magic
tech sky130A
magscale 1 2
timestamp 1665401783
<< metal1 >>
rect 366174 1027828 366180 1027880
rect 366232 1027868 366238 1027880
rect 366542 1027868 366548 1027880
rect 366232 1027840 366548 1027868
rect 366232 1027828 366238 1027840
rect 366542 1027828 366548 1027840
rect 366600 1027828 366606 1027880
rect 366174 1024360 366180 1024412
rect 366232 1024400 366238 1024412
rect 366542 1024400 366548 1024412
rect 366232 1024372 366548 1024400
rect 366232 1024360 366238 1024372
rect 366542 1024360 366548 1024372
rect 366600 1024360 366606 1024412
rect 505002 1007156 505008 1007208
rect 505060 1007196 505066 1007208
rect 513834 1007196 513840 1007208
rect 505060 1007168 513840 1007196
rect 505060 1007156 505066 1007168
rect 513834 1007156 513840 1007168
rect 513892 1007156 513898 1007208
rect 357710 1007088 357716 1007140
rect 357768 1007128 357774 1007140
rect 368934 1007128 368940 1007140
rect 357768 1007100 368940 1007128
rect 357768 1007088 357774 1007100
rect 368934 1007088 368940 1007100
rect 368992 1007088 368998 1007140
rect 505370 1007020 505376 1007072
rect 505428 1007060 505434 1007072
rect 515582 1007060 515588 1007072
rect 505428 1007032 515588 1007060
rect 505428 1007020 505434 1007032
rect 515582 1007020 515588 1007032
rect 515640 1007020 515646 1007072
rect 373258 1006992 373264 1007004
rect 364306 1006964 373264 1006992
rect 357710 1006884 357716 1006936
rect 357768 1006924 357774 1006936
rect 364306 1006924 364334 1006964
rect 373258 1006952 373264 1006964
rect 373316 1006952 373322 1007004
rect 425514 1006952 425520 1007004
rect 425572 1006992 425578 1007004
rect 439682 1006992 439688 1007004
rect 425572 1006964 439688 1006992
rect 425572 1006952 425578 1006964
rect 439682 1006952 439688 1006964
rect 439740 1006952 439746 1007004
rect 520918 1006992 520924 1007004
rect 518866 1006964 520924 1006992
rect 357768 1006896 364334 1006924
rect 357768 1006884 357774 1006896
rect 503346 1006884 503352 1006936
rect 503404 1006924 503410 1006936
rect 518866 1006924 518894 1006964
rect 520918 1006952 520924 1006964
rect 520976 1006952 520982 1007004
rect 551094 1006952 551100 1007004
rect 551152 1006992 551158 1007004
rect 569218 1006992 569224 1007004
rect 551152 1006964 569224 1006992
rect 551152 1006952 551158 1006964
rect 569218 1006952 569224 1006964
rect 569276 1006952 569282 1007004
rect 503404 1006896 518894 1006924
rect 503404 1006884 503410 1006896
rect 427538 1006816 427544 1006868
rect 427596 1006856 427602 1006868
rect 438118 1006856 438124 1006868
rect 427596 1006828 438124 1006856
rect 427596 1006816 427602 1006828
rect 438118 1006816 438124 1006828
rect 438176 1006816 438182 1006868
rect 554130 1006816 554136 1006868
rect 554188 1006856 554194 1006868
rect 559650 1006856 559656 1006868
rect 554188 1006828 559656 1006856
rect 554188 1006816 554194 1006828
rect 559650 1006816 559656 1006828
rect 559708 1006816 559714 1006868
rect 358538 1006748 358544 1006800
rect 358596 1006788 358602 1006800
rect 369118 1006788 369124 1006800
rect 358596 1006760 369124 1006788
rect 358596 1006748 358602 1006760
rect 369118 1006748 369124 1006760
rect 369176 1006748 369182 1006800
rect 400858 1006680 400864 1006732
rect 400916 1006720 400922 1006732
rect 430850 1006720 430856 1006732
rect 400916 1006692 430856 1006720
rect 400916 1006680 400922 1006692
rect 430850 1006680 430856 1006692
rect 430908 1006680 430914 1006732
rect 555970 1006680 555976 1006732
rect 556028 1006720 556034 1006732
rect 566458 1006720 566464 1006732
rect 556028 1006692 566464 1006720
rect 556028 1006680 556034 1006692
rect 566458 1006680 566464 1006692
rect 566516 1006680 566522 1006732
rect 506198 1006612 506204 1006664
rect 506256 1006652 506262 1006664
rect 514018 1006652 514024 1006664
rect 506256 1006624 514024 1006652
rect 506256 1006612 506262 1006624
rect 514018 1006612 514024 1006624
rect 514076 1006612 514082 1006664
rect 94682 1006544 94688 1006596
rect 94740 1006584 94746 1006596
rect 103146 1006584 103152 1006596
rect 94740 1006556 103152 1006584
rect 94740 1006544 94746 1006556
rect 103146 1006544 103152 1006556
rect 103204 1006544 103210 1006596
rect 145558 1006544 145564 1006596
rect 145616 1006584 145622 1006596
rect 153746 1006584 153752 1006596
rect 145616 1006556 153752 1006584
rect 145616 1006544 145622 1006556
rect 153746 1006544 153752 1006556
rect 153804 1006544 153810 1006596
rect 298830 1006544 298836 1006596
rect 298888 1006584 298894 1006596
rect 306926 1006584 306932 1006596
rect 298888 1006556 306932 1006584
rect 298888 1006544 298894 1006556
rect 306926 1006544 306932 1006556
rect 306984 1006544 306990 1006596
rect 429194 1006544 429200 1006596
rect 429252 1006584 429258 1006596
rect 471238 1006584 471244 1006596
rect 429252 1006556 471244 1006584
rect 429252 1006544 429258 1006556
rect 471238 1006544 471244 1006556
rect 471296 1006544 471302 1006596
rect 505370 1006476 505376 1006528
rect 505428 1006516 505434 1006528
rect 516778 1006516 516784 1006528
rect 505428 1006488 516784 1006516
rect 505428 1006476 505434 1006488
rect 516778 1006476 516784 1006488
rect 516836 1006476 516842 1006528
rect 102778 1006408 102784 1006460
rect 102836 1006448 102842 1006460
rect 103974 1006448 103980 1006460
rect 102836 1006420 103980 1006448
rect 102836 1006408 102842 1006420
rect 103974 1006408 103980 1006420
rect 104032 1006408 104038 1006460
rect 145742 1006408 145748 1006460
rect 145800 1006448 145806 1006460
rect 152918 1006448 152924 1006460
rect 145800 1006420 152924 1006448
rect 145800 1006408 145806 1006420
rect 152918 1006408 152924 1006420
rect 152976 1006408 152982 1006460
rect 300302 1006408 300308 1006460
rect 300360 1006448 300366 1006460
rect 307754 1006448 307760 1006460
rect 300360 1006420 307760 1006448
rect 300360 1006408 300366 1006420
rect 307754 1006408 307760 1006420
rect 307812 1006408 307818 1006460
rect 360194 1006408 360200 1006460
rect 360252 1006448 360258 1006460
rect 376018 1006448 376024 1006460
rect 360252 1006420 376024 1006448
rect 360252 1006408 360258 1006420
rect 376018 1006408 376024 1006420
rect 376076 1006408 376082 1006460
rect 553118 1006408 553124 1006460
rect 553176 1006448 553182 1006460
rect 553176 1006420 562364 1006448
rect 553176 1006408 553182 1006420
rect 210418 1006340 210424 1006392
rect 210476 1006380 210482 1006392
rect 228358 1006380 228364 1006392
rect 210476 1006352 228364 1006380
rect 210476 1006340 210482 1006352
rect 228358 1006340 228364 1006352
rect 228416 1006340 228422 1006392
rect 93118 1006272 93124 1006324
rect 93176 1006312 93182 1006324
rect 100294 1006312 100300 1006324
rect 93176 1006284 100300 1006312
rect 93176 1006272 93182 1006284
rect 100294 1006272 100300 1006284
rect 100352 1006272 100358 1006324
rect 144270 1006272 144276 1006324
rect 144328 1006312 144334 1006324
rect 152090 1006312 152096 1006324
rect 144328 1006284 152096 1006312
rect 144328 1006272 144334 1006284
rect 152090 1006272 152096 1006284
rect 152148 1006272 152154 1006324
rect 158254 1006272 158260 1006324
rect 158312 1006312 158318 1006324
rect 175918 1006312 175924 1006324
rect 158312 1006284 175924 1006312
rect 158312 1006272 158318 1006284
rect 175918 1006272 175924 1006284
rect 175976 1006272 175982 1006324
rect 249058 1006272 249064 1006324
rect 249116 1006312 249122 1006324
rect 256142 1006312 256148 1006324
rect 249116 1006284 256148 1006312
rect 249116 1006272 249122 1006284
rect 256142 1006272 256148 1006284
rect 256200 1006272 256206 1006324
rect 299290 1006272 299296 1006324
rect 299348 1006312 299354 1006324
rect 311802 1006312 311808 1006324
rect 299348 1006284 311808 1006312
rect 299348 1006272 299354 1006284
rect 311802 1006272 311808 1006284
rect 311860 1006272 311866 1006324
rect 314654 1006272 314660 1006324
rect 314712 1006312 314718 1006324
rect 319438 1006312 319444 1006324
rect 314712 1006284 319444 1006312
rect 314712 1006272 314718 1006284
rect 319438 1006272 319444 1006284
rect 319496 1006272 319502 1006324
rect 360562 1006272 360568 1006324
rect 360620 1006312 360626 1006324
rect 360620 1006284 365484 1006312
rect 360620 1006272 360626 1006284
rect 208394 1006204 208400 1006256
rect 208452 1006244 208458 1006256
rect 208452 1006216 214604 1006244
rect 208452 1006204 208458 1006216
rect 94498 1006136 94504 1006188
rect 94556 1006176 94562 1006188
rect 101950 1006176 101956 1006188
rect 94556 1006148 101956 1006176
rect 94556 1006136 94562 1006148
rect 101950 1006136 101956 1006148
rect 102008 1006136 102014 1006188
rect 106826 1006136 106832 1006188
rect 106884 1006176 106890 1006188
rect 124858 1006176 124864 1006188
rect 106884 1006148 124864 1006176
rect 106884 1006136 106890 1006148
rect 124858 1006136 124864 1006148
rect 124916 1006136 124922 1006188
rect 144454 1006136 144460 1006188
rect 144512 1006176 144518 1006188
rect 159450 1006176 159456 1006188
rect 144512 1006148 159456 1006176
rect 144512 1006136 144518 1006148
rect 159450 1006136 159456 1006148
rect 159508 1006136 159514 1006188
rect 160278 1006136 160284 1006188
rect 160336 1006176 160342 1006188
rect 164878 1006176 164884 1006188
rect 160336 1006148 164884 1006176
rect 160336 1006136 160342 1006148
rect 164878 1006136 164884 1006148
rect 164936 1006136 164942 1006188
rect 214576 1006108 214604 1006216
rect 247034 1006136 247040 1006188
rect 247092 1006176 247098 1006188
rect 252462 1006176 252468 1006188
rect 247092 1006148 252468 1006176
rect 247092 1006136 247098 1006148
rect 252462 1006136 252468 1006148
rect 252520 1006136 252526 1006188
rect 262674 1006136 262680 1006188
rect 262732 1006176 262738 1006188
rect 278038 1006176 278044 1006188
rect 262732 1006148 278044 1006176
rect 262732 1006136 262738 1006148
rect 278038 1006136 278044 1006148
rect 278096 1006136 278102 1006188
rect 300118 1006136 300124 1006188
rect 300176 1006176 300182 1006188
rect 306098 1006176 306104 1006188
rect 300176 1006148 306104 1006176
rect 300176 1006136 300182 1006148
rect 306098 1006136 306104 1006148
rect 306156 1006136 306162 1006188
rect 365254 1006176 365260 1006188
rect 364720 1006148 365260 1006176
rect 214576 1006080 219434 1006108
rect 93302 1006000 93308 1006052
rect 93360 1006040 93366 1006052
rect 98270 1006040 98276 1006052
rect 93360 1006012 98276 1006040
rect 93360 1006000 93366 1006012
rect 98270 1006000 98276 1006012
rect 98328 1006000 98334 1006052
rect 101398 1006000 101404 1006052
rect 101456 1006040 101462 1006052
rect 103974 1006040 103980 1006052
rect 101456 1006012 103980 1006040
rect 101456 1006000 101462 1006012
rect 103974 1006000 103980 1006012
rect 104032 1006000 104038 1006052
rect 107654 1006000 107660 1006052
rect 107712 1006040 107718 1006052
rect 126238 1006040 126244 1006052
rect 107712 1006012 126244 1006040
rect 107712 1006000 107718 1006012
rect 126238 1006000 126244 1006012
rect 126296 1006000 126302 1006052
rect 148870 1006000 148876 1006052
rect 148928 1006040 148934 1006052
rect 150066 1006040 150072 1006052
rect 148928 1006012 150072 1006040
rect 148928 1006000 148934 1006012
rect 150066 1006000 150072 1006012
rect 150124 1006000 150130 1006052
rect 152642 1006000 152648 1006052
rect 152700 1006040 152706 1006052
rect 155770 1006040 155776 1006052
rect 152700 1006012 155776 1006040
rect 152700 1006000 152706 1006012
rect 155770 1006000 155776 1006012
rect 155828 1006000 155834 1006052
rect 158622 1006000 158628 1006052
rect 158680 1006040 158686 1006052
rect 177298 1006040 177304 1006052
rect 158680 1006012 177304 1006040
rect 158680 1006000 158686 1006012
rect 177298 1006000 177304 1006012
rect 177356 1006000 177362 1006052
rect 198642 1006000 198648 1006052
rect 198700 1006040 198706 1006052
rect 201034 1006040 201040 1006052
rect 198700 1006012 201040 1006040
rect 198700 1006000 198706 1006012
rect 201034 1006000 201040 1006012
rect 201092 1006000 201098 1006052
rect 219406 1006040 219434 1006080
rect 229738 1006040 229744 1006052
rect 219406 1006012 229744 1006040
rect 229738 1006000 229744 1006012
rect 229796 1006000 229802 1006052
rect 249794 1006000 249800 1006052
rect 249852 1006040 249858 1006052
rect 254118 1006040 254124 1006052
rect 249852 1006012 254124 1006040
rect 249852 1006000 249858 1006012
rect 254118 1006000 254124 1006012
rect 254176 1006000 254182 1006052
rect 261846 1006000 261852 1006052
rect 261904 1006040 261910 1006052
rect 280798 1006040 280804 1006052
rect 261904 1006012 280804 1006040
rect 261904 1006000 261910 1006012
rect 280798 1006000 280804 1006012
rect 280856 1006000 280862 1006052
rect 302142 1006000 302148 1006052
rect 302200 1006040 302206 1006052
rect 304074 1006040 304080 1006052
rect 302200 1006012 304080 1006040
rect 302200 1006000 302206 1006012
rect 304074 1006000 304080 1006012
rect 304132 1006000 304138 1006052
rect 314654 1006000 314660 1006052
rect 314712 1006040 314718 1006052
rect 323578 1006040 323584 1006052
rect 314712 1006012 323584 1006040
rect 314712 1006000 314718 1006012
rect 323578 1006000 323584 1006012
rect 323636 1006000 323642 1006052
rect 354582 1006000 354588 1006052
rect 354640 1006040 354646 1006052
rect 354858 1006040 354864 1006052
rect 354640 1006012 354864 1006040
rect 354640 1006000 354646 1006012
rect 354858 1006000 354864 1006012
rect 354916 1006000 354922 1006052
rect 355686 1006000 355692 1006052
rect 355744 1006040 355750 1006052
rect 359550 1006040 359556 1006052
rect 355744 1006012 359556 1006040
rect 355744 1006000 355750 1006012
rect 359550 1006000 359556 1006012
rect 359608 1006000 359614 1006052
rect 361390 1006000 361396 1006052
rect 361448 1006040 361454 1006052
rect 364720 1006040 364748 1006148
rect 365254 1006136 365260 1006148
rect 365312 1006136 365318 1006188
rect 365456 1006176 365484 1006284
rect 369118 1006272 369124 1006324
rect 369176 1006312 369182 1006324
rect 374638 1006312 374644 1006324
rect 369176 1006284 374644 1006312
rect 369176 1006272 369182 1006284
rect 374638 1006272 374644 1006284
rect 374696 1006272 374702 1006324
rect 425146 1006272 425152 1006324
rect 425204 1006312 425210 1006324
rect 443638 1006312 443644 1006324
rect 425204 1006284 443644 1006312
rect 425204 1006272 425210 1006284
rect 443638 1006272 443644 1006284
rect 443696 1006272 443702 1006324
rect 502150 1006272 502156 1006324
rect 502208 1006312 502214 1006324
rect 518158 1006312 518164 1006324
rect 502208 1006284 518164 1006312
rect 502208 1006272 502214 1006284
rect 518158 1006272 518164 1006284
rect 518216 1006272 518222 1006324
rect 556798 1006272 556804 1006324
rect 556856 1006312 556862 1006324
rect 560202 1006312 560208 1006324
rect 556856 1006284 560208 1006312
rect 556856 1006272 556862 1006284
rect 560202 1006272 560208 1006284
rect 560260 1006272 560266 1006324
rect 562336 1006312 562364 1006420
rect 571978 1006312 571984 1006324
rect 562336 1006284 571984 1006312
rect 571978 1006272 571984 1006284
rect 572036 1006272 572042 1006324
rect 371878 1006176 371884 1006188
rect 365456 1006148 371884 1006176
rect 371878 1006136 371884 1006148
rect 371936 1006136 371942 1006188
rect 422018 1006136 422024 1006188
rect 422076 1006176 422082 1006188
rect 423490 1006176 423496 1006188
rect 422076 1006148 423496 1006176
rect 422076 1006136 422082 1006148
rect 423490 1006136 423496 1006148
rect 423548 1006136 423554 1006188
rect 508222 1006136 508228 1006188
rect 508280 1006176 508286 1006188
rect 522298 1006176 522304 1006188
rect 508280 1006148 522304 1006176
rect 508280 1006136 508286 1006148
rect 522298 1006136 522304 1006148
rect 522356 1006136 522362 1006188
rect 557166 1006136 557172 1006188
rect 557224 1006176 557230 1006188
rect 557224 1006148 562364 1006176
rect 557224 1006136 557230 1006148
rect 361448 1006012 364748 1006040
rect 361448 1006000 361454 1006012
rect 365070 1006000 365076 1006052
rect 365128 1006040 365134 1006052
rect 367738 1006040 367744 1006052
rect 365128 1006012 367744 1006040
rect 365128 1006000 365134 1006012
rect 367738 1006000 367744 1006012
rect 367796 1006000 367802 1006052
rect 368934 1006000 368940 1006052
rect 368992 1006040 368998 1006052
rect 378134 1006040 378140 1006052
rect 368992 1006012 378140 1006040
rect 368992 1006000 368998 1006012
rect 378134 1006000 378140 1006012
rect 378192 1006000 378198 1006052
rect 422662 1006000 422668 1006052
rect 422720 1006040 422726 1006052
rect 429838 1006040 429844 1006052
rect 422720 1006012 429844 1006040
rect 422720 1006000 422726 1006012
rect 429838 1006000 429844 1006012
rect 429896 1006000 429902 1006052
rect 430022 1006000 430028 1006052
rect 430080 1006040 430086 1006052
rect 471422 1006040 471428 1006052
rect 430080 1006012 471428 1006040
rect 430080 1006000 430086 1006012
rect 471422 1006000 471428 1006012
rect 471480 1006000 471486 1006052
rect 497918 1006000 497924 1006052
rect 497976 1006040 497982 1006052
rect 498838 1006040 498844 1006052
rect 497976 1006012 498844 1006040
rect 497976 1006000 497982 1006012
rect 498838 1006000 498844 1006012
rect 498896 1006000 498902 1006052
rect 501322 1006000 501328 1006052
rect 501380 1006040 501386 1006052
rect 506474 1006040 506480 1006052
rect 501380 1006012 506480 1006040
rect 501380 1006000 501386 1006012
rect 506474 1006000 506480 1006012
rect 506532 1006000 506538 1006052
rect 509050 1006000 509056 1006052
rect 509108 1006040 509114 1006052
rect 509108 1006012 512316 1006040
rect 509108 1006000 509114 1006012
rect 512288 1005904 512316 1006012
rect 514018 1006000 514024 1006052
rect 514076 1006040 514082 1006052
rect 522482 1006040 522488 1006052
rect 514076 1006012 522488 1006040
rect 514076 1006000 514082 1006012
rect 522482 1006000 522488 1006012
rect 522540 1006000 522546 1006052
rect 562336 1006040 562364 1006148
rect 574738 1006040 574744 1006052
rect 562336 1006012 574744 1006040
rect 574738 1006000 574744 1006012
rect 574796 1006000 574802 1006052
rect 515398 1005904 515404 1005916
rect 512288 1005876 515404 1005904
rect 515398 1005864 515404 1005876
rect 515456 1005864 515462 1005916
rect 432046 1005796 432052 1005848
rect 432104 1005836 432110 1005848
rect 433518 1005836 433524 1005848
rect 432104 1005808 433524 1005836
rect 432104 1005796 432110 1005808
rect 433518 1005796 433524 1005808
rect 433576 1005796 433582 1005848
rect 423490 1005660 423496 1005712
rect 423548 1005700 423554 1005712
rect 446398 1005700 446404 1005712
rect 423548 1005672 446404 1005700
rect 423548 1005660 423554 1005672
rect 446398 1005660 446404 1005672
rect 446456 1005660 446462 1005712
rect 560846 1005660 560852 1005712
rect 560904 1005700 560910 1005712
rect 570598 1005700 570604 1005712
rect 560904 1005672 570604 1005700
rect 560904 1005660 560910 1005672
rect 570598 1005660 570604 1005672
rect 570656 1005660 570662 1005712
rect 428366 1005524 428372 1005576
rect 428424 1005564 428430 1005576
rect 460198 1005564 460204 1005576
rect 428424 1005536 460204 1005564
rect 428424 1005524 428430 1005536
rect 460198 1005524 460204 1005536
rect 460256 1005524 460262 1005576
rect 555142 1005524 555148 1005576
rect 555200 1005564 555206 1005576
rect 567838 1005564 567844 1005576
rect 555200 1005536 567844 1005564
rect 555200 1005524 555206 1005536
rect 567838 1005524 567844 1005536
rect 567896 1005524 567902 1005576
rect 436922 1005388 436928 1005440
rect 436980 1005428 436986 1005440
rect 465718 1005428 465724 1005440
rect 436980 1005400 465724 1005428
rect 436980 1005388 436986 1005400
rect 465718 1005388 465724 1005400
rect 465776 1005388 465782 1005440
rect 553946 1005388 553952 1005440
rect 554004 1005428 554010 1005440
rect 573358 1005428 573364 1005440
rect 554004 1005400 573364 1005428
rect 554004 1005388 554010 1005400
rect 573358 1005388 573364 1005400
rect 573416 1005388 573422 1005440
rect 149882 1005320 149888 1005372
rect 149940 1005360 149946 1005372
rect 152918 1005360 152924 1005372
rect 149940 1005332 152924 1005360
rect 149940 1005320 149946 1005332
rect 152918 1005320 152924 1005332
rect 152976 1005320 152982 1005372
rect 427170 1005320 427176 1005372
rect 427228 1005360 427234 1005372
rect 427228 1005332 436784 1005360
rect 427228 1005320 427234 1005332
rect 195698 1005252 195704 1005304
rect 195756 1005292 195762 1005304
rect 202690 1005292 202696 1005304
rect 195756 1005264 202696 1005292
rect 195756 1005252 195762 1005264
rect 202690 1005252 202696 1005264
rect 202748 1005252 202754 1005304
rect 263042 1005252 263048 1005304
rect 263100 1005292 263106 1005304
rect 279418 1005292 279424 1005304
rect 263100 1005264 279424 1005292
rect 263100 1005252 263106 1005264
rect 279418 1005252 279424 1005264
rect 279476 1005252 279482 1005304
rect 360562 1005252 360568 1005304
rect 360620 1005292 360626 1005304
rect 377398 1005292 377404 1005304
rect 360620 1005264 377404 1005292
rect 360620 1005252 360626 1005264
rect 377398 1005252 377404 1005264
rect 377456 1005252 377462 1005304
rect 436756 1005292 436784 1005332
rect 456058 1005292 456064 1005304
rect 436756 1005264 456064 1005292
rect 456058 1005252 456064 1005264
rect 456116 1005252 456122 1005304
rect 552290 1005252 552296 1005304
rect 552348 1005292 552354 1005304
rect 570782 1005292 570788 1005304
rect 552348 1005264 570788 1005292
rect 552348 1005252 552354 1005264
rect 570782 1005252 570788 1005264
rect 570840 1005252 570846 1005304
rect 430850 1005184 430856 1005236
rect 430908 1005224 430914 1005236
rect 431908 1005224 431914 1005236
rect 430908 1005196 431914 1005224
rect 430908 1005184 430914 1005196
rect 431908 1005184 431914 1005196
rect 431966 1005184 431972 1005236
rect 507026 1005184 507032 1005236
rect 507084 1005224 507090 1005236
rect 509970 1005224 509976 1005236
rect 507084 1005196 509976 1005224
rect 507084 1005184 507090 1005196
rect 509970 1005184 509976 1005196
rect 510028 1005184 510034 1005236
rect 432046 1005116 432052 1005168
rect 432104 1005156 432110 1005168
rect 436922 1005156 436928 1005168
rect 432104 1005128 436928 1005156
rect 432104 1005116 432110 1005128
rect 436922 1005116 436928 1005128
rect 436980 1005116 436986 1005168
rect 209222 1005048 209228 1005100
rect 209280 1005088 209286 1005100
rect 211798 1005088 211804 1005100
rect 209280 1005060 211804 1005088
rect 209280 1005048 209286 1005060
rect 211798 1005048 211804 1005060
rect 211856 1005048 211862 1005100
rect 363414 1005048 363420 1005100
rect 363472 1005088 363478 1005100
rect 366358 1005088 366364 1005100
rect 363472 1005060 366364 1005088
rect 363472 1005048 363478 1005060
rect 366358 1005048 366364 1005060
rect 366416 1005048 366422 1005100
rect 508222 1005048 508228 1005100
rect 508280 1005088 508286 1005100
rect 510890 1005088 510896 1005100
rect 508280 1005060 510896 1005088
rect 508280 1005048 508286 1005060
rect 510890 1005048 510896 1005060
rect 510948 1005048 510954 1005100
rect 432414 1004980 432420 1005032
rect 432472 1005020 432478 1005032
rect 434162 1005020 434168 1005032
rect 432472 1004992 434168 1005020
rect 432472 1004980 432478 1004992
rect 434162 1004980 434168 1004992
rect 434220 1004980 434226 1005032
rect 151078 1004912 151084 1004964
rect 151136 1004952 151142 1004964
rect 153746 1004952 153752 1004964
rect 151136 1004924 153752 1004952
rect 151136 1004912 151142 1004924
rect 153746 1004912 153752 1004924
rect 153804 1004912 153810 1004964
rect 154390 1004912 154396 1004964
rect 154448 1004952 154454 1004964
rect 160646 1004952 160652 1004964
rect 154448 1004924 160652 1004952
rect 154448 1004912 154454 1004924
rect 160646 1004912 160652 1004924
rect 160704 1004912 160710 1004964
rect 207566 1004912 207572 1004964
rect 207624 1004952 207630 1004964
rect 209866 1004952 209872 1004964
rect 207624 1004924 209872 1004952
rect 207624 1004912 207630 1004924
rect 209866 1004912 209872 1004924
rect 209924 1004912 209930 1004964
rect 365070 1004912 365076 1004964
rect 365128 1004952 365134 1004964
rect 370498 1004952 370504 1004964
rect 365128 1004924 370504 1004952
rect 365128 1004912 365134 1004924
rect 370498 1004912 370504 1004924
rect 370556 1004912 370562 1004964
rect 429194 1004912 429200 1004964
rect 429252 1004952 429258 1004964
rect 432230 1004952 432236 1004964
rect 429252 1004924 432236 1004952
rect 429252 1004912 429258 1004924
rect 432230 1004912 432236 1004924
rect 432288 1004912 432294 1004964
rect 507854 1004912 507860 1004964
rect 507912 1004952 507918 1004964
rect 509694 1004952 509700 1004964
rect 507912 1004924 509700 1004952
rect 507912 1004912 507918 1004924
rect 509694 1004912 509700 1004924
rect 509752 1004912 509758 1004964
rect 151262 1004776 151268 1004828
rect 151320 1004816 151326 1004828
rect 154114 1004816 154120 1004828
rect 151320 1004788 154120 1004816
rect 151320 1004776 151326 1004788
rect 154114 1004776 154120 1004788
rect 154172 1004776 154178 1004828
rect 159450 1004776 159456 1004828
rect 159508 1004816 159514 1004828
rect 162118 1004816 162124 1004828
rect 159508 1004788 162124 1004816
rect 159508 1004776 159514 1004788
rect 162118 1004776 162124 1004788
rect 162176 1004776 162182 1004828
rect 313826 1004776 313832 1004828
rect 313884 1004816 313890 1004828
rect 316034 1004816 316040 1004828
rect 313884 1004788 316040 1004816
rect 313884 1004776 313890 1004788
rect 316034 1004776 316040 1004788
rect 316092 1004776 316098 1004828
rect 352834 1004776 352840 1004828
rect 352892 1004816 352898 1004828
rect 355686 1004816 355692 1004828
rect 352892 1004788 355692 1004816
rect 352892 1004776 352898 1004788
rect 355686 1004776 355692 1004788
rect 355744 1004776 355750 1004828
rect 362586 1004776 362592 1004828
rect 362644 1004816 362650 1004828
rect 364978 1004816 364984 1004828
rect 362644 1004788 364984 1004816
rect 362644 1004776 362650 1004788
rect 364978 1004776 364984 1004788
rect 365036 1004776 365042 1004828
rect 431678 1004776 431684 1004828
rect 431736 1004816 431742 1004828
rect 431736 1004788 432092 1004816
rect 431736 1004776 431742 1004788
rect 106182 1004640 106188 1004692
rect 106240 1004680 106246 1004692
rect 108482 1004680 108488 1004692
rect 106240 1004652 108488 1004680
rect 106240 1004640 106246 1004652
rect 108482 1004640 108488 1004652
rect 108540 1004640 108546 1004692
rect 149698 1004640 149704 1004692
rect 149756 1004680 149762 1004692
rect 151722 1004680 151728 1004692
rect 149756 1004652 151728 1004680
rect 149756 1004640 149762 1004652
rect 151722 1004640 151728 1004652
rect 151780 1004640 151786 1004692
rect 160646 1004640 160652 1004692
rect 160704 1004680 160710 1004692
rect 162854 1004680 162860 1004692
rect 160704 1004652 162860 1004680
rect 160704 1004640 160710 1004652
rect 162854 1004640 162860 1004652
rect 162912 1004640 162918 1004692
rect 209222 1004640 209228 1004692
rect 209280 1004680 209286 1004692
rect 211154 1004680 211160 1004692
rect 209280 1004652 211160 1004680
rect 209280 1004640 209286 1004652
rect 211154 1004640 211160 1004652
rect 211212 1004640 211218 1004692
rect 212534 1004640 212540 1004692
rect 212592 1004680 212598 1004692
rect 217318 1004680 217324 1004692
rect 212592 1004652 217324 1004680
rect 212592 1004640 212598 1004652
rect 217318 1004640 217324 1004652
rect 217376 1004640 217382 1004692
rect 250438 1004640 250444 1004692
rect 250496 1004680 250502 1004692
rect 256510 1004680 256516 1004692
rect 250496 1004652 256516 1004680
rect 250496 1004640 250502 1004652
rect 256510 1004640 256516 1004652
rect 256568 1004640 256574 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 364242 1004640 364248 1004692
rect 364300 1004680 364306 1004692
rect 366542 1004680 366548 1004692
rect 364300 1004652 366548 1004680
rect 364300 1004640 364306 1004652
rect 366542 1004640 366548 1004652
rect 366600 1004640 366606 1004692
rect 430022 1004640 430028 1004692
rect 430080 1004680 430086 1004692
rect 431862 1004680 431868 1004692
rect 430080 1004652 431868 1004680
rect 430080 1004640 430086 1004652
rect 431862 1004640 431868 1004652
rect 431920 1004640 431926 1004692
rect 432064 1004680 432092 1004788
rect 498102 1004776 498108 1004828
rect 498160 1004816 498166 1004828
rect 499666 1004816 499672 1004828
rect 498160 1004788 499672 1004816
rect 498160 1004776 498166 1004788
rect 499666 1004776 499672 1004788
rect 499724 1004776 499730 1004828
rect 507394 1004776 507400 1004828
rect 507452 1004816 507458 1004828
rect 509234 1004816 509240 1004828
rect 507452 1004788 509240 1004816
rect 507452 1004776 507458 1004788
rect 509234 1004776 509240 1004788
rect 509292 1004776 509298 1004828
rect 555970 1004776 555976 1004828
rect 556028 1004816 556034 1004828
rect 558178 1004816 558184 1004828
rect 556028 1004788 558184 1004816
rect 556028 1004776 556034 1004788
rect 558178 1004776 558184 1004788
rect 558236 1004776 558242 1004828
rect 433978 1004680 433984 1004692
rect 432064 1004652 433984 1004680
rect 433978 1004640 433984 1004652
rect 434036 1004640 434042 1004692
rect 499482 1004640 499488 1004692
rect 499540 1004680 499546 1004692
rect 500494 1004680 500500 1004692
rect 499540 1004652 500500 1004680
rect 499540 1004640 499546 1004652
rect 500494 1004640 500500 1004652
rect 500552 1004640 500558 1004692
rect 509050 1004640 509056 1004692
rect 509108 1004680 509114 1004692
rect 510706 1004680 510712 1004692
rect 509108 1004652 510712 1004680
rect 509108 1004640 509114 1004652
rect 510706 1004640 510712 1004652
rect 510764 1004640 510770 1004692
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559558 1004680 559564 1004692
rect 557684 1004652 559564 1004680
rect 557684 1004640 557690 1004652
rect 559558 1004640 559564 1004652
rect 559616 1004640 559622 1004692
rect 504542 1004436 504548 1004488
rect 504600 1004476 504606 1004488
rect 510154 1004476 510160 1004488
rect 504600 1004448 510160 1004476
rect 504600 1004436 504606 1004448
rect 510154 1004436 510160 1004448
rect 510212 1004436 510218 1004488
rect 356514 1003892 356520 1003944
rect 356572 1003932 356578 1003944
rect 381446 1003932 381452 1003944
rect 356572 1003904 381452 1003932
rect 356572 1003892 356578 1003904
rect 381446 1003892 381452 1003904
rect 381504 1003892 381510 1003944
rect 422018 1003892 422024 1003944
rect 422076 1003932 422082 1003944
rect 469858 1003932 469864 1003944
rect 422076 1003904 469864 1003932
rect 422076 1003892 422082 1003904
rect 469858 1003892 469864 1003904
rect 469916 1003892 469922 1003944
rect 298646 1003280 298652 1003332
rect 298704 1003320 298710 1003332
rect 331122 1003320 331128 1003332
rect 298704 1003292 331128 1003320
rect 298704 1003280 298710 1003292
rect 331122 1003280 331128 1003292
rect 331180 1003280 331186 1003332
rect 354582 1002804 354588 1002856
rect 354640 1002844 354646 1002856
rect 355134 1002844 355140 1002856
rect 354640 1002816 355140 1002844
rect 354640 1002804 354646 1002816
rect 355134 1002804 355140 1002816
rect 355192 1002804 355198 1002856
rect 456058 1002804 456064 1002856
rect 456116 1002844 456122 1002856
rect 462314 1002844 462320 1002856
rect 456116 1002816 462320 1002844
rect 456116 1002804 456122 1002816
rect 462314 1002804 462320 1002816
rect 462372 1002804 462378 1002856
rect 98638 1002736 98644 1002788
rect 98696 1002776 98702 1002788
rect 101950 1002776 101956 1002788
rect 98696 1002748 101956 1002776
rect 98696 1002736 98702 1002748
rect 101950 1002736 101956 1002748
rect 102008 1002736 102014 1002788
rect 252002 1002736 252008 1002788
rect 252060 1002776 252066 1002788
rect 255314 1002776 255320 1002788
rect 252060 1002748 255320 1002776
rect 252060 1002736 252066 1002748
rect 255314 1002736 255320 1002748
rect 255372 1002736 255378 1002788
rect 424686 1002668 424692 1002720
rect 424744 1002708 424750 1002720
rect 449158 1002708 449164 1002720
rect 424744 1002680 449164 1002708
rect 424744 1002668 424750 1002680
rect 449158 1002668 449164 1002680
rect 449216 1002668 449222 1002720
rect 97258 1002600 97264 1002652
rect 97316 1002640 97322 1002652
rect 100294 1002640 100300 1002652
rect 97316 1002612 100300 1002640
rect 97316 1002600 97322 1002612
rect 100294 1002600 100300 1002612
rect 100352 1002600 100358 1002652
rect 157426 1002600 157432 1002652
rect 157484 1002640 157490 1002652
rect 159358 1002640 159364 1002652
rect 157484 1002612 159364 1002640
rect 157484 1002600 157490 1002612
rect 159358 1002600 159364 1002612
rect 159416 1002600 159422 1002652
rect 560202 1002600 560208 1002652
rect 560260 1002640 560266 1002652
rect 567194 1002640 567200 1002652
rect 560260 1002612 567200 1002640
rect 560260 1002600 560266 1002612
rect 567194 1002600 567200 1002612
rect 567252 1002600 567258 1002652
rect 246758 1002532 246764 1002584
rect 246816 1002572 246822 1002584
rect 255314 1002572 255320 1002584
rect 246816 1002544 255320 1002572
rect 246816 1002532 246822 1002544
rect 255314 1002532 255320 1002544
rect 255372 1002532 255378 1002584
rect 426342 1002532 426348 1002584
rect 426400 1002572 426406 1002584
rect 458082 1002572 458088 1002584
rect 426400 1002544 458088 1002572
rect 426400 1002532 426406 1002544
rect 458082 1002532 458088 1002544
rect 458140 1002532 458146 1002584
rect 98822 1002464 98828 1002516
rect 98880 1002504 98886 1002516
rect 101122 1002504 101128 1002516
rect 98880 1002476 101128 1002504
rect 98880 1002464 98886 1002476
rect 101122 1002464 101128 1002476
rect 101180 1002464 101186 1002516
rect 105998 1002464 106004 1002516
rect 106056 1002504 106062 1002516
rect 109494 1002504 109500 1002516
rect 106056 1002476 109500 1002504
rect 106056 1002464 106062 1002476
rect 109494 1002464 109500 1002476
rect 109552 1002464 109558 1002516
rect 158622 1002464 158628 1002516
rect 158680 1002504 158686 1002516
rect 160186 1002504 160192 1002516
rect 158680 1002476 160192 1002504
rect 158680 1002464 158686 1002476
rect 160186 1002464 160192 1002476
rect 160244 1002464 160250 1002516
rect 261018 1002464 261024 1002516
rect 261076 1002504 261082 1002516
rect 264238 1002504 264244 1002516
rect 261076 1002476 264244 1002504
rect 261076 1002464 261082 1002476
rect 264238 1002464 264244 1002476
rect 264296 1002464 264302 1002516
rect 501690 1002464 501696 1002516
rect 501748 1002504 501754 1002516
rect 504358 1002504 504364 1002516
rect 501748 1002476 504364 1002504
rect 501748 1002464 501754 1002476
rect 504358 1002464 504364 1002476
rect 504416 1002464 504422 1002516
rect 558822 1002464 558828 1002516
rect 558880 1002504 558886 1002516
rect 562318 1002504 562324 1002516
rect 558880 1002476 562324 1002504
rect 558880 1002464 558886 1002476
rect 562318 1002464 562324 1002476
rect 562376 1002464 562382 1002516
rect 96522 1002328 96528 1002380
rect 96580 1002368 96586 1002380
rect 99098 1002368 99104 1002380
rect 96580 1002340 99104 1002368
rect 96580 1002328 96586 1002340
rect 99098 1002328 99104 1002340
rect 99156 1002328 99162 1002380
rect 105630 1002328 105636 1002380
rect 105688 1002368 105694 1002380
rect 107746 1002368 107752 1002380
rect 105688 1002340 107752 1002368
rect 105688 1002328 105694 1002340
rect 107746 1002328 107752 1002340
rect 107804 1002328 107810 1002380
rect 108022 1002328 108028 1002380
rect 108080 1002368 108086 1002380
rect 110414 1002368 110420 1002380
rect 108080 1002340 110420 1002368
rect 108080 1002328 108086 1002340
rect 110414 1002328 110420 1002340
rect 110472 1002328 110478 1002380
rect 144730 1002328 144736 1002380
rect 144788 1002368 144794 1002380
rect 150894 1002368 150900 1002380
rect 144788 1002340 150900 1002368
rect 144788 1002328 144794 1002340
rect 150894 1002328 150900 1002340
rect 150952 1002328 150958 1002380
rect 156598 1002328 156604 1002380
rect 156656 1002368 156662 1002380
rect 158714 1002368 158720 1002380
rect 156656 1002340 158720 1002368
rect 156656 1002328 156662 1002340
rect 158714 1002328 158720 1002340
rect 158772 1002328 158778 1002380
rect 211246 1002328 211252 1002380
rect 211304 1002368 211310 1002380
rect 215938 1002368 215944 1002380
rect 211304 1002340 215944 1002368
rect 211304 1002328 211310 1002340
rect 215938 1002328 215944 1002340
rect 215996 1002328 216002 1002380
rect 500218 1002328 500224 1002380
rect 500276 1002368 500282 1002380
rect 502150 1002368 502156 1002380
rect 500276 1002340 502156 1002368
rect 500276 1002328 500282 1002340
rect 502150 1002328 502156 1002340
rect 502208 1002328 502214 1002380
rect 557994 1002328 558000 1002380
rect 558052 1002368 558058 1002380
rect 560294 1002368 560300 1002380
rect 558052 1002340 560300 1002368
rect 558052 1002328 558058 1002340
rect 560294 1002328 560300 1002340
rect 560352 1002328 560358 1002380
rect 560478 1002328 560484 1002380
rect 560536 1002368 560542 1002380
rect 563054 1002368 563060 1002380
rect 560536 1002340 563060 1002368
rect 560536 1002328 560542 1002340
rect 563054 1002328 563060 1002340
rect 563112 1002328 563118 1002380
rect 99006 1002192 99012 1002244
rect 99064 1002232 99070 1002244
rect 101122 1002232 101128 1002244
rect 99064 1002204 101128 1002232
rect 99064 1002192 99070 1002204
rect 101122 1002192 101128 1002204
rect 101180 1002192 101186 1002244
rect 104802 1002192 104808 1002244
rect 104860 1002232 104866 1002244
rect 106458 1002232 106464 1002244
rect 104860 1002204 106464 1002232
rect 104860 1002192 104866 1002204
rect 106458 1002192 106464 1002204
rect 106516 1002192 106522 1002244
rect 108482 1002192 108488 1002244
rect 108540 1002232 108546 1002244
rect 111058 1002232 111064 1002244
rect 108540 1002204 111064 1002232
rect 108540 1002192 108546 1002204
rect 111058 1002192 111064 1002204
rect 111116 1002192 111122 1002244
rect 148318 1002192 148324 1002244
rect 148376 1002232 148382 1002244
rect 151722 1002232 151728 1002244
rect 148376 1002204 151728 1002232
rect 148376 1002192 148382 1002204
rect 151722 1002192 151728 1002204
rect 151780 1002192 151786 1002244
rect 155770 1002192 155776 1002244
rect 155828 1002232 155834 1002244
rect 157334 1002232 157340 1002244
rect 155828 1002204 157340 1002232
rect 155828 1002192 155834 1002204
rect 157334 1002192 157340 1002204
rect 157392 1002192 157398 1002244
rect 203334 1002192 203340 1002244
rect 203392 1002232 203398 1002244
rect 206370 1002232 206376 1002244
rect 203392 1002204 206376 1002232
rect 203392 1002192 203398 1002204
rect 206370 1002192 206376 1002204
rect 206428 1002192 206434 1002244
rect 210050 1002192 210056 1002244
rect 210108 1002232 210114 1002244
rect 212534 1002232 212540 1002244
rect 210108 1002204 212540 1002232
rect 210108 1002192 210114 1002204
rect 212534 1002192 212540 1002204
rect 212592 1002192 212598 1002244
rect 251818 1002192 251824 1002244
rect 251876 1002232 251882 1002244
rect 254486 1002232 254492 1002244
rect 251876 1002204 254492 1002232
rect 251876 1002192 251882 1002204
rect 254486 1002192 254492 1002204
rect 254544 1002192 254550 1002244
rect 427998 1002192 428004 1002244
rect 428056 1002232 428062 1002244
rect 431126 1002232 431132 1002244
rect 428056 1002204 431132 1002232
rect 428056 1002192 428062 1002204
rect 431126 1002192 431132 1002204
rect 431184 1002192 431190 1002244
rect 500494 1002192 500500 1002244
rect 500552 1002232 500558 1002244
rect 502978 1002232 502984 1002244
rect 500552 1002204 502984 1002232
rect 500552 1002192 500558 1002204
rect 502978 1002192 502984 1002204
rect 503036 1002192 503042 1002244
rect 509878 1002192 509884 1002244
rect 509936 1002232 509942 1002244
rect 512638 1002232 512644 1002244
rect 509936 1002204 512644 1002232
rect 509936 1002192 509942 1002204
rect 512638 1002192 512644 1002204
rect 512696 1002192 512702 1002244
rect 553118 1002192 553124 1002244
rect 553176 1002232 553182 1002244
rect 554314 1002232 554320 1002244
rect 553176 1002204 554320 1002232
rect 553176 1002192 553182 1002204
rect 554314 1002192 554320 1002204
rect 554372 1002192 554378 1002244
rect 560018 1002192 560024 1002244
rect 560076 1002232 560082 1002244
rect 562502 1002232 562508 1002244
rect 560076 1002204 562508 1002232
rect 560076 1002192 560082 1002204
rect 562502 1002192 562508 1002204
rect 562560 1002192 562566 1002244
rect 97442 1002056 97448 1002108
rect 97500 1002096 97506 1002108
rect 99466 1002096 99472 1002108
rect 97500 1002068 99472 1002096
rect 97500 1002056 97506 1002068
rect 99466 1002056 99472 1002068
rect 99524 1002056 99530 1002108
rect 100018 1002056 100024 1002108
rect 100076 1002096 100082 1002108
rect 103146 1002096 103152 1002108
rect 100076 1002068 103152 1002096
rect 100076 1002056 100082 1002068
rect 103146 1002056 103152 1002068
rect 103204 1002056 103210 1002108
rect 106826 1002056 106832 1002108
rect 106884 1002096 106890 1002108
rect 109034 1002096 109040 1002108
rect 106884 1002068 109040 1002096
rect 106884 1002056 106890 1002068
rect 109034 1002056 109040 1002068
rect 109092 1002056 109098 1002108
rect 109678 1002056 109684 1002108
rect 109736 1002096 109742 1002108
rect 111886 1002096 111892 1002108
rect 109736 1002068 111892 1002096
rect 109736 1002056 109742 1002068
rect 111886 1002056 111892 1002068
rect 111944 1002056 111950 1002108
rect 148962 1002056 148968 1002108
rect 149020 1002096 149026 1002108
rect 150894 1002096 150900 1002108
rect 149020 1002068 150900 1002096
rect 149020 1002056 149026 1002068
rect 150894 1002056 150900 1002068
rect 150952 1002056 150958 1002108
rect 155218 1002056 155224 1002108
rect 155276 1002096 155282 1002108
rect 156598 1002096 156604 1002108
rect 155276 1002068 156604 1002096
rect 155276 1002056 155282 1002068
rect 156598 1002056 156604 1002068
rect 156656 1002056 156662 1002108
rect 203702 1002056 203708 1002108
rect 203760 1002096 203766 1002108
rect 205542 1002096 205548 1002108
rect 203760 1002068 205548 1002096
rect 203760 1002056 203766 1002068
rect 205542 1002056 205548 1002068
rect 205600 1002056 205606 1002108
rect 211246 1002056 211252 1002108
rect 211304 1002096 211310 1002108
rect 213178 1002096 213184 1002108
rect 211304 1002068 213184 1002096
rect 211304 1002056 211310 1002068
rect 213178 1002056 213184 1002068
rect 213236 1002056 213242 1002108
rect 253474 1002056 253480 1002108
rect 253532 1002096 253538 1002108
rect 256142 1002096 256148 1002108
rect 253532 1002068 256148 1002096
rect 253532 1002056 253538 1002068
rect 256142 1002056 256148 1002068
rect 256200 1002056 256206 1002108
rect 263502 1002056 263508 1002108
rect 263560 1002096 263566 1002108
rect 265618 1002096 265624 1002108
rect 263560 1002068 265624 1002096
rect 263560 1002056 263566 1002068
rect 265618 1002056 265624 1002068
rect 265676 1002056 265682 1002108
rect 310974 1002056 310980 1002108
rect 311032 1002096 311038 1002108
rect 313274 1002096 313280 1002108
rect 311032 1002068 313280 1002096
rect 311032 1002056 311038 1002068
rect 313274 1002056 313280 1002068
rect 313332 1002056 313338 1002108
rect 355778 1002056 355784 1002108
rect 355836 1002096 355842 1002108
rect 358538 1002096 358544 1002108
rect 355836 1002068 358544 1002096
rect 355836 1002056 355842 1002068
rect 358538 1002056 358544 1002068
rect 358596 1002056 358602 1002108
rect 359734 1002056 359740 1002108
rect 359792 1002096 359798 1002108
rect 362218 1002096 362224 1002108
rect 359792 1002068 362224 1002096
rect 359792 1002056 359798 1002068
rect 362218 1002056 362224 1002068
rect 362276 1002056 362282 1002108
rect 423582 1002056 423588 1002108
rect 423640 1002096 423646 1002108
rect 425146 1002096 425152 1002108
rect 423640 1002068 425152 1002096
rect 423640 1002056 423646 1002068
rect 425146 1002056 425152 1002068
rect 425204 1002056 425210 1002108
rect 428366 1002056 428372 1002108
rect 428424 1002096 428430 1002108
rect 431310 1002096 431316 1002108
rect 428424 1002068 431316 1002096
rect 428424 1002056 428430 1002068
rect 431310 1002056 431316 1002068
rect 431368 1002056 431374 1002108
rect 433334 1002056 433340 1002108
rect 433392 1002096 433398 1002108
rect 435358 1002096 435364 1002108
rect 433392 1002068 435364 1002096
rect 433392 1002056 433398 1002068
rect 435358 1002056 435364 1002068
rect 435416 1002056 435422 1002108
rect 500678 1002056 500684 1002108
rect 500736 1002096 500742 1002108
rect 502518 1002096 502524 1002108
rect 500736 1002068 502524 1002096
rect 500736 1002056 500742 1002068
rect 502518 1002056 502524 1002068
rect 502576 1002056 502582 1002108
rect 510338 1002056 510344 1002108
rect 510396 1002096 510402 1002108
rect 512822 1002096 512828 1002108
rect 510396 1002068 512828 1002096
rect 510396 1002056 510402 1002068
rect 512822 1002056 512828 1002068
rect 512880 1002056 512886 1002108
rect 555142 1002056 555148 1002108
rect 555200 1002096 555206 1002108
rect 556798 1002096 556804 1002108
rect 555200 1002068 556804 1002096
rect 555200 1002056 555206 1002068
rect 556798 1002056 556804 1002068
rect 556856 1002056 556862 1002108
rect 557994 1002056 558000 1002108
rect 558052 1002096 558058 1002108
rect 560662 1002096 560668 1002108
rect 558052 1002068 560668 1002096
rect 558052 1002056 558058 1002068
rect 560662 1002056 560668 1002068
rect 560720 1002056 560726 1002108
rect 560846 1002056 560852 1002108
rect 560904 1002096 560910 1002108
rect 563698 1002096 563704 1002108
rect 560904 1002068 563704 1002096
rect 560904 1002056 560910 1002068
rect 563698 1002056 563704 1002068
rect 563756 1002056 563762 1002108
rect 152458 1001988 152464 1002040
rect 152516 1002028 152522 1002040
rect 154574 1002028 154580 1002040
rect 152516 1002000 154580 1002028
rect 152516 1001988 152522 1002000
rect 154574 1001988 154580 1002000
rect 154632 1001988 154638 1002040
rect 96338 1001920 96344 1001972
rect 96396 1001960 96402 1001972
rect 98270 1001960 98276 1001972
rect 96396 1001932 98276 1001960
rect 96396 1001920 96402 1001932
rect 98270 1001920 98276 1001932
rect 98328 1001920 98334 1001972
rect 100202 1001920 100208 1001972
rect 100260 1001960 100266 1001972
rect 102318 1001960 102324 1001972
rect 100260 1001932 102324 1001960
rect 100260 1001920 100266 1001932
rect 102318 1001920 102324 1001932
rect 102376 1001920 102382 1001972
rect 105998 1001920 106004 1001972
rect 106056 1001960 106062 1001972
rect 108114 1001960 108120 1001972
rect 106056 1001932 108120 1001960
rect 106056 1001920 106062 1001932
rect 108114 1001920 108120 1001932
rect 108172 1001920 108178 1001972
rect 108850 1001920 108856 1001972
rect 108908 1001960 108914 1001972
rect 112070 1001960 112076 1001972
rect 108908 1001932 112076 1001960
rect 108908 1001920 108914 1001932
rect 112070 1001920 112076 1001932
rect 112128 1001920 112134 1001972
rect 147582 1001920 147588 1001972
rect 147640 1001960 147646 1001972
rect 149238 1001960 149244 1001972
rect 147640 1001932 149244 1001960
rect 147640 1001920 147646 1001932
rect 149238 1001920 149244 1001932
rect 149296 1001920 149302 1001972
rect 154942 1001920 154948 1001972
rect 155000 1001960 155006 1001972
rect 155954 1001960 155960 1001972
rect 155000 1001932 155960 1001960
rect 155000 1001920 155006 1001932
rect 155954 1001920 155960 1001932
rect 156012 1001920 156018 1001972
rect 157794 1001920 157800 1001972
rect 157852 1001960 157858 1001972
rect 160370 1001960 160376 1001972
rect 157852 1001932 160376 1001960
rect 157852 1001920 157858 1001932
rect 160370 1001920 160376 1001932
rect 160428 1001920 160434 1001972
rect 195146 1001920 195152 1001972
rect 195204 1001960 195210 1001972
rect 198642 1001960 198648 1001972
rect 195204 1001932 198648 1001960
rect 195204 1001920 195210 1001932
rect 198642 1001920 198648 1001932
rect 198700 1001920 198706 1001972
rect 204898 1001920 204904 1001972
rect 204956 1001960 204962 1001972
rect 206738 1001960 206744 1001972
rect 204956 1001932 206744 1001960
rect 204956 1001920 204962 1001932
rect 206738 1001920 206744 1001932
rect 206796 1001920 206802 1001972
rect 212074 1001920 212080 1001972
rect 212132 1001960 212138 1001972
rect 213914 1001960 213920 1001972
rect 212132 1001932 213920 1001960
rect 212132 1001920 212138 1001932
rect 213914 1001920 213920 1001932
rect 213972 1001920 213978 1001972
rect 261018 1001920 261024 1001972
rect 261076 1001960 261082 1001972
rect 263594 1001960 263600 1001972
rect 261076 1001932 263600 1001960
rect 261076 1001920 261082 1001932
rect 263594 1001920 263600 1001932
rect 263652 1001920 263658 1001972
rect 263870 1001920 263876 1001972
rect 263928 1001960 263934 1001972
rect 266998 1001960 267004 1001972
rect 263928 1001932 267004 1001960
rect 263928 1001920 263934 1001932
rect 266998 1001920 267004 1001932
rect 267056 1001920 267062 1001972
rect 310146 1001920 310152 1001972
rect 310204 1001960 310210 1001972
rect 311894 1001960 311900 1001972
rect 310204 1001932 311900 1001960
rect 310204 1001920 310210 1001932
rect 311894 1001920 311900 1001932
rect 311952 1001920 311958 1001972
rect 312630 1001920 312636 1001972
rect 312688 1001960 312694 1001972
rect 314654 1001960 314660 1001972
rect 312688 1001932 314660 1001960
rect 312688 1001920 312694 1001932
rect 314654 1001920 314660 1001932
rect 314712 1001920 314718 1001972
rect 351822 1001920 351828 1001972
rect 351880 1001960 351886 1001972
rect 354030 1001960 354036 1001972
rect 351880 1001932 354036 1001960
rect 351880 1001920 351886 1001932
rect 354030 1001920 354036 1001932
rect 354088 1001920 354094 1001972
rect 356054 1001920 356060 1001972
rect 356112 1001960 356118 1001972
rect 356514 1001960 356520 1001972
rect 356112 1001932 356520 1001960
rect 356112 1001920 356118 1001932
rect 356514 1001920 356520 1001932
rect 356572 1001920 356578 1001972
rect 357342 1001920 357348 1001972
rect 357400 1001960 357406 1001972
rect 360838 1001960 360844 1001972
rect 357400 1001932 360844 1001960
rect 357400 1001920 357406 1001932
rect 360838 1001920 360844 1001932
rect 360896 1001920 360902 1001972
rect 361390 1001920 361396 1001972
rect 361448 1001960 361454 1001972
rect 363598 1001960 363604 1001972
rect 361448 1001932 363604 1001960
rect 361448 1001920 361454 1001932
rect 363598 1001920 363604 1001932
rect 363656 1001920 363662 1001972
rect 365898 1001920 365904 1001972
rect 365956 1001960 365962 1001972
rect 369118 1001960 369124 1001972
rect 365956 1001932 369124 1001960
rect 365956 1001920 365962 1001932
rect 369118 1001920 369124 1001932
rect 369176 1001920 369182 1001972
rect 419442 1001920 419448 1001972
rect 419500 1001960 419506 1001972
rect 421466 1001960 421472 1001972
rect 419500 1001932 421472 1001960
rect 419500 1001920 419506 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 424318 1001920 424324 1001972
rect 424376 1001960 424382 1001972
rect 425054 1001960 425060 1001972
rect 424376 1001932 425060 1001960
rect 424376 1001920 424382 1001932
rect 425054 1001920 425060 1001932
rect 425112 1001920 425118 1001972
rect 426342 1001920 426348 1001972
rect 426400 1001960 426406 1001972
rect 428458 1001960 428464 1001972
rect 426400 1001932 428464 1001960
rect 426400 1001920 426406 1001932
rect 428458 1001920 428464 1001932
rect 428516 1001920 428522 1001972
rect 432874 1001920 432880 1001972
rect 432932 1001960 432938 1001972
rect 436738 1001960 436744 1001972
rect 432932 1001932 436744 1001960
rect 432932 1001920 432938 1001932
rect 436738 1001920 436744 1001932
rect 436796 1001920 436802 1001972
rect 496722 1001920 496728 1001972
rect 496780 1001960 496786 1001972
rect 498470 1001960 498476 1001972
rect 496780 1001932 498476 1001960
rect 496780 1001920 496786 1001932
rect 498470 1001920 498476 1001932
rect 498528 1001920 498534 1001972
rect 502242 1001920 502248 1001972
rect 502300 1001960 502306 1001972
rect 503346 1001960 503352 1001972
rect 502300 1001932 503352 1001960
rect 502300 1001920 502306 1001932
rect 503346 1001920 503352 1001932
rect 503404 1001920 503410 1001972
rect 504174 1001920 504180 1001972
rect 504232 1001960 504238 1001972
rect 505738 1001960 505744 1001972
rect 504232 1001932 505744 1001960
rect 504232 1001920 504238 1001932
rect 505738 1001920 505744 1001932
rect 505796 1001920 505802 1001972
rect 506198 1001920 506204 1001972
rect 506256 1001960 506262 1001972
rect 507854 1001960 507860 1001972
rect 506256 1001932 507860 1001960
rect 506256 1001920 506262 1001932
rect 507854 1001920 507860 1001932
rect 507912 1001920 507918 1001972
rect 554314 1001920 554320 1001972
rect 554372 1001960 554378 1001972
rect 555418 1001960 555424 1001972
rect 554372 1001932 555424 1001960
rect 554372 1001920 554378 1001932
rect 555418 1001920 555424 1001932
rect 555476 1001920 555482 1001972
rect 558822 1001920 558828 1001972
rect 558880 1001960 558886 1001972
rect 560202 1001960 560208 1001972
rect 558880 1001932 560208 1001960
rect 558880 1001920 558886 1001932
rect 560202 1001920 560208 1001932
rect 560260 1001920 560266 1001972
rect 561674 1001920 561680 1001972
rect 561732 1001960 561738 1001972
rect 565078 1001960 565084 1001972
rect 561732 1001932 565084 1001960
rect 561732 1001920 561738 1001932
rect 565078 1001920 565084 1001932
rect 565136 1001920 565142 1001972
rect 512822 1001376 512828 1001428
rect 512880 1001416 512886 1001428
rect 519538 1001416 519544 1001428
rect 512880 1001388 519544 1001416
rect 512880 1001376 512886 1001388
rect 519538 1001376 519544 1001388
rect 519596 1001376 519602 1001428
rect 246574 1001172 246580 1001224
rect 246632 1001212 246638 1001224
rect 256970 1001212 256976 1001224
rect 246632 1001184 256976 1001212
rect 246632 1001172 246638 1001184
rect 256970 1001172 256976 1001184
rect 257028 1001172 257034 1001224
rect 355778 1001172 355784 1001224
rect 355836 1001212 355842 1001224
rect 378778 1001212 378784 1001224
rect 355836 1001184 378784 1001212
rect 355836 1001172 355842 1001184
rect 378778 1001172 378784 1001184
rect 378836 1001172 378842 1001224
rect 510154 1000900 510160 1000952
rect 510212 1000940 510218 1000952
rect 517238 1000940 517244 1000952
rect 510212 1000912 517244 1000940
rect 510212 1000900 510218 1000912
rect 517238 1000900 517244 1000912
rect 517296 1000900 517302 1000952
rect 92658 999744 92664 999796
rect 92716 999784 92722 999796
rect 99006 999784 99012 999796
rect 92716 999756 99012 999784
rect 92716 999744 92722 999756
rect 99006 999744 99012 999756
rect 99064 999744 99070 999796
rect 195514 999744 195520 999796
rect 195572 999784 195578 999796
rect 209866 999784 209872 999796
rect 195572 999756 209872 999784
rect 195572 999744 195578 999756
rect 209866 999744 209872 999756
rect 209924 999744 209930 999796
rect 591298 999268 591304 999320
rect 591356 999308 591362 999320
rect 616782 999308 616788 999320
rect 591356 999280 616788 999308
rect 591356 999268 591362 999280
rect 616782 999268 616788 999280
rect 616840 999268 616846 999320
rect 298922 999132 298928 999184
rect 298980 999172 298986 999184
rect 305270 999172 305276 999184
rect 298980 999144 305276 999172
rect 298980 999132 298986 999144
rect 305270 999132 305276 999144
rect 305328 999132 305334 999184
rect 378134 999132 378140 999184
rect 378192 999172 378198 999184
rect 383286 999172 383292 999184
rect 378192 999144 383292 999172
rect 378192 999132 378198 999144
rect 383286 999132 383292 999144
rect 383344 999132 383350 999184
rect 458082 999132 458088 999184
rect 458140 999172 458146 999184
rect 458140 999144 460934 999172
rect 458140 999132 458146 999144
rect 373258 999064 373264 999116
rect 373316 999104 373322 999116
rect 375558 999104 375564 999116
rect 373316 999076 375564 999104
rect 373316 999064 373322 999076
rect 375558 999064 375564 999076
rect 375616 999064 375622 999116
rect 446398 999064 446404 999116
rect 446456 999104 446462 999116
rect 452286 999104 452292 999116
rect 446456 999076 452292 999104
rect 446456 999064 446462 999076
rect 452286 999064 452292 999076
rect 452344 999064 452350 999116
rect 460906 998968 460934 999144
rect 591114 999132 591120 999184
rect 591172 999172 591178 999184
rect 625614 999172 625620 999184
rect 591172 999144 625620 999172
rect 591172 999132 591178 999144
rect 625614 999132 625620 999144
rect 625672 999132 625678 999184
rect 516778 999064 516784 999116
rect 516836 999104 516842 999116
rect 523310 999104 523316 999116
rect 516836 999076 523316 999104
rect 516836 999064 516842 999076
rect 523310 999064 523316 999076
rect 523368 999064 523374 999116
rect 472618 998968 472624 998980
rect 460906 998940 472624 998968
rect 472618 998928 472624 998940
rect 472676 998928 472682 998980
rect 513834 998928 513840 998980
rect 513892 998968 513898 998980
rect 523678 998968 523684 998980
rect 513892 998940 523684 998968
rect 513892 998928 513898 998940
rect 523678 998928 523684 998940
rect 523736 998928 523742 998980
rect 428458 998792 428464 998844
rect 428516 998832 428522 998844
rect 466454 998832 466460 998844
rect 428516 998804 466460 998832
rect 428516 998792 428522 998804
rect 466454 998792 466460 998804
rect 466512 998792 466518 998844
rect 504358 998792 504364 998844
rect 504416 998832 504422 998844
rect 516686 998832 516692 998844
rect 504416 998804 516692 998832
rect 504416 998792 504422 998804
rect 516686 998792 516692 998804
rect 516744 998792 516750 998844
rect 378594 998764 378600 998776
rect 373966 998736 378600 998764
rect 196618 998656 196624 998708
rect 196676 998696 196682 998708
rect 204346 998696 204352 998708
rect 196676 998668 204352 998696
rect 196676 998656 196682 998668
rect 204346 998656 204352 998668
rect 204404 998656 204410 998708
rect 199378 998520 199384 998572
rect 199436 998560 199442 998572
rect 203518 998560 203524 998572
rect 199436 998532 203524 998560
rect 199436 998520 199442 998532
rect 203518 998520 203524 998532
rect 203576 998520 203582 998572
rect 303246 998520 303252 998572
rect 303304 998560 303310 998572
rect 308950 998560 308956 998572
rect 303304 998532 308956 998560
rect 303304 998520 303310 998532
rect 308950 998520 308956 998532
rect 309008 998520 309014 998572
rect 355134 998520 355140 998572
rect 355192 998560 355198 998572
rect 373966 998560 373994 998736
rect 378594 998724 378600 998736
rect 378652 998724 378658 998776
rect 431310 998656 431316 998708
rect 431368 998696 431374 998708
rect 472434 998696 472440 998708
rect 431368 998668 472440 998696
rect 431368 998656 431374 998668
rect 472434 998656 472440 998668
rect 472492 998656 472498 998708
rect 499482 998656 499488 998708
rect 499540 998696 499546 998708
rect 510062 998696 510068 998708
rect 499540 998668 510068 998696
rect 499540 998656 499546 998668
rect 510062 998656 510068 998668
rect 510120 998656 510126 998708
rect 377398 998588 377404 998640
rect 377456 998628 377462 998640
rect 383562 998628 383568 998640
rect 377456 998600 383568 998628
rect 377456 998588 377462 998600
rect 383562 998588 383568 998600
rect 383620 998588 383626 998640
rect 355192 998532 373994 998560
rect 355192 998520 355198 998532
rect 425054 998520 425060 998572
rect 425112 998560 425118 998572
rect 472066 998560 472072 998572
rect 425112 998532 472072 998560
rect 425112 998520 425118 998532
rect 472066 998520 472072 998532
rect 472124 998520 472130 998572
rect 506474 998520 506480 998572
rect 506532 998560 506538 998572
rect 524046 998560 524052 998572
rect 506532 998532 524052 998560
rect 506532 998520 506538 998532
rect 524046 998520 524052 998532
rect 524104 998520 524110 998572
rect 200850 998384 200856 998436
rect 200908 998424 200914 998436
rect 203886 998424 203892 998436
rect 200908 998396 203892 998424
rect 200908 998384 200914 998396
rect 203886 998384 203892 998396
rect 203944 998384 203950 998436
rect 247862 998384 247868 998436
rect 247920 998424 247926 998436
rect 258994 998424 259000 998436
rect 247920 998396 259000 998424
rect 247920 998384 247926 998396
rect 258994 998384 259000 998396
rect 259052 998384 259058 998436
rect 304442 998384 304448 998436
rect 304500 998424 304506 998436
rect 307294 998424 307300 998436
rect 304500 998396 307300 998424
rect 304500 998384 304506 998396
rect 307294 998384 307300 998396
rect 307352 998384 307358 998436
rect 356054 998384 356060 998436
rect 356112 998424 356118 998436
rect 383470 998424 383476 998436
rect 356112 998396 383476 998424
rect 356112 998384 356118 998396
rect 383470 998384 383476 998396
rect 383528 998384 383534 998436
rect 423582 998384 423588 998436
rect 423640 998424 423646 998436
rect 472250 998424 472256 998436
rect 423640 998396 472256 998424
rect 423640 998384 423646 998396
rect 472250 998384 472256 998396
rect 472308 998384 472314 998436
rect 500218 998384 500224 998436
rect 500276 998424 500282 998436
rect 523126 998424 523132 998436
rect 500276 998396 523132 998424
rect 500276 998384 500282 998396
rect 523126 998384 523132 998396
rect 523184 998384 523190 998436
rect 616782 998384 616788 998436
rect 616840 998424 616846 998436
rect 625430 998424 625436 998436
rect 616840 998396 625436 998424
rect 616840 998384 616846 998396
rect 625430 998384 625436 998396
rect 625488 998384 625494 998436
rect 196802 998248 196808 998300
rect 196860 998288 196866 998300
rect 202690 998288 202696 998300
rect 196860 998260 202696 998288
rect 196860 998248 196866 998260
rect 202690 998248 202696 998260
rect 202748 998248 202754 998300
rect 302878 998248 302884 998300
rect 302936 998288 302942 998300
rect 306098 998288 306104 998300
rect 302936 998260 306104 998288
rect 302936 998248 302942 998260
rect 306098 998248 306104 998260
rect 306156 998248 306162 998300
rect 443638 998248 443644 998300
rect 443696 998288 443702 998300
rect 446858 998288 446864 998300
rect 443696 998260 446864 998288
rect 443696 998248 443702 998260
rect 446858 998248 446864 998260
rect 446916 998248 446922 998300
rect 510062 998248 510068 998300
rect 510120 998288 510126 998300
rect 520550 998288 520556 998300
rect 510120 998260 520556 998288
rect 510120 998248 510126 998260
rect 520550 998248 520556 998260
rect 520608 998248 520614 998300
rect 254578 998180 254584 998232
rect 254636 998220 254642 998232
rect 257338 998220 257344 998232
rect 254636 998192 257344 998220
rect 254636 998180 254642 998192
rect 257338 998180 257344 998192
rect 257396 998180 257402 998232
rect 198642 998112 198648 998164
rect 198700 998152 198706 998164
rect 200666 998152 200672 998164
rect 198700 998124 200672 998152
rect 198700 998112 198706 998124
rect 200666 998112 200672 998124
rect 200724 998112 200730 998164
rect 202138 998112 202144 998164
rect 202196 998152 202202 998164
rect 204070 998152 204076 998164
rect 202196 998124 204076 998152
rect 202196 998112 202202 998124
rect 204070 998112 204076 998124
rect 204128 998112 204134 998164
rect 247678 998112 247684 998164
rect 247736 998152 247742 998164
rect 253658 998152 253664 998164
rect 247736 998124 253664 998152
rect 247736 998112 247742 998124
rect 253658 998112 253664 998124
rect 253716 998112 253722 998164
rect 305638 998112 305644 998164
rect 305696 998152 305702 998164
rect 308122 998152 308128 998164
rect 305696 998124 308128 998152
rect 305696 998112 305702 998124
rect 308122 998112 308128 998124
rect 308180 998112 308186 998164
rect 143718 998044 143724 998096
rect 143776 998084 143782 998096
rect 146938 998084 146944 998096
rect 143776 998056 146944 998084
rect 143776 998044 143782 998056
rect 146938 998044 146944 998056
rect 146996 998044 147002 998096
rect 255958 998044 255964 998096
rect 256016 998084 256022 998096
rect 258166 998084 258172 998096
rect 256016 998056 258172 998084
rect 256016 998044 256022 998056
rect 258166 998044 258172 998056
rect 258224 998044 258230 998096
rect 260190 998044 260196 998096
rect 260248 998084 260254 998096
rect 262858 998084 262864 998096
rect 260248 998056 262864 998084
rect 260248 998044 260254 998056
rect 262858 998044 262864 998056
rect 262916 998044 262922 998096
rect 92290 997976 92296 998028
rect 92348 998016 92354 998028
rect 94682 998016 94688 998028
rect 92348 997988 94688 998016
rect 92348 997976 92354 997988
rect 94682 997976 94688 997988
rect 94740 997976 94746 998028
rect 200022 997976 200028 998028
rect 200080 998016 200086 998028
rect 201862 998016 201868 998028
rect 200080 997988 201868 998016
rect 200080 997976 200086 997988
rect 201862 997976 201868 997988
rect 201920 997976 201926 998028
rect 250990 997976 250996 998028
rect 251048 998016 251054 998028
rect 253290 998016 253296 998028
rect 251048 997988 253296 998016
rect 251048 997976 251054 997988
rect 253290 997976 253296 997988
rect 253348 997976 253354 998028
rect 304258 997976 304264 998028
rect 304316 998016 304322 998028
rect 306926 998016 306932 998028
rect 304316 997988 306932 998016
rect 304316 997976 304322 997988
rect 306926 997976 306932 997988
rect 306984 997976 306990 998028
rect 308398 997976 308404 998028
rect 308456 998016 308462 998028
rect 310606 998016 310612 998028
rect 308456 997988 310612 998016
rect 308456 997976 308462 997988
rect 310606 997976 310612 997988
rect 310664 997976 310670 998028
rect 549162 997976 549168 998028
rect 549220 998016 549226 998028
rect 551094 998016 551100 998028
rect 549220 997988 551100 998016
rect 549220 997976 549226 997988
rect 551094 997976 551100 997988
rect 551152 997976 551158 998028
rect 202322 997908 202328 997960
rect 202380 997948 202386 997960
rect 204714 997948 204720 997960
rect 202380 997920 204720 997948
rect 202380 997908 202386 997920
rect 204714 997908 204720 997920
rect 204772 997908 204778 997960
rect 257338 997908 257344 997960
rect 257396 997948 257402 997960
rect 258994 997948 259000 997960
rect 257396 997920 259000 997948
rect 257396 997908 257402 997920
rect 258994 997908 259000 997920
rect 259052 997908 259058 997960
rect 259822 997908 259828 997960
rect 259880 997948 259886 997960
rect 262214 997948 262220 997960
rect 259880 997920 262220 997948
rect 259880 997908 259886 997920
rect 262214 997908 262220 997920
rect 262272 997908 262278 997960
rect 143902 997840 143908 997892
rect 143960 997880 143966 997892
rect 151262 997880 151268 997892
rect 143960 997852 151268 997880
rect 143960 997840 143966 997852
rect 151262 997840 151268 997852
rect 151320 997840 151326 997892
rect 249702 997840 249708 997892
rect 249760 997880 249766 997892
rect 252462 997880 252468 997892
rect 249760 997852 252468 997880
rect 249760 997840 249766 997852
rect 252462 997840 252468 997852
rect 252520 997840 252526 997892
rect 303522 997840 303528 997892
rect 303580 997880 303586 997892
rect 304902 997880 304908 997892
rect 303580 997852 304908 997880
rect 303580 997840 303586 997852
rect 304902 997840 304908 997852
rect 304960 997840 304966 997892
rect 307018 997840 307024 997892
rect 307076 997880 307082 997892
rect 308950 997880 308956 997892
rect 307076 997852 308956 997880
rect 307076 997840 307082 997852
rect 308950 997840 308956 997852
rect 309008 997840 309014 997892
rect 547782 997840 547788 997892
rect 547840 997880 547846 997892
rect 550266 997880 550272 997892
rect 547840 997852 550272 997880
rect 547840 997840 547846 997852
rect 550266 997840 550272 997852
rect 550324 997840 550330 997892
rect 550542 997840 550548 997892
rect 550600 997880 550606 997892
rect 553302 997880 553308 997892
rect 550600 997852 553308 997880
rect 550600 997840 550606 997852
rect 553302 997840 553308 997852
rect 553360 997840 553366 997892
rect 200942 997772 200948 997824
rect 201000 997812 201006 997824
rect 203518 997812 203524 997824
rect 201000 997784 203524 997812
rect 201000 997772 201006 997784
rect 203518 997772 203524 997784
rect 203576 997772 203582 997824
rect 258166 997772 258172 997824
rect 258224 997812 258230 997824
rect 259454 997812 259460 997824
rect 258224 997784 259460 997812
rect 258224 997772 258230 997784
rect 259454 997772 259460 997784
rect 259512 997772 259518 997824
rect 260190 997772 260196 997824
rect 260248 997812 260254 997824
rect 260926 997812 260932 997824
rect 260248 997784 260932 997812
rect 260248 997772 260254 997784
rect 260926 997772 260932 997784
rect 260984 997772 260990 997824
rect 378778 997772 378784 997824
rect 378836 997812 378842 997824
rect 383102 997812 383108 997824
rect 378836 997784 383108 997812
rect 378836 997772 378842 997784
rect 383102 997772 383108 997784
rect 383160 997772 383166 997824
rect 488902 997772 488908 997824
rect 488960 997812 488966 997824
rect 493502 997812 493508 997824
rect 488960 997784 493508 997812
rect 488960 997772 488966 997784
rect 493502 997772 493508 997784
rect 493560 997772 493566 997824
rect 520918 997772 520924 997824
rect 520976 997812 520982 997824
rect 523862 997812 523868 997824
rect 520976 997784 523868 997812
rect 520976 997772 520982 997784
rect 523862 997772 523868 997784
rect 523920 997772 523926 997824
rect 592034 997772 592040 997824
rect 592092 997812 592098 997824
rect 625798 997812 625804 997824
rect 592092 997784 625804 997812
rect 592092 997772 592098 997784
rect 625798 997772 625804 997784
rect 625856 997772 625862 997824
rect 144822 997704 144828 997756
rect 144880 997744 144886 997756
rect 152642 997744 152648 997756
rect 144880 997716 152648 997744
rect 144880 997704 144886 997716
rect 152642 997704 152648 997716
rect 152700 997704 152706 997756
rect 247218 997704 247224 997756
rect 247276 997744 247282 997756
rect 254578 997744 254584 997756
rect 247276 997716 254584 997744
rect 247276 997704 247282 997716
rect 254578 997704 254584 997716
rect 254636 997704 254642 997756
rect 299106 997704 299112 997756
rect 299164 997744 299170 997756
rect 310422 997744 310428 997756
rect 299164 997716 310428 997744
rect 299164 997704 299170 997716
rect 310422 997704 310428 997716
rect 310480 997704 310486 997756
rect 363598 997704 363604 997756
rect 363656 997744 363662 997756
rect 372338 997744 372344 997756
rect 363656 997716 372344 997744
rect 363656 997704 363662 997716
rect 372338 997704 372344 997716
rect 372396 997704 372402 997756
rect 431126 997704 431132 997756
rect 431184 997744 431190 997756
rect 439682 997744 439688 997756
rect 431184 997716 439688 997744
rect 431184 997704 431190 997716
rect 439682 997704 439688 997716
rect 439740 997704 439746 997756
rect 515582 997704 515588 997756
rect 515640 997744 515646 997756
rect 516870 997744 516876 997756
rect 515640 997716 516876 997744
rect 515640 997704 515646 997716
rect 516870 997704 516876 997716
rect 516928 997704 516934 997756
rect 164878 997636 164884 997688
rect 164936 997676 164942 997688
rect 170306 997676 170312 997688
rect 164936 997648 170312 997676
rect 164936 997636 164942 997648
rect 170306 997636 170312 997648
rect 170364 997636 170370 997688
rect 566458 997636 566464 997688
rect 566516 997676 566522 997688
rect 623682 997676 623688 997688
rect 566516 997648 623688 997676
rect 566516 997636 566522 997648
rect 623682 997636 623688 997648
rect 623740 997636 623746 997688
rect 438118 997568 438124 997620
rect 438176 997608 438182 997620
rect 439866 997608 439872 997620
rect 438176 997580 439872 997608
rect 438176 997568 438182 997580
rect 439866 997568 439872 997580
rect 439924 997568 439930 997620
rect 573358 997500 573364 997552
rect 573416 997540 573422 997552
rect 573416 997512 581684 997540
rect 573416 997500 573422 997512
rect 553118 997364 553124 997416
rect 553176 997404 553182 997416
rect 581270 997404 581276 997416
rect 553176 997376 581276 997404
rect 553176 997364 553182 997376
rect 581270 997364 581276 997376
rect 581328 997364 581334 997416
rect 581656 997404 581684 997512
rect 581822 997500 581828 997552
rect 581880 997540 581886 997552
rect 591298 997540 591304 997552
rect 581880 997512 591304 997540
rect 581880 997500 581886 997512
rect 591298 997500 591304 997512
rect 591356 997500 591362 997552
rect 590378 997404 590384 997416
rect 581656 997376 590384 997404
rect 590378 997364 590384 997376
rect 590436 997364 590442 997416
rect 319438 997296 319444 997348
rect 319496 997336 319502 997348
rect 332594 997336 332600 997348
rect 319496 997308 332600 997336
rect 319496 997296 319502 997308
rect 332594 997296 332600 997308
rect 332652 997296 332658 997348
rect 97074 997228 97080 997280
rect 97132 997268 97138 997280
rect 98822 997268 98828 997280
rect 97132 997240 98828 997268
rect 97132 997228 97138 997240
rect 98822 997228 98828 997240
rect 98880 997228 98886 997280
rect 331122 997160 331128 997212
rect 331180 997200 331186 997212
rect 357342 997200 357348 997212
rect 331180 997172 357348 997200
rect 331180 997160 331186 997172
rect 357342 997160 357348 997172
rect 357400 997160 357406 997212
rect 569218 997160 569224 997212
rect 569276 997200 569282 997212
rect 620278 997200 620284 997212
rect 569276 997172 620284 997200
rect 569276 997160 569282 997172
rect 620278 997160 620284 997172
rect 620336 997160 620342 997212
rect 318058 997024 318064 997076
rect 318116 997064 318122 997076
rect 349154 997064 349160 997076
rect 318116 997036 349160 997064
rect 318116 997024 318122 997036
rect 349154 997024 349160 997036
rect 349212 997024 349218 997076
rect 360838 997024 360844 997076
rect 360896 997064 360902 997076
rect 380894 997064 380900 997076
rect 360896 997036 380900 997064
rect 360896 997024 360902 997036
rect 380894 997024 380900 997036
rect 380952 997024 380958 997076
rect 558178 997024 558184 997076
rect 558236 997064 558242 997076
rect 617334 997064 617340 997076
rect 558236 997036 617340 997064
rect 558236 997024 558242 997036
rect 617334 997024 617340 997036
rect 617392 997024 617398 997076
rect 106918 996888 106924 996940
rect 106976 996928 106982 996940
rect 111886 996928 111892 996940
rect 106976 996900 111892 996928
rect 106976 996888 106982 996900
rect 111886 996888 111892 996900
rect 111944 996888 111950 996940
rect 570782 996888 570788 996940
rect 570840 996928 570846 996940
rect 581454 996928 581460 996940
rect 570840 996900 581460 996928
rect 570840 996888 570846 996900
rect 581454 996888 581460 996900
rect 581512 996888 581518 996940
rect 592034 996928 592040 996940
rect 581656 996900 592040 996928
rect 574738 996752 574744 996804
rect 574796 996792 574802 996804
rect 581656 996792 581684 996900
rect 592034 996888 592040 996900
rect 592092 996888 592098 996940
rect 574796 996764 581684 996792
rect 574796 996752 574802 996764
rect 581270 996616 581276 996668
rect 581328 996656 581334 996668
rect 590562 996656 590568 996668
rect 581328 996628 590568 996656
rect 581328 996616 581334 996628
rect 590562 996616 590568 996628
rect 590620 996616 590626 996668
rect 200206 996412 200212 996464
rect 200264 996452 200270 996464
rect 203702 996452 203708 996464
rect 200264 996424 203708 996452
rect 200264 996412 200270 996424
rect 203702 996412 203708 996424
rect 203760 996412 203766 996464
rect 421006 996412 421012 996464
rect 421064 996452 421070 996464
rect 426434 996452 426440 996464
rect 421064 996424 426440 996452
rect 421064 996412 421070 996424
rect 426434 996412 426440 996424
rect 426492 996412 426498 996464
rect 92474 996344 92480 996396
rect 92532 996384 92538 996396
rect 121730 996384 121736 996396
rect 92532 996356 121736 996384
rect 92532 996344 92538 996356
rect 121730 996344 121736 996356
rect 121788 996344 121794 996396
rect 555418 996276 555424 996328
rect 555476 996316 555482 996328
rect 591114 996316 591120 996328
rect 555476 996288 591120 996316
rect 555476 996276 555482 996288
rect 591114 996276 591120 996288
rect 591172 996276 591178 996328
rect 551922 996208 551928 996260
rect 551980 996248 551986 996260
rect 554314 996248 554320 996260
rect 551980 996220 554320 996248
rect 551980 996208 551986 996220
rect 554314 996208 554320 996220
rect 554372 996208 554378 996260
rect 109494 996072 109500 996124
rect 109552 996112 109558 996124
rect 158714 996112 158720 996124
rect 109552 996084 158720 996112
rect 109552 996072 109558 996084
rect 158714 996072 158720 996084
rect 158772 996072 158778 996124
rect 159358 996072 159364 996124
rect 159416 996112 159422 996124
rect 208394 996112 208400 996124
rect 159416 996084 208400 996112
rect 159416 996072 159422 996084
rect 208394 996072 208400 996084
rect 208452 996072 208458 996124
rect 229738 996072 229744 996124
rect 229796 996112 229802 996124
rect 262214 996112 262220 996124
rect 229796 996084 262220 996112
rect 229796 996072 229802 996084
rect 262214 996072 262220 996084
rect 262272 996072 262278 996124
rect 278038 996072 278044 996124
rect 278096 996112 278102 996124
rect 316034 996112 316040 996124
rect 278096 996084 316040 996112
rect 278096 996072 278102 996084
rect 316034 996072 316040 996084
rect 316092 996072 316098 996124
rect 366542 996072 366548 996124
rect 366600 996112 366606 996124
rect 433518 996112 433524 996124
rect 366600 996084 433524 996112
rect 366600 996072 366606 996084
rect 433518 996072 433524 996084
rect 433576 996072 433582 996124
rect 433978 996072 433984 996124
rect 434036 996112 434042 996124
rect 510706 996112 510712 996124
rect 434036 996084 510712 996112
rect 434036 996072 434042 996084
rect 510706 996072 510712 996084
rect 510764 996072 510770 996124
rect 522482 996072 522488 996124
rect 522540 996112 522546 996124
rect 560570 996112 560576 996124
rect 522540 996084 560576 996112
rect 522540 996072 522546 996084
rect 560570 996072 560576 996084
rect 560628 996072 560634 996124
rect 567166 996084 621014 996112
rect 111058 995936 111064 995988
rect 111116 995976 111122 995988
rect 144454 995976 144460 995988
rect 111116 995948 144460 995976
rect 111116 995936 111122 995948
rect 144454 995936 144460 995948
rect 144512 995936 144518 995988
rect 162118 995936 162124 995988
rect 162176 995976 162182 995988
rect 210234 995976 210240 995988
rect 162176 995948 210240 995976
rect 162176 995936 162182 995948
rect 210234 995936 210240 995948
rect 210292 995936 210298 995988
rect 228358 995936 228364 995988
rect 228416 995976 228422 995988
rect 263594 995976 263600 995988
rect 228416 995948 263600 995976
rect 228416 995936 228422 995948
rect 263594 995936 263600 995948
rect 263652 995936 263658 995988
rect 264238 995936 264244 995988
rect 264296 995976 264302 995988
rect 299290 995976 299296 995988
rect 264296 995948 299296 995976
rect 264296 995936 264302 995948
rect 299290 995936 299296 995948
rect 299348 995936 299354 995988
rect 365254 995936 365260 995988
rect 365312 995976 365318 995988
rect 432230 995976 432236 995988
rect 365312 995948 432236 995976
rect 365312 995936 365318 995948
rect 432230 995936 432236 995948
rect 432288 995936 432294 995988
rect 434162 995936 434168 995988
rect 434220 995976 434226 995988
rect 510890 995976 510896 995988
rect 434220 995948 510896 995976
rect 434220 995936 434226 995948
rect 510890 995936 510896 995948
rect 510948 995936 510954 995988
rect 522298 995936 522304 995988
rect 522356 995976 522362 995988
rect 563054 995976 563060 995988
rect 522356 995948 563060 995976
rect 522356 995936 522362 995948
rect 563054 995936 563060 995948
rect 563112 995936 563118 995988
rect 124858 995800 124864 995852
rect 124916 995840 124922 995852
rect 160370 995840 160376 995852
rect 124916 995812 160376 995840
rect 124916 995800 124922 995812
rect 160370 995800 160376 995812
rect 160428 995800 160434 995852
rect 175918 995800 175924 995852
rect 175976 995840 175982 995852
rect 211154 995840 211160 995852
rect 175976 995812 211160 995840
rect 175976 995800 175982 995812
rect 211154 995800 211160 995812
rect 211212 995800 211218 995852
rect 213178 995800 213184 995852
rect 213236 995840 213242 995852
rect 261110 995840 261116 995852
rect 213236 995812 261116 995840
rect 213236 995800 213242 995812
rect 261110 995800 261116 995812
rect 261168 995800 261174 995852
rect 280798 995800 280804 995852
rect 280856 995840 280862 995852
rect 314654 995840 314660 995852
rect 280856 995812 314660 995840
rect 280856 995800 280862 995812
rect 314654 995800 314660 995812
rect 314712 995800 314718 995852
rect 364978 995800 364984 995852
rect 365036 995840 365042 995852
rect 432046 995840 432052 995852
rect 365036 995812 432052 995840
rect 365036 995800 365042 995812
rect 432046 995800 432052 995812
rect 432104 995800 432110 995852
rect 471238 995800 471244 995852
rect 471296 995840 471302 995852
rect 507854 995840 507860 995852
rect 471296 995812 507860 995840
rect 471296 995800 471302 995812
rect 507854 995800 507860 995812
rect 507912 995800 507918 995852
rect 509694 995800 509700 995852
rect 509752 995840 509758 995852
rect 554130 995840 554136 995852
rect 509752 995812 554136 995840
rect 509752 995800 509758 995812
rect 554130 995800 554136 995812
rect 554188 995800 554194 995852
rect 554314 995800 554320 995852
rect 554372 995840 554378 995852
rect 567166 995840 567194 996084
rect 554372 995812 567194 995840
rect 620986 995840 621014 996084
rect 625430 995840 625436 995852
rect 620986 995812 625436 995840
rect 554372 995800 554378 995812
rect 625430 995800 625436 995812
rect 625488 995800 625494 995852
rect 195054 995528 195060 995580
rect 195112 995568 195118 995580
rect 200942 995568 200948 995580
rect 195112 995540 200948 995568
rect 195112 995528 195118 995540
rect 200942 995528 200948 995540
rect 201000 995528 201006 995580
rect 246206 995528 246212 995580
rect 246264 995568 246270 995580
rect 252002 995568 252008 995580
rect 246264 995540 252008 995568
rect 246264 995528 246270 995540
rect 252002 995528 252008 995540
rect 252060 995528 252066 995580
rect 298462 995528 298468 995580
rect 298520 995568 298526 995580
rect 304442 995568 304448 995580
rect 298520 995540 304448 995568
rect 298520 995528 298526 995540
rect 304442 995528 304448 995540
rect 304500 995528 304506 995580
rect 323578 995528 323584 995580
rect 323636 995568 323642 995580
rect 364978 995568 364984 995580
rect 323636 995540 364984 995568
rect 323636 995528 323642 995540
rect 364978 995528 364984 995540
rect 365036 995528 365042 995580
rect 366358 995528 366364 995580
rect 366416 995568 366422 995580
rect 366416 995540 373994 995568
rect 366416 995528 366422 995540
rect 177298 995460 177304 995512
rect 177356 995500 177362 995512
rect 177356 995472 180794 995500
rect 177356 995460 177362 995472
rect 126238 995392 126244 995444
rect 126296 995432 126302 995444
rect 160186 995432 160192 995444
rect 126296 995404 160192 995432
rect 126296 995392 126302 995404
rect 160186 995392 160192 995404
rect 160244 995392 160250 995444
rect 180766 995432 180794 995472
rect 212534 995432 212540 995444
rect 180766 995404 212540 995432
rect 212534 995392 212540 995404
rect 212592 995392 212598 995444
rect 262858 995392 262864 995444
rect 262916 995432 262922 995444
rect 313274 995432 313280 995444
rect 262916 995404 313280 995432
rect 262916 995392 262922 995404
rect 313274 995392 313280 995404
rect 313332 995392 313338 995444
rect 88978 995324 88984 995376
rect 89036 995364 89042 995376
rect 92474 995364 92480 995376
rect 89036 995336 92480 995364
rect 89036 995324 89042 995336
rect 92474 995324 92480 995336
rect 92532 995324 92538 995376
rect 373966 995364 373994 995540
rect 472618 995528 472624 995580
rect 472676 995568 472682 995580
rect 473998 995568 474004 995580
rect 472676 995540 474004 995568
rect 472676 995528 472682 995540
rect 473998 995528 474004 995540
rect 474056 995528 474062 995580
rect 493502 995528 493508 995580
rect 493560 995568 493566 995580
rect 511074 995568 511080 995580
rect 493560 995540 511080 995568
rect 493560 995528 493566 995540
rect 511074 995528 511080 995540
rect 511132 995528 511138 995580
rect 523862 995528 523868 995580
rect 523920 995568 523926 995580
rect 525334 995568 525340 995580
rect 523920 995540 525340 995568
rect 523920 995528 523926 995540
rect 525334 995528 525340 995540
rect 525392 995528 525398 995580
rect 625798 995528 625804 995580
rect 625856 995568 625862 995580
rect 627914 995568 627920 995580
rect 625856 995540 627920 995568
rect 625856 995528 625862 995540
rect 627914 995528 627920 995540
rect 627972 995528 627978 995580
rect 475930 995460 475936 995512
rect 475988 995500 475994 995512
rect 478782 995500 478788 995512
rect 475988 995472 478788 995500
rect 475988 995460 475994 995472
rect 478782 995460 478788 995472
rect 478840 995460 478846 995512
rect 630646 995472 630812 995500
rect 472434 995392 472440 995444
rect 472492 995432 472498 995444
rect 474734 995432 474740 995444
rect 472492 995404 474740 995432
rect 472492 995392 472498 995404
rect 474734 995392 474740 995404
rect 474792 995392 474798 995444
rect 509234 995432 509240 995444
rect 480226 995404 509240 995432
rect 400858 995364 400864 995376
rect 373966 995336 400864 995364
rect 400858 995324 400864 995336
rect 400916 995324 400922 995376
rect 402974 995364 402980 995376
rect 402808 995336 402980 995364
rect 142798 995256 142804 995308
rect 142856 995296 142862 995308
rect 149882 995296 149888 995308
rect 142856 995268 149888 995296
rect 142856 995256 142862 995268
rect 149882 995256 149888 995268
rect 149940 995256 149946 995308
rect 194318 995256 194324 995308
rect 194376 995296 194382 995308
rect 195238 995296 195244 995308
rect 194376 995268 195244 995296
rect 194376 995256 194382 995268
rect 195238 995256 195244 995268
rect 195296 995256 195302 995308
rect 211798 995256 211804 995308
rect 211856 995296 211862 995308
rect 211856 995268 234614 995296
rect 211856 995256 211862 995268
rect 180794 995228 180800 995240
rect 180628 995200 180800 995228
rect 77662 995120 77668 995172
rect 77720 995160 77726 995172
rect 100202 995160 100208 995172
rect 77720 995132 100208 995160
rect 77720 995120 77726 995132
rect 100202 995120 100208 995132
rect 100260 995120 100266 995172
rect 137922 995120 137928 995172
rect 137980 995160 137986 995172
rect 144638 995160 144644 995172
rect 137980 995132 144644 995160
rect 137980 995120 137986 995132
rect 144638 995120 144644 995132
rect 144696 995120 144702 995172
rect 77018 994984 77024 995036
rect 77076 995024 77082 995036
rect 102778 995024 102784 995036
rect 77076 994996 102784 995024
rect 77076 994984 77082 994996
rect 102778 994984 102784 994996
rect 102836 994984 102842 995036
rect 128446 994916 128452 994968
rect 128504 994956 128510 994968
rect 157334 994956 157340 994968
rect 128504 994928 157340 994956
rect 128504 994916 128510 994928
rect 157334 994916 157340 994928
rect 157392 994916 157398 994968
rect 180628 994956 180656 995200
rect 180794 995188 180800 995200
rect 180852 995188 180858 995240
rect 234586 995228 234614 995268
rect 244366 995256 244372 995308
rect 244424 995296 244430 995308
rect 260926 995296 260932 995308
rect 244424 995268 260932 995296
rect 244424 995256 244430 995268
rect 260926 995256 260932 995268
rect 260984 995256 260990 995308
rect 291102 995256 291108 995308
rect 291160 995296 291166 995308
rect 302878 995296 302884 995308
rect 291160 995268 302884 995296
rect 291160 995256 291166 995268
rect 302878 995256 302884 995268
rect 302936 995256 302942 995308
rect 244090 995228 244096 995240
rect 234586 995200 244096 995228
rect 244090 995188 244096 995200
rect 244148 995188 244154 995240
rect 194686 995120 194692 995172
rect 194744 995160 194750 995172
rect 199378 995160 199384 995172
rect 194744 995132 199384 995160
rect 194744 995120 194750 995132
rect 199378 995120 199384 995132
rect 199436 995120 199442 995172
rect 293586 995120 293592 995172
rect 293644 995160 293650 995172
rect 298830 995160 298836 995172
rect 293644 995132 298836 995160
rect 293644 995120 293650 995132
rect 298830 995120 298836 995132
rect 298888 995120 298894 995172
rect 234706 995092 234712 995104
rect 234402 995064 234712 995092
rect 180490 994928 180656 994956
rect 78306 994848 78312 994900
rect 78364 994888 78370 994900
rect 104158 994888 104164 994900
rect 78364 994860 104164 994888
rect 78364 994848 78370 994860
rect 104158 994848 104164 994860
rect 104216 994848 104222 994900
rect 132126 994780 132132 994832
rect 132184 994820 132190 994832
rect 145558 994820 145564 994832
rect 132184 994792 145564 994820
rect 132184 994780 132190 994792
rect 145558 994780 145564 994792
rect 145616 994780 145622 994832
rect 155954 994820 155960 994832
rect 151786 994792 155960 994820
rect 80146 994712 80152 994764
rect 80204 994752 80210 994764
rect 101398 994752 101404 994764
rect 80204 994724 101404 994752
rect 80204 994712 80210 994724
rect 101398 994712 101404 994724
rect 101456 994712 101462 994764
rect 132402 994644 132408 994696
rect 132460 994684 132466 994696
rect 149698 994684 149704 994696
rect 132460 994656 149704 994684
rect 132460 994644 132466 994656
rect 149698 994644 149704 994656
rect 149756 994644 149762 994696
rect 81342 994576 81348 994628
rect 81400 994616 81406 994628
rect 98638 994616 98644 994628
rect 81400 994588 98644 994616
rect 81400 994576 81406 994588
rect 98638 994576 98644 994588
rect 98696 994576 98702 994628
rect 131574 994508 131580 994560
rect 131632 994548 131638 994560
rect 151786 994548 151814 994792
rect 155954 994780 155960 994792
rect 156012 994780 156018 994832
rect 131632 994520 151814 994548
rect 180490 994548 180518 994928
rect 183278 994916 183284 994968
rect 183336 994956 183342 994968
rect 205634 994956 205640 994968
rect 183336 994928 205640 994956
rect 183336 994916 183342 994928
rect 205634 994916 205640 994928
rect 205692 994916 205698 994968
rect 229186 994916 229192 994968
rect 229244 994956 229250 994968
rect 234402 994956 234430 995064
rect 234706 995052 234712 995064
rect 234764 995052 234770 995104
rect 398834 995092 398840 995104
rect 393286 995064 398840 995092
rect 358722 994984 358728 995036
rect 358780 995024 358786 995036
rect 393286 995024 393314 995064
rect 398834 995052 398840 995064
rect 398892 995052 398898 995104
rect 358780 994996 393314 995024
rect 358780 994984 358786 994996
rect 229244 994928 234430 994956
rect 229244 994916 229250 994928
rect 234522 994916 234528 994968
rect 234580 994956 234586 994968
rect 259454 994956 259460 994968
rect 234580 994928 259460 994956
rect 234580 994916 234586 994928
rect 259454 994916 259460 994928
rect 259512 994916 259518 994968
rect 286502 994916 286508 994968
rect 286560 994956 286566 994968
rect 300302 994956 300308 994968
rect 286560 994928 300308 994956
rect 286560 994916 286566 994928
rect 300302 994916 300308 994928
rect 300360 994916 300366 994968
rect 396994 994916 397000 994968
rect 397052 994956 397058 994968
rect 402808 994956 402836 995336
rect 402974 995324 402980 995336
rect 403032 995324 403038 995376
rect 471422 995256 471428 995308
rect 471480 995296 471486 995308
rect 480226 995296 480254 995404
rect 509234 995392 509240 995404
rect 509292 995392 509298 995444
rect 509878 995392 509884 995444
rect 509936 995432 509942 995444
rect 560294 995432 560300 995444
rect 509936 995404 560300 995432
rect 509936 995392 509942 995404
rect 560294 995392 560300 995404
rect 560352 995392 560358 995444
rect 620278 995392 620284 995444
rect 620336 995432 620342 995444
rect 630646 995432 630674 995472
rect 620336 995404 630674 995432
rect 620336 995392 620342 995404
rect 630784 995364 630812 995472
rect 639506 995364 639512 995376
rect 630784 995336 639512 995364
rect 639506 995324 639512 995336
rect 639564 995324 639570 995376
rect 471480 995268 480254 995296
rect 471480 995256 471486 995268
rect 505738 995256 505744 995308
rect 505796 995296 505802 995308
rect 532142 995296 532148 995308
rect 505796 995268 532148 995296
rect 505796 995256 505802 995268
rect 532142 995256 532148 995268
rect 532200 995256 532206 995308
rect 567194 995256 567200 995308
rect 567252 995296 567258 995308
rect 630582 995296 630588 995308
rect 567252 995268 630588 995296
rect 567252 995256 567258 995268
rect 630582 995256 630588 995268
rect 630640 995256 630646 995308
rect 489730 995188 489736 995240
rect 489788 995228 489794 995240
rect 489788 995200 489914 995228
rect 489788 995188 489794 995200
rect 472250 995120 472256 995172
rect 472308 995160 472314 995172
rect 477678 995160 477684 995172
rect 472308 995132 477684 995160
rect 472308 995120 472314 995132
rect 477678 995120 477684 995132
rect 477736 995120 477742 995172
rect 397052 994928 402836 994956
rect 397052 994916 397058 994928
rect 429838 994916 429844 994968
rect 429896 994956 429902 994968
rect 489886 994956 489914 995200
rect 523310 995120 523316 995172
rect 523368 995160 523374 995172
rect 526070 995160 526076 995172
rect 523368 995132 526076 995160
rect 523368 995120 523374 995132
rect 526070 995120 526076 995132
rect 526128 995120 526134 995172
rect 526254 995120 526260 995172
rect 526312 995160 526318 995172
rect 529014 995160 529020 995172
rect 526312 995132 529020 995160
rect 526312 995120 526318 995132
rect 529014 995120 529020 995132
rect 529072 995120 529078 995172
rect 556798 995120 556804 995172
rect 556856 995160 556862 995172
rect 640702 995160 640708 995172
rect 556856 995132 640708 995160
rect 556856 995120 556862 995132
rect 640702 995120 640708 995132
rect 640760 995120 640766 995172
rect 534074 995092 534080 995104
rect 532896 995064 534080 995092
rect 500678 994984 500684 995036
rect 500736 995024 500742 995036
rect 528738 995024 528744 995036
rect 500736 994996 528744 995024
rect 500736 994984 500742 994996
rect 528738 994984 528744 994996
rect 528796 994984 528802 995036
rect 429896 994928 489914 994956
rect 429896 994916 429902 994928
rect 359550 994848 359556 994900
rect 359608 994888 359614 994900
rect 393958 994888 393964 994900
rect 359608 994860 393964 994888
rect 359608 994848 359614 994860
rect 393958 994848 393964 994860
rect 394016 994848 394022 994900
rect 520550 994848 520556 994900
rect 520608 994888 520614 994900
rect 532896 994888 532924 995064
rect 534074 995052 534080 995064
rect 534132 995052 534138 995104
rect 550634 994984 550640 995036
rect 550692 995024 550698 995036
rect 635826 995024 635832 995036
rect 550692 994996 635832 995024
rect 550692 994984 550698 994996
rect 635826 994984 635832 994996
rect 635884 994984 635890 995036
rect 638678 995024 638684 995036
rect 636028 994996 638684 995024
rect 533062 994916 533068 994968
rect 533120 994956 533126 994968
rect 537846 994956 537852 994968
rect 533120 994928 537852 994956
rect 533120 994916 533126 994928
rect 537846 994916 537852 994928
rect 537904 994916 537910 994968
rect 520608 994860 532924 994888
rect 520608 994848 520614 994860
rect 550358 994848 550364 994900
rect 550416 994888 550422 994900
rect 625798 994888 625804 994900
rect 550416 994860 625804 994888
rect 550416 994848 550422 994860
rect 625798 994848 625804 994860
rect 625856 994848 625862 994900
rect 630766 994848 630772 994900
rect 630824 994888 630830 994900
rect 636028 994888 636056 994996
rect 638678 994984 638684 994996
rect 638736 994984 638742 995036
rect 640794 994956 640800 994968
rect 640306 994928 640800 994956
rect 630824 994860 636056 994888
rect 630824 994848 630830 994860
rect 638494 994848 638500 994900
rect 638552 994888 638558 994900
rect 640306 994888 640334 994928
rect 640794 994916 640800 994928
rect 640852 994916 640858 994968
rect 638552 994860 640334 994888
rect 638552 994848 638558 994860
rect 180610 994780 180616 994832
rect 180668 994820 180674 994832
rect 192846 994820 192852 994832
rect 180668 994792 192852 994820
rect 180668 994780 180674 994792
rect 192846 994780 192852 994792
rect 192904 994780 192910 994832
rect 195238 994780 195244 994832
rect 195296 994820 195302 994832
rect 207014 994820 207020 994832
rect 195296 994792 207020 994820
rect 195296 994780 195302 994792
rect 207014 994780 207020 994792
rect 207072 994780 207078 994832
rect 231578 994780 231584 994832
rect 231636 994820 231642 994832
rect 255958 994820 255964 994832
rect 231636 994792 255964 994820
rect 231636 994780 231642 994792
rect 255958 994780 255964 994792
rect 256016 994780 256022 994832
rect 305638 994820 305644 994832
rect 289648 994792 305644 994820
rect 180610 994644 180616 994696
rect 180668 994684 180674 994696
rect 204898 994684 204904 994696
rect 180668 994656 204904 994684
rect 180668 994644 180674 994656
rect 204898 994644 204904 994656
rect 204956 994644 204962 994696
rect 232866 994644 232872 994696
rect 232924 994684 232930 994696
rect 257338 994684 257344 994696
rect 232924 994656 257344 994684
rect 232924 994644 232930 994656
rect 257338 994644 257344 994656
rect 257396 994644 257402 994696
rect 285950 994644 285956 994696
rect 286008 994684 286014 994696
rect 289446 994684 289452 994696
rect 286008 994656 289452 994684
rect 286008 994644 286014 994656
rect 289446 994644 289452 994656
rect 289504 994644 289510 994696
rect 195238 994548 195244 994560
rect 180490 994520 195244 994548
rect 131632 994508 131638 994520
rect 195238 994508 195244 994520
rect 195296 994508 195302 994560
rect 229002 994508 229008 994560
rect 229060 994548 229066 994560
rect 239398 994548 239404 994560
rect 229060 994520 239404 994548
rect 229060 994508 229066 994520
rect 239398 994508 239404 994520
rect 239456 994508 239462 994560
rect 283466 994508 283472 994560
rect 283524 994548 283530 994560
rect 289648 994548 289676 994792
rect 305638 994780 305644 994792
rect 305696 994780 305702 994832
rect 460198 994780 460204 994832
rect 460256 994820 460262 994832
rect 485958 994820 485964 994832
rect 460256 994792 485964 994820
rect 460256 994780 460262 994792
rect 485958 994780 485964 994792
rect 486016 994780 486022 994832
rect 486602 994780 486608 994832
rect 486660 994820 486666 994832
rect 489730 994820 489736 994832
rect 486660 994792 489736 994820
rect 486660 994780 486666 994792
rect 489730 994780 489736 994792
rect 489788 994780 489794 994832
rect 371878 994712 371884 994764
rect 371936 994752 371942 994764
rect 388070 994752 388076 994764
rect 371936 994724 388076 994752
rect 371936 994712 371942 994724
rect 388070 994712 388076 994724
rect 388128 994712 388134 994764
rect 388254 994712 388260 994764
rect 388312 994752 388318 994764
rect 393314 994752 393320 994764
rect 388312 994724 393320 994752
rect 388312 994712 388318 994724
rect 393314 994712 393320 994724
rect 393372 994712 393378 994764
rect 502978 994712 502984 994764
rect 503036 994752 503042 994764
rect 538214 994752 538220 994764
rect 503036 994724 538220 994752
rect 503036 994712 503042 994724
rect 538214 994712 538220 994724
rect 538272 994712 538278 994764
rect 571978 994712 571984 994764
rect 572036 994752 572042 994764
rect 635182 994752 635188 994764
rect 572036 994724 635188 994752
rect 572036 994712 572042 994724
rect 635182 994712 635188 994724
rect 635240 994712 635246 994764
rect 311894 994684 311900 994696
rect 283524 994520 289676 994548
rect 291764 994656 311900 994684
rect 283524 994508 283530 994520
rect 81986 994440 81992 994492
rect 82044 994480 82050 994492
rect 93118 994480 93124 994492
rect 82044 994452 93124 994480
rect 82044 994440 82050 994452
rect 93118 994440 93124 994452
rect 93176 994440 93182 994492
rect 192846 994372 192852 994424
rect 192904 994412 192910 994424
rect 202138 994412 202144 994424
rect 192904 994384 202144 994412
rect 192904 994372 192910 994384
rect 202138 994372 202144 994384
rect 202196 994372 202202 994424
rect 207014 994372 207020 994424
rect 207072 994412 207078 994424
rect 213914 994412 213920 994424
rect 207072 994384 213920 994412
rect 207072 994372 207078 994384
rect 213914 994372 213920 994384
rect 213972 994372 213978 994424
rect 232222 994372 232228 994424
rect 232280 994412 232286 994424
rect 250438 994412 250444 994424
rect 232280 994384 250444 994412
rect 232280 994372 232286 994384
rect 250438 994372 250444 994384
rect 250496 994372 250502 994424
rect 282822 994372 282828 994424
rect 282880 994412 282886 994424
rect 291764 994412 291792 994656
rect 311894 994644 311900 994656
rect 311952 994644 311958 994696
rect 469858 994644 469864 994696
rect 469916 994684 469922 994696
rect 481358 994684 481364 994696
rect 469916 994656 481364 994684
rect 469916 994644 469922 994656
rect 481358 994644 481364 994656
rect 481416 994644 481422 994696
rect 362218 994576 362224 994628
rect 362276 994616 362282 994628
rect 393498 994616 393504 994628
rect 362276 994588 393504 994616
rect 362276 994576 362282 994588
rect 393498 994576 393504 994588
rect 393556 994576 393562 994628
rect 502242 994576 502248 994628
rect 502300 994616 502306 994628
rect 539226 994616 539232 994628
rect 502300 994588 539232 994616
rect 502300 994576 502306 994588
rect 539226 994576 539232 994588
rect 539284 994576 539290 994628
rect 625798 994576 625804 994628
rect 625856 994616 625862 994628
rect 637022 994616 637028 994628
rect 625856 994588 637028 994616
rect 625856 994576 625862 994588
rect 637022 994576 637028 994588
rect 637080 994576 637086 994628
rect 282880 994384 291792 994412
rect 291856 994520 296714 994548
rect 282880 994372 282886 994384
rect 140130 994236 140136 994288
rect 140188 994276 140194 994288
rect 186498 994276 186504 994288
rect 140188 994248 186504 994276
rect 140188 994236 140194 994248
rect 186498 994236 186504 994248
rect 186556 994236 186562 994288
rect 191834 994236 191840 994288
rect 191892 994276 191898 994288
rect 251450 994276 251456 994288
rect 191892 994248 251456 994276
rect 191892 994236 191898 994248
rect 251450 994236 251456 994248
rect 251508 994236 251514 994288
rect 284110 994236 284116 994288
rect 284168 994276 284174 994288
rect 291856 994276 291884 994520
rect 296686 994412 296714 994520
rect 301498 994508 301504 994560
rect 301556 994548 301562 994560
rect 309778 994548 309784 994560
rect 301556 994520 309784 994548
rect 301556 994508 301562 994520
rect 309778 994508 309784 994520
rect 309836 994508 309842 994560
rect 563698 994508 563704 994560
rect 563756 994548 563762 994560
rect 624602 994548 624608 994560
rect 563756 994520 624608 994548
rect 563756 994508 563762 994520
rect 624602 994508 624608 994520
rect 624660 994508 624666 994560
rect 380894 994440 380900 994492
rect 380952 994480 380958 994492
rect 388254 994480 388260 994492
rect 380952 994452 388260 994480
rect 380952 994440 380958 994452
rect 388254 994440 388260 994452
rect 388312 994440 388318 994492
rect 397638 994480 397644 994492
rect 388456 994452 397644 994480
rect 308398 994412 308404 994424
rect 296686 994384 308404 994412
rect 308398 994372 308404 994384
rect 308456 994372 308462 994424
rect 388456 994344 388484 994452
rect 397638 994440 397644 994452
rect 397696 994440 397702 994492
rect 402974 994480 402980 994492
rect 402946 994440 402980 994480
rect 403032 994440 403038 994492
rect 497918 994440 497924 994492
rect 497976 994480 497982 994492
rect 538030 994480 538036 994492
rect 497976 994452 538036 994480
rect 497976 994440 497982 994452
rect 538030 994440 538036 994452
rect 538088 994440 538094 994492
rect 383626 994316 388484 994344
rect 284168 994248 291884 994276
rect 284168 994236 284174 994248
rect 357342 994236 357348 994288
rect 357400 994276 357406 994288
rect 381170 994276 381176 994288
rect 357400 994248 381176 994276
rect 357400 994236 357406 994248
rect 381170 994236 381176 994248
rect 381228 994236 381234 994288
rect 184474 994100 184480 994152
rect 184532 994140 184538 994152
rect 196618 994140 196624 994152
rect 184532 994112 196624 994140
rect 184532 994100 184538 994112
rect 196618 994100 196624 994112
rect 196676 994100 196682 994152
rect 239398 994100 239404 994152
rect 239456 994140 239462 994152
rect 249058 994140 249064 994152
rect 239456 994112 249064 994140
rect 239456 994100 239462 994112
rect 249058 994100 249064 994112
rect 249116 994100 249122 994152
rect 265618 994100 265624 994152
rect 265676 994140 265682 994152
rect 267734 994140 267740 994152
rect 265676 994112 267740 994140
rect 265676 994100 265682 994112
rect 267734 994100 267740 994112
rect 267792 994100 267798 994152
rect 289446 994100 289452 994152
rect 289504 994140 289510 994152
rect 301498 994140 301504 994152
rect 289504 994112 301504 994140
rect 289504 994100 289510 994112
rect 301498 994100 301504 994112
rect 301556 994100 301562 994152
rect 378594 994100 378600 994152
rect 378652 994140 378658 994152
rect 383626 994140 383654 994316
rect 388070 994168 388076 994220
rect 388128 994208 388134 994220
rect 402946 994208 402974 994440
rect 549162 994372 549168 994424
rect 549220 994412 549226 994424
rect 667106 994412 667112 994424
rect 549220 994384 667112 994412
rect 549220 994372 549226 994384
rect 667106 994372 667112 994384
rect 667164 994372 667170 994424
rect 426434 994236 426440 994288
rect 426492 994276 426498 994288
rect 446122 994276 446128 994288
rect 426492 994248 446128 994276
rect 426492 994236 426498 994248
rect 446122 994236 446128 994248
rect 446180 994236 446186 994288
rect 547782 994236 547788 994288
rect 547840 994276 547846 994288
rect 666554 994276 666560 994288
rect 547840 994248 666560 994276
rect 547840 994236 547846 994248
rect 666554 994236 666560 994248
rect 666612 994236 666618 994288
rect 388128 994180 402974 994208
rect 388128 994168 388134 994180
rect 378652 994112 383654 994140
rect 378652 994100 378658 994112
rect 240042 993964 240048 994016
rect 240100 994004 240106 994016
rect 246206 994004 246212 994016
rect 240100 993976 246212 994004
rect 240100 993964 240106 993976
rect 246206 993964 246212 993976
rect 246264 993964 246270 994016
rect 496722 993284 496728 993336
rect 496780 993324 496786 993336
rect 666922 993324 666928 993336
rect 496780 993296 666928 993324
rect 496780 993284 496786 993296
rect 666922 993284 666928 993296
rect 666980 993284 666986 993336
rect 280706 993148 280712 993200
rect 280764 993188 280770 993200
rect 316402 993188 316408 993200
rect 280764 993160 316408 993188
rect 280764 993148 280770 993160
rect 316402 993148 316408 993160
rect 316460 993148 316466 993200
rect 351822 993148 351828 993200
rect 351880 993188 351886 993200
rect 665174 993188 665180 993200
rect 351880 993160 665180 993188
rect 351880 993148 351886 993160
rect 665174 993148 665180 993160
rect 665232 993148 665238 993200
rect 51718 993012 51724 993064
rect 51776 993052 51782 993064
rect 107746 993052 107752 993064
rect 51776 993024 107752 993052
rect 51776 993012 51782 993024
rect 107746 993012 107752 993024
rect 107804 993012 107810 993064
rect 147582 993012 147588 993064
rect 147640 993052 147646 993064
rect 649994 993052 650000 993064
rect 147640 993024 650000 993052
rect 147640 993012 147646 993024
rect 649994 993012 650000 993024
rect 650052 993012 650058 993064
rect 46198 992876 46204 992928
rect 46256 992916 46262 992928
rect 108114 992916 108120 992928
rect 46256 992888 108120 992916
rect 46256 992876 46262 992888
rect 108114 992876 108120 992888
rect 108172 992876 108178 992928
rect 148962 992876 148968 992928
rect 149020 992916 149026 992928
rect 651374 992916 651380 992928
rect 149020 992888 651380 992916
rect 149020 992876 149026 992888
rect 651374 992876 651380 992888
rect 651432 992876 651438 992928
rect 512638 991856 512644 991908
rect 512696 991896 512702 991908
rect 527634 991896 527640 991908
rect 512696 991868 527640 991896
rect 512696 991856 512702 991868
rect 527634 991856 527640 991868
rect 527692 991856 527698 991908
rect 266998 991720 267004 991772
rect 267056 991760 267062 991772
rect 284294 991760 284300 991772
rect 267056 991732 284300 991760
rect 267056 991720 267062 991732
rect 284294 991720 284300 991732
rect 284352 991720 284358 991772
rect 367738 991720 367744 991772
rect 367796 991760 367802 991772
rect 415026 991760 415032 991772
rect 367796 991732 415032 991760
rect 367796 991720 367802 991732
rect 415026 991720 415032 991732
rect 415084 991720 415090 991772
rect 419442 991720 419448 991772
rect 419500 991760 419506 991772
rect 668026 991760 668032 991772
rect 419500 991732 668032 991760
rect 419500 991720 419506 991732
rect 668026 991720 668032 991732
rect 668084 991720 668090 991772
rect 73430 991584 73436 991636
rect 73488 991624 73494 991636
rect 112070 991624 112076 991636
rect 73488 991596 112076 991624
rect 73488 991584 73494 991596
rect 112070 991584 112076 991596
rect 112128 991584 112134 991636
rect 200022 991584 200028 991636
rect 200080 991624 200086 991636
rect 651742 991624 651748 991636
rect 200080 991596 651748 991624
rect 200080 991584 200086 991596
rect 651742 991584 651748 991596
rect 651800 991584 651806 991636
rect 50338 991448 50344 991500
rect 50396 991488 50402 991500
rect 110414 991488 110420 991500
rect 50396 991460 110420 991488
rect 50396 991448 50402 991460
rect 110414 991448 110420 991460
rect 110472 991448 110478 991500
rect 138290 991448 138296 991500
rect 138348 991488 138354 991500
rect 162854 991488 162860 991500
rect 138348 991460 162860 991488
rect 138348 991448 138354 991460
rect 162854 991448 162860 991460
rect 162912 991448 162918 991500
rect 198642 991448 198648 991500
rect 198700 991488 198706 991500
rect 650730 991488 650736 991500
rect 198700 991460 650736 991488
rect 198700 991448 198706 991460
rect 650730 991448 650736 991460
rect 650788 991448 650794 991500
rect 562502 990496 562508 990548
rect 562560 990536 562566 990548
rect 672718 990536 672724 990548
rect 562560 990508 672724 990536
rect 562560 990496 562566 990508
rect 672718 990496 672724 990508
rect 672776 990496 672782 990548
rect 435358 990360 435364 990412
rect 435416 990400 435422 990412
rect 463602 990400 463608 990412
rect 435416 990372 463608 990400
rect 435416 990360 435422 990372
rect 463602 990360 463608 990372
rect 463660 990360 463666 990412
rect 498102 990360 498108 990412
rect 498160 990400 498166 990412
rect 666738 990400 666744 990412
rect 498160 990372 666744 990400
rect 498160 990360 498166 990372
rect 666738 990360 666744 990372
rect 666796 990360 666802 990412
rect 303522 990224 303528 990276
rect 303580 990264 303586 990276
rect 665450 990264 665456 990276
rect 303580 990236 665456 990264
rect 303580 990224 303586 990236
rect 665450 990224 665456 990236
rect 665508 990224 665514 990276
rect 48958 990088 48964 990140
rect 49016 990128 49022 990140
rect 109034 990128 109040 990140
rect 49016 990100 109040 990128
rect 49016 990088 49022 990100
rect 109034 990088 109040 990100
rect 109092 990088 109098 990140
rect 249702 990088 249708 990140
rect 249760 990128 249766 990140
rect 648890 990128 648896 990140
rect 249760 990100 648896 990128
rect 249760 990088 249766 990100
rect 648890 990088 648896 990100
rect 648948 990088 648954 990140
rect 422202 988864 422208 988916
rect 422260 988904 422266 988916
rect 668210 988904 668216 988916
rect 422260 988876 668216 988904
rect 422260 988864 422266 988876
rect 668210 988864 668216 988876
rect 668268 988864 668274 988916
rect 250990 988728 250996 988780
rect 251048 988768 251054 988780
rect 650178 988768 650184 988780
rect 251048 988740 650184 988768
rect 251048 988728 251054 988740
rect 650178 988728 650184 988740
rect 650236 988728 650242 988780
rect 559558 987640 559564 987692
rect 559616 987680 559622 987692
rect 669958 987680 669964 987692
rect 559616 987652 669964 987680
rect 559616 987640 559622 987652
rect 669958 987640 669964 987652
rect 670016 987640 670022 987692
rect 352834 987504 352840 987556
rect 352892 987544 352898 987556
rect 668394 987544 668400 987556
rect 352892 987516 668400 987544
rect 352892 987504 352898 987516
rect 668394 987504 668400 987516
rect 668452 987504 668458 987556
rect 96338 987368 96344 987420
rect 96396 987408 96402 987420
rect 650914 987408 650920 987420
rect 96396 987380 650920 987408
rect 96396 987368 96402 987380
rect 650914 987368 650920 987380
rect 650972 987368 650978 987420
rect 203150 986620 203156 986672
rect 203208 986660 203214 986672
rect 207014 986660 207020 986672
rect 203208 986632 207020 986660
rect 203208 986620 203214 986632
rect 207014 986620 207020 986632
rect 207072 986620 207078 986672
rect 217318 986620 217324 986672
rect 217376 986660 217382 986672
rect 219434 986660 219440 986672
rect 217376 986632 219440 986660
rect 217376 986620 217382 986632
rect 219434 986620 219440 986632
rect 219492 986620 219498 986672
rect 570598 986212 570604 986264
rect 570656 986252 570662 986264
rect 592494 986252 592500 986264
rect 570656 986224 592500 986252
rect 570656 986212 570662 986224
rect 592494 986212 592500 986224
rect 592552 986212 592558 986264
rect 370498 986076 370504 986128
rect 370556 986116 370562 986128
rect 397822 986116 397828 986128
rect 370556 986088 397828 986116
rect 370556 986076 370562 986088
rect 397822 986076 397828 986088
rect 397880 986076 397886 986128
rect 463602 986076 463608 986128
rect 463660 986116 463666 986128
rect 478966 986116 478972 986128
rect 463660 986088 478972 986116
rect 463660 986076 463666 986088
rect 478966 986076 478972 986088
rect 479024 986076 479030 986128
rect 519538 986076 519544 986128
rect 519596 986116 519602 986128
rect 543826 986116 543832 986128
rect 519596 986088 543832 986116
rect 519596 986076 519602 986088
rect 543826 986076 543832 986088
rect 543884 986076 543890 986128
rect 565078 986076 565084 986128
rect 565136 986116 565142 986128
rect 608778 986116 608784 986128
rect 565136 986088 608784 986116
rect 565136 986076 565142 986088
rect 608778 986076 608784 986088
rect 608836 986076 608842 986128
rect 89622 985940 89628 985992
rect 89680 985980 89686 985992
rect 106918 985980 106924 985992
rect 89680 985952 106924 985980
rect 89680 985940 89686 985952
rect 106918 985940 106924 985952
rect 106976 985940 106982 985992
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 279418 985940 279424 985992
rect 279476 985980 279482 985992
rect 300486 985980 300492 985992
rect 279476 985952 300492 985980
rect 279476 985940 279482 985952
rect 300486 985940 300492 985952
rect 300544 985940 300550 985992
rect 369118 985940 369124 985992
rect 369176 985980 369182 985992
rect 414106 985980 414112 985992
rect 369176 985952 414112 985980
rect 369176 985940 369182 985952
rect 414106 985940 414112 985952
rect 414164 985940 414170 985992
rect 415026 985940 415032 985992
rect 415084 985980 415090 985992
rect 430298 985980 430304 985992
rect 415084 985952 430304 985980
rect 415084 985940 415090 985952
rect 430298 985940 430304 985952
rect 430356 985940 430362 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 462774 985980 462780 985992
rect 436796 985952 462780 985980
rect 436796 985940 436802 985952
rect 462774 985940 462780 985952
rect 462832 985940 462838 985992
rect 465718 985940 465724 985992
rect 465776 985980 465782 985992
rect 495158 985980 495164 985992
rect 465776 985952 495164 985980
rect 465776 985940 465782 985952
rect 495158 985940 495164 985952
rect 495216 985940 495222 985992
rect 515398 985940 515404 985992
rect 515456 985980 515462 985992
rect 560110 985980 560116 985992
rect 515456 985952 560116 985980
rect 515456 985940 515462 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 562318 985940 562324 985992
rect 562376 985980 562382 985992
rect 658918 985980 658924 985992
rect 562376 985952 658924 985980
rect 562376 985940 562382 985952
rect 658918 985940 658924 985952
rect 658976 985940 658982 985992
rect 560938 984852 560944 984904
rect 560996 984892 561002 984904
rect 660298 984892 660304 984904
rect 560996 984864 660304 984892
rect 560996 984852 561002 984864
rect 660298 984852 660304 984864
rect 660356 984852 660362 984904
rect 302142 984716 302148 984768
rect 302200 984756 302206 984768
rect 665634 984756 665640 984768
rect 302200 984728 665640 984756
rect 302200 984716 302206 984728
rect 665634 984716 665640 984728
rect 665692 984716 665698 984768
rect 96522 984580 96528 984632
rect 96580 984620 96586 984632
rect 650362 984620 650368 984632
rect 96580 984592 650368 984620
rect 96580 984580 96586 984592
rect 650362 984580 650368 984592
rect 650420 984580 650426 984632
rect 55858 975672 55864 975724
rect 55916 975712 55922 975724
rect 62114 975712 62120 975724
rect 55916 975684 62120 975712
rect 55916 975672 55922 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651558 975672 651564 975724
rect 651616 975712 651622 975724
rect 661678 975712 661684 975724
rect 651616 975684 661684 975712
rect 651616 975672 651622 975684
rect 661678 975672 661684 975684
rect 661736 975672 661742 975724
rect 42518 969416 42524 969468
rect 42576 969456 42582 969468
rect 55858 969456 55864 969468
rect 42576 969428 55864 969456
rect 42576 969416 42582 969428
rect 55858 969416 55864 969428
rect 55916 969416 55922 969468
rect 42242 966832 42248 966884
rect 42300 966872 42306 966884
rect 42702 966872 42708 966884
rect 42300 966844 42708 966872
rect 42300 966832 42306 966844
rect 42702 966832 42708 966844
rect 42760 966832 42766 966884
rect 673362 966152 673368 966204
rect 673420 966192 673426 966204
rect 675110 966192 675116 966204
rect 673420 966164 675116 966192
rect 673420 966152 673426 966164
rect 675110 966152 675116 966164
rect 675168 966152 675174 966204
rect 42426 964656 42432 964708
rect 42484 964696 42490 964708
rect 42886 964696 42892 964708
rect 42484 964668 42892 964696
rect 42484 964656 42490 964668
rect 42886 964656 42892 964668
rect 42944 964656 42950 964708
rect 42426 963840 42432 963892
rect 42484 963880 42490 963892
rect 44174 963880 44180 963892
rect 42484 963852 44180 963880
rect 42484 963840 42490 963852
rect 44174 963840 44180 963852
rect 44232 963840 44238 963892
rect 42426 963432 42432 963484
rect 42484 963472 42490 963484
rect 43070 963472 43076 963484
rect 42484 963444 43076 963472
rect 42484 963432 42490 963444
rect 43070 963432 43076 963444
rect 43128 963432 43134 963484
rect 42426 961868 42432 961920
rect 42484 961908 42490 961920
rect 44450 961908 44456 961920
rect 42484 961880 44456 961908
rect 42484 961868 42490 961880
rect 44450 961868 44456 961880
rect 44508 961868 44514 961920
rect 47578 961868 47584 961920
rect 47636 961908 47642 961920
rect 62114 961908 62120 961920
rect 47636 961880 62120 961908
rect 47636 961868 47642 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 651558 961868 651564 961920
rect 651616 961908 651622 961920
rect 663058 961908 663064 961920
rect 651616 961880 663064 961908
rect 651616 961868 651622 961880
rect 663058 961868 663064 961880
rect 663116 961868 663122 961920
rect 674282 961868 674288 961920
rect 674340 961908 674346 961920
rect 675110 961908 675116 961920
rect 674340 961880 675116 961908
rect 674340 961868 674346 961880
rect 675110 961868 675116 961880
rect 675168 961868 675174 961920
rect 42426 959080 42432 959132
rect 42484 959120 42490 959132
rect 43254 959120 43260 959132
rect 42484 959092 43260 959120
rect 42484 959080 42490 959092
rect 43254 959080 43260 959092
rect 43312 959080 43318 959132
rect 42426 958264 42432 958316
rect 42484 958304 42490 958316
rect 44634 958304 44640 958316
rect 42484 958276 44640 958304
rect 42484 958264 42490 958276
rect 44634 958264 44640 958276
rect 44692 958264 44698 958316
rect 674466 957856 674472 957908
rect 674524 957896 674530 957908
rect 675110 957896 675116 957908
rect 674524 957868 675116 957896
rect 674524 957856 674530 957868
rect 675110 957856 675116 957868
rect 675168 957856 675174 957908
rect 660482 957720 660488 957772
rect 660540 957760 660546 957772
rect 660540 957732 675340 957760
rect 660540 957720 660546 957732
rect 675312 957364 675340 957732
rect 675294 957312 675300 957364
rect 675352 957312 675358 957364
rect 673178 956360 673184 956412
rect 673236 956400 673242 956412
rect 675110 956400 675116 956412
rect 673236 956372 675116 956400
rect 673236 956360 673242 956372
rect 675110 956360 675116 956372
rect 675168 956360 675174 956412
rect 35158 951464 35164 951516
rect 35216 951504 35222 951516
rect 41690 951504 41696 951516
rect 35216 951476 41696 951504
rect 35216 951464 35222 951476
rect 41690 951464 41696 951476
rect 41748 951464 41754 951516
rect 675846 949424 675852 949476
rect 675904 949464 675910 949476
rect 678238 949464 678244 949476
rect 675904 949436 678244 949464
rect 675904 949424 675910 949436
rect 678238 949424 678244 949436
rect 678296 949424 678302 949476
rect 675846 948744 675852 948796
rect 675904 948784 675910 948796
rect 682378 948784 682384 948796
rect 675904 948756 682384 948784
rect 675904 948744 675910 948756
rect 682378 948744 682384 948756
rect 682436 948744 682442 948796
rect 651558 948064 651564 948116
rect 651616 948104 651622 948116
rect 671338 948104 671344 948116
rect 651616 948076 671344 948104
rect 651616 948064 651622 948076
rect 671338 948064 671344 948076
rect 671396 948064 671402 948116
rect 43530 945956 43536 946008
rect 43588 945996 43594 946008
rect 62114 945996 62120 946008
rect 43588 945968 62120 945996
rect 43588 945956 43594 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 663058 941808 663064 941860
rect 663116 941848 663122 941860
rect 675478 941848 675484 941860
rect 663116 941820 675484 941848
rect 663116 941808 663122 941820
rect 675478 941808 675484 941820
rect 675536 941808 675542 941860
rect 41322 941468 41328 941520
rect 41380 941508 41386 941520
rect 41690 941508 41696 941520
rect 41380 941480 41696 941508
rect 41380 941468 41386 941480
rect 41690 941468 41696 941480
rect 41748 941468 41754 941520
rect 43622 941332 43628 941384
rect 43680 941372 43686 941384
rect 48958 941372 48964 941384
rect 43680 941344 48964 941372
rect 43680 941332 43686 941344
rect 48958 941332 48964 941344
rect 49016 941332 49022 941384
rect 43438 941196 43444 941248
rect 43496 941236 43502 941248
rect 50338 941236 50344 941248
rect 43496 941208 50344 941236
rect 43496 941196 43502 941208
rect 50338 941196 50344 941208
rect 50396 941196 50402 941248
rect 40954 940108 40960 940160
rect 41012 940148 41018 940160
rect 41690 940148 41696 940160
rect 41012 940120 41696 940148
rect 41012 940108 41018 940120
rect 41690 940108 41696 940120
rect 41748 940108 41754 940160
rect 43438 939768 43444 939820
rect 43496 939808 43502 939820
rect 51718 939808 51724 939820
rect 43496 939780 51724 939808
rect 43496 939768 43502 939780
rect 51718 939768 51724 939780
rect 51776 939768 51782 939820
rect 672718 938680 672724 938732
rect 672776 938720 672782 938732
rect 675478 938720 675484 938732
rect 672776 938692 675484 938720
rect 672776 938680 672782 938692
rect 675478 938680 675484 938692
rect 675536 938680 675542 938732
rect 40954 938544 40960 938596
rect 41012 938584 41018 938596
rect 41506 938584 41512 938596
rect 41012 938556 41512 938584
rect 41012 938544 41018 938556
rect 41506 938544 41512 938556
rect 41564 938544 41570 938596
rect 671338 938544 671344 938596
rect 671396 938584 671402 938596
rect 675294 938584 675300 938596
rect 671396 938556 675300 938584
rect 671396 938544 671402 938556
rect 675294 938544 675300 938556
rect 675352 938544 675358 938596
rect 41138 938408 41144 938460
rect 41196 938448 41202 938460
rect 41506 938448 41512 938460
rect 41196 938420 41512 938448
rect 41196 938408 41202 938420
rect 41506 938408 41512 938420
rect 41564 938408 41570 938460
rect 661678 938408 661684 938460
rect 661736 938448 661742 938460
rect 674926 938448 674932 938460
rect 661736 938420 674932 938448
rect 661736 938408 661742 938420
rect 674926 938408 674932 938420
rect 674984 938408 674990 938460
rect 671522 937524 671528 937576
rect 671580 937564 671586 937576
rect 675478 937564 675484 937576
rect 671580 937536 675484 937564
rect 671580 937524 671586 937536
rect 675478 937524 675484 937536
rect 675536 937524 675542 937576
rect 660298 937320 660304 937372
rect 660356 937360 660362 937372
rect 675478 937360 675484 937372
rect 660356 937332 675484 937360
rect 660356 937320 660362 937332
rect 675478 937320 675484 937332
rect 675536 937320 675542 937372
rect 658918 937184 658924 937236
rect 658976 937224 658982 937236
rect 674926 937224 674932 937236
rect 658976 937196 674932 937224
rect 658976 937184 658982 937196
rect 674926 937184 674932 937196
rect 674984 937184 674990 937236
rect 671154 937048 671160 937100
rect 671212 937088 671218 937100
rect 675294 937088 675300 937100
rect 671212 937060 675300 937088
rect 671212 937048 671218 937060
rect 675294 937048 675300 937060
rect 675352 937048 675358 937100
rect 44634 936980 44640 937032
rect 44692 937020 44698 937032
rect 62114 937020 62120 937032
rect 44692 936992 62120 937020
rect 44692 936980 44698 936992
rect 62114 936980 62120 936992
rect 62172 936980 62178 937032
rect 651558 936980 651564 937032
rect 651616 937020 651622 937032
rect 660482 937020 660488 937032
rect 651616 936992 660488 937020
rect 651616 936980 651622 936992
rect 660482 936980 660488 936992
rect 660540 936980 660546 937032
rect 669958 935892 669964 935944
rect 670016 935932 670022 935944
rect 675478 935932 675484 935944
rect 670016 935904 675484 935932
rect 670016 935892 670022 935904
rect 675478 935892 675484 935904
rect 675536 935892 675542 935944
rect 672074 935756 672080 935808
rect 672132 935796 672138 935808
rect 675478 935796 675484 935808
rect 672132 935768 675484 935796
rect 672132 935756 672138 935768
rect 675478 935756 675484 935768
rect 675536 935756 675542 935808
rect 672442 935620 672448 935672
rect 672500 935660 672506 935672
rect 675294 935660 675300 935672
rect 672500 935632 675300 935660
rect 672500 935620 672506 935632
rect 675294 935620 675300 935632
rect 675352 935620 675358 935672
rect 672994 933308 673000 933360
rect 673052 933348 673058 933360
rect 675478 933348 675484 933360
rect 673052 933320 675484 933348
rect 673052 933308 673058 933320
rect 675478 933308 675484 933320
rect 675536 933308 675542 933360
rect 673362 932968 673368 933020
rect 673420 933008 673426 933020
rect 675478 933008 675484 933020
rect 673420 932980 675484 933008
rect 673420 932968 673426 932980
rect 675478 932968 675484 932980
rect 675536 932968 675542 933020
rect 43438 932900 43444 932952
rect 43496 932940 43502 932952
rect 54478 932940 54484 932952
rect 43496 932912 54484 932940
rect 43496 932900 43502 932912
rect 54478 932900 54484 932912
rect 54536 932900 54542 932952
rect 42794 931540 42800 931592
rect 42852 931580 42858 931592
rect 53098 931580 53104 931592
rect 42852 931552 53104 931580
rect 42852 931540 42858 931552
rect 53098 931540 53104 931552
rect 53156 931540 53162 931592
rect 673178 930112 673184 930164
rect 673236 930152 673242 930164
rect 675478 930152 675484 930164
rect 673236 930124 675484 930152
rect 673236 930112 673242 930124
rect 675478 930112 675484 930124
rect 675536 930112 675542 930164
rect 678238 930044 678244 930096
rect 678296 930084 678302 930096
rect 683114 930084 683120 930096
rect 678296 930056 683120 930084
rect 678296 930044 678302 930056
rect 683114 930044 683120 930056
rect 683172 930044 683178 930096
rect 669774 928752 669780 928804
rect 669832 928792 669838 928804
rect 675478 928792 675484 928804
rect 669832 928764 675484 928792
rect 669832 928752 669838 928764
rect 675478 928752 675484 928764
rect 675536 928752 675542 928804
rect 670602 927392 670608 927444
rect 670660 927432 670666 927444
rect 675478 927432 675484 927444
rect 670660 927404 675484 927432
rect 670660 927392 670666 927404
rect 675478 927392 675484 927404
rect 675536 927392 675542 927444
rect 47578 923244 47584 923296
rect 47636 923284 47642 923296
rect 62114 923284 62120 923296
rect 47636 923256 62120 923284
rect 47636 923244 47642 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651558 921816 651564 921868
rect 651616 921856 651622 921868
rect 661678 921856 661684 921868
rect 651616 921828 661684 921856
rect 651616 921816 651622 921828
rect 661678 921816 661684 921828
rect 661736 921816 661742 921868
rect 50338 909440 50344 909492
rect 50396 909480 50402 909492
rect 62114 909480 62120 909492
rect 50396 909452 62120 909480
rect 50396 909440 50402 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 651558 909440 651564 909492
rect 651616 909480 651622 909492
rect 664438 909480 664444 909492
rect 651616 909452 664444 909480
rect 651616 909440 651622 909452
rect 664438 909440 664444 909452
rect 664496 909440 664502 909492
rect 46198 896996 46204 897048
rect 46256 897036 46262 897048
rect 62114 897036 62120 897048
rect 46256 897008 62120 897036
rect 46256 896996 46262 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651558 895636 651564 895688
rect 651616 895676 651622 895688
rect 663058 895676 663064 895688
rect 651616 895648 663064 895676
rect 651616 895636 651622 895648
rect 663058 895636 663064 895648
rect 663116 895636 663122 895688
rect 42426 884688 42432 884740
rect 42484 884728 42490 884740
rect 62114 884728 62120 884740
rect 42484 884700 62120 884728
rect 42484 884688 42490 884700
rect 62114 884688 62120 884700
rect 62172 884688 62178 884740
rect 652386 881832 652392 881884
rect 652444 881872 652450 881884
rect 671338 881872 671344 881884
rect 652444 881844 671344 881872
rect 652444 881832 652450 881844
rect 671338 881832 671344 881844
rect 671396 881832 671402 881884
rect 669590 879044 669596 879096
rect 669648 879084 669654 879096
rect 675294 879084 675300 879096
rect 669648 879056 675300 879084
rect 669648 879044 669654 879056
rect 675294 879044 675300 879056
rect 675352 879044 675358 879096
rect 43438 870816 43444 870868
rect 43496 870856 43502 870868
rect 62114 870856 62120 870868
rect 43496 870828 62120 870856
rect 43496 870816 43502 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 651558 869388 651564 869440
rect 651616 869428 651622 869440
rect 658918 869428 658924 869440
rect 651616 869400 658924 869428
rect 651616 869388 651622 869400
rect 658918 869388 658924 869400
rect 658976 869388 658982 869440
rect 672994 869388 673000 869440
rect 673052 869428 673058 869440
rect 675110 869428 675116 869440
rect 673052 869400 675116 869428
rect 673052 869388 673058 869400
rect 675110 869388 675116 869400
rect 675168 869388 675174 869440
rect 671338 868980 671344 869032
rect 671396 869020 671402 869032
rect 675018 869020 675024 869032
rect 671396 868992 675024 869020
rect 671396 868980 671402 868992
rect 675018 868980 675024 868992
rect 675076 868980 675082 869032
rect 674650 868028 674656 868080
rect 674708 868068 674714 868080
rect 675110 868068 675116 868080
rect 674708 868040 675116 868068
rect 674708 868028 674714 868040
rect 675110 868028 675116 868040
rect 675168 868028 675174 868080
rect 670970 866804 670976 866856
rect 671028 866844 671034 866856
rect 675110 866844 675116 866856
rect 671028 866816 675116 866844
rect 671028 866804 671034 866816
rect 675110 866804 675116 866816
rect 675168 866804 675174 866856
rect 669222 866668 669228 866720
rect 669280 866708 669286 866720
rect 669280 866680 675064 866708
rect 669280 866668 669286 866680
rect 675036 866448 675064 866680
rect 675018 866396 675024 866448
rect 675076 866396 675082 866448
rect 674466 864628 674472 864680
rect 674524 864668 674530 864680
rect 675294 864668 675300 864680
rect 674524 864640 675300 864668
rect 674524 864628 674530 864640
rect 675294 864628 675300 864640
rect 675352 864628 675358 864680
rect 673362 862860 673368 862912
rect 673420 862900 673426 862912
rect 675110 862900 675116 862912
rect 673420 862872 675116 862900
rect 673420 862860 673426 862872
rect 675110 862860 675116 862872
rect 675168 862860 675174 862912
rect 51902 858372 51908 858424
rect 51960 858412 51966 858424
rect 62114 858412 62120 858424
rect 51960 858384 62120 858412
rect 51960 858372 51966 858384
rect 62114 858372 62120 858384
rect 62172 858372 62178 858424
rect 651558 855584 651564 855636
rect 651616 855624 651622 855636
rect 671338 855624 671344 855636
rect 651616 855596 671344 855624
rect 651616 855584 651622 855596
rect 671338 855584 671344 855596
rect 671396 855584 671402 855636
rect 44818 844568 44824 844620
rect 44876 844608 44882 844620
rect 62114 844608 62120 844620
rect 44876 844580 62120 844608
rect 44876 844568 44882 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 651558 841780 651564 841832
rect 651616 841820 651622 841832
rect 659102 841820 659108 841832
rect 651616 841792 659108 841820
rect 651616 841780 651622 841792
rect 659102 841780 659108 841792
rect 659160 841780 659166 841832
rect 55858 832124 55864 832176
rect 55916 832164 55922 832176
rect 62114 832164 62120 832176
rect 55916 832136 62120 832164
rect 55916 832124 55922 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651558 829404 651564 829456
rect 651616 829444 651622 829456
rect 660298 829444 660304 829456
rect 651616 829416 660304 829444
rect 651616 829404 651622 829416
rect 660298 829404 660304 829416
rect 660356 829404 660362 829456
rect 51718 818320 51724 818372
rect 51776 818360 51782 818372
rect 62114 818360 62120 818372
rect 51776 818332 62120 818360
rect 51776 818320 51782 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 35802 817096 35808 817148
rect 35860 817136 35866 817148
rect 40678 817136 40684 817148
rect 35860 817108 40684 817136
rect 35860 817096 35866 817108
rect 40678 817096 40684 817108
rect 40736 817096 40742 817148
rect 35618 816960 35624 817012
rect 35676 817000 35682 817012
rect 39942 817000 39948 817012
rect 35676 816972 39948 817000
rect 35676 816960 35682 816972
rect 39942 816960 39948 816972
rect 40000 816960 40006 817012
rect 35618 816008 35624 816060
rect 35676 816048 35682 816060
rect 41690 816048 41696 816060
rect 35676 816020 41696 816048
rect 35676 816008 35682 816020
rect 41690 816008 41696 816020
rect 41748 816008 41754 816060
rect 35434 815872 35440 815924
rect 35492 815912 35498 815924
rect 41690 815912 41696 815924
rect 35492 815884 41696 815912
rect 35492 815872 35498 815884
rect 41690 815872 41696 815884
rect 41748 815872 41754 815924
rect 35802 815736 35808 815788
rect 35860 815776 35866 815788
rect 41322 815776 41328 815788
rect 35860 815748 41328 815776
rect 35860 815736 35866 815748
rect 41322 815736 41328 815748
rect 41380 815736 41386 815788
rect 35250 815600 35256 815652
rect 35308 815640 35314 815652
rect 41690 815640 41696 815652
rect 35308 815612 41696 815640
rect 35308 815600 35314 815612
rect 41690 815600 41696 815612
rect 41748 815600 41754 815652
rect 42150 815600 42156 815652
rect 42208 815640 42214 815652
rect 50338 815640 50344 815652
rect 42208 815612 50344 815640
rect 42208 815600 42214 815612
rect 50338 815600 50344 815612
rect 50396 815600 50402 815652
rect 651558 815600 651564 815652
rect 651616 815640 651622 815652
rect 661862 815640 661868 815652
rect 651616 815612 661868 815640
rect 651616 815600 651622 815612
rect 661862 815600 661868 815612
rect 661920 815600 661926 815652
rect 41690 814756 41696 814768
rect 38626 814728 41696 814756
rect 35802 814648 35808 814700
rect 35860 814688 35866 814700
rect 38626 814688 38654 814728
rect 41690 814716 41696 814728
rect 41748 814716 41754 814768
rect 35860 814660 38654 814688
rect 35860 814648 35866 814660
rect 35618 814376 35624 814428
rect 35676 814416 35682 814428
rect 40310 814416 40316 814428
rect 35676 814388 40316 814416
rect 35676 814376 35682 814388
rect 40310 814376 40316 814388
rect 40368 814376 40374 814428
rect 35434 814240 35440 814292
rect 35492 814280 35498 814292
rect 41690 814280 41696 814292
rect 35492 814252 41696 814280
rect 35492 814240 35498 814252
rect 41690 814240 41696 814252
rect 41748 814240 41754 814292
rect 42058 814240 42064 814292
rect 42116 814280 42122 814292
rect 44174 814280 44180 814292
rect 42116 814252 44180 814280
rect 42116 814240 42122 814252
rect 44174 814240 44180 814252
rect 44232 814240 44238 814292
rect 41138 812948 41144 813000
rect 41196 812988 41202 813000
rect 41506 812988 41512 813000
rect 41196 812960 41512 812988
rect 41196 812948 41202 812960
rect 41506 812948 41512 812960
rect 41564 812948 41570 813000
rect 41322 811588 41328 811640
rect 41380 811628 41386 811640
rect 41690 811628 41696 811640
rect 41380 811600 41696 811628
rect 41380 811588 41386 811600
rect 41690 811588 41696 811600
rect 41748 811588 41754 811640
rect 43622 807440 43628 807492
rect 43680 807480 43686 807492
rect 48958 807480 48964 807492
rect 43680 807452 48964 807480
rect 43680 807440 43686 807452
rect 48958 807440 48964 807452
rect 49016 807440 49022 807492
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 651558 803224 651564 803276
rect 651616 803264 651622 803276
rect 663242 803264 663248 803276
rect 651616 803236 663248 803264
rect 651616 803224 651622 803236
rect 663242 803224 663248 803236
rect 663300 803224 663306 803276
rect 32398 802544 32404 802596
rect 32456 802584 32462 802596
rect 41690 802584 41696 802596
rect 32456 802556 41696 802584
rect 32456 802544 32462 802556
rect 41690 802544 41696 802556
rect 41748 802544 41754 802596
rect 31662 802272 31668 802324
rect 31720 802312 31726 802324
rect 39758 802312 39764 802324
rect 31720 802284 39764 802312
rect 31720 802272 31726 802284
rect 39758 802272 39764 802284
rect 39816 802272 39822 802324
rect 36538 801728 36544 801780
rect 36596 801768 36602 801780
rect 39850 801768 39856 801780
rect 36596 801740 39856 801768
rect 36596 801728 36602 801740
rect 39850 801728 39856 801740
rect 39908 801728 39914 801780
rect 33778 800912 33784 800964
rect 33836 800952 33842 800964
rect 40034 800952 40040 800964
rect 33836 800924 40040 800952
rect 33836 800912 33842 800924
rect 40034 800912 40040 800924
rect 40092 800912 40098 800964
rect 43622 799008 43628 799060
rect 43680 799048 43686 799060
rect 47578 799048 47584 799060
rect 43680 799020 47584 799048
rect 43680 799008 43686 799020
rect 47578 799008 47584 799020
rect 47636 799008 47642 799060
rect 47762 793568 47768 793620
rect 47820 793608 47826 793620
rect 62114 793608 62120 793620
rect 47820 793580 62120 793608
rect 47820 793568 47826 793580
rect 62114 793568 62120 793580
rect 62172 793568 62178 793620
rect 42242 792548 42248 792600
rect 42300 792588 42306 792600
rect 43070 792588 43076 792600
rect 42300 792560 43076 792588
rect 42300 792548 42306 792560
rect 43070 792548 43076 792560
rect 43128 792548 43134 792600
rect 42702 790236 42708 790288
rect 42760 790236 42766 790288
rect 42150 789964 42156 790016
rect 42208 790004 42214 790016
rect 42720 790004 42748 790236
rect 42208 789976 42748 790004
rect 42208 789964 42214 789976
rect 651558 789352 651564 789404
rect 651616 789392 651622 789404
rect 662046 789392 662052 789404
rect 651616 789364 662052 789392
rect 651616 789352 651622 789364
rect 662046 789352 662052 789364
rect 662104 789352 662110 789404
rect 670234 789352 670240 789404
rect 670292 789392 670298 789404
rect 675110 789392 675116 789404
rect 670292 789364 675116 789392
rect 670292 789352 670298 789364
rect 675110 789352 675116 789364
rect 675168 789352 675174 789404
rect 670786 787992 670792 788044
rect 670844 788032 670850 788044
rect 675110 788032 675116 788044
rect 670844 788004 675116 788032
rect 670844 787992 670850 788004
rect 675110 787992 675116 788004
rect 675168 787992 675174 788044
rect 674282 784116 674288 784168
rect 674340 784156 674346 784168
rect 675110 784156 675116 784168
rect 674340 784128 675116 784156
rect 674340 784116 674346 784128
rect 675110 784116 675116 784128
rect 675168 784116 675174 784168
rect 672258 782620 672264 782672
rect 672316 782660 672322 782672
rect 675110 782660 675116 782672
rect 672316 782632 675116 782660
rect 672316 782620 672322 782632
rect 675110 782620 675116 782632
rect 675168 782620 675174 782672
rect 668762 782484 668768 782536
rect 668820 782524 668826 782536
rect 675294 782524 675300 782536
rect 668820 782496 675300 782524
rect 668820 782484 668826 782496
rect 675294 782484 675300 782496
rect 675352 782484 675358 782536
rect 56226 780036 56232 780088
rect 56284 780076 56290 780088
rect 62114 780076 62120 780088
rect 56284 780048 62120 780076
rect 56284 780036 56290 780048
rect 62114 780036 62120 780048
rect 62172 780036 62178 780088
rect 673638 779764 673644 779816
rect 673696 779804 673702 779816
rect 675110 779804 675116 779816
rect 673696 779776 675116 779804
rect 673696 779764 673702 779776
rect 675110 779764 675116 779776
rect 675168 779764 675174 779816
rect 673822 779084 673828 779136
rect 673880 779124 673886 779136
rect 675110 779124 675116 779136
rect 673880 779096 675116 779124
rect 673880 779084 673886 779096
rect 675110 779084 675116 779096
rect 675168 779084 675174 779136
rect 660298 778948 660304 779000
rect 660356 778988 660362 779000
rect 675110 778988 675116 779000
rect 660356 778960 675116 778988
rect 660356 778948 660362 778960
rect 675110 778948 675116 778960
rect 675168 778948 675174 779000
rect 672810 778336 672816 778388
rect 672868 778376 672874 778388
rect 675294 778376 675300 778388
rect 672868 778348 675300 778376
rect 672868 778336 672874 778348
rect 675294 778336 675300 778348
rect 675352 778336 675358 778388
rect 674190 776976 674196 777028
rect 674248 777016 674254 777028
rect 675294 777016 675300 777028
rect 674248 776988 675300 777016
rect 674248 776976 674254 776988
rect 675294 776976 675300 776988
rect 675352 776976 675358 777028
rect 674834 775888 674840 775940
rect 674892 775928 674898 775940
rect 675202 775928 675208 775940
rect 674892 775900 675208 775928
rect 674892 775888 674898 775900
rect 675202 775888 675208 775900
rect 675260 775888 675266 775940
rect 675018 775752 675024 775804
rect 675076 775752 675082 775804
rect 651558 775548 651564 775600
rect 651616 775588 651622 775600
rect 660482 775588 660488 775600
rect 651616 775560 660488 775588
rect 651616 775548 651622 775560
rect 660482 775548 660488 775560
rect 660540 775548 660546 775600
rect 674834 775548 674840 775600
rect 674892 775588 674898 775600
rect 675036 775588 675064 775752
rect 674892 775560 675064 775588
rect 674892 775548 674898 775560
rect 35802 774324 35808 774376
rect 35860 774364 35866 774376
rect 39758 774364 39764 774376
rect 35860 774336 39764 774364
rect 35860 774324 35866 774336
rect 39758 774324 39764 774336
rect 39816 774324 39822 774376
rect 35526 773372 35532 773424
rect 35584 773412 35590 773424
rect 40862 773412 40868 773424
rect 35584 773384 40868 773412
rect 35584 773372 35590 773384
rect 40862 773372 40868 773384
rect 40920 773372 40926 773424
rect 35802 773276 35808 773288
rect 35636 773248 35808 773276
rect 35636 773004 35664 773248
rect 35802 773236 35808 773248
rect 35860 773236 35866 773288
rect 35802 773100 35808 773152
rect 35860 773140 35866 773152
rect 41690 773140 41696 773152
rect 35860 773112 41696 773140
rect 35860 773100 35866 773112
rect 41690 773100 41696 773112
rect 41748 773100 41754 773152
rect 42058 773100 42064 773152
rect 42116 773140 42122 773152
rect 44450 773140 44456 773152
rect 42116 773112 44456 773140
rect 42116 773100 42122 773112
rect 44450 773100 44456 773112
rect 44508 773100 44514 773152
rect 41690 773004 41696 773016
rect 35636 772976 41696 773004
rect 41690 772964 41696 772976
rect 41748 772964 41754 773016
rect 42058 772964 42064 773016
rect 42116 773004 42122 773016
rect 55858 773004 55864 773016
rect 42116 772976 55864 773004
rect 42116 772964 42122 772976
rect 55858 772964 55864 772976
rect 55916 772964 55922 773016
rect 35342 772828 35348 772880
rect 35400 772868 35406 772880
rect 51902 772868 51908 772880
rect 35400 772840 41736 772868
rect 35400 772828 35406 772840
rect 41708 772744 41736 772840
rect 42076 772840 51908 772868
rect 42076 772744 42104 772840
rect 51902 772828 51908 772840
rect 51960 772828 51966 772880
rect 41690 772692 41696 772744
rect 41748 772692 41754 772744
rect 42058 772692 42064 772744
rect 42116 772692 42122 772744
rect 676030 772216 676036 772268
rect 676088 772256 676094 772268
rect 683298 772256 683304 772268
rect 676088 772228 683304 772256
rect 676088 772216 676094 772228
rect 683298 772216 683304 772228
rect 683356 772216 683362 772268
rect 675846 772080 675852 772132
rect 675904 772120 675910 772132
rect 684126 772120 684132 772132
rect 675904 772092 684132 772120
rect 675904 772080 675910 772092
rect 684126 772080 684132 772092
rect 684184 772080 684190 772132
rect 35526 771672 35532 771724
rect 35584 771712 35590 771724
rect 39850 771712 39856 771724
rect 35584 771684 39856 771712
rect 35584 771672 35590 771684
rect 39850 771672 39856 771684
rect 39908 771672 39914 771724
rect 35802 771536 35808 771588
rect 35860 771576 35866 771588
rect 41690 771576 41696 771588
rect 35860 771548 41696 771576
rect 35860 771536 35866 771548
rect 41690 771536 41696 771548
rect 41748 771536 41754 771588
rect 42058 771536 42064 771588
rect 42116 771576 42122 771588
rect 42886 771576 42892 771588
rect 42116 771548 42892 771576
rect 42116 771536 42122 771548
rect 42886 771536 42892 771548
rect 42944 771536 42950 771588
rect 35342 771400 35348 771452
rect 35400 771440 35406 771452
rect 41690 771440 41696 771452
rect 35400 771412 41696 771440
rect 35400 771400 35406 771412
rect 41690 771400 41696 771412
rect 41748 771400 41754 771452
rect 42058 771400 42064 771452
rect 42116 771440 42122 771452
rect 44174 771440 44180 771452
rect 42116 771412 44180 771440
rect 42116 771400 42122 771412
rect 44174 771400 44180 771412
rect 44232 771400 44238 771452
rect 35802 770448 35808 770500
rect 35860 770488 35866 770500
rect 39850 770488 39856 770500
rect 35860 770460 39856 770488
rect 35860 770448 35866 770460
rect 39850 770448 39856 770460
rect 39908 770448 39914 770500
rect 41690 770284 41696 770296
rect 41386 770256 41696 770284
rect 35618 770176 35624 770228
rect 35676 770216 35682 770228
rect 41386 770216 41414 770256
rect 41690 770244 41696 770256
rect 41748 770244 41754 770296
rect 42058 770244 42064 770296
rect 42116 770284 42122 770296
rect 43254 770284 43260 770296
rect 42116 770256 43260 770284
rect 42116 770244 42122 770256
rect 43254 770244 43260 770256
rect 43312 770244 43318 770296
rect 35676 770188 41414 770216
rect 35676 770176 35682 770188
rect 35802 770040 35808 770092
rect 35860 770080 35866 770092
rect 41690 770080 41696 770092
rect 35860 770052 41696 770080
rect 35860 770040 35866 770052
rect 41690 770040 41696 770052
rect 41748 770040 41754 770092
rect 42058 770040 42064 770092
rect 42116 770080 42122 770092
rect 44634 770080 44640 770092
rect 42116 770052 44640 770080
rect 42116 770040 42122 770052
rect 44634 770040 44640 770052
rect 44692 770040 44698 770092
rect 35802 768816 35808 768868
rect 35860 768856 35866 768868
rect 39298 768856 39304 768868
rect 35860 768828 39304 768856
rect 35860 768816 35866 768828
rect 39298 768816 39304 768828
rect 39356 768816 39362 768868
rect 35618 768680 35624 768732
rect 35676 768720 35682 768732
rect 41322 768720 41328 768732
rect 35676 768692 41328 768720
rect 35676 768680 35682 768692
rect 41322 768680 41328 768692
rect 41380 768680 41386 768732
rect 35802 767592 35808 767644
rect 35860 767632 35866 767644
rect 40034 767632 40040 767644
rect 35860 767604 40040 767632
rect 35860 767592 35866 767604
rect 40034 767592 40040 767604
rect 40092 767592 40098 767644
rect 35618 767456 35624 767508
rect 35676 767496 35682 767508
rect 36538 767496 36544 767508
rect 35676 767468 36544 767496
rect 35676 767456 35682 767468
rect 36538 767456 36544 767468
rect 36596 767456 36602 767508
rect 43622 767320 43628 767372
rect 43680 767360 43686 767372
rect 62114 767360 62120 767372
rect 43680 767332 62120 767360
rect 43680 767320 43686 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 674926 766368 674932 766420
rect 674984 766408 674990 766420
rect 675386 766408 675392 766420
rect 674984 766380 675392 766408
rect 674984 766368 674990 766380
rect 675386 766368 675392 766380
rect 675444 766368 675450 766420
rect 35802 766300 35808 766352
rect 35860 766340 35866 766352
rect 35860 766300 35894 766340
rect 35866 766204 35894 766300
rect 39758 766204 39764 766216
rect 35866 766176 39764 766204
rect 39758 766164 39764 766176
rect 39816 766164 39822 766216
rect 41690 766000 41696 766012
rect 41386 765972 41696 766000
rect 35802 765892 35808 765944
rect 35860 765932 35866 765944
rect 41386 765932 41414 765972
rect 41690 765960 41696 765972
rect 41748 765960 41754 766012
rect 35860 765904 41414 765932
rect 35860 765892 35866 765904
rect 42058 765892 42064 765944
rect 42116 765932 42122 765944
rect 44450 765932 44456 765944
rect 42116 765904 44456 765932
rect 42116 765892 42122 765904
rect 44450 765892 44456 765904
rect 44508 765892 44514 765944
rect 40034 765144 40040 765196
rect 40092 765184 40098 765196
rect 41690 765184 41696 765196
rect 40092 765156 41696 765184
rect 40092 765144 40098 765156
rect 41690 765144 41696 765156
rect 41748 765144 41754 765196
rect 42058 765008 42064 765060
rect 42116 765048 42122 765060
rect 42518 765048 42524 765060
rect 42116 765020 42524 765048
rect 42116 765008 42122 765020
rect 42518 765008 42524 765020
rect 42576 765008 42582 765060
rect 35802 764668 35808 764720
rect 35860 764708 35866 764720
rect 39114 764708 39120 764720
rect 35860 764680 39120 764708
rect 35860 764668 35866 764680
rect 39114 764668 39120 764680
rect 39172 764668 39178 764720
rect 35802 763308 35808 763360
rect 35860 763348 35866 763360
rect 37918 763348 37924 763360
rect 35860 763320 37924 763348
rect 35860 763308 35866 763320
rect 37918 763308 37924 763320
rect 37976 763308 37982 763360
rect 41690 763280 41696 763292
rect 38626 763252 41696 763280
rect 35618 763172 35624 763224
rect 35676 763212 35682 763224
rect 38626 763212 38654 763252
rect 41690 763240 41696 763252
rect 41748 763240 41754 763292
rect 651558 763240 651564 763292
rect 651616 763280 651622 763292
rect 651616 763252 654134 763280
rect 651616 763240 651622 763252
rect 35676 763184 38654 763212
rect 654106 763212 654134 763252
rect 660298 763212 660304 763224
rect 654106 763184 660304 763212
rect 35676 763172 35682 763184
rect 660298 763172 660304 763184
rect 660356 763172 660362 763224
rect 35802 761880 35808 761932
rect 35860 761920 35866 761932
rect 40218 761920 40224 761932
rect 35860 761892 40224 761920
rect 35860 761880 35866 761892
rect 40218 761880 40224 761892
rect 40276 761880 40282 761932
rect 664438 760860 664444 760912
rect 664496 760900 664502 760912
rect 675478 760900 675484 760912
rect 664496 760872 675484 760900
rect 664496 760860 664502 760872
rect 675478 760860 675484 760872
rect 675536 760860 675542 760912
rect 661678 760520 661684 760572
rect 661736 760560 661742 760572
rect 675294 760560 675300 760572
rect 661736 760532 675300 760560
rect 661736 760520 661742 760532
rect 675294 760520 675300 760532
rect 675352 760520 675358 760572
rect 663058 760384 663064 760436
rect 663116 760424 663122 760436
rect 675478 760424 675484 760436
rect 663116 760396 675484 760424
rect 663116 760384 663122 760396
rect 675478 760384 675484 760396
rect 675536 760384 675542 760436
rect 671522 760248 671528 760300
rect 671580 760288 671586 760300
rect 675294 760288 675300 760300
rect 671580 760260 675300 760288
rect 671580 760248 671586 760260
rect 675294 760248 675300 760260
rect 675352 760248 675358 760300
rect 671522 759840 671528 759892
rect 671580 759880 671586 759892
rect 675478 759880 675484 759892
rect 671580 759852 675484 759880
rect 671580 759840 671586 759852
rect 675478 759840 675484 759852
rect 675536 759840 675542 759892
rect 671154 759500 671160 759552
rect 671212 759540 671218 759552
rect 675478 759540 675484 759552
rect 671212 759512 675484 759540
rect 671212 759500 671218 759512
rect 675478 759500 675484 759512
rect 675536 759500 675542 759552
rect 36538 759024 36544 759076
rect 36596 759064 36602 759076
rect 39942 759064 39948 759076
rect 36596 759036 39948 759064
rect 36596 759024 36602 759036
rect 39942 759024 39948 759036
rect 40000 759024 40006 759076
rect 671154 759024 671160 759076
rect 671212 759064 671218 759076
rect 675478 759064 675484 759076
rect 671212 759036 675484 759064
rect 671212 759024 671218 759036
rect 675478 759024 675484 759036
rect 675536 759024 675542 759076
rect 672074 758684 672080 758736
rect 672132 758724 672138 758736
rect 675478 758724 675484 758736
rect 672132 758696 675484 758724
rect 672132 758684 672138 758696
rect 675478 758684 675484 758696
rect 675536 758684 675542 758736
rect 673178 758208 673184 758260
rect 673236 758248 673242 758260
rect 675478 758248 675484 758260
rect 673236 758220 675484 758248
rect 673236 758208 673242 758220
rect 675478 758208 675484 758220
rect 675536 758208 675542 758260
rect 35158 758140 35164 758192
rect 35216 758180 35222 758192
rect 41690 758180 41696 758192
rect 35216 758152 41696 758180
rect 35216 758140 35222 758152
rect 41690 758140 41696 758152
rect 41748 758140 41754 758192
rect 42426 758140 42432 758192
rect 42484 758140 42490 758192
rect 37918 757732 37924 757784
rect 37976 757772 37982 757784
rect 41598 757772 41604 757784
rect 37976 757744 41604 757772
rect 37976 757732 37982 757744
rect 41598 757732 41604 757744
rect 41656 757732 41662 757784
rect 42444 757648 42472 758140
rect 672442 757868 672448 757920
rect 672500 757908 672506 757920
rect 675478 757908 675484 757920
rect 672500 757880 675484 757908
rect 672500 757868 672506 757880
rect 675478 757868 675484 757880
rect 675536 757868 675542 757920
rect 42426 757596 42432 757648
rect 42484 757596 42490 757648
rect 672074 757392 672080 757444
rect 672132 757432 672138 757444
rect 675478 757432 675484 757444
rect 672132 757404 675484 757432
rect 672132 757392 672138 757404
rect 675478 757392 675484 757404
rect 675536 757392 675542 757444
rect 674006 756236 674012 756288
rect 674064 756276 674070 756288
rect 675110 756276 675116 756288
rect 674064 756248 675116 756276
rect 674064 756236 674070 756248
rect 675110 756236 675116 756248
rect 675168 756236 675174 756288
rect 673362 755012 673368 755064
rect 673420 755052 673426 755064
rect 675478 755052 675484 755064
rect 673420 755024 675484 755052
rect 673420 755012 673426 755024
rect 675478 755012 675484 755024
rect 675536 755012 675542 755064
rect 44450 754916 44456 754928
rect 42260 754888 44456 754916
rect 42260 754316 42288 754888
rect 44450 754876 44456 754888
rect 44508 754876 44514 754928
rect 669590 754604 669596 754656
rect 669648 754644 669654 754656
rect 675478 754644 675484 754656
rect 669648 754616 675484 754644
rect 669648 754604 669654 754616
rect 675478 754604 675484 754616
rect 675536 754604 675542 754656
rect 42242 754264 42248 754316
rect 42300 754264 42306 754316
rect 672626 754196 672632 754248
rect 672684 754236 672690 754248
rect 675478 754236 675484 754248
rect 672684 754208 675484 754236
rect 672684 754196 672690 754208
rect 675478 754196 675484 754208
rect 675536 754196 675542 754248
rect 43438 753516 43444 753568
rect 43496 753556 43502 753568
rect 45002 753556 45008 753568
rect 43496 753528 45008 753556
rect 43496 753516 43502 753528
rect 45002 753516 45008 753528
rect 45060 753516 45066 753568
rect 50706 753516 50712 753568
rect 50764 753556 50770 753568
rect 62114 753556 62120 753568
rect 50764 753528 62120 753556
rect 50764 753516 50770 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 670970 753380 670976 753432
rect 671028 753420 671034 753432
rect 675478 753420 675484 753432
rect 671028 753392 675484 753420
rect 671028 753380 671034 753392
rect 675478 753380 675484 753392
rect 675536 753380 675542 753432
rect 672994 752156 673000 752208
rect 673052 752196 673058 752208
rect 675478 752196 675484 752208
rect 673052 752168 675484 752196
rect 673052 752156 673058 752168
rect 675478 752156 675484 752168
rect 675536 752156 675542 752208
rect 671798 751748 671804 751800
rect 671856 751788 671862 751800
rect 675478 751788 675484 751800
rect 671856 751760 675484 751788
rect 671856 751748 671862 751760
rect 675478 751748 675484 751760
rect 675536 751748 675542 751800
rect 675846 750932 675852 750984
rect 675904 750972 675910 750984
rect 683114 750972 683120 750984
rect 675904 750944 683120 750972
rect 675904 750932 675910 750944
rect 683114 750932 683120 750944
rect 683172 750932 683178 750984
rect 669590 750048 669596 750100
rect 669648 750088 669654 750100
rect 675478 750088 675484 750100
rect 669648 750060 675484 750088
rect 669648 750048 669654 750060
rect 675478 750048 675484 750060
rect 675536 750048 675542 750100
rect 651558 749368 651564 749420
rect 651616 749408 651622 749420
rect 664438 749408 664444 749420
rect 651616 749380 664444 749408
rect 651616 749368 651622 749380
rect 664438 749368 664444 749380
rect 664496 749368 664502 749420
rect 42426 749300 42432 749352
rect 42484 749340 42490 749352
rect 43254 749340 43260 749352
rect 42484 749312 43260 749340
rect 42484 749300 42490 749312
rect 43254 749300 43260 749312
rect 43312 749300 43318 749352
rect 669222 743656 669228 743708
rect 669280 743696 669286 743708
rect 675110 743696 675116 743708
rect 669280 743668 675116 743696
rect 669280 743656 669286 743668
rect 675110 743656 675116 743668
rect 675168 743656 675174 743708
rect 671890 742772 671896 742824
rect 671948 742812 671954 742824
rect 675294 742812 675300 742824
rect 671948 742784 675300 742812
rect 671948 742772 671954 742784
rect 675294 742772 675300 742784
rect 675352 742772 675358 742824
rect 666370 742432 666376 742484
rect 666428 742472 666434 742484
rect 675294 742472 675300 742484
rect 666428 742444 675300 742472
rect 666428 742432 666434 742444
rect 675294 742432 675300 742444
rect 675352 742432 675358 742484
rect 674834 741616 674840 741668
rect 674892 741656 674898 741668
rect 675478 741656 675484 741668
rect 674892 741628 675484 741656
rect 674892 741616 674898 741628
rect 675478 741616 675484 741628
rect 675536 741616 675542 741668
rect 56042 741072 56048 741124
rect 56100 741112 56106 741124
rect 62114 741112 62120 741124
rect 56100 741084 62120 741112
rect 56100 741072 56106 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 674466 739712 674472 739764
rect 674524 739752 674530 739764
rect 675110 739752 675116 739764
rect 674524 739724 675116 739752
rect 674524 739712 674530 739724
rect 675110 739712 675116 739724
rect 675168 739712 675174 739764
rect 674006 738624 674012 738676
rect 674064 738664 674070 738676
rect 675386 738664 675392 738676
rect 674064 738636 675392 738664
rect 674064 738624 674070 738636
rect 675386 738624 675392 738636
rect 675444 738624 675450 738676
rect 651558 735564 651564 735616
rect 651616 735604 651622 735616
rect 663058 735604 663064 735616
rect 651616 735576 663064 735604
rect 651616 735564 651622 735576
rect 663058 735564 663064 735576
rect 663116 735564 663122 735616
rect 670786 734952 670792 735004
rect 670844 734992 670850 735004
rect 675294 734992 675300 735004
rect 670844 734964 675300 734992
rect 670844 734952 670850 734964
rect 675294 734952 675300 734964
rect 675352 734952 675358 735004
rect 660482 734816 660488 734868
rect 660540 734856 660546 734868
rect 675294 734856 675300 734868
rect 660540 734828 675300 734856
rect 660540 734816 660546 734828
rect 675294 734816 675300 734828
rect 675352 734816 675358 734868
rect 667658 732776 667664 732828
rect 667716 732816 667722 732828
rect 675110 732816 675116 732828
rect 667716 732788 675116 732816
rect 667716 732776 667722 732788
rect 675110 732776 675116 732788
rect 675168 732776 675174 732828
rect 43438 731144 43444 731196
rect 43496 731184 43502 731196
rect 50338 731184 50344 731196
rect 43496 731156 50344 731184
rect 43496 731144 43502 731156
rect 50338 731144 50344 731156
rect 50396 731144 50402 731196
rect 43254 730124 43260 730176
rect 43312 730164 43318 730176
rect 43312 730136 51074 730164
rect 43312 730124 43318 730136
rect 51046 730096 51074 730136
rect 56226 730096 56232 730108
rect 51046 730068 56232 730096
rect 56226 730056 56232 730068
rect 56284 730056 56290 730108
rect 41322 728628 41328 728680
rect 41380 728668 41386 728680
rect 41690 728668 41696 728680
rect 41380 728640 41696 728668
rect 41380 728628 41386 728640
rect 41690 728628 41696 728640
rect 41748 728628 41754 728680
rect 42058 728628 42064 728680
rect 42116 728668 42122 728680
rect 45002 728668 45008 728680
rect 42116 728640 45008 728668
rect 42116 728628 42122 728640
rect 45002 728628 45008 728640
rect 45060 728628 45066 728680
rect 670418 728628 670424 728680
rect 670476 728668 670482 728680
rect 675110 728668 675116 728680
rect 670476 728640 675116 728668
rect 670476 728628 670482 728640
rect 675110 728628 675116 728640
rect 675168 728628 675174 728680
rect 41046 727404 41052 727456
rect 41104 727444 41110 727456
rect 41690 727444 41696 727456
rect 41104 727416 41696 727444
rect 41104 727404 41110 727416
rect 41690 727404 41696 727416
rect 41748 727404 41754 727456
rect 42058 727404 42064 727456
rect 42116 727444 42122 727456
rect 43070 727444 43076 727456
rect 42116 727416 43076 727444
rect 42116 727404 42122 727416
rect 43070 727404 43076 727416
rect 43128 727404 43134 727456
rect 40862 727268 40868 727320
rect 40920 727308 40926 727320
rect 41690 727308 41696 727320
rect 40920 727280 41696 727308
rect 40920 727268 40926 727280
rect 41690 727268 41696 727280
rect 41748 727268 41754 727320
rect 42058 727268 42064 727320
rect 42116 727308 42122 727320
rect 44266 727308 44272 727320
rect 42116 727280 44272 727308
rect 42116 727268 42122 727280
rect 44266 727268 44272 727280
rect 44324 727268 44330 727320
rect 51902 727268 51908 727320
rect 51960 727308 51966 727320
rect 62114 727308 62120 727320
rect 51960 727280 62120 727308
rect 51960 727268 51966 727280
rect 62114 727268 62120 727280
rect 62172 727268 62178 727320
rect 675846 726792 675852 726844
rect 675904 726832 675910 726844
rect 684218 726832 684224 726844
rect 675904 726804 684224 726832
rect 675904 726792 675910 726804
rect 684218 726792 684224 726804
rect 684276 726792 684282 726844
rect 676030 726520 676036 726572
rect 676088 726560 676094 726572
rect 683206 726560 683212 726572
rect 676088 726532 683212 726560
rect 676088 726520 676094 726532
rect 683206 726520 683212 726532
rect 683264 726520 683270 726572
rect 41322 726316 41328 726368
rect 41380 726356 41386 726368
rect 41598 726356 41604 726368
rect 41380 726328 41604 726356
rect 41380 726316 41386 726328
rect 41598 726316 41604 726328
rect 41656 726316 41662 726368
rect 651558 723120 651564 723172
rect 651616 723160 651622 723172
rect 659286 723160 659292 723172
rect 651616 723132 659292 723160
rect 651616 723120 651622 723132
rect 659286 723120 659292 723132
rect 659344 723120 659350 723172
rect 31754 720264 31760 720316
rect 31812 720304 31818 720316
rect 40034 720304 40040 720316
rect 31812 720276 40040 720304
rect 31812 720264 31818 720276
rect 40034 720264 40040 720276
rect 40092 720264 40098 720316
rect 42334 719108 42340 719160
rect 42392 719148 42398 719160
rect 55858 719148 55864 719160
rect 42392 719120 55864 719148
rect 42392 719108 42398 719120
rect 55858 719108 55864 719120
rect 55916 719108 55922 719160
rect 671338 716524 671344 716576
rect 671396 716564 671402 716576
rect 675478 716564 675484 716576
rect 671396 716536 675484 716564
rect 671396 716524 671402 716536
rect 675478 716524 675484 716536
rect 675536 716524 675542 716576
rect 37918 716048 37924 716100
rect 37976 716088 37982 716100
rect 40310 716088 40316 716100
rect 37976 716060 40316 716088
rect 37976 716048 37982 716060
rect 40310 716048 40316 716060
rect 40368 716048 40374 716100
rect 35158 715640 35164 715692
rect 35216 715680 35222 715692
rect 41322 715680 41328 715692
rect 35216 715652 41328 715680
rect 35216 715640 35222 715652
rect 41322 715640 41328 715652
rect 41380 715640 41386 715692
rect 33778 715368 33784 715420
rect 33836 715408 33842 715420
rect 41690 715408 41696 715420
rect 33836 715380 41696 715408
rect 33836 715368 33842 715380
rect 41690 715368 41696 715380
rect 41748 715368 41754 715420
rect 671522 715300 671528 715352
rect 671580 715340 671586 715352
rect 675110 715340 675116 715352
rect 671580 715312 675116 715340
rect 671580 715300 671586 715312
rect 675110 715300 675116 715312
rect 675168 715300 675174 715352
rect 42058 715232 42064 715284
rect 42116 715272 42122 715284
rect 42702 715272 42708 715284
rect 42116 715244 42708 715272
rect 42116 715232 42122 715244
rect 42702 715232 42708 715244
rect 42760 715232 42766 715284
rect 659102 715096 659108 715148
rect 659160 715136 659166 715148
rect 675478 715136 675484 715148
rect 659160 715108 675484 715136
rect 659160 715096 659166 715108
rect 675478 715096 675484 715108
rect 675536 715096 675542 715148
rect 658918 714960 658924 715012
rect 658976 715000 658982 715012
rect 675294 715000 675300 715012
rect 658976 714972 675300 715000
rect 658976 714960 658982 714972
rect 675294 714960 675300 714972
rect 675352 714960 675358 715012
rect 50522 714824 50528 714876
rect 50580 714864 50586 714876
rect 62114 714864 62120 714876
rect 50580 714836 62120 714864
rect 50580 714824 50586 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 671522 714824 671528 714876
rect 671580 714864 671586 714876
rect 675478 714864 675484 714876
rect 671580 714836 675484 714864
rect 671580 714824 671586 714836
rect 675478 714824 675484 714836
rect 675536 714824 675542 714876
rect 40034 714484 40040 714536
rect 40092 714524 40098 714536
rect 41690 714524 41696 714536
rect 40092 714496 41696 714524
rect 40092 714484 40098 714496
rect 41690 714484 41696 714496
rect 41748 714484 41754 714536
rect 671154 714484 671160 714536
rect 671212 714524 671218 714536
rect 675478 714524 675484 714536
rect 671212 714496 675484 714524
rect 671212 714484 671218 714496
rect 675478 714484 675484 714496
rect 675536 714484 675542 714536
rect 672994 714008 673000 714060
rect 673052 714048 673058 714060
rect 675478 714048 675484 714060
rect 673052 714020 675484 714048
rect 673052 714008 673058 714020
rect 675478 714008 675484 714020
rect 675536 714008 675542 714060
rect 673178 713668 673184 713720
rect 673236 713708 673242 713720
rect 675478 713708 675484 713720
rect 673236 713680 675484 713708
rect 673236 713668 673242 713680
rect 675478 713668 675484 713680
rect 675536 713668 675542 713720
rect 671154 713192 671160 713244
rect 671212 713232 671218 713244
rect 675478 713232 675484 713244
rect 671212 713204 675484 713232
rect 671212 713192 671218 713204
rect 675478 713192 675484 713204
rect 675536 713192 675542 713244
rect 672074 712852 672080 712904
rect 672132 712892 672138 712904
rect 675478 712892 675484 712904
rect 672132 712864 675484 712892
rect 672132 712852 672138 712864
rect 675478 712852 675484 712864
rect 675536 712852 675542 712904
rect 671338 712376 671344 712428
rect 671396 712416 671402 712428
rect 675478 712416 675484 712428
rect 671396 712388 675484 712416
rect 671396 712376 671402 712388
rect 675478 712376 675484 712388
rect 675536 712376 675542 712428
rect 42886 712240 42892 712292
rect 42944 712280 42950 712292
rect 51718 712280 51724 712292
rect 42944 712252 51724 712280
rect 42944 712240 42950 712252
rect 51718 712240 51724 712252
rect 51776 712240 51782 712292
rect 676214 712036 676220 712088
rect 676272 712076 676278 712088
rect 677502 712076 677508 712088
rect 676272 712048 677508 712076
rect 676272 712036 676278 712048
rect 677502 712036 677508 712048
rect 677560 712036 677566 712088
rect 676030 711832 676036 711884
rect 676088 711872 676094 711884
rect 676766 711872 676772 711884
rect 676088 711844 676772 711872
rect 676088 711832 676094 711844
rect 676766 711832 676772 711844
rect 676824 711832 676830 711884
rect 670970 711220 670976 711272
rect 671028 711260 671034 711272
rect 675478 711260 675484 711272
rect 671028 711232 675484 711260
rect 671028 711220 671034 711232
rect 675478 711220 675484 711232
rect 675536 711220 675542 711272
rect 42242 710948 42248 711000
rect 42300 710988 42306 711000
rect 42886 710988 42892 711000
rect 42300 710960 42892 710988
rect 42300 710948 42306 710960
rect 42886 710948 42892 710960
rect 42944 710948 42950 711000
rect 668578 709724 668584 709776
rect 668636 709764 668642 709776
rect 675478 709764 675484 709776
rect 668636 709736 675484 709764
rect 668636 709724 668642 709736
rect 675478 709724 675484 709736
rect 675536 709724 675542 709776
rect 670234 709588 670240 709640
rect 670292 709628 670298 709640
rect 675478 709628 675484 709640
rect 670292 709600 675484 709628
rect 670292 709588 670298 709600
rect 675478 709588 675484 709600
rect 675536 709588 675542 709640
rect 44174 709356 44180 709368
rect 42352 709328 44180 709356
rect 42352 708416 42380 709328
rect 44174 709316 44180 709328
rect 44232 709316 44238 709368
rect 651558 709316 651564 709368
rect 651616 709356 651622 709368
rect 658918 709356 658924 709368
rect 651616 709328 658924 709356
rect 651616 709316 651622 709328
rect 658918 709316 658924 709328
rect 658976 709316 658982 709368
rect 668762 709316 668768 709368
rect 668820 709356 668826 709368
rect 675294 709356 675300 709368
rect 668820 709328 675300 709356
rect 668820 709316 668826 709328
rect 675294 709316 675300 709328
rect 675352 709316 675358 709368
rect 42334 708364 42340 708416
rect 42392 708364 42398 708416
rect 673822 707956 673828 708008
rect 673880 707996 673886 708008
rect 675478 707996 675484 708008
rect 673880 707968 675484 707996
rect 673880 707956 673886 707968
rect 675478 707956 675484 707968
rect 675536 707956 675542 708008
rect 43070 707752 43076 707804
rect 43128 707792 43134 707804
rect 43438 707792 43444 707804
rect 43128 707764 43444 707792
rect 43128 707752 43134 707764
rect 43438 707752 43444 707764
rect 43496 707752 43502 707804
rect 672350 707548 672356 707600
rect 672408 707588 672414 707600
rect 675478 707588 675484 707600
rect 672408 707560 675484 707588
rect 672408 707548 672414 707560
rect 675478 707548 675484 707560
rect 675536 707548 675542 707600
rect 673638 707140 673644 707192
rect 673696 707180 673702 707192
rect 675478 707180 675484 707192
rect 673696 707152 675484 707180
rect 673696 707140 673702 707152
rect 675478 707140 675484 707152
rect 675536 707140 675542 707192
rect 672810 706732 672816 706784
rect 672868 706772 672874 706784
rect 675478 706772 675484 706784
rect 672868 706744 675484 706772
rect 672868 706732 672874 706744
rect 675478 706732 675484 706744
rect 675536 706732 675542 706784
rect 675846 705168 675852 705220
rect 675904 705208 675910 705220
rect 683114 705208 683120 705220
rect 675904 705180 683120 705208
rect 675904 705168 675910 705180
rect 683114 705168 683120 705180
rect 683172 705168 683178 705220
rect 669958 705032 669964 705084
rect 670016 705072 670022 705084
rect 675478 705072 675484 705084
rect 670016 705044 675484 705072
rect 670016 705032 670022 705044
rect 675478 705032 675484 705044
rect 675536 705032 675542 705084
rect 42242 702108 42248 702160
rect 42300 702108 42306 702160
rect 42260 701888 42288 702108
rect 42242 701836 42248 701888
rect 42300 701836 42306 701888
rect 51718 701020 51724 701072
rect 51776 701060 51782 701072
rect 62114 701060 62120 701072
rect 51776 701032 62120 701060
rect 51776 701020 51782 701032
rect 62114 701020 62120 701032
rect 62172 701020 62178 701072
rect 668762 699660 668768 699712
rect 668820 699700 668826 699712
rect 675110 699700 675116 699712
rect 668820 699672 675116 699700
rect 668820 699660 668826 699672
rect 675110 699660 675116 699672
rect 675168 699660 675174 699712
rect 651558 696940 651564 696992
rect 651616 696980 651622 696992
rect 664622 696980 664628 696992
rect 651616 696952 664628 696980
rect 651616 696940 651622 696952
rect 664622 696940 664628 696952
rect 664680 696940 664686 696992
rect 673638 694152 673644 694204
rect 673696 694192 673702 694204
rect 675110 694192 675116 694204
rect 673696 694164 675116 694192
rect 673696 694152 673702 694164
rect 675110 694152 675116 694164
rect 675168 694152 675174 694204
rect 673822 693336 673828 693388
rect 673880 693376 673886 693388
rect 675110 693376 675116 693388
rect 673880 693348 675116 693376
rect 673880 693336 673886 693348
rect 675110 693336 675116 693348
rect 675168 693336 675174 693388
rect 674650 692996 674656 693048
rect 674708 693036 674714 693048
rect 675386 693036 675392 693048
rect 674708 693008 675392 693036
rect 674708 692996 674714 693008
rect 675386 692996 675392 693008
rect 675444 692996 675450 693048
rect 666094 692860 666100 692912
rect 666152 692900 666158 692912
rect 675110 692900 675116 692912
rect 666152 692872 675116 692900
rect 666152 692860 666158 692872
rect 675110 692860 675116 692872
rect 675168 692860 675174 692912
rect 672810 690004 672816 690056
rect 672868 690044 672874 690056
rect 675110 690044 675116 690056
rect 672868 690016 675116 690044
rect 672868 690004 672874 690016
rect 675110 690004 675116 690016
rect 675168 690004 675174 690056
rect 659286 689256 659292 689308
rect 659344 689296 659350 689308
rect 674926 689296 674932 689308
rect 659344 689268 674932 689296
rect 659344 689256 659350 689268
rect 674926 689256 674932 689268
rect 674984 689256 674990 689308
rect 43806 688644 43812 688696
rect 43864 688684 43870 688696
rect 62114 688684 62120 688696
rect 43864 688656 62120 688684
rect 43864 688644 43870 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 674190 687896 674196 687948
rect 674248 687936 674254 687948
rect 675294 687936 675300 687948
rect 674248 687908 675300 687936
rect 674248 687896 674254 687908
rect 675294 687896 675300 687908
rect 675352 687896 675358 687948
rect 43438 687692 43444 687744
rect 43496 687732 43502 687744
rect 50706 687732 50712 687744
rect 43496 687704 50712 687732
rect 43496 687692 43502 687704
rect 50706 687692 50712 687704
rect 50764 687692 50770 687744
rect 671246 687420 671252 687472
rect 671304 687460 671310 687472
rect 675110 687460 675116 687472
rect 671304 687432 675116 687460
rect 671304 687420 671310 687432
rect 675110 687420 675116 687432
rect 675168 687420 675174 687472
rect 43254 687352 43260 687404
rect 43312 687392 43318 687404
rect 51902 687392 51908 687404
rect 43312 687364 51908 687392
rect 43312 687352 43318 687364
rect 51902 687352 51908 687364
rect 51960 687352 51966 687404
rect 40954 687216 40960 687268
rect 41012 687256 41018 687268
rect 41690 687256 41696 687268
rect 41012 687228 41696 687256
rect 41012 687216 41018 687228
rect 41690 687216 41696 687228
rect 41748 687216 41754 687268
rect 42058 687216 42064 687268
rect 42116 687256 42122 687268
rect 56042 687256 56048 687268
rect 42116 687228 56048 687256
rect 42116 687216 42122 687228
rect 56042 687216 56048 687228
rect 56100 687216 56106 687268
rect 41690 686100 41696 686112
rect 41386 686072 41696 686100
rect 41138 685992 41144 686044
rect 41196 686032 41202 686044
rect 41386 686032 41414 686072
rect 41690 686060 41696 686072
rect 41748 686060 41754 686112
rect 42058 686060 42064 686112
rect 42116 686100 42122 686112
rect 44450 686100 44456 686112
rect 42116 686072 44456 686100
rect 42116 686060 42122 686072
rect 44450 686060 44456 686072
rect 44508 686060 44514 686112
rect 41196 686004 41414 686032
rect 41196 685992 41202 686004
rect 41322 685856 41328 685908
rect 41380 685896 41386 685908
rect 41690 685896 41696 685908
rect 41380 685868 41696 685896
rect 41380 685856 41386 685868
rect 41690 685856 41696 685868
rect 41748 685856 41754 685908
rect 42058 685856 42064 685908
rect 42116 685896 42122 685908
rect 45002 685896 45008 685908
rect 42116 685868 45008 685896
rect 42116 685856 42122 685868
rect 45002 685856 45008 685868
rect 45060 685856 45066 685908
rect 669406 685856 669412 685908
rect 669464 685896 669470 685908
rect 669464 685868 675340 685896
rect 669464 685856 669470 685868
rect 675312 685568 675340 685868
rect 675294 685516 675300 685568
rect 675352 685516 675358 685568
rect 40862 684768 40868 684820
rect 40920 684768 40926 684820
rect 40880 684536 40908 684768
rect 41690 684740 41696 684752
rect 41386 684712 41696 684740
rect 41138 684632 41144 684684
rect 41196 684672 41202 684684
rect 41386 684672 41414 684712
rect 41690 684700 41696 684712
rect 41748 684700 41754 684752
rect 42058 684700 42064 684752
rect 42116 684740 42122 684752
rect 42886 684740 42892 684752
rect 42116 684712 42892 684740
rect 42116 684700 42122 684712
rect 42886 684700 42892 684712
rect 42944 684700 42950 684752
rect 41196 684644 41414 684672
rect 41196 684632 41202 684644
rect 41690 684536 41696 684548
rect 40880 684508 41696 684536
rect 41690 684496 41696 684508
rect 41748 684496 41754 684548
rect 42058 684496 42064 684548
rect 42116 684536 42122 684548
rect 44266 684536 44272 684548
rect 42116 684508 44272 684536
rect 42116 684496 42122 684508
rect 44266 684496 44272 684508
rect 44324 684496 44330 684548
rect 41322 683476 41328 683528
rect 41380 683516 41386 683528
rect 41690 683516 41696 683528
rect 41380 683488 41696 683516
rect 41380 683476 41386 683488
rect 41690 683476 41696 683488
rect 41748 683476 41754 683528
rect 651558 683136 651564 683188
rect 651616 683176 651622 683188
rect 659102 683176 659108 683188
rect 651616 683148 659108 683176
rect 651616 683136 651622 683148
rect 659102 683136 659108 683148
rect 659160 683136 659166 683188
rect 675846 682388 675852 682440
rect 675904 682428 675910 682440
rect 683390 682428 683396 682440
rect 675904 682400 683396 682428
rect 675904 682388 675910 682400
rect 683390 682388 683396 682400
rect 683448 682388 683454 682440
rect 40770 679328 40776 679380
rect 40828 679368 40834 679380
rect 41322 679368 41328 679380
rect 40828 679340 41328 679368
rect 40828 679328 40834 679340
rect 41322 679328 41328 679340
rect 41380 679328 41386 679380
rect 40586 679192 40592 679244
rect 40644 679232 40650 679244
rect 41690 679232 41696 679244
rect 40644 679204 41696 679232
rect 40644 679192 40650 679204
rect 41690 679192 41696 679204
rect 41748 679192 41754 679244
rect 43990 676404 43996 676456
rect 44048 676444 44054 676456
rect 50338 676444 50344 676456
rect 44048 676416 50344 676444
rect 44048 676404 44054 676416
rect 50338 676404 50344 676416
rect 50396 676404 50402 676456
rect 47762 674840 47768 674892
rect 47820 674880 47826 674892
rect 62114 674880 62120 674892
rect 47820 674852 62120 674880
rect 47820 674840 47826 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 33778 672732 33784 672784
rect 33836 672772 33842 672784
rect 39482 672772 39488 672784
rect 33836 672744 39488 672772
rect 33836 672732 33842 672744
rect 39482 672732 39488 672744
rect 39540 672732 39546 672784
rect 36538 672052 36544 672104
rect 36596 672092 36602 672104
rect 41690 672092 41696 672104
rect 36596 672064 41696 672092
rect 36596 672052 36602 672064
rect 41690 672052 41696 672064
rect 41748 672052 41754 672104
rect 37918 671236 37924 671288
rect 37976 671276 37982 671288
rect 40034 671276 40040 671288
rect 37976 671248 40040 671276
rect 37976 671236 37982 671248
rect 40034 671236 40040 671248
rect 40092 671236 40098 671288
rect 663242 670828 663248 670880
rect 663300 670868 663306 670880
rect 675294 670868 675300 670880
rect 663300 670840 675300 670868
rect 663300 670828 663306 670840
rect 675294 670828 675300 670840
rect 675352 670828 675358 670880
rect 661862 670692 661868 670744
rect 661920 670732 661926 670744
rect 675478 670732 675484 670744
rect 661920 670704 675484 670732
rect 661920 670692 661926 670704
rect 675478 670692 675484 670704
rect 675536 670692 675542 670744
rect 672994 669740 673000 669792
rect 673052 669780 673058 669792
rect 674834 669780 674840 669792
rect 673052 669752 674840 669780
rect 673052 669740 673058 669752
rect 674834 669740 674840 669752
rect 674892 669740 674898 669792
rect 671522 669604 671528 669656
rect 671580 669644 671586 669656
rect 675294 669644 675300 669656
rect 671580 669616 675300 669644
rect 671580 669604 671586 669616
rect 675294 669604 675300 669616
rect 675352 669604 675358 669656
rect 671614 669468 671620 669520
rect 671672 669508 671678 669520
rect 675478 669508 675484 669520
rect 671672 669480 675484 669508
rect 671672 669468 671678 669480
rect 675478 669468 675484 669480
rect 675536 669468 675542 669520
rect 651558 669332 651564 669384
rect 651616 669372 651622 669384
rect 661862 669372 661868 669384
rect 651616 669344 661868 669372
rect 651616 669332 651622 669344
rect 661862 669332 661868 669344
rect 661920 669332 661926 669384
rect 662046 669332 662052 669384
rect 662104 669372 662110 669384
rect 675478 669372 675484 669384
rect 662104 669344 675484 669372
rect 662104 669332 662110 669344
rect 675478 669332 675484 669344
rect 675536 669332 675542 669384
rect 671062 668516 671068 668568
rect 671120 668556 671126 668568
rect 675478 668556 675484 668568
rect 671120 668528 675484 668556
rect 671120 668516 671126 668528
rect 675478 668516 675484 668528
rect 675536 668516 675542 668568
rect 671062 668380 671068 668432
rect 671120 668420 671126 668432
rect 675294 668420 675300 668432
rect 671120 668392 675300 668420
rect 671120 668380 671126 668392
rect 675294 668380 675300 668392
rect 675352 668380 675358 668432
rect 672350 668040 672356 668092
rect 672408 668080 672414 668092
rect 675478 668080 675484 668092
rect 672408 668052 675484 668080
rect 672408 668040 672414 668052
rect 675478 668040 675484 668052
rect 675536 668040 675542 668092
rect 45186 667944 45192 667956
rect 42260 667916 45192 667944
rect 42260 667820 42288 667916
rect 45186 667904 45192 667916
rect 45244 667904 45250 667956
rect 42242 667768 42248 667820
rect 42300 667768 42306 667820
rect 671430 667700 671436 667752
rect 671488 667740 671494 667752
rect 675478 667740 675484 667752
rect 671488 667712 675484 667740
rect 671488 667700 671494 667712
rect 675478 667700 675484 667712
rect 675536 667700 675542 667752
rect 673270 667224 673276 667276
rect 673328 667264 673334 667276
rect 675478 667264 675484 667276
rect 673328 667236 675484 667264
rect 673328 667224 673334 667236
rect 675478 667224 675484 667236
rect 675536 667224 675542 667276
rect 44634 666584 44640 666596
rect 42260 666556 44640 666584
rect 42260 666052 42288 666556
rect 44634 666544 44640 666556
rect 44692 666544 44698 666596
rect 671982 666068 671988 666120
rect 672040 666108 672046 666120
rect 675478 666108 675484 666120
rect 672040 666080 675484 666108
rect 672040 666068 672046 666080
rect 675478 666068 675484 666080
rect 675536 666068 675542 666120
rect 42242 666000 42248 666052
rect 42300 666000 42306 666052
rect 667658 665320 667664 665372
rect 667716 665360 667722 665372
rect 675294 665360 675300 665372
rect 667716 665332 675300 665360
rect 667716 665320 667722 665332
rect 675294 665320 675300 665332
rect 675352 665320 675358 665372
rect 666370 665184 666376 665236
rect 666428 665224 666434 665236
rect 675478 665224 675484 665236
rect 666428 665196 675484 665224
rect 666428 665184 666434 665196
rect 675478 665184 675484 665196
rect 675536 665184 675542 665236
rect 670418 664844 670424 664896
rect 670476 664884 670482 664896
rect 675478 664884 675484 664896
rect 670476 664856 675484 664884
rect 670476 664844 670482 664856
rect 675478 664844 675484 664856
rect 675536 664844 675542 664896
rect 669222 663756 669228 663808
rect 669280 663796 669286 663808
rect 675478 663796 675484 663808
rect 669280 663768 675484 663796
rect 669280 663756 669286 663768
rect 675478 663756 675484 663768
rect 675536 663756 675542 663808
rect 42518 663280 42524 663332
rect 42576 663280 42582 663332
rect 42334 663212 42340 663264
rect 42392 663212 42398 663264
rect 42352 662708 42380 663212
rect 42536 662992 42564 663280
rect 673454 663212 673460 663264
rect 673512 663252 673518 663264
rect 675478 663252 675484 663264
rect 673512 663224 675484 663252
rect 673512 663212 673518 663224
rect 675478 663212 675484 663224
rect 675536 663212 675542 663264
rect 42702 663008 42708 663060
rect 42760 663048 42766 663060
rect 43438 663048 43444 663060
rect 42760 663020 43444 663048
rect 42760 663008 42766 663020
rect 43438 663008 43444 663020
rect 43496 663008 43502 663060
rect 42518 662940 42524 662992
rect 42576 662940 42582 662992
rect 672534 662804 672540 662856
rect 672592 662844 672598 662856
rect 675478 662844 675484 662856
rect 672592 662816 675484 662844
rect 672592 662804 672598 662816
rect 675478 662804 675484 662816
rect 675536 662804 675542 662856
rect 42518 662708 42524 662720
rect 42352 662680 42524 662708
rect 42518 662668 42524 662680
rect 42576 662668 42582 662720
rect 43438 662396 43444 662448
rect 43496 662436 43502 662448
rect 62114 662436 62120 662448
rect 43496 662408 62120 662436
rect 43496 662396 43502 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 670786 661988 670792 662040
rect 670844 662028 670850 662040
rect 675478 662028 675484 662040
rect 670844 662000 675484 662028
rect 670844 661988 670850 662000
rect 675478 661988 675484 662000
rect 675536 661988 675542 662040
rect 671798 661580 671804 661632
rect 671856 661620 671862 661632
rect 675478 661620 675484 661632
rect 671856 661592 675484 661620
rect 671856 661580 671862 661592
rect 675478 661580 675484 661592
rect 675536 661580 675542 661632
rect 670786 661104 670792 661156
rect 670844 661144 670850 661156
rect 675478 661144 675484 661156
rect 670844 661116 675484 661144
rect 670844 661104 670850 661116
rect 675478 661104 675484 661116
rect 675536 661104 675542 661156
rect 42150 660492 42156 660544
rect 42208 660532 42214 660544
rect 42702 660532 42708 660544
rect 42208 660504 42708 660532
rect 42208 660492 42214 660504
rect 42702 660492 42708 660504
rect 42760 660492 42766 660544
rect 670970 659948 670976 660000
rect 671028 659988 671034 660000
rect 675478 659988 675484 660000
rect 671028 659960 675484 659988
rect 671028 659948 671034 659960
rect 675478 659948 675484 659960
rect 675536 659948 675542 660000
rect 675846 659812 675852 659864
rect 675904 659852 675910 659864
rect 683114 659852 683120 659864
rect 675904 659824 683120 659852
rect 675904 659812 675910 659824
rect 683114 659812 683120 659824
rect 683172 659812 683178 659864
rect 42058 657364 42064 657416
rect 42116 657404 42122 657416
rect 42610 657404 42616 657416
rect 42116 657376 42616 657404
rect 42116 657364 42122 657376
rect 42610 657364 42616 657376
rect 42668 657364 42674 657416
rect 651558 656888 651564 656940
rect 651616 656928 651622 656940
rect 661678 656928 661684 656940
rect 651616 656900 661684 656928
rect 651616 656888 651622 656900
rect 661678 656888 661684 656900
rect 661736 656888 661742 656940
rect 664990 654100 664996 654152
rect 665048 654140 665054 654152
rect 675294 654140 675300 654152
rect 665048 654112 675300 654140
rect 665048 654100 665054 654112
rect 675294 654100 675300 654112
rect 675352 654100 675358 654152
rect 671890 651380 671896 651432
rect 671948 651420 671954 651432
rect 675294 651420 675300 651432
rect 671948 651392 675300 651420
rect 671948 651380 671954 651392
rect 675294 651380 675300 651392
rect 675352 651380 675358 651432
rect 674834 649176 674840 649188
rect 669286 649148 674840 649176
rect 668946 649068 668952 649120
rect 669004 649108 669010 649120
rect 669286 649108 669314 649148
rect 674834 649136 674840 649148
rect 674892 649136 674898 649188
rect 669004 649080 669314 649108
rect 669004 649068 669010 649080
rect 51902 647844 51908 647896
rect 51960 647884 51966 647896
rect 62114 647884 62120 647896
rect 51960 647856 62120 647884
rect 51960 647844 51966 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 669222 647708 669228 647760
rect 669280 647748 669286 647760
rect 675386 647748 675392 647760
rect 669280 647720 675392 647748
rect 669280 647708 669286 647720
rect 675386 647708 675392 647720
rect 675444 647708 675450 647760
rect 35802 644716 35808 644768
rect 35860 644756 35866 644768
rect 39390 644756 39396 644768
rect 35860 644728 39396 644756
rect 35860 644716 35866 644728
rect 39390 644716 39396 644728
rect 39448 644716 39454 644768
rect 35526 644444 35532 644496
rect 35584 644484 35590 644496
rect 39758 644484 39764 644496
rect 35584 644456 39764 644484
rect 35584 644444 35590 644456
rect 39758 644444 39764 644456
rect 39816 644444 39822 644496
rect 670234 644444 670240 644496
rect 670292 644484 670298 644496
rect 674834 644484 674840 644496
rect 670292 644456 674840 644484
rect 670292 644444 670298 644456
rect 674834 644444 674840 644456
rect 674892 644444 674898 644496
rect 661862 643696 661868 643748
rect 661920 643736 661926 643748
rect 661920 643708 666554 643736
rect 661920 643696 661926 643708
rect 666526 643668 666554 643708
rect 675294 643668 675300 643680
rect 666526 643640 675300 643668
rect 675294 643628 675300 643640
rect 675352 643628 675358 643680
rect 35802 643492 35808 643544
rect 35860 643532 35866 643544
rect 39666 643532 39672 643544
rect 35860 643504 39672 643532
rect 35860 643492 35866 643504
rect 39666 643492 39672 643504
rect 39724 643492 39730 643544
rect 41690 643328 41696 643340
rect 41386 643300 41696 643328
rect 35526 643220 35532 643272
rect 35584 643260 35590 643272
rect 41386 643260 41414 643300
rect 41690 643288 41696 643300
rect 41748 643288 41754 643340
rect 42058 643288 42064 643340
rect 42116 643328 42122 643340
rect 44450 643328 44456 643340
rect 42116 643300 44456 643328
rect 42116 643288 42122 643300
rect 44450 643288 44456 643300
rect 44508 643288 44514 643340
rect 35584 643232 41414 643260
rect 35584 643220 35590 643232
rect 35342 643084 35348 643136
rect 35400 643124 35406 643136
rect 41690 643124 41696 643136
rect 35400 643096 41696 643124
rect 35400 643084 35406 643096
rect 41690 643084 41696 643096
rect 41748 643084 41754 643136
rect 42058 643084 42064 643136
rect 42116 643124 42122 643136
rect 51718 643124 51724 643136
rect 42116 643096 51724 643124
rect 42116 643084 42122 643096
rect 51718 643084 51724 643096
rect 51776 643084 51782 643136
rect 651558 643084 651564 643136
rect 651616 643124 651622 643136
rect 663242 643124 663248 643136
rect 651616 643096 663248 643124
rect 651616 643084 651622 643096
rect 663242 643084 663248 643096
rect 663300 643084 663306 643136
rect 38930 642240 38936 642252
rect 38626 642212 38936 642240
rect 35802 642132 35808 642184
rect 35860 642172 35866 642184
rect 38626 642172 38654 642212
rect 38930 642200 38936 642212
rect 38988 642200 38994 642252
rect 35860 642144 38654 642172
rect 35860 642132 35866 642144
rect 39574 642036 39580 642048
rect 36004 642008 39580 642036
rect 35434 641860 35440 641912
rect 35492 641900 35498 641912
rect 36004 641900 36032 642008
rect 39574 641996 39580 642008
rect 39632 641996 39638 642048
rect 35492 641872 36032 641900
rect 35492 641860 35498 641872
rect 666278 641860 666284 641912
rect 666336 641900 666342 641912
rect 674834 641900 674840 641912
rect 666336 641872 674840 641900
rect 666336 641860 666342 641872
rect 674834 641860 674840 641872
rect 674892 641860 674898 641912
rect 35618 641724 35624 641776
rect 35676 641764 35682 641776
rect 41690 641764 41696 641776
rect 35676 641736 41696 641764
rect 35676 641724 35682 641736
rect 41690 641724 41696 641736
rect 41748 641724 41754 641776
rect 42058 641724 42064 641776
rect 42116 641764 42122 641776
rect 44174 641764 44180 641776
rect 42116 641736 44180 641764
rect 42116 641724 42122 641736
rect 44174 641724 44180 641736
rect 44232 641724 44238 641776
rect 665910 641724 665916 641776
rect 665968 641764 665974 641776
rect 670418 641764 670424 641776
rect 665968 641736 670424 641764
rect 665968 641724 665974 641736
rect 670418 641724 670424 641736
rect 670476 641724 670482 641776
rect 670418 641248 670424 641300
rect 670476 641288 670482 641300
rect 675294 641288 675300 641300
rect 670476 641260 675300 641288
rect 670476 641248 670482 641260
rect 675294 641248 675300 641260
rect 675352 641248 675358 641300
rect 35802 640772 35808 640824
rect 35860 640812 35866 640824
rect 35860 640772 35894 640812
rect 35866 640744 35894 640772
rect 39666 640744 39672 640756
rect 35866 640716 39672 640744
rect 39666 640704 39672 640716
rect 39724 640704 39730 640756
rect 673638 640568 673644 640620
rect 673696 640568 673702 640620
rect 673822 640568 673828 640620
rect 673880 640568 673886 640620
rect 35618 640432 35624 640484
rect 35676 640472 35682 640484
rect 39850 640472 39856 640484
rect 35676 640444 39856 640472
rect 35676 640432 35682 640444
rect 39850 640432 39856 640444
rect 39908 640432 39914 640484
rect 673656 640348 673684 640568
rect 673840 640348 673868 640568
rect 35802 640296 35808 640348
rect 35860 640336 35866 640348
rect 41690 640336 41696 640348
rect 35860 640308 41696 640336
rect 35860 640296 35866 640308
rect 41690 640296 41696 640308
rect 41748 640296 41754 640348
rect 42058 640296 42064 640348
rect 42116 640336 42122 640348
rect 43070 640336 43076 640348
rect 42116 640308 43076 640336
rect 42116 640296 42122 640308
rect 43070 640296 43076 640308
rect 43128 640296 43134 640348
rect 673638 640296 673644 640348
rect 673696 640296 673702 640348
rect 673822 640296 673828 640348
rect 673880 640296 673886 640348
rect 35802 639072 35808 639124
rect 35860 639112 35866 639124
rect 40218 639112 40224 639124
rect 35860 639084 40224 639112
rect 35860 639072 35866 639084
rect 40218 639072 40224 639084
rect 40276 639072 40282 639124
rect 35526 638936 35532 638988
rect 35584 638976 35590 638988
rect 40034 638976 40040 638988
rect 35584 638948 40040 638976
rect 35584 638936 35590 638948
rect 40034 638936 40040 638948
rect 40092 638936 40098 638988
rect 35342 638188 35348 638240
rect 35400 638228 35406 638240
rect 41690 638228 41696 638240
rect 35400 638200 41696 638228
rect 35400 638188 35406 638200
rect 41690 638188 41696 638200
rect 41748 638188 41754 638240
rect 35526 637916 35532 637968
rect 35584 637956 35590 637968
rect 40954 637956 40960 637968
rect 35584 637928 40960 637956
rect 35584 637916 35590 637928
rect 40954 637916 40960 637928
rect 41012 637916 41018 637968
rect 35802 637712 35808 637764
rect 35860 637752 35866 637764
rect 41506 637752 41512 637764
rect 35860 637724 41512 637752
rect 35860 637712 35866 637724
rect 41506 637712 41512 637724
rect 41564 637712 41570 637764
rect 676030 637508 676036 637560
rect 676088 637548 676094 637560
rect 682378 637548 682384 637560
rect 676088 637520 682384 637548
rect 676088 637508 676094 637520
rect 682378 637508 682384 637520
rect 682436 637508 682442 637560
rect 676030 636828 676036 636880
rect 676088 636868 676094 636880
rect 683298 636868 683304 636880
rect 676088 636840 683304 636868
rect 676088 636828 676094 636840
rect 683298 636828 683304 636840
rect 683356 636828 683362 636880
rect 35802 636352 35808 636404
rect 35860 636392 35866 636404
rect 40678 636392 40684 636404
rect 35860 636364 40684 636392
rect 35860 636352 35866 636364
rect 40678 636352 40684 636364
rect 40736 636352 40742 636404
rect 49142 636216 49148 636268
rect 49200 636256 49206 636268
rect 62114 636256 62120 636268
rect 49200 636228 62120 636256
rect 49200 636216 49206 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 35802 635060 35808 635112
rect 35860 635100 35866 635112
rect 39574 635100 39580 635112
rect 35860 635072 39580 635100
rect 35860 635060 35866 635072
rect 39574 635060 39580 635072
rect 39632 635060 39638 635112
rect 35618 634788 35624 634840
rect 35676 634828 35682 634840
rect 40494 634828 40500 634840
rect 35676 634800 40500 634828
rect 35676 634788 35682 634800
rect 40494 634788 40500 634800
rect 40552 634788 40558 634840
rect 35802 633836 35808 633888
rect 35860 633876 35866 633888
rect 35860 633836 35894 633876
rect 35866 633740 35894 633836
rect 41690 633740 41696 633752
rect 35866 633712 41696 633740
rect 41690 633700 41696 633712
rect 41748 633700 41754 633752
rect 42058 633700 42064 633752
rect 42116 633740 42122 633752
rect 53282 633740 53288 633752
rect 42116 633712 53288 633740
rect 42116 633700 42122 633712
rect 53282 633700 53288 633712
rect 53340 633700 53346 633752
rect 51718 633604 51724 633616
rect 48286 633576 51724 633604
rect 35802 633496 35808 633548
rect 35860 633536 35866 633548
rect 41690 633536 41696 633548
rect 35860 633508 41696 633536
rect 35860 633496 35866 633508
rect 41690 633496 41696 633508
rect 41748 633496 41754 633548
rect 42058 633496 42064 633548
rect 42116 633536 42122 633548
rect 48286 633536 48314 633576
rect 51718 633564 51724 633576
rect 51776 633564 51782 633616
rect 675846 633564 675852 633616
rect 675904 633604 675910 633616
rect 682562 633604 682568 633616
rect 675904 633576 682568 633604
rect 675904 633564 675910 633576
rect 682562 633564 682568 633576
rect 682620 633564 682626 633616
rect 42116 633508 48314 633536
rect 42116 633496 42122 633508
rect 33778 630028 33784 630080
rect 33836 630068 33842 630080
rect 41690 630068 41696 630080
rect 33836 630040 41696 630068
rect 33836 630028 33842 630040
rect 41690 630028 41696 630040
rect 41748 630028 41754 630080
rect 42058 629960 42064 630012
rect 42116 630000 42122 630012
rect 42702 630000 42708 630012
rect 42116 629972 42708 630000
rect 42116 629960 42122 629972
rect 42702 629960 42708 629972
rect 42760 629960 42766 630012
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41690 629932 41696 629944
rect 32456 629904 41696 629932
rect 32456 629892 32462 629904
rect 41690 629892 41696 629904
rect 41748 629892 41754 629944
rect 651558 629280 651564 629332
rect 651616 629320 651622 629332
rect 661862 629320 661868 629332
rect 651616 629292 661868 629320
rect 651616 629280 651622 629292
rect 661862 629280 661868 629292
rect 661920 629280 661926 629332
rect 42886 626628 42892 626680
rect 42944 626668 42950 626680
rect 50522 626668 50528 626680
rect 42944 626640 50528 626668
rect 42944 626628 42950 626640
rect 50522 626628 50528 626640
rect 50580 626628 50586 626680
rect 664438 625676 664444 625728
rect 664496 625716 664502 625728
rect 675478 625716 675484 625728
rect 664496 625688 675484 625716
rect 664496 625676 664502 625688
rect 675478 625676 675484 625688
rect 675536 625676 675542 625728
rect 663058 625404 663064 625456
rect 663116 625444 663122 625456
rect 663116 625416 663794 625444
rect 663116 625404 663122 625416
rect 42518 625336 42524 625388
rect 42576 625336 42582 625388
rect 42242 625132 42248 625184
rect 42300 625172 42306 625184
rect 42536 625172 42564 625336
rect 663766 625308 663794 625416
rect 675478 625308 675484 625320
rect 663766 625280 675484 625308
rect 675478 625268 675484 625280
rect 675536 625268 675542 625320
rect 42300 625144 42564 625172
rect 42300 625132 42306 625144
rect 660298 625132 660304 625184
rect 660356 625172 660362 625184
rect 675110 625172 675116 625184
rect 660356 625144 675116 625172
rect 660356 625132 660362 625144
rect 675110 625132 675116 625144
rect 675168 625132 675174 625184
rect 671522 624928 671528 624980
rect 671580 624968 671586 624980
rect 675478 624968 675484 624980
rect 671580 624940 675484 624968
rect 671580 624928 671586 624940
rect 675478 624928 675484 624940
rect 675536 624928 675542 624980
rect 42334 624656 42340 624708
rect 42392 624696 42398 624708
rect 43806 624696 43812 624708
rect 42392 624668 43812 624696
rect 42392 624656 42398 624668
rect 43806 624656 43812 624668
rect 43864 624656 43870 624708
rect 672902 624656 672908 624708
rect 672960 624696 672966 624708
rect 675478 624696 675484 624708
rect 672960 624668 675484 624696
rect 672960 624656 672966 624668
rect 675478 624656 675484 624668
rect 675536 624656 675542 624708
rect 671154 624316 671160 624368
rect 671212 624356 671218 624368
rect 675478 624356 675484 624368
rect 671212 624328 675484 624356
rect 671212 624316 671218 624328
rect 675478 624316 675484 624328
rect 675536 624316 675542 624368
rect 47762 623772 47768 623824
rect 47820 623812 47826 623824
rect 62114 623812 62120 623824
rect 47820 623784 62120 623812
rect 47820 623772 47826 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 672350 623500 672356 623552
rect 672408 623540 672414 623552
rect 675478 623540 675484 623552
rect 672408 623512 675484 623540
rect 672408 623500 672414 623512
rect 675478 623500 675484 623512
rect 675536 623500 675542 623552
rect 671522 623024 671528 623076
rect 671580 623064 671586 623076
rect 675478 623064 675484 623076
rect 671580 623036 675484 623064
rect 671580 623024 671586 623036
rect 675478 623024 675484 623036
rect 675536 623024 675542 623076
rect 673454 622888 673460 622940
rect 673512 622888 673518 622940
rect 673472 622736 673500 622888
rect 673454 622684 673460 622736
rect 673512 622684 673518 622736
rect 673638 622684 673644 622736
rect 673696 622724 673702 622736
rect 675478 622724 675484 622736
rect 673696 622696 675484 622724
rect 673696 622684 673702 622696
rect 675478 622684 675484 622696
rect 675536 622684 675542 622736
rect 672074 622208 672080 622260
rect 672132 622248 672138 622260
rect 675478 622248 675484 622260
rect 672132 622220 675484 622248
rect 672132 622208 672138 622220
rect 675478 622208 675484 622220
rect 675536 622208 675542 622260
rect 669406 619828 669412 619880
rect 669464 619868 669470 619880
rect 675018 619868 675024 619880
rect 669464 619840 675024 619868
rect 669464 619828 669470 619840
rect 675018 619828 675024 619840
rect 675076 619828 675082 619880
rect 666094 619624 666100 619676
rect 666152 619664 666158 619676
rect 675478 619664 675484 619676
rect 666152 619636 675484 619664
rect 666152 619624 666158 619636
rect 675478 619624 675484 619636
rect 675536 619624 675542 619676
rect 673086 619080 673092 619132
rect 673144 619120 673150 619132
rect 674834 619120 674840 619132
rect 673144 619092 674840 619120
rect 673144 619080 673150 619092
rect 674834 619080 674840 619092
rect 674892 619080 674898 619132
rect 42610 618876 42616 618928
rect 42668 618916 42674 618928
rect 43622 618916 43628 618928
rect 42668 618888 43628 618916
rect 42668 618876 42674 618888
rect 43622 618876 43628 618888
rect 43680 618876 43686 618928
rect 668762 618264 668768 618316
rect 668820 618304 668826 618316
rect 675478 618304 675484 618316
rect 668820 618276 675484 618304
rect 668820 618264 668826 618276
rect 675478 618264 675484 618276
rect 675536 618264 675542 618316
rect 671338 618128 671344 618180
rect 671396 618168 671402 618180
rect 675478 618168 675484 618180
rect 671396 618140 675484 618168
rect 671396 618128 671402 618140
rect 675478 618128 675484 618140
rect 675536 618128 675542 618180
rect 673270 616972 673276 617024
rect 673328 617012 673334 617024
rect 675478 617012 675484 617024
rect 673328 616984 675484 617012
rect 673328 616972 673334 616984
rect 675478 616972 675484 616984
rect 675536 616972 675542 617024
rect 651558 616836 651564 616888
rect 651616 616876 651622 616888
rect 660482 616876 660488 616888
rect 651616 616848 660488 616876
rect 651616 616836 651622 616848
rect 660482 616836 660488 616848
rect 660540 616836 660546 616888
rect 668578 616768 668584 616820
rect 668636 616808 668642 616820
rect 669774 616808 669780 616820
rect 668636 616780 669780 616808
rect 668636 616768 668642 616780
rect 669774 616768 669780 616780
rect 669832 616768 669838 616820
rect 672718 616564 672724 616616
rect 672776 616604 672782 616616
rect 675478 616604 675484 616616
rect 672776 616576 675484 616604
rect 672776 616564 672782 616576
rect 675478 616564 675484 616576
rect 675536 616564 675542 616616
rect 670418 616088 670424 616140
rect 670476 616128 670482 616140
rect 675478 616128 675484 616140
rect 670476 616100 675484 616128
rect 670476 616088 670482 616100
rect 675478 616088 675484 616100
rect 675536 616088 675542 616140
rect 42242 615680 42248 615732
rect 42300 615680 42306 615732
rect 42260 615528 42288 615680
rect 675846 615612 675852 615664
rect 675904 615652 675910 615664
rect 683114 615652 683120 615664
rect 675904 615624 683120 615652
rect 675904 615612 675910 615624
rect 683114 615612 683120 615624
rect 683172 615612 683178 615664
rect 42242 615476 42248 615528
rect 42300 615476 42306 615528
rect 672166 614864 672172 614916
rect 672224 614904 672230 614916
rect 675478 614904 675484 614916
rect 672224 614876 675484 614904
rect 672224 614864 672230 614876
rect 675478 614864 675484 614876
rect 675536 614864 675542 614916
rect 42150 613572 42156 613624
rect 42208 613612 42214 613624
rect 44358 613612 44364 613624
rect 42208 613584 44364 613612
rect 42208 613572 42214 613584
rect 44358 613572 44364 613584
rect 44416 613572 44422 613624
rect 43622 609220 43628 609272
rect 43680 609260 43686 609272
rect 62114 609260 62120 609272
rect 43680 609232 62120 609260
rect 43680 609220 43686 609232
rect 62114 609220 62120 609232
rect 62172 609220 62178 609272
rect 675202 608852 675208 608864
rect 663766 608824 675208 608852
rect 663518 608608 663524 608660
rect 663576 608648 663582 608660
rect 663766 608648 663794 608824
rect 675202 608812 675208 608824
rect 675260 608812 675266 608864
rect 663576 608620 663794 608648
rect 663576 608608 663582 608620
rect 670326 607112 670332 607164
rect 670384 607112 670390 607164
rect 670142 606840 670148 606892
rect 670200 606880 670206 606892
rect 670344 606880 670372 607112
rect 670200 606852 670372 606880
rect 670200 606840 670206 606852
rect 674282 604324 674288 604376
rect 674340 604364 674346 604376
rect 675294 604364 675300 604376
rect 674340 604336 675300 604364
rect 674340 604324 674346 604336
rect 675294 604324 675300 604336
rect 675352 604324 675358 604376
rect 673638 603440 673644 603492
rect 673696 603480 673702 603492
rect 675386 603480 675392 603492
rect 673696 603452 675392 603480
rect 673696 603440 673702 603452
rect 675386 603440 675392 603452
rect 675444 603440 675450 603492
rect 652570 603100 652576 603152
rect 652628 603140 652634 603152
rect 660298 603140 660304 603152
rect 652628 603112 660304 603140
rect 652628 603100 652634 603112
rect 660298 603100 660304 603112
rect 660356 603100 660362 603152
rect 667842 603100 667848 603152
rect 667900 603140 667906 603152
rect 674834 603140 674840 603152
rect 667900 603112 674840 603140
rect 667900 603100 667906 603112
rect 674834 603100 674840 603112
rect 674892 603100 674898 603152
rect 35802 601672 35808 601724
rect 35860 601712 35866 601724
rect 41690 601712 41696 601724
rect 35860 601684 41696 601712
rect 35860 601672 35866 601684
rect 41690 601672 41696 601684
rect 41748 601672 41754 601724
rect 42058 601672 42064 601724
rect 42116 601712 42122 601724
rect 49142 601712 49148 601724
rect 42116 601684 49148 601712
rect 42116 601672 42122 601684
rect 49142 601672 49148 601684
rect 49200 601672 49206 601724
rect 670418 601672 670424 601724
rect 670476 601712 670482 601724
rect 675294 601712 675300 601724
rect 670476 601684 675300 601712
rect 670476 601672 670482 601684
rect 675294 601672 675300 601684
rect 675352 601672 675358 601724
rect 43806 600380 43812 600432
rect 43864 600420 43870 600432
rect 43864 600392 51074 600420
rect 43864 600380 43870 600392
rect 51046 600352 51074 600392
rect 51902 600352 51908 600364
rect 51046 600324 51908 600352
rect 51902 600312 51908 600324
rect 51960 600312 51966 600364
rect 660482 599564 660488 599616
rect 660540 599604 660546 599616
rect 675294 599604 675300 599616
rect 660540 599576 675300 599604
rect 660540 599564 660546 599576
rect 675294 599564 675300 599576
rect 675352 599564 675358 599616
rect 41322 598952 41328 599004
rect 41380 598992 41386 599004
rect 41690 598992 41696 599004
rect 41380 598964 41696 598992
rect 41380 598952 41386 598964
rect 41690 598952 41696 598964
rect 41748 598952 41754 599004
rect 42058 598952 42064 599004
rect 42116 598992 42122 599004
rect 44450 598992 44456 599004
rect 42116 598964 44456 598992
rect 42116 598952 42122 598964
rect 44450 598952 44456 598964
rect 44508 598952 44514 599004
rect 41690 597904 41696 597916
rect 41386 597876 41696 597904
rect 41046 597796 41052 597848
rect 41104 597836 41110 597848
rect 41386 597836 41414 597876
rect 41690 597864 41696 597876
rect 41748 597864 41754 597916
rect 42058 597864 42064 597916
rect 42116 597904 42122 597916
rect 42886 597904 42892 597916
rect 42116 597876 42892 597904
rect 42116 597864 42122 597876
rect 42886 597864 42892 597876
rect 42944 597864 42950 597916
rect 41104 597808 41414 597836
rect 41104 597796 41110 597808
rect 41690 597768 41696 597780
rect 41524 597740 41696 597768
rect 40862 597660 40868 597712
rect 40920 597700 40926 597712
rect 41524 597700 41552 597740
rect 41690 597728 41696 597740
rect 41748 597728 41754 597780
rect 42058 597728 42064 597780
rect 42116 597768 42122 597780
rect 43162 597768 43168 597780
rect 42116 597740 43168 597768
rect 42116 597728 42122 597740
rect 43162 597728 43168 597740
rect 43220 597728 43226 597780
rect 40920 597672 41552 597700
rect 40920 597660 40926 597672
rect 41322 597524 41328 597576
rect 41380 597564 41386 597576
rect 41690 597564 41696 597576
rect 41380 597536 41696 597564
rect 41380 597524 41386 597536
rect 41690 597524 41696 597536
rect 41748 597524 41754 597576
rect 42058 597524 42064 597576
rect 42116 597564 42122 597576
rect 43806 597564 43812 597576
rect 42116 597536 43812 597564
rect 42116 597524 42122 597536
rect 43806 597524 43812 597536
rect 43864 597524 43870 597576
rect 49142 597524 49148 597576
rect 49200 597564 49206 597576
rect 62114 597564 62120 597576
rect 49200 597536 62120 597564
rect 49200 597524 49206 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 666094 596164 666100 596216
rect 666152 596204 666158 596216
rect 674742 596204 674748 596216
rect 666152 596176 674748 596204
rect 666152 596164 666158 596176
rect 674742 596164 674748 596176
rect 674800 596164 674806 596216
rect 41138 595892 41144 595944
rect 41196 595932 41202 595944
rect 41690 595932 41696 595944
rect 41196 595904 41696 595932
rect 41196 595892 41202 595904
rect 41690 595892 41696 595904
rect 41748 595892 41754 595944
rect 668762 595212 668768 595264
rect 668820 595252 668826 595264
rect 675294 595252 675300 595264
rect 668820 595224 675300 595252
rect 668820 595212 668826 595224
rect 675294 595212 675300 595224
rect 675352 595212 675358 595264
rect 674742 595008 674748 595060
rect 674800 595048 674806 595060
rect 675294 595048 675300 595060
rect 674800 595020 675300 595048
rect 674800 595008 674806 595020
rect 675294 595008 675300 595020
rect 675352 595008 675358 595060
rect 40770 592832 40776 592884
rect 40828 592872 40834 592884
rect 41690 592872 41696 592884
rect 40828 592844 41696 592872
rect 40828 592832 40834 592844
rect 41690 592832 41696 592844
rect 41748 592832 41754 592884
rect 675846 592628 675852 592680
rect 675904 592668 675910 592680
rect 683298 592668 683304 592680
rect 675904 592640 683304 592668
rect 675904 592628 675910 592640
rect 683298 592628 683304 592640
rect 683356 592628 683362 592680
rect 675846 592492 675852 592544
rect 675904 592532 675910 592544
rect 678238 592532 678244 592544
rect 675904 592504 678244 592532
rect 675904 592492 675910 592504
rect 678238 592492 678244 592504
rect 678296 592492 678302 592544
rect 42058 591880 42064 591932
rect 42116 591920 42122 591932
rect 42426 591920 42432 591932
rect 42116 591892 42432 591920
rect 42116 591880 42122 591892
rect 42426 591880 42432 591892
rect 42484 591880 42490 591932
rect 675846 591404 675852 591456
rect 675904 591444 675910 591456
rect 683482 591444 683488 591456
rect 675904 591416 683488 591444
rect 675904 591404 675910 591416
rect 683482 591404 683488 591416
rect 683540 591404 683546 591456
rect 675846 591268 675852 591320
rect 675904 591308 675910 591320
rect 684126 591308 684132 591320
rect 675904 591280 684132 591308
rect 675904 591268 675910 591280
rect 684126 591268 684132 591280
rect 684184 591268 684190 591320
rect 43254 590792 43260 590844
rect 43312 590832 43318 590844
rect 50522 590832 50528 590844
rect 43312 590804 50528 590832
rect 43312 590792 43318 590804
rect 50522 590792 50528 590804
rect 50580 590792 50586 590844
rect 651558 590656 651564 590708
rect 651616 590696 651622 590708
rect 664438 590696 664444 590708
rect 651616 590668 664444 590696
rect 651616 590656 651622 590668
rect 664438 590656 664444 590668
rect 664496 590656 664502 590708
rect 668762 589228 668768 589280
rect 668820 589268 668826 589280
rect 669406 589268 669412 589280
rect 668820 589240 669412 589268
rect 668820 589228 668826 589240
rect 669406 589228 669412 589240
rect 669464 589228 669470 589280
rect 33042 587120 33048 587172
rect 33100 587160 33106 587172
rect 39574 587160 39580 587172
rect 33100 587132 39580 587160
rect 33100 587120 33106 587132
rect 39574 587120 39580 587132
rect 39632 587120 39638 587172
rect 36538 586372 36544 586424
rect 36596 586412 36602 586424
rect 39574 586412 39580 586424
rect 36596 586384 39580 586412
rect 36596 586372 36602 586384
rect 39574 586372 39580 586384
rect 39632 586372 39638 586424
rect 35158 585896 35164 585948
rect 35216 585936 35222 585948
rect 40494 585936 40500 585948
rect 35216 585908 40500 585936
rect 35216 585896 35222 585908
rect 40494 585896 40500 585908
rect 40552 585896 40558 585948
rect 31018 585556 31024 585608
rect 31076 585596 31082 585608
rect 39666 585596 39672 585608
rect 31076 585568 39672 585596
rect 31076 585556 31082 585568
rect 39666 585556 39672 585568
rect 39724 585556 39730 585608
rect 51902 583720 51908 583772
rect 51960 583760 51966 583772
rect 62114 583760 62120 583772
rect 51960 583732 62120 583760
rect 51960 583720 51966 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 43162 581000 43168 581052
rect 43220 581040 43226 581052
rect 44634 581040 44640 581052
rect 43220 581012 44640 581040
rect 43220 581000 43226 581012
rect 44634 581000 44640 581012
rect 44692 581000 44698 581052
rect 664622 581000 664628 581052
rect 664680 581040 664686 581052
rect 675478 581040 675484 581052
rect 664680 581012 675484 581040
rect 664680 581000 664686 581012
rect 675478 581000 675484 581012
rect 675536 581000 675542 581052
rect 672994 579980 673000 580032
rect 673052 580020 673058 580032
rect 675478 580020 675484 580032
rect 673052 579992 675484 580020
rect 673052 579980 673058 579992
rect 675478 579980 675484 579992
rect 675536 579980 675542 580032
rect 658918 579776 658924 579828
rect 658976 579816 658982 579828
rect 674926 579816 674932 579828
rect 658976 579788 674932 579816
rect 658976 579776 658982 579788
rect 674926 579776 674932 579788
rect 674984 579776 674990 579828
rect 659102 579640 659108 579692
rect 659160 579680 659166 579692
rect 675294 579680 675300 579692
rect 659160 579652 675300 579680
rect 659160 579640 659166 579652
rect 675294 579640 675300 579652
rect 675352 579640 675358 579692
rect 673270 578484 673276 578536
rect 673328 578524 673334 578536
rect 675294 578524 675300 578536
rect 673328 578496 675300 578524
rect 673328 578484 673334 578496
rect 675294 578484 675300 578496
rect 675352 578484 675358 578536
rect 42242 578416 42248 578468
rect 42300 578416 42306 578468
rect 42260 577856 42288 578416
rect 673086 578348 673092 578400
rect 673144 578388 673150 578400
rect 675478 578388 675484 578400
rect 673144 578360 675484 578388
rect 673144 578348 673150 578360
rect 675478 578348 675484 578360
rect 675536 578348 675542 578400
rect 672902 578212 672908 578264
rect 672960 578252 672966 578264
rect 674926 578252 674932 578264
rect 672960 578224 674932 578252
rect 672960 578212 672966 578224
rect 674926 578212 674932 578224
rect 674984 578212 674990 578264
rect 42242 577804 42248 577856
rect 42300 577804 42306 577856
rect 673454 577600 673460 577652
rect 673512 577640 673518 577652
rect 675478 577640 675484 577652
rect 673512 577612 675484 577640
rect 673512 577600 673518 577612
rect 675478 577600 675484 577612
rect 675536 577600 675542 577652
rect 671338 577260 671344 577312
rect 671396 577300 671402 577312
rect 675294 577300 675300 577312
rect 671396 577272 675300 577300
rect 671396 577260 671402 577272
rect 675294 577260 675300 577272
rect 675352 577260 675358 577312
rect 671982 577124 671988 577176
rect 672040 577164 672046 577176
rect 675478 577164 675484 577176
rect 672040 577136 675484 577164
rect 672040 577124 672046 577136
rect 675478 577124 675484 577136
rect 675536 577124 675542 577176
rect 671522 576988 671528 577040
rect 671580 577028 671586 577040
rect 673362 577028 673368 577040
rect 671580 577000 673368 577028
rect 671580 576988 671586 577000
rect 673362 576988 673368 577000
rect 673420 576988 673426 577040
rect 675478 576960 675484 576972
rect 673564 576932 675484 576960
rect 651558 576852 651564 576904
rect 651616 576892 651622 576904
rect 659286 576892 659292 576904
rect 651616 576864 659292 576892
rect 651616 576852 651622 576864
rect 659286 576852 659292 576864
rect 659344 576852 659350 576904
rect 671154 576852 671160 576904
rect 671212 576892 671218 576904
rect 673564 576892 673592 576932
rect 675478 576920 675484 576932
rect 675536 576920 675542 576972
rect 671212 576864 673592 576892
rect 671212 576852 671218 576864
rect 671890 575492 671896 575544
rect 671948 575532 671954 575544
rect 675478 575532 675484 575544
rect 671948 575504 675484 575532
rect 671948 575492 671954 575504
rect 675478 575492 675484 575504
rect 675536 575492 675542 575544
rect 672534 574336 672540 574388
rect 672592 574376 672598 574388
rect 675478 574376 675484 574388
rect 672592 574348 675484 574376
rect 672592 574336 672598 574348
rect 675478 574336 675484 574348
rect 675536 574336 675542 574388
rect 666278 574200 666284 574252
rect 666336 574240 666342 574252
rect 675294 574240 675300 574252
rect 666336 574212 675300 574240
rect 666336 574200 666342 574212
rect 675294 574200 675300 574212
rect 675352 574200 675358 574252
rect 664990 574064 664996 574116
rect 665048 574104 665054 574116
rect 675478 574104 675484 574116
rect 665048 574076 675484 574104
rect 665048 574064 665054 574076
rect 675478 574064 675484 574076
rect 675536 574064 675542 574116
rect 42150 573452 42156 573504
rect 42208 573492 42214 573504
rect 42610 573492 42616 573504
rect 42208 573464 42616 573492
rect 42208 573452 42214 573464
rect 42610 573452 42616 573464
rect 42668 573452 42674 573504
rect 670234 572840 670240 572892
rect 670292 572880 670298 572892
rect 675478 572880 675484 572892
rect 670292 572852 675484 572880
rect 670292 572840 670298 572852
rect 675478 572840 675484 572852
rect 675536 572840 675542 572892
rect 668854 572704 668860 572756
rect 668912 572744 668918 572756
rect 675294 572744 675300 572756
rect 668912 572716 675300 572744
rect 668912 572704 668918 572716
rect 675294 572704 675300 572716
rect 675352 572704 675358 572756
rect 43438 571344 43444 571396
rect 43496 571384 43502 571396
rect 62114 571384 62120 571396
rect 43496 571356 62120 571384
rect 43496 571344 43502 571356
rect 62114 571344 62120 571356
rect 62172 571344 62178 571396
rect 671706 571208 671712 571260
rect 671764 571248 671770 571260
rect 675294 571248 675300 571260
rect 671764 571220 675300 571248
rect 671764 571208 671770 571220
rect 675294 571208 675300 571220
rect 675352 571208 675358 571260
rect 675846 570052 675852 570104
rect 675904 570092 675910 570104
rect 683114 570092 683120 570104
rect 675904 570064 683120 570092
rect 675904 570052 675910 570064
rect 683114 570052 683120 570064
rect 683172 570052 683178 570104
rect 665910 569984 665916 570036
rect 665968 570024 665974 570036
rect 675478 570024 675484 570036
rect 665968 569996 675484 570024
rect 665968 569984 665974 569996
rect 675478 569984 675484 569996
rect 675536 569984 675542 570036
rect 671338 569576 671344 569628
rect 671396 569616 671402 569628
rect 675478 569616 675484 569628
rect 671396 569588 675484 569616
rect 671396 569576 671402 569588
rect 675478 569576 675484 569588
rect 675536 569576 675542 569628
rect 675846 565156 675852 565208
rect 675904 565196 675910 565208
rect 676214 565196 676220 565208
rect 675904 565168 676220 565196
rect 675904 565156 675910 565168
rect 676214 565156 676220 565168
rect 676272 565156 676278 565208
rect 664990 564544 664996 564596
rect 665048 564584 665054 564596
rect 675294 564584 675300 564596
rect 665048 564556 675300 564584
rect 665048 564544 665054 564556
rect 675294 564544 675300 564556
rect 675352 564544 675358 564596
rect 663702 564408 663708 564460
rect 663760 564448 663766 564460
rect 675478 564448 675484 564460
rect 663760 564420 675484 564448
rect 663760 564408 663766 564420
rect 675478 564408 675484 564420
rect 675536 564408 675542 564460
rect 652386 563048 652392 563100
rect 652444 563088 652450 563100
rect 658918 563088 658924 563100
rect 652444 563060 658924 563088
rect 652444 563048 652450 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 674650 558220 674656 558272
rect 674708 558260 674714 558272
rect 675386 558260 675392 558272
rect 674708 558232 675392 558260
rect 674708 558220 674714 558232
rect 675386 558220 675392 558232
rect 675444 558220 675450 558272
rect 43438 557812 43444 557864
rect 43496 557852 43502 557864
rect 49142 557852 49148 557864
rect 43496 557824 49148 557852
rect 43496 557812 43502 557824
rect 49142 557812 49148 557824
rect 49200 557812 49206 557864
rect 673270 557676 673276 557728
rect 673328 557716 673334 557728
rect 675294 557716 675300 557728
rect 673328 557688 675300 557716
rect 673328 557676 673334 557688
rect 675294 557676 675300 557688
rect 675352 557676 675358 557728
rect 43254 557540 43260 557592
rect 43312 557580 43318 557592
rect 51902 557580 51908 557592
rect 43312 557552 51908 557580
rect 43312 557540 43318 557552
rect 51902 557540 51908 557552
rect 51960 557540 51966 557592
rect 54846 557540 54852 557592
rect 54904 557580 54910 557592
rect 62114 557580 62120 557592
rect 54904 557552 62120 557580
rect 54904 557540 54910 557552
rect 62114 557540 62120 557552
rect 62172 557540 62178 557592
rect 666370 557540 666376 557592
rect 666428 557580 666434 557592
rect 675294 557580 675300 557592
rect 666428 557552 675300 557580
rect 666428 557540 666434 557552
rect 675294 557540 675300 557552
rect 675352 557540 675358 557592
rect 40862 554888 40868 554940
rect 40920 554928 40926 554940
rect 41690 554928 41696 554940
rect 40920 554900 41696 554928
rect 40920 554888 40926 554900
rect 41690 554888 41696 554900
rect 41748 554888 41754 554940
rect 42058 554888 42064 554940
rect 42116 554928 42122 554940
rect 42794 554928 42800 554940
rect 42116 554900 42800 554928
rect 42116 554888 42122 554900
rect 42794 554888 42800 554900
rect 42852 554888 42858 554940
rect 40586 554752 40592 554804
rect 40644 554792 40650 554804
rect 41690 554792 41696 554804
rect 40644 554764 41696 554792
rect 40644 554752 40650 554764
rect 41690 554752 41696 554764
rect 41748 554752 41754 554804
rect 42058 554752 42064 554804
rect 42116 554792 42122 554804
rect 44358 554792 44364 554804
rect 42116 554764 44364 554792
rect 42116 554752 42122 554764
rect 44358 554752 44364 554764
rect 44416 554752 44422 554804
rect 671798 554752 671804 554804
rect 671856 554792 671862 554804
rect 675110 554792 675116 554804
rect 671856 554764 675116 554792
rect 671856 554752 671862 554764
rect 675110 554752 675116 554764
rect 675168 554752 675174 554804
rect 673454 554140 673460 554192
rect 673512 554180 673518 554192
rect 675110 554180 675116 554192
rect 673512 554152 675116 554180
rect 673512 554140 673518 554152
rect 675110 554140 675116 554152
rect 675168 554140 675174 554192
rect 658918 554004 658924 554056
rect 658976 554044 658982 554056
rect 675110 554044 675116 554056
rect 658976 554016 675116 554044
rect 658976 554004 658982 554016
rect 675110 554004 675116 554016
rect 675168 554004 675174 554056
rect 42058 550672 42064 550724
rect 42116 550712 42122 550724
rect 43162 550712 43168 550724
rect 42116 550684 43168 550712
rect 42116 550672 42122 550684
rect 43162 550672 43168 550684
rect 43220 550672 43226 550724
rect 651558 550604 651564 550656
rect 651616 550644 651622 550656
rect 658918 550644 658924 550656
rect 651616 550616 658924 550644
rect 651616 550604 651622 550616
rect 658918 550604 658924 550616
rect 658976 550604 658982 550656
rect 40034 550400 40040 550452
rect 40092 550440 40098 550452
rect 41690 550440 41696 550452
rect 40092 550412 41696 550440
rect 40092 550400 40098 550412
rect 41690 550400 41696 550412
rect 41748 550400 41754 550452
rect 42058 550332 42064 550384
rect 42116 550372 42122 550384
rect 42518 550372 42524 550384
rect 42116 550344 42524 550372
rect 42116 550332 42122 550344
rect 42518 550332 42524 550344
rect 42576 550332 42582 550384
rect 674466 549720 674472 549772
rect 674524 549760 674530 549772
rect 675294 549760 675300 549772
rect 674524 549732 675300 549760
rect 674524 549720 674530 549732
rect 675294 549720 675300 549732
rect 675352 549720 675358 549772
rect 41138 548088 41144 548140
rect 41196 548128 41202 548140
rect 41690 548128 41696 548140
rect 41196 548100 41696 548128
rect 41196 548088 41202 548100
rect 41690 548088 41696 548100
rect 41748 548088 41754 548140
rect 43438 547884 43444 547936
rect 43496 547924 43502 547936
rect 56042 547924 56048 547936
rect 43496 547896 56048 547924
rect 43496 547884 43502 547896
rect 56042 547884 56048 547896
rect 56100 547884 56106 547936
rect 31754 547408 31760 547460
rect 31812 547448 31818 547460
rect 38470 547448 38476 547460
rect 31812 547420 38476 547448
rect 31812 547408 31818 547420
rect 38470 547408 38476 547420
rect 38528 547408 38534 547460
rect 675938 546796 675944 546848
rect 675996 546836 676002 546848
rect 680998 546836 681004 546848
rect 675996 546808 681004 546836
rect 675996 546796 676002 546808
rect 680998 546796 681004 546808
rect 681056 546796 681062 546848
rect 43438 546524 43444 546576
rect 43496 546564 43502 546576
rect 49142 546564 49148 546576
rect 43496 546536 49148 546564
rect 43496 546524 43502 546536
rect 49142 546524 49148 546536
rect 49200 546524 49206 546576
rect 676122 545708 676128 545760
rect 676180 545748 676186 545760
rect 683206 545748 683212 545760
rect 676180 545720 683212 545748
rect 676180 545708 676186 545720
rect 683206 545708 683212 545720
rect 683264 545708 683270 545760
rect 674466 545436 674472 545488
rect 674524 545476 674530 545488
rect 675018 545476 675024 545488
rect 674524 545448 675024 545476
rect 674524 545436 674530 545448
rect 675018 545436 675024 545448
rect 675076 545436 675082 545488
rect 43438 545096 43444 545148
rect 43496 545136 43502 545148
rect 62114 545136 62120 545148
rect 43496 545108 62120 545136
rect 43496 545096 43502 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 34422 544348 34428 544400
rect 34480 544388 34486 544400
rect 39482 544388 39488 544400
rect 34480 544360 39488 544388
rect 34480 544348 34486 544360
rect 39482 544348 39488 544360
rect 39540 544348 39546 544400
rect 38470 542172 38476 542224
rect 38528 542212 38534 542224
rect 39758 542212 39764 542224
rect 38528 542184 39764 542212
rect 38528 542172 38534 542184
rect 39758 542172 39764 542184
rect 39816 542172 39822 542224
rect 42702 540676 42708 540728
rect 42760 540716 42766 540728
rect 43622 540716 43628 540728
rect 42760 540688 43628 540716
rect 42760 540676 42766 540688
rect 43622 540676 43628 540688
rect 43680 540676 43686 540728
rect 42426 537616 42432 537668
rect 42484 537656 42490 537668
rect 44082 537656 44088 537668
rect 42484 537628 44088 537656
rect 42484 537616 42490 537628
rect 44082 537616 44088 537628
rect 44140 537616 44146 537668
rect 651558 536800 651564 536852
rect 651616 536840 651622 536852
rect 663058 536840 663064 536852
rect 651616 536812 663064 536840
rect 651616 536800 651622 536812
rect 663058 536800 663064 536812
rect 663116 536800 663122 536852
rect 42702 536596 42708 536648
rect 42760 536636 42766 536648
rect 45370 536636 45376 536648
rect 42760 536608 45376 536636
rect 42760 536596 42766 536608
rect 45370 536596 45376 536608
rect 45428 536596 45434 536648
rect 675478 535684 675484 535696
rect 663766 535656 675484 535684
rect 663242 535576 663248 535628
rect 663300 535616 663306 535628
rect 663766 535616 663794 535656
rect 675478 535644 675484 535656
rect 675536 535644 675542 535696
rect 663300 535588 663794 535616
rect 663300 535576 663306 535588
rect 661678 535440 661684 535492
rect 661736 535480 661742 535492
rect 675478 535480 675484 535492
rect 661736 535452 675484 535480
rect 661736 535440 661742 535452
rect 675478 535440 675484 535452
rect 675536 535440 675542 535492
rect 42334 535236 42340 535288
rect 42392 535276 42398 535288
rect 43898 535276 43904 535288
rect 42392 535248 43904 535276
rect 42392 535236 42398 535248
rect 43898 535236 43904 535248
rect 43956 535236 43962 535288
rect 673086 534556 673092 534608
rect 673144 534596 673150 534608
rect 674926 534596 674932 534608
rect 673144 534568 674932 534596
rect 673144 534556 673150 534568
rect 674926 534556 674932 534568
rect 674984 534556 674990 534608
rect 675478 534460 675484 534472
rect 673564 534432 675484 534460
rect 672902 534352 672908 534404
rect 672960 534392 672966 534404
rect 673564 534392 673592 534432
rect 675478 534420 675484 534432
rect 675536 534420 675542 534472
rect 672960 534364 673592 534392
rect 672960 534352 672966 534364
rect 661862 534216 661868 534268
rect 661920 534256 661926 534268
rect 674466 534256 674472 534268
rect 661920 534228 674472 534256
rect 661920 534216 661926 534228
rect 674466 534216 674472 534228
rect 674524 534216 674530 534268
rect 672994 534080 673000 534132
rect 673052 534120 673058 534132
rect 675478 534120 675484 534132
rect 673052 534092 675484 534120
rect 673052 534080 673058 534092
rect 675478 534080 675484 534092
rect 675536 534080 675542 534132
rect 42426 533400 42432 533452
rect 42484 533440 42490 533452
rect 43070 533440 43076 533452
rect 42484 533412 43076 533440
rect 42484 533400 42490 533412
rect 43070 533400 43076 533412
rect 43128 533400 43134 533452
rect 671522 533332 671528 533384
rect 671580 533372 671586 533384
rect 675478 533372 675484 533384
rect 671580 533344 675484 533372
rect 671580 533332 671586 533344
rect 675478 533332 675484 533344
rect 675536 533332 675542 533384
rect 672534 532720 672540 532772
rect 672592 532760 672598 532772
rect 675478 532760 675484 532772
rect 672592 532732 675484 532760
rect 672592 532720 672598 532732
rect 675478 532720 675484 532732
rect 675536 532720 675542 532772
rect 42702 532652 42708 532704
rect 42760 532692 42766 532704
rect 45186 532692 45192 532704
rect 42760 532664 45192 532692
rect 42760 532652 42766 532664
rect 45186 532652 45192 532664
rect 45244 532652 45250 532704
rect 671154 532516 671160 532568
rect 671212 532556 671218 532568
rect 675478 532556 675484 532568
rect 671212 532528 675484 532556
rect 671212 532516 671218 532528
rect 675478 532516 675484 532528
rect 675536 532516 675542 532568
rect 663518 531428 663524 531480
rect 663576 531468 663582 531480
rect 663576 531440 663794 531468
rect 663576 531428 663582 531440
rect 663766 531400 663794 531440
rect 675478 531400 675484 531412
rect 663766 531372 675484 531400
rect 675478 531360 675484 531372
rect 675536 531360 675542 531412
rect 667842 530068 667848 530120
rect 667900 530108 667906 530120
rect 675478 530108 675484 530120
rect 667900 530080 675484 530108
rect 667900 530068 667906 530080
rect 675478 530068 675484 530080
rect 675536 530068 675542 530120
rect 669038 529932 669044 529984
rect 669096 529972 669102 529984
rect 674926 529972 674932 529984
rect 669096 529944 674932 529972
rect 669096 529932 669102 529944
rect 674926 529932 674932 529944
rect 674984 529932 674990 529984
rect 42518 529048 42524 529100
rect 42576 529088 42582 529100
rect 43254 529088 43260 529100
rect 42576 529060 43260 529088
rect 42576 529048 42582 529060
rect 43254 529048 43260 529060
rect 43312 529048 43318 529100
rect 666094 528572 666100 528624
rect 666152 528612 666158 528624
rect 675478 528612 675484 528624
rect 666152 528584 675484 528612
rect 666152 528572 666158 528584
rect 675478 528572 675484 528584
rect 675536 528572 675542 528624
rect 673638 528436 673644 528488
rect 673696 528476 673702 528488
rect 675478 528476 675484 528488
rect 673696 528448 675484 528476
rect 673696 528436 673702 528448
rect 675478 528436 675484 528448
rect 675536 528436 675542 528488
rect 673822 528028 673828 528080
rect 673880 528068 673886 528080
rect 675478 528068 675484 528080
rect 673880 528040 675484 528068
rect 673880 528028 673886 528040
rect 675478 528028 675484 528040
rect 675536 528028 675542 528080
rect 670418 526804 670424 526856
rect 670476 526844 670482 526856
rect 675478 526844 675484 526856
rect 670476 526816 675484 526844
rect 670476 526804 670482 526816
rect 675478 526804 675484 526816
rect 675536 526804 675542 526856
rect 672718 526396 672724 526448
rect 672776 526436 672782 526448
rect 675478 526436 675484 526448
rect 672776 526408 675484 526436
rect 672776 526396 672782 526408
rect 675478 526396 675484 526408
rect 675536 526396 675542 526448
rect 673730 525784 673736 525836
rect 673788 525824 673794 525836
rect 675478 525824 675484 525836
rect 673788 525796 675484 525824
rect 673788 525784 673794 525796
rect 675478 525784 675484 525796
rect 675536 525784 675542 525836
rect 680998 525716 681004 525768
rect 681056 525756 681062 525768
rect 683114 525756 683120 525768
rect 681056 525728 683120 525756
rect 681056 525716 681062 525728
rect 683114 525716 683120 525728
rect 683172 525716 683178 525768
rect 43254 523676 43260 523728
rect 43312 523716 43318 523728
rect 62758 523716 62764 523728
rect 43312 523688 62764 523716
rect 43312 523676 43318 523688
rect 62758 523676 62764 523688
rect 62816 523676 62822 523728
rect 651558 522996 651564 523048
rect 651616 523036 651622 523048
rect 661678 523036 661684 523048
rect 651616 523008 661684 523036
rect 651616 522996 651622 523008
rect 661678 522996 661684 523008
rect 661736 522996 661742 523048
rect 42058 518916 42064 518968
rect 42116 518956 42122 518968
rect 62114 518956 62120 518968
rect 42116 518928 62120 518956
rect 42116 518916 42122 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 651558 510620 651564 510672
rect 651616 510660 651622 510672
rect 660482 510660 660488 510672
rect 651616 510632 660488 510660
rect 651616 510620 651622 510632
rect 660482 510620 660488 510632
rect 660540 510620 660546 510672
rect 52086 506472 52092 506524
rect 52144 506512 52150 506524
rect 62114 506512 62120 506524
rect 52144 506484 62120 506512
rect 52144 506472 52150 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 676030 503480 676036 503532
rect 676088 503520 676094 503532
rect 679618 503520 679624 503532
rect 676088 503492 679624 503520
rect 676088 503480 676094 503492
rect 679618 503480 679624 503492
rect 679676 503480 679682 503532
rect 676030 498244 676036 498296
rect 676088 498284 676094 498296
rect 679802 498284 679808 498296
rect 676088 498256 679808 498284
rect 676088 498244 676094 498256
rect 679802 498244 679808 498256
rect 679860 498244 679866 498296
rect 651558 496816 651564 496868
rect 651616 496856 651622 496868
rect 659102 496856 659108 496868
rect 651616 496828 659108 496856
rect 651616 496816 651622 496828
rect 659102 496816 659108 496828
rect 659160 496816 659166 496868
rect 43622 491920 43628 491972
rect 43680 491960 43686 491972
rect 62114 491960 62120 491972
rect 43680 491932 62120 491960
rect 43680 491920 43686 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 664438 491580 664444 491632
rect 664496 491620 664502 491632
rect 675294 491620 675300 491632
rect 664496 491592 675300 491620
rect 664496 491580 664502 491592
rect 675294 491580 675300 491592
rect 675352 491580 675358 491632
rect 660298 491444 660304 491496
rect 660356 491484 660362 491496
rect 675478 491484 675484 491496
rect 660356 491456 675484 491484
rect 660356 491444 660362 491456
rect 675478 491444 675484 491456
rect 675536 491444 675542 491496
rect 659286 491308 659292 491360
rect 659344 491348 659350 491360
rect 675478 491348 675484 491360
rect 659344 491320 675484 491348
rect 659344 491308 659350 491320
rect 675478 491308 675484 491320
rect 675536 491308 675542 491360
rect 676214 490152 676220 490204
rect 676272 490192 676278 490204
rect 677410 490192 677416 490204
rect 676272 490164 677416 490192
rect 676272 490152 676278 490164
rect 677410 490152 677416 490164
rect 677468 490152 677474 490204
rect 672994 490016 673000 490068
rect 673052 490056 673058 490068
rect 675478 490056 675484 490068
rect 673052 490028 675484 490056
rect 673052 490016 673058 490028
rect 675478 490016 675484 490028
rect 675536 490016 675542 490068
rect 672534 488656 672540 488708
rect 672592 488696 672598 488708
rect 675478 488696 675484 488708
rect 672592 488668 675484 488696
rect 672592 488656 672598 488668
rect 675478 488656 675484 488668
rect 675536 488656 675542 488708
rect 676214 488520 676220 488572
rect 676272 488560 676278 488572
rect 677226 488560 677232 488572
rect 676272 488532 677232 488560
rect 676272 488520 676278 488532
rect 677226 488520 677232 488532
rect 677284 488520 677290 488572
rect 666370 485936 666376 485988
rect 666428 485976 666434 485988
rect 675478 485976 675484 485988
rect 666428 485948 675484 485976
rect 666428 485936 666434 485948
rect 675478 485936 675484 485948
rect 675536 485936 675542 485988
rect 663702 485800 663708 485852
rect 663760 485840 663766 485852
rect 675294 485840 675300 485852
rect 663760 485812 675300 485840
rect 663760 485800 663766 485812
rect 675294 485800 675300 485812
rect 675352 485800 675358 485852
rect 670234 485596 670240 485648
rect 670292 485636 670298 485648
rect 675478 485636 675484 485648
rect 670292 485608 675484 485636
rect 670292 485596 670298 485608
rect 675478 485596 675484 485608
rect 675536 485596 675542 485648
rect 651558 484440 651564 484492
rect 651616 484480 651622 484492
rect 651616 484452 654134 484480
rect 651616 484440 651622 484452
rect 654106 484412 654134 484452
rect 664806 484412 664812 484424
rect 654106 484384 664812 484412
rect 664806 484372 664812 484384
rect 664864 484372 664870 484424
rect 664990 484372 664996 484424
rect 665048 484412 665054 484424
rect 675478 484412 675484 484424
rect 665048 484384 675484 484412
rect 665048 484372 665054 484384
rect 675478 484372 675484 484384
rect 675536 484372 675542 484424
rect 673454 483556 673460 483608
rect 673512 483596 673518 483608
rect 675478 483596 675484 483608
rect 673512 483568 675484 483596
rect 673512 483556 673518 483568
rect 675478 483556 675484 483568
rect 675536 483556 675542 483608
rect 673270 483148 673276 483200
rect 673328 483188 673334 483200
rect 675478 483188 675484 483200
rect 673328 483160 675484 483188
rect 673328 483148 673334 483160
rect 675478 483148 675484 483160
rect 675536 483148 675542 483200
rect 671798 482740 671804 482792
rect 671856 482780 671862 482792
rect 675478 482780 675484 482792
rect 671856 482752 675484 482780
rect 671856 482740 671862 482752
rect 675478 482740 675484 482752
rect 675536 482740 675542 482792
rect 671982 482332 671988 482384
rect 672040 482372 672046 482384
rect 675478 482372 675484 482384
rect 672040 482344 675484 482372
rect 672040 482332 672046 482344
rect 675478 482332 675484 482344
rect 675536 482332 675542 482384
rect 674098 481856 674104 481908
rect 674156 481896 674162 481908
rect 675478 481896 675484 481908
rect 674156 481868 675484 481896
rect 674156 481856 674162 481868
rect 675478 481856 675484 481868
rect 675536 481856 675542 481908
rect 671522 480632 671528 480684
rect 671580 480672 671586 480684
rect 675478 480672 675484 480684
rect 671580 480644 675484 480672
rect 671580 480632 671586 480644
rect 675478 480632 675484 480644
rect 675536 480632 675542 480684
rect 47946 480224 47952 480276
rect 48004 480264 48010 480276
rect 62114 480264 62120 480276
rect 48004 480236 62120 480264
rect 48004 480224 48010 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 651558 470568 651564 470620
rect 651616 470608 651622 470620
rect 661862 470608 661868 470620
rect 651616 470580 661868 470608
rect 651616 470568 651622 470580
rect 661862 470568 661868 470580
rect 661920 470568 661926 470620
rect 49326 466420 49332 466472
rect 49384 466460 49390 466472
rect 62114 466460 62120 466472
rect 49384 466432 62120 466460
rect 49384 466420 49390 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 651558 456764 651564 456816
rect 651616 456804 651622 456816
rect 663242 456804 663248 456816
rect 651616 456776 663248 456804
rect 651616 456764 651622 456776
rect 663242 456764 663248 456776
rect 663300 456764 663306 456816
rect 55030 454044 55036 454096
rect 55088 454084 55094 454096
rect 62114 454084 62120 454096
rect 55088 454056 62120 454084
rect 55088 454044 55094 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 651558 444456 651564 444508
rect 651616 444496 651622 444508
rect 651616 444468 654134 444496
rect 651616 444456 651622 444468
rect 654106 444428 654134 444468
rect 660666 444428 660672 444440
rect 654106 444400 660672 444428
rect 660666 444388 660672 444400
rect 660724 444388 660730 444440
rect 50706 440240 50712 440292
rect 50764 440280 50770 440292
rect 62114 440280 62120 440292
rect 50764 440252 62120 440280
rect 50764 440240 50770 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 651558 430584 651564 430636
rect 651616 430624 651622 430636
rect 660298 430624 660304 430636
rect 651616 430596 660304 430624
rect 651616 430584 651622 430596
rect 660298 430584 660304 430596
rect 660356 430584 660362 430636
rect 41322 429564 41328 429616
rect 41380 429604 41386 429616
rect 41690 429604 41696 429616
rect 41380 429576 41696 429604
rect 41380 429564 41386 429576
rect 41690 429564 41696 429576
rect 41748 429564 41754 429616
rect 41322 429428 41328 429480
rect 41380 429468 41386 429480
rect 41690 429468 41696 429480
rect 41380 429440 41696 429468
rect 41380 429428 41386 429440
rect 41690 429428 41696 429440
rect 41748 429428 41754 429480
rect 42058 429428 42064 429480
rect 42116 429468 42122 429480
rect 43254 429468 43260 429480
rect 42116 429440 43260 429468
rect 42116 429428 42122 429440
rect 43254 429428 43260 429440
rect 43312 429428 43318 429480
rect 41138 429292 41144 429344
rect 41196 429332 41202 429344
rect 41690 429332 41696 429344
rect 41196 429304 41696 429332
rect 41196 429292 41202 429304
rect 41690 429292 41696 429304
rect 41748 429292 41754 429344
rect 42058 429292 42064 429344
rect 42116 429332 42122 429344
rect 43438 429332 43444 429344
rect 42116 429304 43444 429332
rect 42116 429292 42122 429304
rect 43438 429292 43444 429304
rect 43496 429292 43502 429344
rect 40954 429156 40960 429208
rect 41012 429196 41018 429208
rect 41690 429196 41696 429208
rect 41012 429168 41696 429196
rect 41012 429156 41018 429168
rect 41690 429156 41696 429168
rect 41748 429156 41754 429208
rect 42058 429156 42064 429208
rect 42116 429196 42122 429208
rect 44542 429196 44548 429208
rect 42116 429168 44548 429196
rect 42116 429156 42122 429168
rect 44542 429156 44548 429168
rect 44600 429156 44606 429208
rect 42058 428408 42064 428460
rect 42116 428448 42122 428460
rect 42886 428448 42892 428460
rect 42116 428420 42892 428448
rect 42116 428408 42122 428420
rect 42886 428408 42892 428420
rect 42944 428408 42950 428460
rect 41690 428040 41696 428052
rect 41386 428012 41696 428040
rect 41386 427984 41414 428012
rect 41690 428000 41696 428012
rect 41748 428000 41754 428052
rect 41322 427932 41328 427984
rect 41380 427944 41414 427984
rect 41380 427932 41386 427944
rect 41138 427796 41144 427848
rect 41196 427836 41202 427848
rect 41690 427836 41696 427848
rect 41196 427808 41696 427836
rect 41196 427796 41202 427808
rect 41690 427796 41696 427808
rect 41748 427796 41754 427848
rect 42058 427796 42064 427848
rect 42116 427836 42122 427848
rect 44266 427836 44272 427848
rect 42116 427808 44272 427836
rect 42116 427796 42122 427808
rect 44266 427796 44272 427808
rect 44324 427796 44330 427848
rect 46566 427796 46572 427848
rect 46624 427836 46630 427848
rect 62114 427836 62120 427848
rect 46624 427808 62120 427836
rect 46624 427796 46630 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 41690 426680 41696 426692
rect 41386 426652 41696 426680
rect 41138 426572 41144 426624
rect 41196 426612 41202 426624
rect 41386 426612 41414 426652
rect 41690 426640 41696 426652
rect 41748 426640 41754 426692
rect 42058 426640 42064 426692
rect 42116 426680 42122 426692
rect 43806 426680 43812 426692
rect 42116 426652 43812 426680
rect 42116 426640 42122 426652
rect 43806 426640 43812 426652
rect 43864 426640 43870 426692
rect 41196 426584 41414 426612
rect 41196 426572 41202 426584
rect 40954 426436 40960 426488
rect 41012 426476 41018 426488
rect 41690 426476 41696 426488
rect 41012 426448 41696 426476
rect 41012 426436 41018 426448
rect 41690 426436 41696 426448
rect 41748 426436 41754 426488
rect 42058 426436 42064 426488
rect 42116 426476 42122 426488
rect 44266 426476 44272 426488
rect 42116 426448 44272 426476
rect 42116 426436 42122 426448
rect 44266 426436 44272 426448
rect 44324 426436 44330 426488
rect 41322 424328 41328 424380
rect 41380 424368 41386 424380
rect 41690 424368 41696 424380
rect 41380 424340 41696 424368
rect 41380 424328 41386 424340
rect 41690 424328 41696 424340
rect 41748 424328 41754 424380
rect 42426 419500 42432 419552
rect 42484 419540 42490 419552
rect 51902 419540 51908 419552
rect 42484 419512 51908 419540
rect 42484 419500 42490 419512
rect 51902 419500 51908 419512
rect 51960 419500 51966 419552
rect 45738 418140 45744 418192
rect 45796 418180 45802 418192
rect 54662 418180 54668 418192
rect 45796 418152 54668 418180
rect 45796 418140 45802 418152
rect 54662 418140 54668 418152
rect 54720 418140 54726 418192
rect 651558 416780 651564 416832
rect 651616 416820 651622 416832
rect 664438 416820 664444 416832
rect 651616 416792 664444 416820
rect 651616 416780 651622 416792
rect 664438 416780 664444 416792
rect 664496 416780 664502 416832
rect 56226 415420 56232 415472
rect 56284 415460 56290 415472
rect 62114 415460 62120 415472
rect 56284 415432 62120 415460
rect 56284 415420 56290 415432
rect 62114 415420 62120 415432
rect 62172 415420 62178 415472
rect 42242 409776 42248 409828
rect 42300 409816 42306 409828
rect 43438 409816 43444 409828
rect 42300 409788 43444 409816
rect 42300 409776 42306 409788
rect 43438 409776 43444 409788
rect 43496 409776 43502 409828
rect 42426 408416 42432 408468
rect 42484 408456 42490 408468
rect 54846 408456 54852 408468
rect 42484 408428 54852 408456
rect 42484 408416 42490 408428
rect 54846 408416 54852 408428
rect 54904 408416 54910 408468
rect 42426 408280 42432 408332
rect 42484 408320 42490 408332
rect 45370 408320 45376 408332
rect 42484 408292 45376 408320
rect 42484 408280 42490 408292
rect 45370 408280 45376 408292
rect 45428 408280 45434 408332
rect 42426 407056 42432 407108
rect 42484 407096 42490 407108
rect 43070 407096 43076 407108
rect 42484 407068 43076 407096
rect 42484 407056 42490 407068
rect 43070 407056 43076 407068
rect 43128 407056 43134 407108
rect 42334 405968 42340 406020
rect 42392 406008 42398 406020
rect 45554 406008 45560 406020
rect 42392 405980 45560 406008
rect 42392 405968 42398 405980
rect 45554 405968 45560 405980
rect 45612 405968 45618 406020
rect 651558 404336 651564 404388
rect 651616 404376 651622 404388
rect 659286 404376 659292 404388
rect 651616 404348 659292 404376
rect 651616 404336 651622 404348
rect 659286 404336 659292 404348
rect 659344 404336 659350 404388
rect 669314 403384 669320 403436
rect 669372 403424 669378 403436
rect 675294 403424 675300 403436
rect 669372 403396 675300 403424
rect 669372 403384 669378 403396
rect 675294 403384 675300 403396
rect 675352 403384 675358 403436
rect 663058 403248 663064 403300
rect 663116 403288 663122 403300
rect 675478 403288 675484 403300
rect 663116 403260 675484 403288
rect 663116 403248 663122 403260
rect 675478 403248 675484 403260
rect 675536 403248 675542 403300
rect 661678 403112 661684 403164
rect 661736 403152 661742 403164
rect 661736 403124 669452 403152
rect 661736 403112 661742 403124
rect 669424 403084 669452 403124
rect 675478 403084 675484 403096
rect 669424 403056 675484 403084
rect 675478 403044 675484 403056
rect 675536 403044 675542 403096
rect 658918 402976 658924 403028
rect 658976 403016 658982 403028
rect 658976 402988 669314 403016
rect 658976 402976 658982 402988
rect 669286 402960 669314 402988
rect 42242 402908 42248 402960
rect 42300 402948 42306 402960
rect 43806 402948 43812 402960
rect 42300 402920 43812 402948
rect 42300 402908 42306 402920
rect 43806 402908 43812 402920
rect 43864 402908 43870 402960
rect 669286 402920 669320 402960
rect 669314 402908 669320 402920
rect 669372 402908 669378 402960
rect 42426 402500 42432 402552
rect 42484 402540 42490 402552
rect 45186 402540 45192 402552
rect 42484 402512 45192 402540
rect 42484 402500 42490 402512
rect 45186 402500 45192 402512
rect 45244 402500 45250 402552
rect 43438 401616 43444 401668
rect 43496 401656 43502 401668
rect 62114 401656 62120 401668
rect 43496 401628 62120 401656
rect 43496 401616 43502 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 672810 400528 672816 400580
rect 672868 400568 672874 400580
rect 675478 400568 675484 400580
rect 672868 400540 675484 400568
rect 672868 400528 672874 400540
rect 675478 400528 675484 400540
rect 675536 400528 675542 400580
rect 42426 400120 42432 400172
rect 42484 400160 42490 400172
rect 43990 400160 43996 400172
rect 42484 400132 43996 400160
rect 42484 400120 42490 400132
rect 43990 400120 43996 400132
rect 44048 400120 44054 400172
rect 673178 399712 673184 399764
rect 673236 399752 673242 399764
rect 675478 399752 675484 399764
rect 673236 399724 675484 399752
rect 673236 399712 673242 399724
rect 675478 399712 675484 399724
rect 675536 399712 675542 399764
rect 671154 397264 671160 397316
rect 671212 397304 671218 397316
rect 675478 397304 675484 397316
rect 671212 397276 675484 397304
rect 671212 397264 671218 397276
rect 675478 397264 675484 397276
rect 675536 397264 675542 397316
rect 670418 396040 670424 396092
rect 670476 396080 670482 396092
rect 675478 396080 675484 396092
rect 670476 396052 675484 396080
rect 670476 396040 670482 396052
rect 675478 396040 675484 396052
rect 675536 396040 675542 396092
rect 673914 395632 673920 395684
rect 673972 395672 673978 395684
rect 675478 395672 675484 395684
rect 673972 395644 675484 395672
rect 673972 395632 673978 395644
rect 675478 395632 675484 395644
rect 675536 395632 675542 395684
rect 673362 394408 673368 394460
rect 673420 394448 673426 394460
rect 675478 394448 675484 394460
rect 673420 394420 675484 394448
rect 673420 394408 673426 394420
rect 675478 394408 675484 394420
rect 675536 394408 675542 394460
rect 672534 394136 672540 394188
rect 672592 394176 672598 394188
rect 672902 394176 672908 394188
rect 672592 394148 672908 394176
rect 672592 394136 672598 394148
rect 672902 394136 672908 394148
rect 672960 394136 672966 394188
rect 672994 394000 673000 394052
rect 673052 394040 673058 394052
rect 675478 394040 675484 394052
rect 673052 394012 675484 394040
rect 673052 394000 673058 394012
rect 675478 394000 675484 394012
rect 675536 394000 675542 394052
rect 671614 392368 671620 392420
rect 671672 392408 671678 392420
rect 675478 392408 675484 392420
rect 671672 392380 675484 392408
rect 671672 392368 671678 392380
rect 675478 392368 675484 392380
rect 675536 392368 675542 392420
rect 675846 392096 675852 392148
rect 675904 392136 675910 392148
rect 683114 392136 683120 392148
rect 675904 392108 683120 392136
rect 675904 392096 675910 392108
rect 683114 392096 683120 392108
rect 683172 392096 683178 392148
rect 651558 390532 651564 390584
rect 651616 390572 651622 390584
rect 661678 390572 661684 390584
rect 651616 390544 661684 390572
rect 651616 390532 651622 390544
rect 661678 390532 661684 390544
rect 661736 390532 661742 390584
rect 48130 389240 48136 389292
rect 48188 389280 48194 389292
rect 62114 389280 62120 389292
rect 48188 389252 62120 389280
rect 48188 389240 48194 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 35802 387540 35808 387592
rect 35860 387580 35866 387592
rect 41690 387580 41696 387592
rect 35860 387552 41696 387580
rect 35860 387540 35866 387552
rect 41690 387540 41696 387552
rect 41748 387540 41754 387592
rect 42058 387472 42064 387524
rect 42116 387512 42122 387524
rect 49326 387512 49332 387524
rect 42116 387484 49332 387512
rect 42116 387472 42122 387484
rect 49326 387472 49332 387484
rect 49384 387472 49390 387524
rect 35618 386792 35624 386844
rect 35676 386832 35682 386844
rect 39942 386832 39948 386844
rect 35676 386804 39948 386832
rect 35676 386792 35682 386804
rect 39942 386792 39948 386804
rect 40000 386792 40006 386844
rect 40126 386696 40132 386708
rect 38626 386668 40132 386696
rect 38626 386628 38654 386668
rect 40126 386656 40132 386668
rect 40184 386656 40190 386708
rect 36004 386600 38654 386628
rect 35802 386520 35808 386572
rect 35860 386560 35866 386572
rect 36004 386560 36032 386600
rect 35860 386532 36032 386560
rect 35860 386520 35866 386532
rect 41690 386492 41696 386504
rect 40696 386464 41696 386492
rect 35434 386384 35440 386436
rect 35492 386424 35498 386436
rect 40696 386424 40724 386464
rect 41690 386452 41696 386464
rect 41748 386452 41754 386504
rect 42058 386452 42064 386504
rect 42116 386492 42122 386504
rect 47946 386492 47952 386504
rect 42116 386464 47952 386492
rect 42116 386452 42122 386464
rect 47946 386452 47952 386464
rect 48004 386452 48010 386504
rect 35492 386396 40724 386424
rect 35492 386384 35498 386396
rect 35802 385432 35808 385484
rect 35860 385472 35866 385484
rect 40126 385472 40132 385484
rect 35860 385444 40132 385472
rect 35860 385432 35866 385444
rect 40126 385432 40132 385444
rect 40184 385432 40190 385484
rect 41690 385268 41696 385280
rect 41386 385240 41696 385268
rect 35526 385160 35532 385212
rect 35584 385200 35590 385212
rect 41386 385200 41414 385240
rect 41690 385228 41696 385240
rect 41748 385228 41754 385280
rect 42058 385228 42064 385280
rect 42116 385268 42122 385280
rect 42886 385268 42892 385280
rect 42116 385240 42892 385268
rect 42116 385228 42122 385240
rect 42886 385228 42892 385240
rect 42944 385228 42950 385280
rect 35584 385172 41414 385200
rect 35584 385160 35590 385172
rect 35342 385024 35348 385076
rect 35400 385064 35406 385076
rect 41690 385064 41696 385076
rect 35400 385036 41696 385064
rect 35400 385024 35406 385036
rect 41690 385024 41696 385036
rect 41748 385024 41754 385076
rect 42058 385024 42064 385076
rect 42116 385064 42122 385076
rect 45370 385064 45376 385076
rect 42116 385036 45376 385064
rect 42116 385024 42122 385036
rect 45370 385024 45376 385036
rect 45428 385024 45434 385076
rect 674926 384752 674932 384804
rect 674984 384792 674990 384804
rect 675478 384792 675484 384804
rect 674984 384764 675484 384792
rect 674984 384752 674990 384764
rect 675478 384752 675484 384764
rect 675536 384752 675542 384804
rect 35802 384072 35808 384124
rect 35860 384112 35866 384124
rect 39758 384112 39764 384124
rect 35860 384084 39764 384112
rect 35860 384072 35866 384084
rect 39758 384072 39764 384084
rect 39816 384072 39822 384124
rect 39942 383908 39948 383920
rect 36004 383880 39948 383908
rect 35618 383800 35624 383852
rect 35676 383840 35682 383852
rect 36004 383840 36032 383880
rect 39942 383868 39948 383880
rect 40000 383868 40006 383920
rect 35676 383812 36032 383840
rect 35676 383800 35682 383812
rect 42058 383732 42064 383784
rect 42116 383772 42122 383784
rect 44542 383772 44548 383784
rect 42116 383744 44548 383772
rect 42116 383732 42122 383744
rect 44542 383732 44548 383744
rect 44600 383732 44606 383784
rect 35802 383664 35808 383716
rect 35860 383704 35866 383716
rect 41690 383704 41696 383716
rect 35860 383676 41696 383704
rect 35860 383664 35866 383676
rect 41690 383664 41696 383676
rect 41748 383664 41754 383716
rect 35802 382644 35808 382696
rect 35860 382684 35866 382696
rect 41690 382684 41696 382696
rect 35860 382656 41696 382684
rect 35860 382644 35866 382656
rect 41690 382644 41696 382656
rect 41748 382644 41754 382696
rect 35618 382508 35624 382560
rect 35676 382548 35682 382560
rect 40218 382548 40224 382560
rect 35676 382520 40224 382548
rect 35676 382508 35682 382520
rect 40218 382508 40224 382520
rect 40276 382508 40282 382560
rect 35434 382372 35440 382424
rect 35492 382412 35498 382424
rect 40034 382412 40040 382424
rect 35492 382384 40040 382412
rect 35492 382372 35498 382384
rect 40034 382372 40040 382384
rect 40092 382372 40098 382424
rect 35250 382236 35256 382288
rect 35308 382276 35314 382288
rect 39022 382276 39028 382288
rect 35308 382248 39028 382276
rect 35308 382236 35314 382248
rect 39022 382236 39028 382248
rect 39080 382236 39086 382288
rect 35802 381148 35808 381200
rect 35860 381188 35866 381200
rect 41414 381188 41420 381200
rect 35860 381160 41420 381188
rect 35860 381148 35866 381160
rect 41414 381148 41420 381160
rect 41472 381148 41478 381200
rect 35618 381012 35624 381064
rect 35676 381052 35682 381064
rect 40034 381052 40040 381064
rect 35676 381024 40040 381052
rect 35676 381012 35682 381024
rect 40034 381012 40040 381024
rect 40092 381012 40098 381064
rect 35802 379924 35808 379976
rect 35860 379964 35866 379976
rect 41506 379964 41512 379976
rect 35860 379936 41512 379964
rect 35860 379924 35866 379936
rect 41506 379924 41512 379936
rect 41564 379924 41570 379976
rect 35618 379652 35624 379704
rect 35676 379692 35682 379704
rect 39942 379692 39948 379704
rect 35676 379664 39948 379692
rect 35676 379652 35682 379664
rect 39942 379652 39948 379664
rect 40000 379652 40006 379704
rect 35802 379516 35808 379568
rect 35860 379556 35866 379568
rect 39574 379556 39580 379568
rect 35860 379528 39580 379556
rect 35860 379516 35866 379528
rect 39574 379516 39580 379528
rect 39632 379516 39638 379568
rect 670418 379448 670424 379500
rect 670476 379488 670482 379500
rect 675110 379488 675116 379500
rect 670476 379460 675116 379488
rect 670476 379448 670482 379460
rect 675110 379448 675116 379460
rect 675168 379448 675174 379500
rect 35802 378292 35808 378344
rect 35860 378332 35866 378344
rect 41230 378332 41236 378344
rect 35860 378304 41236 378332
rect 35860 378292 35866 378304
rect 41230 378292 41236 378304
rect 41288 378292 41294 378344
rect 651558 378156 651564 378208
rect 651616 378196 651622 378208
rect 663058 378196 663064 378208
rect 651616 378168 663064 378196
rect 651616 378156 651622 378168
rect 663058 378156 663064 378168
rect 663116 378156 663122 378208
rect 673362 377816 673368 377868
rect 673420 377856 673426 377868
rect 675294 377856 675300 377868
rect 673420 377828 675300 377856
rect 673420 377816 673426 377828
rect 675294 377816 675300 377828
rect 675352 377816 675358 377868
rect 35618 377000 35624 377052
rect 35676 377040 35682 377052
rect 35676 377012 38654 377040
rect 35676 377000 35682 377012
rect 38626 376972 38654 377012
rect 41690 376972 41696 376984
rect 38626 376944 41696 376972
rect 41690 376932 41696 376944
rect 41748 376932 41754 376984
rect 42058 376796 42064 376848
rect 42116 376836 42122 376848
rect 42116 376808 51074 376836
rect 42116 376796 42122 376808
rect 35802 376728 35808 376780
rect 35860 376768 35866 376780
rect 41690 376768 41696 376780
rect 35860 376740 41696 376768
rect 35860 376728 35866 376740
rect 41690 376728 41696 376740
rect 41748 376728 41754 376780
rect 51046 376768 51074 376808
rect 53466 376768 53472 376780
rect 51046 376740 53472 376768
rect 53466 376728 53472 376740
rect 53524 376728 53530 376780
rect 672994 376592 673000 376644
rect 673052 376632 673058 376644
rect 675110 376632 675116 376644
rect 673052 376604 675116 376632
rect 673052 376592 673058 376604
rect 675110 376592 675116 376604
rect 675168 376592 675174 376644
rect 28810 375844 28816 375896
rect 28868 375884 28874 375896
rect 33778 375884 33784 375896
rect 28868 375856 33784 375884
rect 28868 375844 28874 375856
rect 33778 375844 33784 375856
rect 33836 375844 33842 375896
rect 35802 375572 35808 375624
rect 35860 375612 35866 375624
rect 41690 375612 41696 375624
rect 35860 375584 41696 375612
rect 35860 375572 35866 375584
rect 41690 375572 41696 375584
rect 41748 375572 41754 375624
rect 42058 375504 42064 375556
rect 42116 375544 42122 375556
rect 52270 375544 52276 375556
rect 42116 375516 52276 375544
rect 42116 375504 42122 375516
rect 52270 375504 52276 375516
rect 52328 375504 52334 375556
rect 49326 375368 49332 375420
rect 49384 375408 49390 375420
rect 62114 375408 62120 375420
rect 49384 375380 62120 375408
rect 49384 375368 49390 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 33778 373260 33784 373312
rect 33836 373300 33842 373312
rect 41690 373300 41696 373312
rect 33836 373272 41696 373300
rect 33836 373260 33842 373272
rect 41690 373260 41696 373272
rect 41748 373260 41754 373312
rect 672810 372512 672816 372564
rect 672868 372552 672874 372564
rect 675294 372552 675300 372564
rect 672868 372524 675300 372552
rect 672868 372512 672874 372524
rect 675294 372512 675300 372524
rect 675352 372512 675358 372564
rect 32398 371832 32404 371884
rect 32456 371872 32462 371884
rect 41690 371872 41696 371884
rect 32456 371844 41696 371872
rect 32456 371832 32462 371844
rect 41690 371832 41696 371844
rect 41748 371832 41754 371884
rect 42058 371696 42064 371748
rect 42116 371736 42122 371748
rect 42610 371736 42616 371748
rect 42116 371708 42616 371736
rect 42116 371696 42122 371708
rect 42610 371696 42616 371708
rect 42668 371696 42674 371748
rect 42242 365644 42248 365696
rect 42300 365684 42306 365696
rect 45186 365684 45192 365696
rect 42300 365656 45192 365684
rect 42300 365644 42306 365656
rect 45186 365644 45192 365656
rect 45244 365644 45250 365696
rect 651558 364352 651564 364404
rect 651616 364392 651622 364404
rect 664622 364392 664628 364404
rect 651616 364364 664628 364392
rect 651616 364352 651622 364364
rect 664622 364352 664628 364364
rect 664680 364352 664686 364404
rect 42334 364216 42340 364268
rect 42392 364256 42398 364268
rect 52086 364256 52092 364268
rect 42392 364228 52092 364256
rect 42392 364216 42398 364228
rect 52086 364216 52092 364228
rect 52144 364216 52150 364268
rect 42334 364080 42340 364132
rect 42392 364120 42398 364132
rect 43806 364120 43812 364132
rect 42392 364092 43812 364120
rect 42392 364080 42398 364092
rect 43806 364080 43812 364092
rect 43864 364080 43870 364132
rect 42426 360136 42432 360188
rect 42484 360176 42490 360188
rect 44358 360176 44364 360188
rect 42484 360148 44364 360176
rect 42484 360136 42490 360148
rect 44358 360136 44364 360148
rect 44416 360136 44422 360188
rect 42150 359932 42156 359984
rect 42208 359972 42214 359984
rect 43254 359972 43260 359984
rect 42208 359944 43260 359972
rect 42208 359932 42214 359944
rect 43254 359932 43260 359944
rect 43312 359932 43318 359984
rect 675294 357864 675300 357876
rect 663766 357836 675300 357864
rect 659102 357688 659108 357740
rect 659160 357728 659166 357740
rect 663766 357728 663794 357836
rect 675294 357824 675300 357836
rect 675352 357824 675358 357876
rect 659160 357700 663794 357728
rect 659160 357688 659166 357700
rect 664806 357552 664812 357604
rect 664864 357592 664870 357604
rect 675478 357592 675484 357604
rect 664864 357564 675484 357592
rect 664864 357552 664870 357564
rect 675478 357552 675484 357564
rect 675536 357552 675542 357604
rect 660482 357416 660488 357468
rect 660540 357456 660546 357468
rect 675110 357456 675116 357468
rect 660540 357428 675116 357456
rect 660540 357416 660546 357428
rect 675110 357416 675116 357428
rect 675168 357416 675174 357468
rect 673914 357008 673920 357060
rect 673972 357048 673978 357060
rect 675478 357048 675484 357060
rect 673972 357020 675484 357048
rect 673972 357008 673978 357020
rect 675478 357008 675484 357020
rect 675536 357008 675542 357060
rect 50890 356668 50896 356720
rect 50948 356708 50954 356720
rect 62114 356708 62120 356720
rect 50948 356680 62120 356708
rect 50948 356668 50954 356680
rect 62114 356668 62120 356680
rect 62172 356668 62178 356720
rect 42426 355988 42432 356040
rect 42484 356028 42490 356040
rect 42978 356028 42984 356040
rect 42484 356000 42984 356028
rect 42484 355988 42490 356000
rect 42978 355988 42984 356000
rect 43036 355988 43042 356040
rect 672442 355852 672448 355904
rect 672500 355892 672506 355904
rect 675478 355892 675484 355904
rect 672500 355864 675484 355892
rect 672500 355852 672506 355864
rect 675478 355852 675484 355864
rect 675536 355852 675542 355904
rect 672442 355376 672448 355428
rect 672500 355416 672506 355428
rect 675478 355416 675484 355428
rect 672500 355388 675484 355416
rect 672500 355376 672506 355388
rect 675478 355376 675484 355388
rect 675536 355376 675542 355428
rect 673178 355036 673184 355088
rect 673236 355076 673242 355088
rect 675478 355076 675484 355088
rect 673236 355048 675484 355076
rect 673236 355036 673242 355048
rect 675478 355036 675484 355048
rect 675536 355036 675542 355088
rect 673178 354560 673184 354612
rect 673236 354600 673242 354612
rect 675478 354600 675484 354612
rect 673236 354572 675484 354600
rect 673236 354560 673242 354572
rect 675478 354560 675484 354572
rect 675536 354560 675542 354612
rect 667842 353608 667848 353660
rect 667900 353648 667906 353660
rect 675478 353648 675484 353660
rect 667900 353620 675484 353648
rect 667900 353608 667906 353620
rect 675478 353608 675484 353620
rect 675536 353608 675542 353660
rect 671798 353336 671804 353388
rect 671856 353376 671862 353388
rect 675478 353376 675484 353388
rect 671856 353348 675484 353376
rect 671856 353336 671862 353348
rect 675478 353336 675484 353348
rect 675536 353336 675542 353388
rect 670418 352520 670424 352572
rect 670476 352560 670482 352572
rect 675478 352560 675484 352572
rect 670476 352532 675484 352560
rect 670476 352520 670482 352532
rect 675478 352520 675484 352532
rect 675536 352520 675542 352572
rect 673362 350072 673368 350124
rect 673420 350112 673426 350124
rect 675478 350112 675484 350124
rect 673420 350084 675484 350112
rect 673420 350072 673426 350084
rect 675478 350072 675484 350084
rect 675536 350072 675542 350124
rect 673546 349664 673552 349716
rect 673604 349704 673610 349716
rect 675478 349704 675484 349716
rect 673604 349676 675484 349704
rect 673604 349664 673610 349676
rect 675478 349664 675484 349676
rect 675536 349664 675542 349716
rect 669774 349256 669780 349308
rect 669832 349296 669838 349308
rect 675478 349296 675484 349308
rect 669832 349268 675484 349296
rect 669832 349256 669838 349268
rect 675478 349256 675484 349268
rect 675536 349256 675542 349308
rect 672994 348848 673000 348900
rect 673052 348888 673058 348900
rect 675478 348888 675484 348900
rect 673052 348860 675484 348888
rect 673052 348848 673058 348860
rect 675478 348848 675484 348860
rect 675536 348848 675542 348900
rect 671154 348440 671160 348492
rect 671212 348480 671218 348492
rect 675478 348480 675484 348492
rect 671212 348452 675484 348480
rect 671212 348440 671218 348452
rect 675478 348440 675484 348452
rect 675536 348440 675542 348492
rect 675846 347896 675852 347948
rect 675904 347936 675910 347948
rect 676582 347936 676588 347948
rect 675904 347908 676588 347936
rect 675904 347896 675910 347908
rect 676582 347896 676588 347908
rect 676640 347896 676646 347948
rect 672350 347216 672356 347268
rect 672408 347256 672414 347268
rect 675478 347256 675484 347268
rect 672408 347228 675484 347256
rect 672408 347216 672414 347228
rect 675478 347216 675484 347228
rect 675536 347216 675542 347268
rect 45186 347012 45192 347064
rect 45244 347052 45250 347064
rect 62114 347052 62120 347064
rect 45244 347024 62120 347052
rect 45244 347012 45250 347024
rect 62114 347012 62120 347024
rect 62172 347012 62178 347064
rect 675846 346400 675852 346452
rect 675904 346440 675910 346452
rect 683114 346440 683120 346452
rect 675904 346412 683120 346440
rect 675904 346400 675910 346412
rect 683114 346400 683120 346412
rect 683172 346400 683178 346452
rect 35802 344020 35808 344072
rect 35860 344060 35866 344072
rect 39206 344060 39212 344072
rect 35860 344032 39212 344060
rect 35860 344020 35866 344032
rect 39206 344020 39212 344032
rect 39264 344020 39270 344072
rect 41690 343856 41696 343868
rect 41386 343828 41696 343856
rect 35802 343748 35808 343800
rect 35860 343788 35866 343800
rect 41386 343788 41414 343828
rect 41690 343816 41696 343828
rect 41748 343816 41754 343868
rect 42058 343816 42064 343868
rect 42116 343856 42122 343868
rect 50706 343856 50712 343868
rect 42116 343828 50712 343856
rect 42116 343816 42122 343828
rect 50706 343816 50712 343828
rect 50764 343816 50770 343868
rect 35860 343760 41414 343788
rect 35860 343748 35866 343760
rect 35618 343612 35624 343664
rect 35676 343652 35682 343664
rect 41690 343652 41696 343664
rect 35676 343624 41696 343652
rect 35676 343612 35682 343624
rect 41690 343612 41696 343624
rect 41748 343612 41754 343664
rect 42058 343612 42064 343664
rect 42116 343652 42122 343664
rect 56226 343652 56232 343664
rect 42116 343624 56232 343652
rect 42116 343612 42122 343624
rect 56226 343612 56232 343624
rect 56284 343612 56290 343664
rect 35802 342660 35808 342712
rect 35860 342700 35866 342712
rect 40310 342700 40316 342712
rect 35860 342672 40316 342700
rect 35860 342660 35866 342672
rect 40310 342660 40316 342672
rect 40368 342660 40374 342712
rect 35618 342388 35624 342440
rect 35676 342428 35682 342440
rect 40034 342428 40040 342440
rect 35676 342400 40040 342428
rect 35676 342388 35682 342400
rect 40034 342388 40040 342400
rect 40092 342388 40098 342440
rect 35618 342252 35624 342304
rect 35676 342292 35682 342304
rect 41690 342292 41696 342304
rect 35676 342264 41696 342292
rect 35676 342252 35682 342264
rect 41690 342252 41696 342264
rect 41748 342252 41754 342304
rect 42058 342252 42064 342304
rect 42116 342292 42122 342304
rect 44634 342292 44640 342304
rect 42116 342264 44640 342292
rect 42116 342252 42122 342264
rect 44634 342252 44640 342264
rect 44692 342252 44698 342304
rect 35802 341436 35808 341488
rect 35860 341476 35866 341488
rect 41690 341476 41696 341488
rect 35860 341448 41696 341476
rect 35860 341436 35866 341448
rect 41690 341436 41696 341448
rect 41748 341436 41754 341488
rect 42058 341368 42064 341420
rect 42116 341408 42122 341420
rect 42886 341408 42892 341420
rect 42116 341380 42892 341408
rect 42116 341368 42122 341380
rect 42886 341368 42892 341380
rect 42944 341368 42950 341420
rect 41690 341272 41696 341284
rect 41386 341244 41696 341272
rect 35342 341164 35348 341216
rect 35400 341204 35406 341216
rect 41386 341204 41414 341244
rect 41690 341232 41696 341244
rect 41748 341232 41754 341284
rect 42058 341232 42064 341284
rect 42116 341272 42122 341284
rect 42702 341272 42708 341284
rect 42116 341244 42708 341272
rect 42116 341232 42122 341244
rect 42702 341232 42708 341244
rect 42760 341232 42766 341284
rect 35400 341176 41414 341204
rect 35400 341164 35406 341176
rect 35802 341028 35808 341080
rect 35860 341068 35866 341080
rect 41690 341068 41696 341080
rect 35860 341040 41696 341068
rect 35860 341028 35866 341040
rect 41690 341028 41696 341040
rect 41748 341028 41754 341080
rect 42058 341028 42064 341080
rect 42116 341068 42122 341080
rect 43622 341068 43628 341080
rect 42116 341040 43628 341068
rect 42116 341028 42122 341040
rect 43622 341028 43628 341040
rect 43680 341028 43686 341080
rect 35618 340892 35624 340944
rect 35676 340932 35682 340944
rect 41690 340932 41696 340944
rect 35676 340904 41696 340932
rect 35676 340892 35682 340904
rect 41690 340892 41696 340904
rect 41748 340892 41754 340944
rect 42058 340892 42064 340944
rect 42116 340932 42122 340944
rect 44450 340932 44456 340944
rect 42116 340904 44456 340932
rect 42116 340892 42122 340904
rect 44450 340892 44456 340904
rect 44508 340892 44514 340944
rect 35802 339600 35808 339652
rect 35860 339640 35866 339652
rect 41414 339640 41420 339652
rect 35860 339612 41420 339640
rect 35860 339600 35866 339612
rect 41414 339600 41420 339612
rect 41472 339600 41478 339652
rect 35802 338376 35808 338428
rect 35860 338416 35866 338428
rect 41690 338416 41696 338428
rect 35860 338388 41696 338416
rect 35860 338376 35866 338388
rect 41690 338376 41696 338388
rect 41748 338376 41754 338428
rect 35618 338104 35624 338156
rect 35676 338144 35682 338156
rect 41506 338144 41512 338156
rect 35676 338116 41512 338144
rect 35676 338104 35682 338116
rect 41506 338104 41512 338116
rect 41564 338104 41570 338156
rect 652202 338104 652208 338156
rect 652260 338144 652266 338156
rect 667382 338144 667388 338156
rect 652260 338116 667388 338144
rect 652260 338104 652266 338116
rect 667382 338104 667388 338116
rect 667440 338104 667446 338156
rect 671798 338036 671804 338088
rect 671856 338076 671862 338088
rect 675110 338076 675116 338088
rect 671856 338048 675116 338076
rect 671856 338036 671862 338048
rect 675110 338036 675116 338048
rect 675168 338036 675174 338088
rect 674466 337900 674472 337952
rect 674524 337940 674530 337952
rect 675110 337940 675116 337952
rect 674524 337912 675116 337940
rect 674524 337900 674530 337912
rect 675110 337900 675116 337912
rect 675168 337900 675174 337952
rect 35802 337084 35808 337136
rect 35860 337124 35866 337136
rect 39850 337124 39856 337136
rect 35860 337096 39856 337124
rect 35860 337084 35866 337096
rect 39850 337084 39856 337096
rect 39908 337084 39914 337136
rect 35802 336880 35808 336932
rect 35860 336920 35866 336932
rect 40310 336920 40316 336932
rect 35860 336892 40316 336920
rect 35860 336880 35866 336892
rect 40310 336880 40316 336892
rect 40368 336880 40374 336932
rect 35526 336744 35532 336796
rect 35584 336784 35590 336796
rect 41690 336784 41696 336796
rect 35584 336756 41696 336784
rect 35584 336744 35590 336756
rect 41690 336744 41696 336756
rect 41748 336744 41754 336796
rect 42058 336744 42064 336796
rect 42116 336784 42122 336796
rect 43622 336784 43628 336796
rect 42116 336756 43628 336784
rect 42116 336744 42122 336756
rect 43622 336744 43628 336756
rect 43680 336744 43686 336796
rect 46566 336744 46572 336796
rect 46624 336784 46630 336796
rect 62114 336784 62120 336796
rect 46624 336756 62120 336784
rect 46624 336744 46630 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 673362 335996 673368 336048
rect 673420 336036 673426 336048
rect 674926 336036 674932 336048
rect 673420 336008 674932 336036
rect 673420 335996 673426 336008
rect 674926 335996 674932 336008
rect 674984 335996 674990 336048
rect 673546 335860 673552 335912
rect 673604 335900 673610 335912
rect 675386 335900 675392 335912
rect 673604 335872 675392 335900
rect 673604 335860 673610 335872
rect 675386 335860 675392 335872
rect 675444 335860 675450 335912
rect 35802 335588 35808 335640
rect 35860 335628 35866 335640
rect 40862 335628 40868 335640
rect 35860 335600 40868 335628
rect 35860 335588 35866 335600
rect 40862 335588 40868 335600
rect 40920 335588 40926 335640
rect 35618 335316 35624 335368
rect 35676 335356 35682 335368
rect 40218 335356 40224 335368
rect 35676 335328 40224 335356
rect 35676 335316 35682 335328
rect 40218 335316 40224 335328
rect 40276 335316 40282 335368
rect 35618 334364 35624 334416
rect 35676 334404 35682 334416
rect 40310 334404 40316 334416
rect 35676 334376 40316 334404
rect 35676 334364 35682 334376
rect 40310 334364 40316 334376
rect 40368 334364 40374 334416
rect 35434 334092 35440 334144
rect 35492 334132 35498 334144
rect 40126 334132 40132 334144
rect 35492 334104 40132 334132
rect 35492 334092 35498 334104
rect 40126 334092 40132 334104
rect 40184 334092 40190 334144
rect 35802 333956 35808 334008
rect 35860 333996 35866 334008
rect 41690 333996 41696 334008
rect 35860 333968 41696 333996
rect 35860 333956 35866 333968
rect 41690 333956 41696 333968
rect 41748 333956 41754 334008
rect 42058 333956 42064 334008
rect 42116 333996 42122 334008
rect 50706 333996 50712 334008
rect 42116 333968 50712 333996
rect 42116 333956 42122 333968
rect 50706 333956 50712 333968
rect 50764 333956 50770 334008
rect 670418 333888 670424 333940
rect 670476 333928 670482 333940
rect 675110 333928 675116 333940
rect 670476 333900 675116 333928
rect 670476 333888 670482 333900
rect 675110 333888 675116 333900
rect 675168 333888 675174 333940
rect 35802 333004 35808 333056
rect 35860 333044 35866 333056
rect 35860 333004 35894 333044
rect 35866 332908 35894 333004
rect 39298 332908 39304 332920
rect 35866 332880 39304 332908
rect 39298 332868 39304 332880
rect 39356 332868 39362 332920
rect 35802 332596 35808 332648
rect 35860 332636 35866 332648
rect 41690 332636 41696 332648
rect 35860 332608 41696 332636
rect 35860 332596 35866 332608
rect 41690 332596 41696 332608
rect 41748 332596 41754 332648
rect 42058 332596 42064 332648
rect 42116 332636 42122 332648
rect 56226 332636 56232 332648
rect 42116 332608 56232 332636
rect 42116 332596 42122 332608
rect 56226 332596 56232 332608
rect 56284 332596 56290 332648
rect 669774 332596 669780 332648
rect 669832 332636 669838 332648
rect 675110 332636 675116 332648
rect 669832 332608 675116 332636
rect 669832 332596 669838 332608
rect 675110 332596 675116 332608
rect 675168 332596 675174 332648
rect 672994 331712 673000 331764
rect 673052 331752 673058 331764
rect 675110 331752 675116 331764
rect 673052 331724 675116 331752
rect 673052 331712 673058 331724
rect 675110 331712 675116 331724
rect 675168 331712 675174 331764
rect 42426 327020 42432 327072
rect 42484 327060 42490 327072
rect 45830 327060 45836 327072
rect 42484 327032 45836 327060
rect 42484 327020 42490 327032
rect 45830 327020 45836 327032
rect 45888 327020 45894 327072
rect 670234 325592 670240 325644
rect 670292 325632 670298 325644
rect 675110 325632 675116 325644
rect 670292 325604 675116 325632
rect 670292 325592 670298 325604
rect 675110 325592 675116 325604
rect 675168 325592 675174 325644
rect 667842 325456 667848 325508
rect 667900 325496 667906 325508
rect 674926 325496 674932 325508
rect 667900 325468 674932 325496
rect 667900 325456 667906 325468
rect 674926 325456 674932 325468
rect 674984 325456 674990 325508
rect 42426 325320 42432 325372
rect 42484 325360 42490 325372
rect 44634 325360 44640 325372
rect 42484 325332 44640 325360
rect 42484 325320 42490 325332
rect 44634 325320 44640 325332
rect 44692 325320 44698 325372
rect 651558 324300 651564 324352
rect 651616 324340 651622 324352
rect 673546 324340 673552 324352
rect 651616 324312 673552 324340
rect 651616 324300 651622 324312
rect 673546 324300 673552 324312
rect 673604 324300 673610 324352
rect 42426 321512 42432 321564
rect 42484 321552 42490 321564
rect 55030 321552 55036 321564
rect 42484 321524 55036 321552
rect 42484 321512 42490 321524
rect 55030 321512 55036 321524
rect 55088 321512 55094 321564
rect 42426 321240 42432 321292
rect 42484 321280 42490 321292
rect 43990 321280 43996 321292
rect 42484 321252 43996 321280
rect 42484 321240 42490 321252
rect 43990 321240 43996 321252
rect 44048 321240 44054 321292
rect 42242 319948 42248 320000
rect 42300 319988 42306 320000
rect 45370 319988 45376 320000
rect 42300 319960 45376 319988
rect 42300 319948 42306 319960
rect 45370 319948 45376 319960
rect 45428 319948 45434 320000
rect 42426 319132 42432 319184
rect 42484 319172 42490 319184
rect 46014 319172 46020 319184
rect 42484 319144 46020 319172
rect 42484 319132 42490 319144
rect 46014 319132 46020 319144
rect 46072 319132 46078 319184
rect 42610 318724 42616 318776
rect 42668 318764 42674 318776
rect 46750 318764 46756 318776
rect 42668 318736 46756 318764
rect 42668 318724 42674 318736
rect 46750 318724 46756 318736
rect 46808 318724 46814 318776
rect 42426 317364 42432 317416
rect 42484 317404 42490 317416
rect 43070 317404 43076 317416
rect 42484 317376 43076 317404
rect 42484 317364 42490 317376
rect 43070 317364 43076 317376
rect 43128 317364 43134 317416
rect 42426 316888 42432 316940
rect 42484 316928 42490 316940
rect 43806 316928 43812 316940
rect 42484 316900 43812 316928
rect 42484 316888 42490 316900
rect 43806 316888 43812 316900
rect 43864 316888 43870 316940
rect 42426 315868 42432 315920
rect 42484 315908 42490 315920
rect 43622 315908 43628 315920
rect 42484 315880 43628 315908
rect 42484 315868 42490 315880
rect 43622 315868 43628 315880
rect 43680 315868 43686 315920
rect 43806 313896 43812 313948
rect 43864 313936 43870 313948
rect 62758 313936 62764 313948
rect 43864 313908 62764 313936
rect 43864 313896 43870 313908
rect 62758 313896 62764 313908
rect 62816 313896 62822 313948
rect 663242 313420 663248 313472
rect 663300 313460 663306 313472
rect 675478 313460 675484 313472
rect 663300 313432 675484 313460
rect 663300 313420 663306 313432
rect 675478 313420 675484 313432
rect 675536 313420 675542 313472
rect 661862 313284 661868 313336
rect 661920 313324 661926 313336
rect 675478 313324 675484 313336
rect 661920 313296 675484 313324
rect 661920 313284 661926 313296
rect 675478 313284 675484 313296
rect 675536 313284 675542 313336
rect 673914 312468 673920 312520
rect 673972 312508 673978 312520
rect 675478 312508 675484 312520
rect 673972 312480 675484 312508
rect 673972 312468 673978 312480
rect 675478 312468 675484 312480
rect 675536 312468 675542 312520
rect 660666 311992 660672 312044
rect 660724 312032 660730 312044
rect 675294 312032 675300 312044
rect 660724 312004 675300 312032
rect 660724 311992 660730 312004
rect 675294 311992 675300 312004
rect 675352 311992 675358 312044
rect 664254 311856 664260 311908
rect 664312 311896 664318 311908
rect 675478 311896 675484 311908
rect 664312 311868 675484 311896
rect 664312 311856 664318 311868
rect 675478 311856 675484 311868
rect 675536 311856 675542 311908
rect 666370 310700 666376 310752
rect 666428 310740 666434 310752
rect 675478 310740 675484 310752
rect 666428 310712 675484 310740
rect 666428 310700 666434 310712
rect 675478 310700 675484 310712
rect 675536 310700 675542 310752
rect 651558 310496 651564 310548
rect 651616 310536 651622 310548
rect 667198 310536 667204 310548
rect 651616 310508 667204 310536
rect 651616 310496 651622 310508
rect 667198 310496 667204 310508
rect 667256 310496 667262 310548
rect 42426 310428 42432 310480
rect 42484 310468 42490 310480
rect 45554 310468 45560 310480
rect 42484 310440 45560 310468
rect 42484 310428 42490 310440
rect 45554 310428 45560 310440
rect 45612 310428 45618 310480
rect 670418 310360 670424 310412
rect 670476 310400 670482 310412
rect 675478 310400 675484 310412
rect 670476 310372 675484 310400
rect 670476 310360 670482 310372
rect 675478 310360 675484 310372
rect 675536 310360 675542 310412
rect 673178 310020 673184 310072
rect 673236 310060 673242 310072
rect 675478 310060 675484 310072
rect 673236 310032 675484 310060
rect 673236 310020 673242 310032
rect 675478 310020 675484 310032
rect 675536 310020 675542 310072
rect 664990 309136 664996 309188
rect 665048 309176 665054 309188
rect 675478 309176 675484 309188
rect 665048 309148 675484 309176
rect 665048 309136 665054 309148
rect 675478 309136 675484 309148
rect 675536 309136 675542 309188
rect 673270 305464 673276 305516
rect 673328 305504 673334 305516
rect 675478 305504 675484 305516
rect 673328 305476 675484 305504
rect 673328 305464 673334 305476
rect 675478 305464 675484 305476
rect 675536 305464 675542 305516
rect 673086 303832 673092 303884
rect 673144 303872 673150 303884
rect 675478 303872 675484 303884
rect 673144 303844 675484 303872
rect 673144 303832 673150 303844
rect 675478 303832 675484 303844
rect 675536 303832 675542 303884
rect 672810 303424 672816 303476
rect 672868 303464 672874 303476
rect 675478 303464 675484 303476
rect 672868 303436 675484 303464
rect 672868 303424 672874 303436
rect 675478 303424 675484 303436
rect 675536 303424 675542 303476
rect 670234 302200 670240 302252
rect 670292 302240 670298 302252
rect 675478 302240 675484 302252
rect 670292 302212 675484 302240
rect 670292 302200 670298 302212
rect 675478 302200 675484 302212
rect 675536 302200 675542 302252
rect 680354 302200 680360 302252
rect 680412 302240 680418 302252
rect 683114 302240 683120 302252
rect 680412 302212 683120 302240
rect 680412 302200 680418 302212
rect 683114 302200 683120 302212
rect 683172 302200 683178 302252
rect 43622 301248 43628 301300
rect 43680 301288 43686 301300
rect 50890 301288 50896 301300
rect 43680 301260 50896 301288
rect 43680 301248 43686 301260
rect 50890 301248 50896 301260
rect 50948 301248 50954 301300
rect 43070 300976 43076 301028
rect 43128 301016 43134 301028
rect 49326 301016 49332 301028
rect 43128 300988 49332 301016
rect 43128 300976 43134 300988
rect 49326 300976 49332 300988
rect 49384 300976 49390 301028
rect 41690 299724 41696 299736
rect 41386 299696 41696 299724
rect 41138 299616 41144 299668
rect 41196 299656 41202 299668
rect 41386 299656 41414 299696
rect 41690 299684 41696 299696
rect 41748 299684 41754 299736
rect 42058 299684 42064 299736
rect 42116 299724 42122 299736
rect 43254 299724 43260 299736
rect 42116 299696 43260 299724
rect 42116 299684 42122 299696
rect 43254 299684 43260 299696
rect 43312 299684 43318 299736
rect 41196 299628 41414 299656
rect 41196 299616 41202 299628
rect 40954 299480 40960 299532
rect 41012 299520 41018 299532
rect 41690 299520 41696 299532
rect 41012 299492 41696 299520
rect 41012 299480 41018 299492
rect 41690 299480 41696 299492
rect 41748 299480 41754 299532
rect 42058 299480 42064 299532
rect 42116 299520 42122 299532
rect 48130 299520 48136 299532
rect 42116 299492 48136 299520
rect 42116 299480 42122 299492
rect 48130 299480 48136 299492
rect 48188 299480 48194 299532
rect 41690 298364 41696 298376
rect 41386 298336 41696 298364
rect 40954 298256 40960 298308
rect 41012 298256 41018 298308
rect 41138 298256 41144 298308
rect 41196 298296 41202 298308
rect 41386 298296 41414 298336
rect 41690 298324 41696 298336
rect 41748 298324 41754 298376
rect 42058 298324 42064 298376
rect 42116 298364 42122 298376
rect 42886 298364 42892 298376
rect 42116 298336 42892 298364
rect 42116 298324 42122 298336
rect 42886 298324 42892 298336
rect 42944 298324 42950 298376
rect 41196 298268 41414 298296
rect 41196 298256 41202 298268
rect 40972 298160 41000 298256
rect 42058 298188 42064 298240
rect 42116 298228 42122 298240
rect 44450 298228 44456 298240
rect 42116 298200 44456 298228
rect 42116 298188 42122 298200
rect 44450 298188 44456 298200
rect 44508 298188 44514 298240
rect 41690 298160 41696 298172
rect 40972 298132 41696 298160
rect 41690 298120 41696 298132
rect 41748 298120 41754 298172
rect 49326 298120 49332 298172
rect 49384 298160 49390 298172
rect 62114 298160 62120 298172
rect 49384 298132 62120 298160
rect 49384 298120 49390 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 41690 296936 41696 296948
rect 41386 296908 41696 296936
rect 41138 296828 41144 296880
rect 41196 296868 41202 296880
rect 41386 296868 41414 296908
rect 41690 296896 41696 296908
rect 41748 296896 41754 296948
rect 42058 296896 42064 296948
rect 42116 296936 42122 296948
rect 44174 296936 44180 296948
rect 42116 296908 44180 296936
rect 42116 296896 42122 296908
rect 44174 296896 44180 296908
rect 44232 296896 44238 296948
rect 675846 296896 675852 296948
rect 675904 296936 675910 296948
rect 680998 296936 681004 296948
rect 675904 296908 681004 296936
rect 675904 296896 675910 296908
rect 680998 296896 681004 296908
rect 681056 296896 681062 296948
rect 41196 296840 41414 296868
rect 41196 296828 41202 296840
rect 40954 296692 40960 296744
rect 41012 296732 41018 296744
rect 41690 296732 41696 296744
rect 41012 296704 41696 296732
rect 41012 296692 41018 296704
rect 41690 296692 41696 296704
rect 41748 296692 41754 296744
rect 42058 296692 42064 296744
rect 42116 296732 42122 296744
rect 44542 296732 44548 296744
rect 42116 296704 44548 296732
rect 42116 296692 42122 296704
rect 44542 296692 44548 296704
rect 44600 296692 44606 296744
rect 675478 296352 675484 296404
rect 675536 296352 675542 296404
rect 675496 295928 675524 296352
rect 675478 295876 675484 295928
rect 675536 295876 675542 295928
rect 41322 293972 41328 294024
rect 41380 294012 41386 294024
rect 41690 294012 41696 294024
rect 41380 293984 41696 294012
rect 41380 293972 41386 293984
rect 41690 293972 41696 293984
rect 41748 293972 41754 294024
rect 42058 293972 42064 294024
rect 42116 294012 42122 294024
rect 47210 294012 47216 294024
rect 42116 293984 47216 294012
rect 42116 293972 42122 293984
rect 47210 293972 47216 293984
rect 47268 293972 47274 294024
rect 40494 292544 40500 292596
rect 40552 292584 40558 292596
rect 41598 292584 41604 292596
rect 40552 292556 41604 292584
rect 40552 292544 40558 292556
rect 41598 292544 41604 292556
rect 41656 292544 41662 292596
rect 674466 292272 674472 292324
rect 674524 292312 674530 292324
rect 675110 292312 675116 292324
rect 674524 292284 675116 292312
rect 674524 292272 674530 292284
rect 675110 292272 675116 292284
rect 675168 292272 675174 292324
rect 41138 291184 41144 291236
rect 41196 291224 41202 291236
rect 41690 291224 41696 291236
rect 41196 291196 41696 291224
rect 41196 291184 41202 291196
rect 41690 291184 41696 291196
rect 41748 291184 41754 291236
rect 42058 291184 42064 291236
rect 42116 291224 42122 291236
rect 43990 291224 43996 291236
rect 42116 291196 43996 291224
rect 42116 291184 42122 291196
rect 43990 291184 43996 291196
rect 44048 291184 44054 291236
rect 43622 290300 43628 290352
rect 43680 290340 43686 290352
rect 49510 290340 49516 290352
rect 43680 290312 49516 290340
rect 43680 290300 43686 290312
rect 49510 290300 49516 290312
rect 49568 290300 49574 290352
rect 42058 290028 42064 290080
rect 42116 290068 42122 290080
rect 42116 290040 51074 290068
rect 42116 290028 42122 290040
rect 51046 290000 51074 290040
rect 59998 290000 60004 290012
rect 51046 289972 60004 290000
rect 59998 289960 60004 289972
rect 60056 289960 60062 290012
rect 40954 289824 40960 289876
rect 41012 289864 41018 289876
rect 41690 289864 41696 289876
rect 41012 289836 41696 289864
rect 41012 289824 41018 289836
rect 41690 289824 41696 289836
rect 41748 289824 41754 289876
rect 42058 289824 42064 289876
rect 42116 289864 42122 289876
rect 64138 289864 64144 289876
rect 42116 289836 64144 289864
rect 42116 289824 42122 289836
rect 64138 289824 64144 289836
rect 64196 289824 64202 289876
rect 41138 289076 41144 289128
rect 41196 289116 41202 289128
rect 41690 289116 41696 289128
rect 41196 289088 41696 289116
rect 41196 289076 41202 289088
rect 41690 289076 41696 289088
rect 41748 289076 41754 289128
rect 37918 284996 37924 285048
rect 37976 285036 37982 285048
rect 41690 285036 41696 285048
rect 37976 285008 41696 285036
rect 37976 284996 37982 285008
rect 41690 284996 41696 285008
rect 41748 284996 41754 285048
rect 43622 284316 43628 284368
rect 43680 284356 43686 284368
rect 62114 284356 62120 284368
rect 43680 284328 62120 284356
rect 43680 284316 43686 284328
rect 62114 284316 62120 284328
rect 62172 284316 62178 284368
rect 651558 284316 651564 284368
rect 651616 284356 651622 284368
rect 664806 284356 664812 284368
rect 651616 284328 664812 284356
rect 651616 284316 651622 284328
rect 664806 284316 664812 284328
rect 664864 284316 664870 284368
rect 42426 281460 42432 281512
rect 42484 281500 42490 281512
rect 43438 281500 43444 281512
rect 42484 281472 43444 281500
rect 42484 281460 42490 281472
rect 43438 281460 43444 281472
rect 43496 281460 43502 281512
rect 42426 280100 42432 280152
rect 42484 280140 42490 280152
rect 42978 280140 42984 280152
rect 42484 280112 42984 280140
rect 42484 280100 42490 280112
rect 42978 280100 42984 280112
rect 43036 280100 43042 280152
rect 406930 278672 406936 278724
rect 406988 278712 406994 278724
rect 499574 278712 499580 278724
rect 406988 278684 499580 278712
rect 406988 278672 406994 278684
rect 499574 278672 499580 278684
rect 499632 278672 499638 278724
rect 437198 278536 437204 278588
rect 437256 278576 437262 278588
rect 546678 278576 546684 278588
rect 437256 278548 546684 278576
rect 437256 278536 437262 278548
rect 546678 278536 546684 278548
rect 546736 278536 546742 278588
rect 48958 278400 48964 278452
rect 49016 278440 49022 278452
rect 644658 278440 644664 278452
rect 49016 278412 644664 278440
rect 49016 278400 49022 278412
rect 644658 278400 644664 278412
rect 644716 278400 644722 278452
rect 64138 278264 64144 278316
rect 64196 278304 64202 278316
rect 661034 278304 661040 278316
rect 64196 278276 661040 278304
rect 64196 278264 64202 278276
rect 661034 278264 661040 278276
rect 661092 278264 661098 278316
rect 56226 278128 56232 278180
rect 56284 278168 56290 278180
rect 658274 278168 658280 278180
rect 56284 278140 658280 278168
rect 56284 278128 56290 278140
rect 658274 278128 658280 278140
rect 658332 278128 658338 278180
rect 49510 277992 49516 278044
rect 49568 278032 49574 278044
rect 659654 278032 659660 278044
rect 49568 278004 659660 278032
rect 49568 277992 49574 278004
rect 659654 277992 659660 278004
rect 659712 277992 659718 278044
rect 424686 277788 424692 277840
rect 424744 277828 424750 277840
rect 527726 277828 527732 277840
rect 424744 277800 527732 277828
rect 424744 277788 424750 277800
rect 527726 277788 527732 277800
rect 527784 277788 527790 277840
rect 413738 277652 413744 277704
rect 413796 277692 413802 277704
rect 510062 277692 510068 277704
rect 413796 277664 510068 277692
rect 413796 277652 413802 277664
rect 510062 277652 510068 277664
rect 510120 277652 510126 277704
rect 422202 277516 422208 277568
rect 422260 277556 422266 277568
rect 524506 277556 524512 277568
rect 422260 277528 524512 277556
rect 422260 277516 422266 277528
rect 524506 277516 524512 277528
rect 524564 277516 524570 277568
rect 467650 277380 467656 277432
rect 467708 277420 467714 277432
rect 570966 277420 570972 277432
rect 467708 277392 570972 277420
rect 467708 277380 467714 277392
rect 570966 277380 570972 277392
rect 571024 277380 571030 277432
rect 42334 277176 42340 277228
rect 42392 277216 42398 277228
rect 44082 277216 44088 277228
rect 42392 277188 44088 277216
rect 42392 277176 42398 277188
rect 44082 277176 44088 277188
rect 44140 277176 44146 277228
rect 457438 277176 457444 277228
rect 457496 277216 457502 277228
rect 563514 277216 563520 277228
rect 457496 277188 563520 277216
rect 457496 277176 457502 277188
rect 563514 277176 563520 277188
rect 563572 277176 563578 277228
rect 42334 277040 42340 277092
rect 42392 277080 42398 277092
rect 43990 277080 43996 277092
rect 42392 277052 43996 277080
rect 42392 277040 42398 277052
rect 43990 277040 43996 277052
rect 44048 277040 44054 277092
rect 409414 277040 409420 277092
rect 409472 277080 409478 277092
rect 499482 277080 499488 277092
rect 409472 277052 499488 277080
rect 409472 277040 409478 277052
rect 499482 277040 499488 277052
rect 499540 277040 499546 277092
rect 499758 277040 499764 277092
rect 499816 277080 499822 277092
rect 509050 277080 509056 277092
rect 499816 277052 509056 277080
rect 499816 277040 499822 277052
rect 509050 277040 509056 277052
rect 509108 277040 509114 277092
rect 509234 277040 509240 277092
rect 509292 277080 509298 277092
rect 601418 277080 601424 277092
rect 509292 277052 601424 277080
rect 509292 277040 509298 277052
rect 601418 277040 601424 277052
rect 601476 277040 601482 277092
rect 380710 276904 380716 276956
rect 380768 276944 380774 276956
rect 457162 276944 457168 276956
rect 380768 276916 457168 276944
rect 380768 276904 380774 276916
rect 457162 276904 457168 276916
rect 457220 276904 457226 276956
rect 472986 276904 472992 276956
rect 473044 276944 473050 276956
rect 606110 276944 606116 276956
rect 473044 276916 606116 276944
rect 473044 276904 473050 276916
rect 606110 276904 606116 276916
rect 606168 276904 606174 276956
rect 387334 276768 387340 276820
rect 387392 276808 387398 276820
rect 467834 276808 467840 276820
rect 387392 276780 467840 276808
rect 387392 276768 387398 276780
rect 467834 276768 467840 276780
rect 467892 276768 467898 276820
rect 469030 276768 469036 276820
rect 469088 276808 469094 276820
rect 599026 276808 599032 276820
rect 469088 276780 599032 276808
rect 469088 276768 469094 276780
rect 599026 276768 599032 276780
rect 599084 276768 599090 276820
rect 52270 276632 52276 276684
rect 52328 276672 52334 276684
rect 655514 276672 655520 276684
rect 52328 276644 655520 276672
rect 52328 276632 52334 276644
rect 655514 276632 655520 276644
rect 655572 276632 655578 276684
rect 402422 276496 402428 276548
rect 402480 276536 402486 276548
rect 492214 276536 492220 276548
rect 402480 276508 492220 276536
rect 402480 276496 402486 276508
rect 492214 276496 492220 276508
rect 492272 276496 492278 276548
rect 493318 276496 493324 276548
rect 493376 276536 493382 276548
rect 499390 276536 499396 276548
rect 493376 276508 499396 276536
rect 493376 276496 493382 276508
rect 499390 276496 499396 276508
rect 499448 276496 499454 276548
rect 499528 276496 499534 276548
rect 499586 276536 499592 276548
rect 616782 276536 616788 276548
rect 499586 276508 616788 276536
rect 499586 276496 499592 276508
rect 616782 276496 616788 276508
rect 616840 276496 616846 276548
rect 420362 276360 420368 276412
rect 420420 276400 420426 276412
rect 521010 276400 521016 276412
rect 420420 276372 521016 276400
rect 420420 276360 420426 276372
rect 521010 276360 521016 276372
rect 521068 276360 521074 276412
rect 442902 276224 442908 276276
rect 442960 276264 442966 276276
rect 557626 276264 557632 276276
rect 442960 276236 557632 276264
rect 442960 276224 442966 276236
rect 557626 276224 557632 276236
rect 557684 276224 557690 276276
rect 410886 276088 410892 276140
rect 410944 276128 410950 276140
rect 410944 276100 411392 276128
rect 410944 276088 410950 276100
rect 110782 275952 110788 276004
rect 110840 275992 110846 276004
rect 156690 275992 156696 276004
rect 110840 275964 156696 275992
rect 110840 275952 110846 275964
rect 156690 275952 156696 275964
rect 156748 275952 156754 276004
rect 171042 275952 171048 276004
rect 171100 275992 171106 276004
rect 171100 275964 174676 275992
rect 171100 275952 171106 275964
rect 107194 275816 107200 275868
rect 107252 275856 107258 275868
rect 153838 275856 153844 275868
rect 107252 275828 153844 275856
rect 107252 275816 107258 275828
rect 153838 275816 153844 275828
rect 153896 275816 153902 275868
rect 160462 275816 160468 275868
rect 160520 275856 160526 275868
rect 174446 275856 174452 275868
rect 160520 275828 174452 275856
rect 160520 275816 160526 275828
rect 174446 275816 174452 275828
rect 174504 275816 174510 275868
rect 174648 275856 174676 275964
rect 175826 275952 175832 276004
rect 175884 275992 175890 276004
rect 177850 275992 177856 276004
rect 175884 275964 177856 275992
rect 175884 275952 175890 275964
rect 177850 275952 177856 275964
rect 177908 275952 177914 276004
rect 317138 275952 317144 276004
rect 317196 275992 317202 276004
rect 319990 275992 319996 276004
rect 317196 275964 319996 275992
rect 317196 275952 317202 275964
rect 319990 275952 319996 275964
rect 320048 275952 320054 276004
rect 331214 275952 331220 276004
rect 331272 275992 331278 276004
rect 340138 275992 340144 276004
rect 331272 275964 340144 275992
rect 331272 275952 331278 275964
rect 340138 275952 340144 275964
rect 340196 275952 340202 276004
rect 342254 275952 342260 276004
rect 342312 275992 342318 276004
rect 350718 275992 350724 276004
rect 342312 275964 350724 275992
rect 342312 275952 342318 275964
rect 350718 275952 350724 275964
rect 350776 275952 350782 276004
rect 355318 275952 355324 276004
rect 355376 275992 355382 276004
rect 369670 275992 369676 276004
rect 355376 275964 369676 275992
rect 355376 275952 355382 275964
rect 369670 275952 369676 275964
rect 369728 275952 369734 276004
rect 369946 275952 369952 276004
rect 370004 275992 370010 276004
rect 407482 275992 407488 276004
rect 370004 275964 407488 275992
rect 370004 275952 370010 275964
rect 407482 275952 407488 275964
rect 407540 275952 407546 276004
rect 408218 275952 408224 276004
rect 408276 275992 408282 276004
rect 411364 275992 411392 276100
rect 436554 276088 436560 276140
rect 436612 276128 436618 276140
rect 436612 276100 436968 276128
rect 436612 276088 436618 276100
rect 421650 275992 421656 276004
rect 408276 275964 411300 275992
rect 411364 275964 421656 275992
rect 408276 275952 408282 275964
rect 175918 275856 175924 275868
rect 174648 275828 175924 275856
rect 175918 275816 175924 275828
rect 175976 275816 175982 275868
rect 305086 275816 305092 275868
rect 305144 275856 305150 275868
rect 316494 275856 316500 275868
rect 305144 275828 316500 275856
rect 305144 275816 305150 275828
rect 316494 275816 316500 275828
rect 316552 275816 316558 275868
rect 317322 275816 317328 275868
rect 317380 275856 317386 275868
rect 336550 275856 336556 275868
rect 317380 275828 336556 275856
rect 317380 275816 317386 275828
rect 336550 275816 336556 275828
rect 336608 275816 336614 275868
rect 343818 275816 343824 275868
rect 343876 275856 343882 275868
rect 354306 275856 354312 275868
rect 343876 275828 354312 275856
rect 343876 275816 343882 275828
rect 354306 275816 354312 275828
rect 354364 275816 354370 275868
rect 356882 275816 356888 275868
rect 356940 275856 356946 275868
rect 399202 275856 399208 275868
rect 356940 275828 399208 275856
rect 356940 275816 356946 275828
rect 399202 275816 399208 275828
rect 399260 275816 399266 275868
rect 400214 275816 400220 275868
rect 400272 275856 400278 275868
rect 411070 275856 411076 275868
rect 400272 275828 411076 275856
rect 400272 275816 400278 275828
rect 411070 275816 411076 275828
rect 411128 275816 411134 275868
rect 411272 275856 411300 275964
rect 421650 275952 421656 275964
rect 421708 275952 421714 276004
rect 421834 275952 421840 276004
rect 421892 275992 421898 276004
rect 425238 275992 425244 276004
rect 421892 275964 425244 275992
rect 421892 275952 421898 275964
rect 425238 275952 425244 275964
rect 425296 275952 425302 276004
rect 426066 275952 426072 276004
rect 426124 275992 426130 276004
rect 436738 275992 436744 276004
rect 426124 275964 436744 275992
rect 426124 275952 426130 275964
rect 436738 275952 436744 275964
rect 436796 275952 436802 276004
rect 436940 275992 436968 276100
rect 450722 276088 450728 276140
rect 450780 276128 450786 276140
rect 531222 276128 531228 276140
rect 450780 276100 531228 276128
rect 450780 276088 450786 276100
rect 531222 276088 531228 276100
rect 531280 276088 531286 276140
rect 465718 275992 465724 276004
rect 436940 275964 465724 275992
rect 465718 275952 465724 275964
rect 465776 275952 465782 276004
rect 465902 275952 465908 276004
rect 465960 275992 465966 276004
rect 466638 275992 466644 276004
rect 465960 275964 466644 275992
rect 465960 275952 465966 275964
rect 466638 275952 466644 275964
rect 466696 275952 466702 276004
rect 467098 275952 467104 276004
rect 467156 275992 467162 276004
rect 475562 275992 475568 276004
rect 467156 275964 475568 275992
rect 467156 275952 467162 275964
rect 475562 275952 475568 275964
rect 475620 275952 475626 276004
rect 475746 275952 475752 276004
rect 475804 275992 475810 276004
rect 480162 275992 480168 276004
rect 475804 275964 480168 275992
rect 475804 275952 475810 275964
rect 480162 275952 480168 275964
rect 480220 275952 480226 276004
rect 480346 275952 480352 276004
rect 480404 275992 480410 276004
rect 484302 275992 484308 276004
rect 480404 275964 484308 275992
rect 480404 275952 480410 275964
rect 484302 275952 484308 275964
rect 484360 275952 484366 276004
rect 485774 275952 485780 276004
rect 485832 275992 485838 276004
rect 489730 275992 489736 276004
rect 485832 275964 489736 275992
rect 485832 275952 485838 275964
rect 489730 275952 489736 275964
rect 489788 275952 489794 276004
rect 489914 275952 489920 276004
rect 489972 275992 489978 276004
rect 494974 275992 494980 276004
rect 489972 275964 494980 275992
rect 489972 275952 489978 275964
rect 494974 275952 494980 275964
rect 495032 275952 495038 276004
rect 495342 275952 495348 276004
rect 495400 275992 495406 276004
rect 504358 275992 504364 276004
rect 495400 275964 504364 275992
rect 495400 275952 495406 275964
rect 504358 275952 504364 275964
rect 504416 275952 504422 276004
rect 504726 275952 504732 276004
rect 504784 275992 504790 276004
rect 504784 275964 508912 275992
rect 504784 275952 504790 275964
rect 501782 275856 501788 275868
rect 411272 275828 501788 275856
rect 501782 275816 501788 275828
rect 501840 275816 501846 275868
rect 501966 275816 501972 275868
rect 502024 275856 502030 275868
rect 508682 275856 508688 275868
rect 502024 275828 508688 275856
rect 502024 275816 502030 275828
rect 508682 275816 508688 275828
rect 508740 275816 508746 275868
rect 508884 275856 508912 275964
rect 509050 275952 509056 276004
rect 509108 275992 509114 276004
rect 511994 275992 512000 276004
rect 509108 275964 512000 275992
rect 509108 275952 509114 275964
rect 511994 275952 512000 275964
rect 512052 275952 512058 276004
rect 512178 275952 512184 276004
rect 512236 275992 512242 276004
rect 516226 275992 516232 276004
rect 512236 275964 516232 275992
rect 512236 275952 512242 275964
rect 516226 275952 516232 275964
rect 516284 275952 516290 276004
rect 523678 275952 523684 276004
rect 523736 275992 523742 276004
rect 533338 275992 533344 276004
rect 523736 275964 533344 275992
rect 523736 275952 523742 275964
rect 533338 275952 533344 275964
rect 533396 275952 533402 276004
rect 616782 275952 616788 276004
rect 616840 275992 616846 276004
rect 635642 275992 635648 276004
rect 616840 275964 635648 275992
rect 616840 275952 616846 275964
rect 635642 275952 635648 275964
rect 635700 275952 635706 276004
rect 574186 275856 574192 275868
rect 508884 275828 574192 275856
rect 574186 275816 574192 275828
rect 574244 275816 574250 275868
rect 103698 275680 103704 275732
rect 103756 275720 103762 275732
rect 160554 275720 160560 275732
rect 103756 275692 160560 275720
rect 103756 275680 103762 275692
rect 160554 275680 160560 275692
rect 160612 275680 160618 275732
rect 174630 275680 174636 275732
rect 174688 275720 174694 275732
rect 197538 275720 197544 275732
rect 174688 275692 197544 275720
rect 174688 275680 174694 275692
rect 197538 275680 197544 275692
rect 197596 275680 197602 275732
rect 199470 275680 199476 275732
rect 199528 275720 199534 275732
rect 210878 275720 210884 275732
rect 199528 275692 210884 275720
rect 199528 275680 199534 275692
rect 210878 275680 210884 275692
rect 210936 275680 210942 275732
rect 297266 275680 297272 275732
rect 297324 275720 297330 275732
rect 311710 275720 311716 275732
rect 297324 275692 311716 275720
rect 297324 275680 297330 275692
rect 311710 275680 311716 275692
rect 311768 275680 311774 275732
rect 319990 275680 319996 275732
rect 320048 275720 320054 275732
rect 343634 275720 343640 275732
rect 320048 275692 343640 275720
rect 320048 275680 320054 275692
rect 343634 275680 343640 275692
rect 343692 275680 343698 275732
rect 345382 275680 345388 275732
rect 345440 275720 345446 275732
rect 370866 275720 370872 275732
rect 345440 275692 370872 275720
rect 345440 275680 345446 275692
rect 370866 275680 370872 275692
rect 370924 275680 370930 275732
rect 374178 275680 374184 275732
rect 374236 275720 374242 275732
rect 393314 275720 393320 275732
rect 374236 275692 393320 275720
rect 374236 275680 374242 275692
rect 393314 275680 393320 275692
rect 393372 275680 393378 275732
rect 395430 275680 395436 275732
rect 395488 275720 395494 275732
rect 399662 275720 399668 275732
rect 395488 275692 399668 275720
rect 395488 275680 395494 275692
rect 399662 275680 399668 275692
rect 399720 275680 399726 275732
rect 399846 275680 399852 275732
rect 399904 275720 399910 275732
rect 400582 275720 400588 275732
rect 399904 275692 400588 275720
rect 399904 275680 399910 275692
rect 400582 275680 400588 275692
rect 400640 275680 400646 275732
rect 400766 275680 400772 275732
rect 400824 275720 400830 275732
rect 480806 275720 480812 275732
rect 400824 275692 480812 275720
rect 400824 275680 400830 275692
rect 480806 275680 480812 275692
rect 480864 275680 480870 275732
rect 480990 275680 480996 275732
rect 481048 275720 481054 275732
rect 487890 275720 487896 275732
rect 481048 275692 487896 275720
rect 481048 275680 481054 275692
rect 487890 275680 487896 275692
rect 487948 275680 487954 275732
rect 488074 275680 488080 275732
rect 488132 275720 488138 275732
rect 489868 275720 489874 275732
rect 488132 275692 489874 275720
rect 488132 275680 488138 275692
rect 489868 275680 489874 275692
rect 489926 275680 489932 275732
rect 490006 275680 490012 275732
rect 490064 275720 490070 275732
rect 604914 275720 604920 275732
rect 490064 275692 604920 275720
rect 490064 275680 490070 275692
rect 604914 275680 604920 275692
rect 604972 275680 604978 275732
rect 610066 275680 610072 275732
rect 610124 275720 610130 275732
rect 614390 275720 614396 275732
rect 610124 275692 614396 275720
rect 610124 275680 610130 275692
rect 614390 275680 614396 275692
rect 614448 275680 614454 275732
rect 74074 275544 74080 275596
rect 74132 275584 74138 275596
rect 77754 275584 77760 275596
rect 74132 275556 77760 275584
rect 74132 275544 74138 275556
rect 77754 275544 77760 275556
rect 77812 275544 77818 275596
rect 85942 275544 85948 275596
rect 86000 275584 86006 275596
rect 149054 275584 149060 275596
rect 86000 275556 149060 275584
rect 86000 275544 86006 275556
rect 149054 275544 149060 275556
rect 149112 275544 149118 275596
rect 149790 275544 149796 275596
rect 149848 275584 149854 275596
rect 179966 275584 179972 275596
rect 149848 275556 179972 275584
rect 149848 275544 149854 275556
rect 179966 275544 179972 275556
rect 180024 275544 180030 275596
rect 181714 275544 181720 275596
rect 181772 275584 181778 275596
rect 207014 275584 207020 275596
rect 181772 275556 207020 275584
rect 181772 275544 181778 275556
rect 207014 275544 207020 275556
rect 207072 275544 207078 275596
rect 282914 275544 282920 275596
rect 282972 275584 282978 275596
rect 285766 275584 285772 275596
rect 282972 275556 285772 275584
rect 282972 275544 282978 275556
rect 285766 275544 285772 275556
rect 285824 275544 285830 275596
rect 302510 275544 302516 275596
rect 302568 275584 302574 275596
rect 318794 275584 318800 275596
rect 302568 275556 318800 275584
rect 302568 275544 302574 275556
rect 318794 275544 318800 275556
rect 318852 275544 318858 275596
rect 329190 275544 329196 275596
rect 329248 275584 329254 275596
rect 374362 275584 374368 275596
rect 329248 275556 374368 275584
rect 329248 275544 329254 275556
rect 374362 275544 374368 275556
rect 374420 275544 374426 275596
rect 374638 275544 374644 275596
rect 374696 275584 374702 275596
rect 379146 275584 379152 275596
rect 374696 275556 379152 275584
rect 374696 275544 374702 275556
rect 379146 275544 379152 275556
rect 379204 275544 379210 275596
rect 380894 275544 380900 275596
rect 380952 275584 380958 275596
rect 386414 275584 386420 275596
rect 380952 275556 386420 275584
rect 380952 275544 380958 275556
rect 386414 275544 386420 275556
rect 386472 275544 386478 275596
rect 391566 275544 391572 275596
rect 391624 275584 391630 275596
rect 473446 275584 473452 275596
rect 391624 275556 473452 275584
rect 391624 275544 391630 275556
rect 473446 275544 473452 275556
rect 473504 275544 473510 275596
rect 473998 275544 474004 275596
rect 474056 275584 474062 275596
rect 475194 275584 475200 275596
rect 474056 275556 475200 275584
rect 474056 275544 474062 275556
rect 475194 275544 475200 275556
rect 475252 275544 475258 275596
rect 475378 275544 475384 275596
rect 475436 275584 475442 275596
rect 475436 275556 494836 275584
rect 475436 275544 475442 275556
rect 213914 275516 213920 275528
rect 209746 275488 213920 275516
rect 68186 275408 68192 275460
rect 68244 275448 68250 275460
rect 135254 275448 135260 275460
rect 68244 275420 135260 275448
rect 68244 275408 68250 275420
rect 135254 275408 135260 275420
rect 135312 275408 135318 275460
rect 136818 275408 136824 275460
rect 136876 275448 136882 275460
rect 152734 275448 152740 275460
rect 136876 275420 152740 275448
rect 136876 275408 136882 275420
rect 152734 275408 152740 275420
rect 152792 275408 152798 275460
rect 153286 275408 153292 275460
rect 153344 275448 153350 275460
rect 185578 275448 185584 275460
rect 153344 275420 185584 275448
rect 153344 275408 153350 275420
rect 185578 275408 185584 275420
rect 185636 275408 185642 275460
rect 188798 275408 188804 275460
rect 188856 275448 188862 275460
rect 209746 275448 209774 275488
rect 213914 275476 213920 275488
rect 213972 275476 213978 275528
rect 188856 275420 209774 275448
rect 188856 275408 188862 275420
rect 236086 275408 236092 275460
rect 236144 275448 236150 275460
rect 242250 275448 242256 275460
rect 236144 275420 242256 275448
rect 236144 275408 236150 275420
rect 242250 275408 242256 275420
rect 242308 275408 242314 275460
rect 285674 275408 285680 275460
rect 285732 275448 285738 275460
rect 303430 275448 303436 275460
rect 285732 275420 303436 275448
rect 285732 275408 285738 275420
rect 303430 275408 303436 275420
rect 303488 275408 303494 275460
rect 311066 275408 311072 275460
rect 311124 275448 311130 275460
rect 329466 275448 329472 275460
rect 311124 275420 329472 275448
rect 311124 275408 311130 275420
rect 329466 275408 329472 275420
rect 329524 275408 329530 275460
rect 333606 275408 333612 275460
rect 333664 275448 333670 275460
rect 381538 275448 381544 275460
rect 333664 275420 381544 275448
rect 333664 275408 333670 275420
rect 381538 275408 381544 275420
rect 381596 275408 381602 275460
rect 382642 275408 382648 275460
rect 382700 275448 382706 275460
rect 388622 275448 388628 275460
rect 382700 275420 388628 275448
rect 382700 275408 382706 275420
rect 388622 275408 388628 275420
rect 388680 275408 388686 275460
rect 392118 275448 392124 275460
rect 389146 275420 392124 275448
rect 210050 275340 210056 275392
rect 210108 275380 210114 275392
rect 226426 275380 226432 275392
rect 210108 275352 226432 275380
rect 210108 275340 210114 275352
rect 226426 275340 226432 275352
rect 226484 275340 226490 275392
rect 70578 275272 70584 275324
rect 70636 275312 70642 275324
rect 139302 275312 139308 275324
rect 70636 275284 139308 275312
rect 70636 275272 70642 275284
rect 139302 275272 139308 275284
rect 139360 275272 139366 275324
rect 152182 275272 152188 275324
rect 152240 275312 152246 275324
rect 162578 275312 162584 275324
rect 152240 275284 162584 275312
rect 152240 275272 152246 275284
rect 162578 275272 162584 275284
rect 162636 275272 162642 275324
rect 167546 275272 167552 275324
rect 167604 275312 167610 275324
rect 200022 275312 200028 275324
rect 167604 275284 200028 275312
rect 167604 275272 167610 275284
rect 200022 275272 200028 275284
rect 200080 275272 200086 275324
rect 227806 275272 227812 275324
rect 227864 275312 227870 275324
rect 237374 275312 237380 275324
rect 227864 275284 237380 275312
rect 227864 275272 227870 275284
rect 237374 275272 237380 275284
rect 237432 275272 237438 275324
rect 238478 275272 238484 275324
rect 238536 275312 238542 275324
rect 243722 275312 243728 275324
rect 238536 275284 243728 275312
rect 238536 275272 238542 275284
rect 243722 275272 243728 275284
rect 243780 275272 243786 275324
rect 265894 275272 265900 275324
rect 265952 275312 265958 275324
rect 271506 275312 271512 275324
rect 265952 275284 271512 275312
rect 265952 275272 265958 275284
rect 271506 275272 271512 275284
rect 271564 275272 271570 275324
rect 278406 275272 278412 275324
rect 278464 275312 278470 275324
rect 292850 275312 292856 275324
rect 278464 275284 292856 275312
rect 278464 275272 278470 275284
rect 292850 275272 292856 275284
rect 292908 275272 292914 275324
rect 295334 275272 295340 275324
rect 295392 275312 295398 275324
rect 299934 275312 299940 275324
rect 295392 275284 299940 275312
rect 295392 275272 295398 275284
rect 299934 275272 299940 275284
rect 299992 275272 299998 275324
rect 301130 275272 301136 275324
rect 301188 275312 301194 275324
rect 322382 275312 322388 275324
rect 301188 275284 322388 275312
rect 301188 275272 301194 275284
rect 322382 275272 322388 275284
rect 322440 275272 322446 275324
rect 322566 275272 322572 275324
rect 322624 275312 322630 275324
rect 333054 275312 333060 275324
rect 322624 275284 333060 275312
rect 322624 275272 322630 275284
rect 333054 275272 333060 275284
rect 333112 275272 333118 275324
rect 340230 275272 340236 275324
rect 340288 275312 340294 275324
rect 389146 275312 389174 275420
rect 392118 275408 392124 275420
rect 392176 275408 392182 275460
rect 396718 275408 396724 275460
rect 396776 275448 396782 275460
rect 400398 275448 400404 275460
rect 396776 275420 400404 275448
rect 396776 275408 396782 275420
rect 400398 275408 400404 275420
rect 400456 275408 400462 275460
rect 400582 275408 400588 275460
rect 400640 275448 400646 275460
rect 480162 275448 480168 275460
rect 400640 275420 480168 275448
rect 400640 275408 400646 275420
rect 480162 275408 480168 275420
rect 480220 275408 480226 275460
rect 480346 275408 480352 275460
rect 480404 275448 480410 275460
rect 484854 275448 484860 275460
rect 480404 275420 484860 275448
rect 480404 275408 480410 275420
rect 484854 275408 484860 275420
rect 484912 275408 484918 275460
rect 485038 275408 485044 275460
rect 485096 275448 485102 275460
rect 485096 275420 494560 275448
rect 485096 275408 485102 275420
rect 494532 275380 494560 275420
rect 494532 275352 494744 275380
rect 340288 275284 389174 275312
rect 340288 275272 340294 275284
rect 391934 275272 391940 275324
rect 391992 275312 391998 275324
rect 396902 275312 396908 275324
rect 391992 275284 396908 275312
rect 391992 275272 391998 275284
rect 396902 275272 396908 275284
rect 396960 275272 396966 275324
rect 397454 275272 397460 275324
rect 397512 275312 397518 275324
rect 397512 275284 414704 275312
rect 397512 275272 397518 275284
rect 211246 275204 211252 275256
rect 211304 275244 211310 275256
rect 212442 275244 212448 275256
rect 211304 275216 212448 275244
rect 211304 275204 211310 275216
rect 212442 275204 212448 275216
rect 212500 275204 212506 275256
rect 113174 275136 113180 275188
rect 113232 275176 113238 275188
rect 142982 275176 142988 275188
rect 113232 275148 142988 275176
rect 113232 275136 113238 275148
rect 142982 275136 142988 275148
rect 143040 275136 143046 275188
rect 156874 275136 156880 275188
rect 156932 275176 156938 275188
rect 166166 275176 166172 275188
rect 156932 275148 166172 275176
rect 156932 275136 156938 275148
rect 166166 275136 166172 275148
rect 166224 275136 166230 275188
rect 245562 275136 245568 275188
rect 245620 275176 245626 275188
rect 246298 275176 246304 275188
rect 245620 275148 246304 275176
rect 245620 275136 245626 275148
rect 246298 275136 246304 275148
rect 246356 275136 246362 275188
rect 350534 275136 350540 275188
rect 350592 275176 350598 275188
rect 357894 275176 357900 275188
rect 350592 275148 357900 275176
rect 350592 275136 350598 275148
rect 357894 275136 357900 275148
rect 357952 275136 357958 275188
rect 365622 275136 365628 275188
rect 365680 275176 365686 275188
rect 375558 275176 375564 275188
rect 365680 275148 375564 275176
rect 365680 275136 365686 275148
rect 375558 275136 375564 275148
rect 375616 275136 375622 275188
rect 386414 275136 386420 275188
rect 386472 275176 386478 275188
rect 414382 275176 414388 275188
rect 386472 275148 414388 275176
rect 386472 275136 386478 275148
rect 414382 275136 414388 275148
rect 414440 275136 414446 275188
rect 414676 275176 414704 275284
rect 415210 275272 415216 275324
rect 415268 275312 415274 275324
rect 418338 275312 418344 275324
rect 415268 275284 418344 275312
rect 415268 275272 415274 275284
rect 418338 275272 418344 275284
rect 418396 275272 418402 275324
rect 418522 275272 418528 275324
rect 418580 275312 418586 275324
rect 421834 275312 421840 275324
rect 418580 275284 421840 275312
rect 418580 275272 418586 275284
rect 421834 275272 421840 275284
rect 421892 275272 421898 275324
rect 422018 275272 422024 275324
rect 422076 275312 422082 275324
rect 422938 275312 422944 275324
rect 422076 275284 422944 275312
rect 422076 275272 422082 275284
rect 422938 275272 422944 275284
rect 422996 275272 423002 275324
rect 465534 275312 465540 275324
rect 423140 275284 465540 275312
rect 423140 275176 423168 275284
rect 465534 275272 465540 275284
rect 465592 275272 465598 275324
rect 465718 275272 465724 275324
rect 465776 275312 465782 275324
rect 475378 275312 475384 275324
rect 465776 275284 475384 275312
rect 465776 275272 465782 275284
rect 475378 275272 475384 275284
rect 475436 275272 475442 275324
rect 475562 275272 475568 275324
rect 475620 275312 475626 275324
rect 475620 275284 490052 275312
rect 475620 275272 475626 275284
rect 414676 275148 423168 275176
rect 423306 275136 423312 275188
rect 423364 275176 423370 275188
rect 427078 275176 427084 275188
rect 423364 275148 427084 275176
rect 423364 275136 423370 275148
rect 427078 275136 427084 275148
rect 427136 275136 427142 275188
rect 427262 275136 427268 275188
rect 427320 275176 427326 275188
rect 431126 275176 431132 275188
rect 427320 275148 431132 275176
rect 427320 275136 427326 275148
rect 431126 275136 431132 275148
rect 431184 275136 431190 275188
rect 431310 275136 431316 275188
rect 431368 275176 431374 275188
rect 436554 275176 436560 275188
rect 431368 275148 436560 275176
rect 431368 275136 431374 275148
rect 436554 275136 436560 275148
rect 436612 275136 436618 275188
rect 436738 275136 436744 275188
rect 436796 275176 436802 275188
rect 485038 275176 485044 275188
rect 436796 275148 485044 275176
rect 436796 275136 436802 275148
rect 485038 275136 485044 275148
rect 485096 275136 485102 275188
rect 485222 275136 485228 275188
rect 485280 275176 485286 275188
rect 489868 275176 489874 275188
rect 485280 275148 489874 275176
rect 485280 275136 485286 275148
rect 489868 275136 489874 275148
rect 489926 275136 489932 275188
rect 490024 275176 490052 275284
rect 494514 275176 494520 275188
rect 490024 275148 494520 275176
rect 494514 275136 494520 275148
rect 494572 275136 494578 275188
rect 494716 275176 494744 275352
rect 494808 275312 494836 275556
rect 494974 275544 494980 275596
rect 495032 275584 495038 275596
rect 611998 275584 612004 275596
rect 495032 275556 612004 275584
rect 495032 275544 495038 275556
rect 611998 275544 612004 275556
rect 612056 275544 612062 275596
rect 494974 275408 494980 275460
rect 495032 275448 495038 275460
rect 498562 275448 498568 275460
rect 495032 275420 498568 275448
rect 495032 275408 495038 275420
rect 498562 275408 498568 275420
rect 498620 275408 498626 275460
rect 498746 275408 498752 275460
rect 498804 275448 498810 275460
rect 498804 275420 502196 275448
rect 498804 275408 498810 275420
rect 501966 275312 501972 275324
rect 494808 275284 501972 275312
rect 501966 275272 501972 275284
rect 502024 275272 502030 275324
rect 502168 275312 502196 275420
rect 504358 275408 504364 275460
rect 504416 275448 504422 275460
rect 640426 275448 640432 275460
rect 504416 275420 640432 275448
rect 504416 275408 504422 275420
rect 640426 275408 640432 275420
rect 640484 275408 640490 275460
rect 648522 275312 648528 275324
rect 502168 275284 648528 275312
rect 648522 275272 648528 275284
rect 648580 275272 648586 275324
rect 523494 275176 523500 275188
rect 494716 275148 523500 275176
rect 523494 275136 523500 275148
rect 523552 275136 523558 275188
rect 537570 275176 537576 275188
rect 523696 275148 537576 275176
rect 194686 275068 194692 275120
rect 194744 275108 194750 275120
rect 195882 275108 195888 275120
rect 194744 275080 195888 275108
rect 194744 275068 194750 275080
rect 195882 275068 195888 275080
rect 195940 275068 195946 275120
rect 378778 275068 378784 275120
rect 378836 275108 378842 275120
rect 386230 275108 386236 275120
rect 378836 275080 386236 275108
rect 378836 275068 378842 275080
rect 386230 275068 386236 275080
rect 386288 275068 386294 275120
rect 142706 275000 142712 275052
rect 142764 275040 142770 275052
rect 169754 275040 169760 275052
rect 142764 275012 169760 275040
rect 142764 275000 142770 275012
rect 169754 275000 169760 275012
rect 169812 275000 169818 275052
rect 249058 275000 249064 275052
rect 249116 275040 249122 275052
rect 250346 275040 250352 275052
rect 249116 275012 250352 275040
rect 249116 275000 249122 275012
rect 250346 275000 250352 275012
rect 250404 275000 250410 275052
rect 386414 275000 386420 275052
rect 386472 275040 386478 275052
rect 414566 275040 414572 275052
rect 386472 275012 414572 275040
rect 386472 275000 386478 275012
rect 414566 275000 414572 275012
rect 414624 275000 414630 275052
rect 415486 275000 415492 275052
rect 415544 275040 415550 275052
rect 501782 275040 501788 275052
rect 415544 275012 501788 275040
rect 415544 275000 415550 275012
rect 501782 275000 501788 275012
rect 501840 275000 501846 275052
rect 501966 275000 501972 275052
rect 502024 275040 502030 275052
rect 523696 275040 523724 275148
rect 537570 275136 537576 275148
rect 537628 275136 537634 275188
rect 537754 275136 537760 275188
rect 537812 275176 537818 275188
rect 552934 275176 552940 275188
rect 537812 275148 552940 275176
rect 537812 275136 537818 275148
rect 552934 275136 552940 275148
rect 552992 275136 552998 275188
rect 556154 275136 556160 275188
rect 556212 275176 556218 275188
rect 565906 275176 565912 275188
rect 556212 275148 565912 275176
rect 556212 275136 556218 275148
rect 565906 275136 565912 275148
rect 565964 275136 565970 275188
rect 570966 275136 570972 275188
rect 571024 275176 571030 275188
rect 596082 275176 596088 275188
rect 571024 275148 596088 275176
rect 571024 275136 571030 275148
rect 596082 275136 596088 275148
rect 596140 275136 596146 275188
rect 597462 275136 597468 275188
rect 597520 275176 597526 275188
rect 610802 275176 610808 275188
rect 597520 275148 610808 275176
rect 597520 275136 597526 275148
rect 610802 275136 610808 275148
rect 610860 275136 610866 275188
rect 633342 275040 633348 275052
rect 502024 275012 523724 275040
rect 528526 275012 633348 275040
rect 502024 275000 502030 275012
rect 71774 274932 71780 274984
rect 71832 274972 71838 274984
rect 73798 274972 73804 274984
rect 71832 274944 73804 274972
rect 71832 274932 71838 274944
rect 73798 274932 73804 274944
rect 73856 274932 73862 274984
rect 81250 274932 81256 274984
rect 81308 274972 81314 274984
rect 86218 274972 86224 274984
rect 81308 274944 86224 274972
rect 81308 274932 81314 274944
rect 86218 274932 86224 274944
rect 86276 274932 86282 274984
rect 186406 274932 186412 274984
rect 186464 274972 186470 274984
rect 188062 274972 188068 274984
rect 186464 274944 188068 274972
rect 186464 274932 186470 274944
rect 188062 274932 188068 274944
rect 188120 274932 188126 274984
rect 207750 274932 207756 274984
rect 207808 274972 207814 274984
rect 208394 274972 208400 274984
rect 207808 274944 208400 274972
rect 207808 274932 207814 274944
rect 208394 274932 208400 274944
rect 208452 274932 208458 274984
rect 135622 274864 135628 274916
rect 135680 274904 135686 274916
rect 158714 274904 158720 274916
rect 135680 274876 158720 274904
rect 135680 274864 135686 274876
rect 158714 274864 158720 274876
rect 158772 274864 158778 274916
rect 376110 274864 376116 274916
rect 376168 274904 376174 274916
rect 403986 274904 403992 274916
rect 376168 274876 403992 274904
rect 376168 274864 376174 274876
rect 403986 274864 403992 274876
rect 404044 274864 404050 274916
rect 404170 274864 404176 274916
rect 404228 274904 404234 274916
rect 412266 274904 412272 274916
rect 404228 274876 412272 274904
rect 404228 274864 404234 274876
rect 412266 274864 412272 274876
rect 412324 274864 412330 274916
rect 414382 274864 414388 274916
rect 414440 274904 414446 274916
rect 418154 274904 418160 274916
rect 414440 274876 418160 274904
rect 414440 274864 414446 274876
rect 418154 274864 418160 274876
rect 418212 274864 418218 274916
rect 418338 274864 418344 274916
rect 418396 274904 418402 274916
rect 421926 274904 421932 274916
rect 418396 274876 421932 274904
rect 418396 274864 418402 274876
rect 421926 274864 421932 274876
rect 421984 274864 421990 274916
rect 422294 274864 422300 274916
rect 422352 274904 422358 274916
rect 422352 274876 423076 274904
rect 422352 274864 422358 274876
rect 214834 274796 214840 274848
rect 214892 274836 214898 274848
rect 221734 274836 221740 274848
rect 214892 274808 221740 274836
rect 214892 274796 214898 274808
rect 221734 274796 221740 274808
rect 221792 274796 221798 274848
rect 338850 274728 338856 274780
rect 338908 274768 338914 274780
rect 344830 274768 344836 274780
rect 338908 274740 344836 274768
rect 338908 274728 338914 274740
rect 344830 274728 344836 274740
rect 344888 274728 344894 274780
rect 353386 274728 353392 274780
rect 353444 274768 353450 274780
rect 355502 274768 355508 274780
rect 353444 274740 355508 274768
rect 353444 274728 353450 274740
rect 355502 274728 355508 274740
rect 355560 274728 355566 274780
rect 358722 274728 358728 274780
rect 358780 274768 358786 274780
rect 364978 274768 364984 274780
rect 358780 274740 364984 274768
rect 358780 274728 358786 274740
rect 364978 274728 364984 274740
rect 365036 274728 365042 274780
rect 365438 274728 365444 274780
rect 365496 274768 365502 274780
rect 382642 274768 382648 274780
rect 365496 274740 382648 274768
rect 365496 274728 365502 274740
rect 382642 274728 382648 274740
rect 382700 274728 382706 274780
rect 382826 274728 382832 274780
rect 382884 274768 382890 274780
rect 386414 274768 386420 274780
rect 382884 274740 386420 274768
rect 382884 274728 382890 274740
rect 386414 274728 386420 274740
rect 386472 274728 386478 274780
rect 388070 274728 388076 274780
rect 388128 274768 388134 274780
rect 408678 274768 408684 274780
rect 388128 274740 408684 274768
rect 388128 274728 388134 274740
rect 408678 274728 408684 274740
rect 408736 274728 408742 274780
rect 411254 274728 411260 274780
rect 411312 274768 411318 274780
rect 415762 274768 415768 274780
rect 411312 274740 415768 274768
rect 411312 274728 411318 274740
rect 415762 274728 415768 274740
rect 415820 274728 415826 274780
rect 417970 274728 417976 274780
rect 418028 274768 418034 274780
rect 422662 274768 422668 274780
rect 418028 274740 422668 274768
rect 418028 274728 418034 274740
rect 422662 274728 422668 274740
rect 422720 274728 422726 274780
rect 423048 274768 423076 274876
rect 423214 274864 423220 274916
rect 423272 274904 423278 274916
rect 509188 274904 509194 274916
rect 423272 274876 509194 274904
rect 423272 274864 423278 274876
rect 509188 274864 509194 274876
rect 509246 274864 509252 274916
rect 509326 274864 509332 274916
rect 509384 274904 509390 274916
rect 513926 274904 513932 274916
rect 509384 274876 513932 274904
rect 509384 274864 509390 274876
rect 513926 274864 513932 274876
rect 513984 274864 513990 274916
rect 514110 274864 514116 274916
rect 514168 274904 514174 274916
rect 528526 274904 528554 275012
rect 633342 275000 633348 275012
rect 633400 275000 633406 275052
rect 514168 274876 528554 274904
rect 514168 274864 514174 274876
rect 531222 274864 531228 274916
rect 531280 274904 531286 274916
rect 570690 274904 570696 274916
rect 531280 274876 570696 274904
rect 531280 274864 531286 274876
rect 570690 274864 570696 274876
rect 570748 274864 570754 274916
rect 619634 274796 619640 274848
rect 619692 274836 619698 274848
rect 623866 274836 623872 274848
rect 619692 274808 623872 274836
rect 619692 274796 619698 274808
rect 623866 274796 623872 274808
rect 623924 274796 623930 274848
rect 523310 274768 523316 274780
rect 423048 274740 523316 274768
rect 523310 274728 523316 274740
rect 523368 274728 523374 274780
rect 523494 274728 523500 274780
rect 523552 274768 523558 274780
rect 530486 274768 530492 274780
rect 523552 274740 530492 274768
rect 523552 274728 523558 274740
rect 530486 274728 530492 274740
rect 530544 274728 530550 274780
rect 533338 274728 533344 274780
rect 533396 274768 533402 274780
rect 549346 274768 549352 274780
rect 533396 274740 549352 274768
rect 533396 274728 533402 274740
rect 549346 274728 549352 274740
rect 549404 274728 549410 274780
rect 552842 274728 552848 274780
rect 552900 274768 552906 274780
rect 556430 274768 556436 274780
rect 552900 274740 556436 274768
rect 552900 274728 552906 274740
rect 556430 274728 556436 274740
rect 556488 274728 556494 274780
rect 89530 274660 89536 274712
rect 89588 274700 89594 274712
rect 92474 274700 92480 274712
rect 89588 274672 92480 274700
rect 89588 274660 89594 274672
rect 92474 274660 92480 274672
rect 92532 274660 92538 274712
rect 161566 274660 161572 274712
rect 161624 274700 161630 274712
rect 163682 274700 163688 274712
rect 161624 274672 163688 274700
rect 161624 274660 161630 274672
rect 163682 274660 163688 274672
rect 163740 274660 163746 274712
rect 163958 274660 163964 274712
rect 164016 274700 164022 274712
rect 167638 274700 167644 274712
rect 164016 274672 167644 274700
rect 164016 274660 164022 274672
rect 167638 274660 167644 274672
rect 167696 274660 167702 274712
rect 178126 274660 178132 274712
rect 178184 274700 178190 274712
rect 179322 274700 179328 274712
rect 178184 274672 179328 274700
rect 178184 274660 178190 274672
rect 179322 274660 179328 274672
rect 179380 274660 179386 274712
rect 185210 274660 185216 274712
rect 185268 274700 185274 274712
rect 186958 274700 186964 274712
rect 185268 274672 186964 274700
rect 185268 274660 185274 274672
rect 186958 274660 186964 274672
rect 187016 274660 187022 274712
rect 241974 274660 241980 274712
rect 242032 274700 242038 274712
rect 246022 274700 246028 274712
rect 242032 274672 246028 274700
rect 242032 274660 242038 274672
rect 246022 274660 246028 274672
rect 246080 274660 246086 274712
rect 246758 274660 246764 274712
rect 246816 274700 246822 274712
rect 248874 274700 248880 274712
rect 246816 274672 248880 274700
rect 246816 274660 246822 274672
rect 248874 274660 248880 274672
rect 248932 274660 248938 274712
rect 271138 274660 271144 274712
rect 271196 274700 271202 274712
rect 276290 274700 276296 274712
rect 271196 274672 276296 274700
rect 271196 274660 271202 274672
rect 276290 274660 276296 274672
rect 276348 274660 276354 274712
rect 276658 274660 276664 274712
rect 276716 274700 276722 274712
rect 278682 274700 278688 274712
rect 276716 274672 278688 274700
rect 276716 274660 276722 274672
rect 278682 274660 278688 274672
rect 278740 274660 278746 274712
rect 280706 274660 280712 274712
rect 280764 274700 280770 274712
rect 283374 274700 283380 274712
rect 280764 274672 283380 274700
rect 280764 274660 280770 274672
rect 283374 274660 283380 274672
rect 283432 274660 283438 274712
rect 293218 274660 293224 274712
rect 293276 274700 293282 274712
rect 294046 274700 294052 274712
rect 293276 274672 294052 274700
rect 293276 274660 293282 274672
rect 294046 274660 294052 274672
rect 294104 274660 294110 274712
rect 319622 274660 319628 274712
rect 319680 274700 319686 274712
rect 327074 274700 327080 274712
rect 319680 274672 327080 274700
rect 319680 274660 319686 274672
rect 327074 274660 327080 274672
rect 327132 274660 327138 274712
rect 614758 274660 614764 274712
rect 614816 274700 614822 274712
rect 616598 274700 616604 274712
rect 614816 274672 616604 274700
rect 614816 274660 614822 274672
rect 616598 274660 616604 274672
rect 616656 274660 616662 274712
rect 618898 274660 618904 274712
rect 618956 274700 618962 274712
rect 620278 274700 620284 274712
rect 618956 274672 620284 274700
rect 618956 274660 618962 274672
rect 620278 274660 620284 274672
rect 620336 274660 620342 274712
rect 643738 274660 643744 274712
rect 643796 274700 643802 274712
rect 645118 274700 645124 274712
rect 643796 274672 645124 274700
rect 643796 274660 643802 274672
rect 645118 274660 645124 274672
rect 645176 274660 645182 274712
rect 42242 274592 42248 274644
rect 42300 274632 42306 274644
rect 47026 274632 47032 274644
rect 42300 274604 47032 274632
rect 42300 274592 42306 274604
rect 47026 274592 47032 274604
rect 47084 274592 47090 274644
rect 119338 274632 119344 274644
rect 103486 274604 119344 274632
rect 96614 274456 96620 274508
rect 96672 274496 96678 274508
rect 103486 274496 103514 274604
rect 119338 274592 119344 274604
rect 119396 274592 119402 274644
rect 120258 274592 120264 274644
rect 120316 274632 120322 274644
rect 161428 274632 161434 274644
rect 120316 274604 161434 274632
rect 120316 274592 120322 274604
rect 161428 274592 161434 274604
rect 161486 274592 161492 274644
rect 329650 274592 329656 274644
rect 329708 274632 329714 274644
rect 365622 274632 365628 274644
rect 329708 274604 365628 274632
rect 329708 274592 329714 274604
rect 365622 274592 365628 274604
rect 365680 274592 365686 274644
rect 390278 274592 390284 274644
rect 390336 274632 390342 274644
rect 470226 274632 470232 274644
rect 390336 274604 470232 274632
rect 390336 274592 390342 274604
rect 470226 274592 470232 274604
rect 470284 274592 470290 274644
rect 470410 274592 470416 274644
rect 470468 274632 470474 274644
rect 475378 274632 475384 274644
rect 470468 274604 475384 274632
rect 470468 274592 470474 274604
rect 475378 274592 475384 274604
rect 475436 274592 475442 274644
rect 475562 274592 475568 274644
rect 475620 274632 475626 274644
rect 479610 274632 479616 274644
rect 475620 274604 479616 274632
rect 475620 274592 475626 274604
rect 479610 274592 479616 274604
rect 479668 274592 479674 274644
rect 479794 274592 479800 274644
rect 479852 274632 479858 274644
rect 597462 274632 597468 274644
rect 479852 274604 597468 274632
rect 479852 274592 479858 274604
rect 597462 274592 597468 274604
rect 597520 274592 597526 274644
rect 96672 274468 103514 274496
rect 96672 274456 96678 274468
rect 119062 274456 119068 274508
rect 119120 274496 119126 274508
rect 168466 274496 168472 274508
rect 119120 274468 168472 274496
rect 119120 274456 119126 274468
rect 168466 274456 168472 274468
rect 168524 274456 168530 274508
rect 169754 274456 169760 274508
rect 169812 274496 169818 274508
rect 185118 274496 185124 274508
rect 169812 274468 185124 274496
rect 169812 274456 169818 274468
rect 185118 274456 185124 274468
rect 185176 274456 185182 274508
rect 294598 274456 294604 274508
rect 294656 274496 294662 274508
rect 307018 274496 307024 274508
rect 294656 274468 307024 274496
rect 294656 274456 294662 274468
rect 307018 274456 307024 274468
rect 307076 274456 307082 274508
rect 318702 274456 318708 274508
rect 318760 274496 318766 274508
rect 350534 274496 350540 274508
rect 318760 274468 350540 274496
rect 318760 274456 318766 274468
rect 350534 274456 350540 274468
rect 350592 274456 350598 274508
rect 351822 274456 351828 274508
rect 351880 274496 351886 274508
rect 400214 274496 400220 274508
rect 351880 274468 400220 274496
rect 351880 274456 351886 274468
rect 400214 274456 400220 274468
rect 400272 274456 400278 274508
rect 401318 274456 401324 274508
rect 401376 274496 401382 274508
rect 489914 274496 489920 274508
rect 401376 274468 489920 274496
rect 401376 274456 401382 274468
rect 489914 274456 489920 274468
rect 489972 274456 489978 274508
rect 490098 274456 490104 274508
rect 490156 274496 490162 274508
rect 494882 274496 494888 274508
rect 490156 274468 494888 274496
rect 490156 274456 490162 274468
rect 494882 274456 494888 274468
rect 494940 274456 494946 274508
rect 495066 274456 495072 274508
rect 495124 274496 495130 274508
rect 496998 274496 497004 274508
rect 495124 274468 497004 274496
rect 495124 274456 495130 274468
rect 496998 274456 497004 274468
rect 497056 274456 497062 274508
rect 497182 274456 497188 274508
rect 497240 274496 497246 274508
rect 617978 274496 617984 274508
rect 497240 274468 617984 274496
rect 497240 274456 497246 274468
rect 617978 274456 617984 274468
rect 618036 274456 618042 274508
rect 111978 274320 111984 274372
rect 112036 274360 112042 274372
rect 164234 274360 164240 274372
rect 112036 274332 164240 274360
rect 112036 274320 112042 274332
rect 164234 274320 164240 274332
rect 164292 274320 164298 274372
rect 177850 274320 177856 274372
rect 177908 274360 177914 274372
rect 204254 274360 204260 274372
rect 177908 274332 204260 274360
rect 177908 274320 177914 274332
rect 204254 274320 204260 274332
rect 204312 274320 204318 274372
rect 302878 274320 302884 274372
rect 302936 274360 302942 274372
rect 317690 274360 317696 274372
rect 302936 274332 317696 274360
rect 302936 274320 302942 274332
rect 317690 274320 317696 274332
rect 317748 274320 317754 274372
rect 336550 274320 336556 274372
rect 336608 274360 336614 274372
rect 378778 274360 378784 274372
rect 336608 274332 378784 274360
rect 336608 274320 336614 274332
rect 378778 274320 378784 274332
rect 378836 274320 378842 274372
rect 393222 274320 393228 274372
rect 393280 274360 393286 274372
rect 476114 274360 476120 274372
rect 393280 274332 476120 274360
rect 393280 274320 393286 274332
rect 476114 274320 476120 274332
rect 476172 274320 476178 274372
rect 478598 274320 478604 274372
rect 478656 274360 478662 274372
rect 610066 274360 610072 274372
rect 478656 274332 610072 274360
rect 478656 274320 478662 274332
rect 610066 274320 610072 274332
rect 610124 274320 610130 274372
rect 102502 274184 102508 274236
rect 102560 274224 102566 274236
rect 157886 274224 157892 274236
rect 102560 274196 157892 274224
rect 102560 274184 102566 274196
rect 157886 274184 157892 274196
rect 157944 274184 157950 274236
rect 166350 274184 166356 274236
rect 166408 274224 166414 274236
rect 198918 274224 198924 274236
rect 166408 274196 198924 274224
rect 166408 274184 166414 274196
rect 198918 274184 198924 274196
rect 198976 274184 198982 274236
rect 200574 274184 200580 274236
rect 200632 274224 200638 274236
rect 213178 274224 213184 274236
rect 200632 274196 213184 274224
rect 200632 274184 200638 274196
rect 213178 274184 213184 274196
rect 213236 274184 213242 274236
rect 283926 274184 283932 274236
rect 283984 274224 283990 274236
rect 302326 274224 302332 274236
rect 283984 274196 302332 274224
rect 283984 274184 283990 274196
rect 302326 274184 302332 274196
rect 302384 274184 302390 274236
rect 307570 274184 307576 274236
rect 307628 274224 307634 274236
rect 331214 274224 331220 274236
rect 307628 274196 331220 274224
rect 307628 274184 307634 274196
rect 331214 274184 331220 274196
rect 331272 274184 331278 274236
rect 343542 274184 343548 274236
rect 343600 274224 343606 274236
rect 391934 274224 391940 274236
rect 343600 274196 391940 274224
rect 343600 274184 343606 274196
rect 391934 274184 391940 274196
rect 391992 274184 391998 274236
rect 394326 274184 394332 274236
rect 394384 274224 394390 274236
rect 475194 274224 475200 274236
rect 394384 274196 475200 274224
rect 394384 274184 394390 274196
rect 475194 274184 475200 274196
rect 475252 274184 475258 274236
rect 475378 274184 475384 274236
rect 475436 274224 475442 274236
rect 485038 274224 485044 274236
rect 475436 274196 485044 274224
rect 475436 274184 475442 274196
rect 485038 274184 485044 274196
rect 485096 274184 485102 274236
rect 485222 274184 485228 274236
rect 485280 274224 485286 274236
rect 489730 274224 489736 274236
rect 485280 274196 489736 274224
rect 485280 274184 485286 274196
rect 489730 274184 489736 274196
rect 489788 274184 489794 274236
rect 489914 274184 489920 274236
rect 489972 274224 489978 274236
rect 621474 274224 621480 274236
rect 489972 274196 621480 274224
rect 489972 274184 489978 274196
rect 621474 274184 621480 274196
rect 621532 274184 621538 274236
rect 234890 274116 234896 274168
rect 234948 274156 234954 274168
rect 239490 274156 239496 274168
rect 234948 274128 239496 274156
rect 234948 274116 234954 274128
rect 239490 274116 239496 274128
rect 239548 274116 239554 274168
rect 77570 274048 77576 274100
rect 77628 274088 77634 274100
rect 143626 274088 143632 274100
rect 77628 274060 143632 274088
rect 77628 274048 77634 274060
rect 143626 274048 143632 274060
rect 143684 274048 143690 274100
rect 158070 274048 158076 274100
rect 158128 274088 158134 274100
rect 193306 274088 193312 274100
rect 158128 274060 193312 274088
rect 158128 274048 158134 274060
rect 193306 274048 193312 274060
rect 193364 274048 193370 274100
rect 198274 274048 198280 274100
rect 198332 274088 198338 274100
rect 218698 274088 218704 274100
rect 198332 274060 218704 274088
rect 198332 274048 198338 274060
rect 218698 274048 218704 274060
rect 218756 274048 218762 274100
rect 279878 274048 279884 274100
rect 279936 274088 279942 274100
rect 295150 274088 295156 274100
rect 279936 274060 295156 274088
rect 279936 274048 279942 274060
rect 295150 274048 295156 274060
rect 295208 274048 295214 274100
rect 300118 274048 300124 274100
rect 300176 274088 300182 274100
rect 325970 274088 325976 274100
rect 300176 274060 325976 274088
rect 300176 274048 300182 274060
rect 325970 274048 325976 274060
rect 326028 274048 326034 274100
rect 371878 274048 371884 274100
rect 371936 274088 371942 274100
rect 395706 274088 395712 274100
rect 371936 274060 395712 274088
rect 371936 274048 371942 274060
rect 395706 274048 395712 274060
rect 395764 274048 395770 274100
rect 397270 274048 397276 274100
rect 397328 274088 397334 274100
rect 483198 274088 483204 274100
rect 397328 274060 483204 274088
rect 397328 274048 397334 274060
rect 483198 274048 483204 274060
rect 483256 274048 483262 274100
rect 486694 274088 486700 274100
rect 483492 274060 486700 274088
rect 72970 273912 72976 273964
rect 73028 273952 73034 273964
rect 140958 273952 140964 273964
rect 73028 273924 140964 273952
rect 73028 273912 73034 273924
rect 140958 273912 140964 273924
rect 141016 273912 141022 273964
rect 141510 273912 141516 273964
rect 141568 273952 141574 273964
rect 183738 273952 183744 273964
rect 141568 273924 183744 273952
rect 141568 273912 141574 273924
rect 183738 273912 183744 273924
rect 183796 273912 183802 273964
rect 184106 273912 184112 273964
rect 184164 273952 184170 273964
rect 206278 273952 206284 273964
rect 184164 273924 206284 273952
rect 184164 273912 184170 273924
rect 206278 273912 206284 273924
rect 206336 273912 206342 273964
rect 206554 273912 206560 273964
rect 206612 273952 206618 273964
rect 223850 273952 223856 273964
rect 206612 273924 223856 273952
rect 206612 273912 206618 273924
rect 223850 273912 223856 273924
rect 223908 273912 223914 273964
rect 224218 273912 224224 273964
rect 224276 273952 224282 273964
rect 234890 273952 234896 273964
rect 224276 273924 234896 273952
rect 224276 273912 224282 273924
rect 234890 273912 234896 273924
rect 234948 273912 234954 273964
rect 274358 273912 274364 273964
rect 274416 273952 274422 273964
rect 286870 273952 286876 273964
rect 274416 273924 286876 273952
rect 274416 273912 274422 273924
rect 286870 273912 286876 273924
rect 286928 273912 286934 273964
rect 288066 273912 288072 273964
rect 288124 273952 288130 273964
rect 309410 273952 309416 273964
rect 288124 273924 309416 273952
rect 288124 273912 288130 273924
rect 309410 273912 309416 273924
rect 309468 273912 309474 273964
rect 314470 273912 314476 273964
rect 314528 273952 314534 273964
rect 342254 273952 342260 273964
rect 314528 273924 342260 273952
rect 314528 273912 314534 273924
rect 342254 273912 342260 273924
rect 342312 273912 342318 273964
rect 344646 273912 344652 273964
rect 344704 273952 344710 273964
rect 396718 273952 396724 273964
rect 344704 273924 396724 273952
rect 344704 273912 344710 273924
rect 396718 273912 396724 273924
rect 396776 273912 396782 273964
rect 398742 273912 398748 273964
rect 398800 273952 398806 273964
rect 483492 273952 483520 274060
rect 486694 274048 486700 274060
rect 486752 274048 486758 274100
rect 487062 274048 487068 274100
rect 487120 274088 487126 274100
rect 487120 274060 494744 274088
rect 487120 274048 487126 274060
rect 398800 273924 483520 273952
rect 398800 273912 398806 273924
rect 485038 273912 485044 273964
rect 485096 273952 485102 273964
rect 494514 273952 494520 273964
rect 485096 273924 494520 273952
rect 485096 273912 485102 273924
rect 494514 273912 494520 273924
rect 494572 273912 494578 273964
rect 494716 273952 494744 274060
rect 494882 274048 494888 274100
rect 494940 274088 494946 274100
rect 625062 274088 625068 274100
rect 494940 274060 625068 274088
rect 494940 274048 494946 274060
rect 625062 274048 625068 274060
rect 625120 274048 625126 274100
rect 628558 273952 628564 273964
rect 494716 273924 628564 273952
rect 628558 273912 628564 273924
rect 628616 273912 628622 273964
rect 632698 273912 632704 273964
rect 632756 273952 632762 273964
rect 643922 273952 643928 273964
rect 632756 273924 643928 273952
rect 632756 273912 632762 273924
rect 643922 273912 643928 273924
rect 643980 273912 643986 273964
rect 130838 273776 130844 273828
rect 130896 273816 130902 273828
rect 176746 273816 176752 273828
rect 130896 273788 176752 273816
rect 130896 273776 130902 273788
rect 176746 273776 176752 273788
rect 176804 273776 176810 273828
rect 322750 273776 322756 273828
rect 322808 273816 322814 273828
rect 358722 273816 358728 273828
rect 322808 273788 358728 273816
rect 322808 273776 322814 273788
rect 358722 273776 358728 273788
rect 358780 273776 358786 273828
rect 367002 273776 367008 273828
rect 367060 273816 367066 273828
rect 435910 273816 435916 273828
rect 367060 273788 435916 273816
rect 367060 273776 367066 273788
rect 435910 273776 435916 273788
rect 435968 273776 435974 273828
rect 446490 273816 446496 273828
rect 441586 273788 446496 273816
rect 124950 273640 124956 273692
rect 125008 273680 125014 273692
rect 149698 273680 149704 273692
rect 125008 273652 149704 273680
rect 125008 273640 125014 273652
rect 149698 273640 149704 273652
rect 149756 273640 149762 273692
rect 161474 273640 161480 273692
rect 161532 273680 161538 273692
rect 169938 273680 169944 273692
rect 161532 273652 169944 273680
rect 161532 273640 161538 273652
rect 169938 273640 169944 273652
rect 169996 273640 170002 273692
rect 374362 273640 374368 273692
rect 374420 273680 374426 273692
rect 420546 273680 420552 273692
rect 374420 273652 420552 273680
rect 374420 273640 374426 273652
rect 420546 273640 420552 273652
rect 420604 273640 420610 273692
rect 422662 273640 422668 273692
rect 422720 273680 422726 273692
rect 441586 273680 441614 273788
rect 446490 273776 446496 273788
rect 446548 273776 446554 273828
rect 448146 273776 448152 273828
rect 448204 273816 448210 273828
rect 448204 273788 460934 273816
rect 448204 273776 448210 273788
rect 422720 273652 441614 273680
rect 422720 273640 422726 273652
rect 446398 273640 446404 273692
rect 446456 273680 446462 273692
rect 460750 273680 460756 273692
rect 446456 273652 460756 273680
rect 446456 273640 446462 273652
rect 460750 273640 460756 273652
rect 460808 273640 460814 273692
rect 460906 273680 460934 273788
rect 461026 273776 461032 273828
rect 461084 273816 461090 273828
rect 569494 273816 569500 273828
rect 461084 273788 569500 273816
rect 461084 273776 461090 273788
rect 569494 273776 569500 273788
rect 569552 273776 569558 273828
rect 556154 273680 556160 273692
rect 460906 273652 556160 273680
rect 556154 273640 556160 273652
rect 556212 273640 556218 273692
rect 358078 273504 358084 273556
rect 358136 273544 358142 273556
rect 389726 273544 389732 273556
rect 358136 273516 389732 273544
rect 358136 273504 358142 273516
rect 389726 273504 389732 273516
rect 389784 273504 389790 273556
rect 394786 273504 394792 273556
rect 394844 273544 394850 273556
rect 397454 273544 397460 273556
rect 394844 273516 397460 273544
rect 394844 273504 394850 273516
rect 397454 273504 397460 273516
rect 397512 273504 397518 273556
rect 405182 273504 405188 273556
rect 405240 273544 405246 273556
rect 494330 273544 494336 273556
rect 405240 273516 494336 273544
rect 405240 273504 405246 273516
rect 494330 273504 494336 273516
rect 494388 273504 494394 273556
rect 494514 273504 494520 273556
rect 494572 273544 494578 273556
rect 529290 273544 529296 273556
rect 494572 273516 529296 273544
rect 494572 273504 494578 273516
rect 529290 273504 529296 273516
rect 529348 273504 529354 273556
rect 332502 273368 332508 273420
rect 332560 273408 332566 273420
rect 374638 273408 374644 273420
rect 332560 273380 374644 273408
rect 332560 273368 332566 273380
rect 374638 273368 374644 273380
rect 374696 273368 374702 273420
rect 378962 273368 378968 273420
rect 379020 273408 379026 273420
rect 409874 273408 409880 273420
rect 379020 273380 409880 273408
rect 379020 273368 379026 273380
rect 409874 273368 409880 273380
rect 409932 273368 409938 273420
rect 416406 273368 416412 273420
rect 416464 273408 416470 273420
rect 515122 273408 515128 273420
rect 416464 273380 515128 273408
rect 416464 273368 416470 273380
rect 515122 273368 515128 273380
rect 515180 273368 515186 273420
rect 414658 273300 414664 273352
rect 414716 273340 414722 273352
rect 414716 273312 415900 273340
rect 414716 273300 414722 273312
rect 353938 273232 353944 273284
rect 353996 273272 354002 273284
rect 382366 273272 382372 273284
rect 353996 273244 382372 273272
rect 353996 273232 354002 273244
rect 382366 273232 382372 273244
rect 382424 273232 382430 273284
rect 385954 273232 385960 273284
rect 386012 273272 386018 273284
rect 394786 273272 394792 273284
rect 386012 273244 394792 273272
rect 386012 273232 386018 273244
rect 394786 273232 394792 273244
rect 394844 273232 394850 273284
rect 42426 273164 42432 273216
rect 42484 273204 42490 273216
rect 45370 273204 45376 273216
rect 42484 273176 45376 273204
rect 42484 273164 42490 273176
rect 45370 273164 45376 273176
rect 45428 273164 45434 273216
rect 127342 273164 127348 273216
rect 127400 273204 127406 273216
rect 174630 273204 174636 273216
rect 127400 273176 174636 273204
rect 127400 273164 127406 273176
rect 174630 273164 174636 273176
rect 174688 273164 174694 273216
rect 326982 273164 326988 273216
rect 327040 273204 327046 273216
rect 345382 273204 345388 273216
rect 327040 273176 345388 273204
rect 327040 273164 327046 273176
rect 345382 273164 345388 273176
rect 345440 273164 345446 273216
rect 394970 273164 394976 273216
rect 395028 273204 395034 273216
rect 415670 273204 415676 273216
rect 395028 273176 415676 273204
rect 395028 273164 395034 273176
rect 415670 273164 415676 273176
rect 415728 273164 415734 273216
rect 415872 273204 415900 273312
rect 432046 273232 432052 273284
rect 432104 273272 432110 273284
rect 446398 273272 446404 273284
rect 432104 273244 446404 273272
rect 432104 273232 432110 273244
rect 446398 273232 446404 273244
rect 446456 273232 446462 273284
rect 431862 273204 431868 273216
rect 415872 273176 431868 273204
rect 431862 273164 431868 273176
rect 431920 273164 431926 273216
rect 450998 273164 451004 273216
rect 451056 273204 451062 273216
rect 568298 273204 568304 273216
rect 451056 273176 568304 273204
rect 451056 273164 451062 273176
rect 568298 273164 568304 273176
rect 568356 273164 568362 273216
rect 121362 273028 121368 273080
rect 121420 273068 121426 273080
rect 171594 273068 171600 273080
rect 121420 273040 171600 273068
rect 121420 273028 121426 273040
rect 171594 273028 171600 273040
rect 171652 273028 171658 273080
rect 174446 273028 174452 273080
rect 174504 273068 174510 273080
rect 196158 273068 196164 273080
rect 174504 273040 196164 273068
rect 174504 273028 174510 273040
rect 196158 273028 196164 273040
rect 196216 273028 196222 273080
rect 317506 273028 317512 273080
rect 317564 273068 317570 273080
rect 343818 273068 343824 273080
rect 317564 273040 343824 273068
rect 317564 273028 317570 273040
rect 343818 273028 343824 273040
rect 343876 273028 343882 273080
rect 345474 273028 345480 273080
rect 345532 273068 345538 273080
rect 372062 273068 372068 273080
rect 345532 273040 372068 273068
rect 345532 273028 345538 273040
rect 372062 273028 372068 273040
rect 372120 273028 372126 273080
rect 372430 273028 372436 273080
rect 372488 273068 372494 273080
rect 443822 273068 443828 273080
rect 372488 273040 443828 273068
rect 372488 273028 372494 273040
rect 443822 273028 443828 273040
rect 443880 273028 443886 273080
rect 444006 273028 444012 273080
rect 444064 273068 444070 273080
rect 450538 273068 450544 273080
rect 444064 273040 450544 273068
rect 444064 273028 444070 273040
rect 450538 273028 450544 273040
rect 450596 273028 450602 273080
rect 451274 273068 451280 273080
rect 450924 273040 451280 273068
rect 109586 272892 109592 272944
rect 109644 272932 109650 272944
rect 163406 272932 163412 272944
rect 109644 272904 163412 272932
rect 109644 272892 109650 272904
rect 163406 272892 163412 272904
rect 163464 272892 163470 272944
rect 180794 272892 180800 272944
rect 180852 272932 180858 272944
rect 207474 272932 207480 272944
rect 180852 272904 207480 272932
rect 180852 272892 180858 272904
rect 207474 272892 207480 272904
rect 207532 272892 207538 272944
rect 295058 272892 295064 272944
rect 295116 272932 295122 272944
rect 302510 272932 302516 272944
rect 295116 272904 302516 272932
rect 295116 272892 295122 272904
rect 302510 272892 302516 272904
rect 302568 272892 302574 272944
rect 310054 272892 310060 272944
rect 310112 272932 310118 272944
rect 319990 272932 319996 272944
rect 310112 272904 319996 272932
rect 310112 272892 310118 272904
rect 319990 272892 319996 272904
rect 320048 272892 320054 272944
rect 321462 272892 321468 272944
rect 321520 272932 321526 272944
rect 361390 272932 361396 272944
rect 321520 272904 361396 272932
rect 321520 272892 321526 272904
rect 361390 272892 361396 272904
rect 361448 272892 361454 272944
rect 376570 272892 376576 272944
rect 376628 272932 376634 272944
rect 450924 272932 450952 273040
rect 451274 273028 451280 273040
rect 451332 273028 451338 273080
rect 454034 273028 454040 273080
rect 454092 273068 454098 273080
rect 458174 273068 458180 273080
rect 454092 273040 458180 273068
rect 454092 273028 454098 273040
rect 458174 273028 458180 273040
rect 458232 273028 458238 273080
rect 461394 273028 461400 273080
rect 461452 273068 461458 273080
rect 571794 273068 571800 273080
rect 461452 273040 571800 273068
rect 461452 273028 461458 273040
rect 571794 273028 571800 273040
rect 571852 273028 571858 273080
rect 571978 273028 571984 273080
rect 572036 273068 572042 273080
rect 608502 273068 608508 273080
rect 572036 273040 608508 273068
rect 572036 273028 572042 273040
rect 608502 273028 608508 273040
rect 608560 273028 608566 273080
rect 376628 272904 450952 272932
rect 376628 272892 376634 272904
rect 451090 272892 451096 272944
rect 451148 272932 451154 272944
rect 451148 272904 454540 272932
rect 451148 272892 451154 272904
rect 97718 272756 97724 272808
rect 97776 272796 97782 272808
rect 155402 272796 155408 272808
rect 97776 272768 155408 272796
rect 97776 272756 97782 272768
rect 155402 272756 155408 272768
rect 155460 272756 155466 272808
rect 168650 272756 168656 272808
rect 168708 272796 168714 272808
rect 198734 272796 198740 272808
rect 168708 272768 198740 272796
rect 168708 272756 168714 272768
rect 198734 272756 198740 272768
rect 198792 272756 198798 272808
rect 298738 272756 298744 272808
rect 298796 272796 298802 272808
rect 310514 272796 310520 272808
rect 298796 272768 310520 272796
rect 298796 272756 298802 272768
rect 310514 272756 310520 272768
rect 310572 272756 310578 272808
rect 324038 272756 324044 272808
rect 324096 272796 324102 272808
rect 366082 272796 366088 272808
rect 324096 272768 366088 272796
rect 324096 272756 324102 272768
rect 366082 272756 366088 272768
rect 366140 272756 366146 272808
rect 371786 272756 371792 272808
rect 371844 272796 371850 272808
rect 377950 272796 377956 272808
rect 371844 272768 377956 272796
rect 371844 272756 371850 272768
rect 377950 272756 377956 272768
rect 378008 272756 378014 272808
rect 378134 272756 378140 272808
rect 378192 272796 378198 272808
rect 437382 272796 437388 272808
rect 378192 272768 437388 272796
rect 378192 272756 378198 272768
rect 437382 272756 437388 272768
rect 437440 272756 437446 272808
rect 437566 272756 437572 272808
rect 437624 272796 437630 272808
rect 441614 272796 441620 272808
rect 437624 272768 441620 272796
rect 437624 272756 437630 272768
rect 441614 272756 441620 272768
rect 441672 272756 441678 272808
rect 442258 272756 442264 272808
rect 442316 272796 442322 272808
rect 454034 272796 454040 272808
rect 442316 272768 454040 272796
rect 442316 272756 442322 272768
rect 454034 272756 454040 272768
rect 454092 272756 454098 272808
rect 454512 272796 454540 272904
rect 454678 272892 454684 272944
rect 454736 272932 454742 272944
rect 575382 272932 575388 272944
rect 454736 272904 575388 272932
rect 454736 272892 454742 272904
rect 575382 272892 575388 272904
rect 575440 272892 575446 272944
rect 564710 272796 564716 272808
rect 454512 272768 564716 272796
rect 564710 272756 564716 272768
rect 564768 272756 564774 272808
rect 578878 272756 578884 272808
rect 578936 272796 578942 272808
rect 636838 272796 636844 272808
rect 578936 272768 636844 272796
rect 578936 272756 578942 272768
rect 636838 272756 636844 272768
rect 636896 272756 636902 272808
rect 91830 272620 91836 272672
rect 91888 272660 91894 272672
rect 152366 272660 152372 272672
rect 91888 272632 152372 272660
rect 91888 272620 91894 272632
rect 152366 272620 152372 272632
rect 152424 272620 152430 272672
rect 159266 272620 159272 272672
rect 159324 272660 159330 272672
rect 194778 272660 194784 272672
rect 159324 272632 194784 272660
rect 159324 272620 159330 272632
rect 194778 272620 194784 272632
rect 194836 272620 194842 272672
rect 195698 272620 195704 272672
rect 195756 272660 195762 272672
rect 217226 272660 217232 272672
rect 195756 272632 217232 272660
rect 195756 272620 195762 272632
rect 217226 272620 217232 272632
rect 217284 272620 217290 272672
rect 217410 272620 217416 272672
rect 217468 272660 217474 272672
rect 230658 272660 230664 272672
rect 217468 272632 230664 272660
rect 217468 272620 217474 272632
rect 230658 272620 230664 272632
rect 230716 272620 230722 272672
rect 286870 272620 286876 272672
rect 286928 272660 286934 272672
rect 305822 272660 305828 272672
rect 286928 272632 305828 272660
rect 286928 272620 286934 272632
rect 305822 272620 305828 272632
rect 305880 272620 305886 272672
rect 306282 272620 306288 272672
rect 306340 272660 306346 272672
rect 317322 272660 317328 272672
rect 306340 272632 317328 272660
rect 306340 272620 306346 272632
rect 317322 272620 317328 272632
rect 317380 272620 317386 272672
rect 325510 272620 325516 272672
rect 325568 272660 325574 272672
rect 368474 272660 368480 272672
rect 325568 272632 368480 272660
rect 325568 272620 325574 272632
rect 368474 272620 368480 272632
rect 368532 272620 368538 272672
rect 369762 272620 369768 272672
rect 369820 272660 369826 272672
rect 436922 272660 436928 272672
rect 369820 272632 436928 272660
rect 369820 272620 369826 272632
rect 436922 272620 436928 272632
rect 436980 272620 436986 272672
rect 437106 272620 437112 272672
rect 437164 272660 437170 272672
rect 455966 272660 455972 272672
rect 437164 272632 455972 272660
rect 437164 272620 437170 272632
rect 455966 272620 455972 272632
rect 456024 272620 456030 272672
rect 461394 272660 461400 272672
rect 456168 272632 461400 272660
rect 239674 272552 239680 272604
rect 239732 272592 239738 272604
rect 244550 272592 244556 272604
rect 239732 272564 244556 272592
rect 239732 272552 239738 272564
rect 244550 272552 244556 272564
rect 244608 272552 244614 272604
rect 77754 272484 77760 272536
rect 77812 272524 77818 272536
rect 142154 272524 142160 272536
rect 77812 272496 142160 272524
rect 77812 272484 77818 272496
rect 142154 272484 142160 272496
rect 142212 272484 142218 272536
rect 154482 272484 154488 272536
rect 154540 272524 154546 272536
rect 190730 272524 190736 272536
rect 154540 272496 190736 272524
rect 154540 272484 154546 272496
rect 190730 272484 190736 272496
rect 190788 272484 190794 272536
rect 197078 272484 197084 272536
rect 197136 272524 197142 272536
rect 218054 272524 218060 272536
rect 197136 272496 218060 272524
rect 197136 272484 197142 272496
rect 218054 272484 218060 272496
rect 218112 272484 218118 272536
rect 218330 272484 218336 272536
rect 218388 272524 218394 272536
rect 231210 272524 231216 272536
rect 218388 272496 231216 272524
rect 218388 272484 218394 272496
rect 231210 272484 231216 272496
rect 231268 272484 231274 272536
rect 231394 272484 231400 272536
rect 231452 272524 231458 272536
rect 239306 272524 239312 272536
rect 231452 272496 239312 272524
rect 231452 272484 231458 272496
rect 239306 272484 239312 272496
rect 239364 272484 239370 272536
rect 271690 272484 271696 272536
rect 271748 272524 271754 272536
rect 280982 272524 280988 272536
rect 271748 272496 280988 272524
rect 271748 272484 271754 272496
rect 280982 272484 280988 272496
rect 281040 272484 281046 272536
rect 282178 272484 282184 272536
rect 282236 272524 282242 272536
rect 297542 272524 297548 272536
rect 282236 272496 297548 272524
rect 282236 272484 282242 272496
rect 297542 272484 297548 272496
rect 297600 272484 297606 272536
rect 303430 272484 303436 272536
rect 303488 272524 303494 272536
rect 322566 272524 322572 272536
rect 303488 272496 322572 272524
rect 303488 272484 303494 272496
rect 322566 272484 322572 272496
rect 322624 272484 322630 272536
rect 333238 272484 333244 272536
rect 333296 272524 333302 272536
rect 371786 272524 371792 272536
rect 333296 272496 371792 272524
rect 333296 272484 333302 272496
rect 371786 272484 371792 272496
rect 371844 272484 371850 272536
rect 371970 272484 371976 272536
rect 372028 272524 372034 272536
rect 374178 272524 374184 272536
rect 372028 272496 374184 272524
rect 372028 272484 372034 272496
rect 374178 272484 374184 272496
rect 374236 272484 374242 272536
rect 375006 272484 375012 272536
rect 375064 272524 375070 272536
rect 378134 272524 378140 272536
rect 375064 272496 378140 272524
rect 375064 272484 375070 272496
rect 378134 272484 378140 272496
rect 378192 272484 378198 272536
rect 384298 272484 384304 272536
rect 384356 272524 384362 272536
rect 388254 272524 388260 272536
rect 384356 272496 388260 272524
rect 384356 272484 384362 272496
rect 388254 272484 388260 272496
rect 388312 272484 388318 272536
rect 388438 272484 388444 272536
rect 388496 272524 388502 272536
rect 454218 272524 454224 272536
rect 388496 272496 454224 272524
rect 388496 272484 388502 272496
rect 454218 272484 454224 272496
rect 454276 272484 454282 272536
rect 454402 272484 454408 272536
rect 454460 272524 454466 272536
rect 456168 272524 456196 272632
rect 461394 272620 461400 272632
rect 461452 272620 461458 272672
rect 578510 272660 578516 272672
rect 461596 272632 578516 272660
rect 454460 272496 456196 272524
rect 454460 272484 454466 272496
rect 456518 272484 456524 272536
rect 456576 272524 456582 272536
rect 461596 272524 461624 272632
rect 578510 272620 578516 272632
rect 578568 272620 578574 272672
rect 456576 272496 461624 272524
rect 456576 272484 456582 272496
rect 461762 272484 461768 272536
rect 461820 272524 461826 272536
rect 466270 272524 466276 272536
rect 461820 272496 466276 272524
rect 461820 272484 461826 272496
rect 466270 272484 466276 272496
rect 466328 272484 466334 272536
rect 466454 272484 466460 272536
rect 466512 272524 466518 272536
rect 582466 272524 582472 272536
rect 466512 272496 582472 272524
rect 466512 272484 466518 272496
rect 582466 272484 582472 272496
rect 582524 272484 582530 272536
rect 585778 272484 585784 272536
rect 585836 272524 585842 272536
rect 622670 272524 622676 272536
rect 585836 272496 622676 272524
rect 585836 272484 585842 272496
rect 622670 272484 622676 272496
rect 622728 272484 622734 272536
rect 93026 272348 93032 272400
rect 93084 272388 93090 272400
rect 137554 272388 137560 272400
rect 93084 272360 137560 272388
rect 93084 272348 93090 272360
rect 137554 272348 137560 272360
rect 137612 272348 137618 272400
rect 137922 272348 137928 272400
rect 137980 272388 137986 272400
rect 181162 272388 181168 272400
rect 137980 272360 181168 272388
rect 137980 272348 137986 272360
rect 181162 272348 181168 272360
rect 181220 272348 181226 272400
rect 364242 272348 364248 272400
rect 364300 272388 364306 272400
rect 424502 272388 424508 272400
rect 364300 272360 424508 272388
rect 364300 272348 364306 272360
rect 424502 272348 424508 272360
rect 424560 272348 424566 272400
rect 442258 272388 442264 272400
rect 424796 272360 442264 272388
rect 116670 272212 116676 272264
rect 116728 272252 116734 272264
rect 159634 272252 159640 272264
rect 116728 272224 159640 272252
rect 116728 272212 116734 272224
rect 159634 272212 159640 272224
rect 159692 272212 159698 272264
rect 362770 272212 362776 272264
rect 362828 272252 362834 272264
rect 405366 272252 405372 272264
rect 362828 272224 405372 272252
rect 362828 272212 362834 272224
rect 405366 272212 405372 272224
rect 405424 272212 405430 272264
rect 424796 272252 424824 272360
rect 442258 272348 442264 272360
rect 442316 272348 442322 272400
rect 442442 272348 442448 272400
rect 442500 272388 442506 272400
rect 444006 272388 444012 272400
rect 442500 272360 444012 272388
rect 442500 272348 442506 272360
rect 444006 272348 444012 272360
rect 444064 272348 444070 272400
rect 444190 272348 444196 272400
rect 444248 272388 444254 272400
rect 475654 272388 475660 272400
rect 444248 272360 475660 272388
rect 444248 272348 444254 272360
rect 475654 272348 475660 272360
rect 475712 272348 475718 272400
rect 476022 272348 476028 272400
rect 476080 272388 476086 272400
rect 480070 272388 480076 272400
rect 476080 272360 480076 272388
rect 476080 272348 476086 272360
rect 480070 272348 480076 272360
rect 480128 272348 480134 272400
rect 480208 272348 480214 272400
rect 480266 272388 480272 272400
rect 487614 272388 487620 272400
rect 480266 272360 487620 272388
rect 480266 272348 480272 272360
rect 487614 272348 487620 272360
rect 487672 272348 487678 272400
rect 490650 272348 490656 272400
rect 490708 272388 490714 272400
rect 499022 272388 499028 272400
rect 490708 272360 499028 272388
rect 490708 272348 490714 272360
rect 499022 272348 499028 272360
rect 499080 272348 499086 272400
rect 499390 272348 499396 272400
rect 499448 272388 499454 272400
rect 551554 272388 551560 272400
rect 499448 272360 551560 272388
rect 499448 272348 499454 272360
rect 551554 272348 551560 272360
rect 551612 272348 551618 272400
rect 552658 272348 552664 272400
rect 552716 272388 552722 272400
rect 586054 272388 586060 272400
rect 552716 272360 586060 272388
rect 552716 272348 552722 272360
rect 586054 272348 586060 272360
rect 586112 272348 586118 272400
rect 405568 272224 424824 272252
rect 340690 272076 340696 272128
rect 340748 272116 340754 272128
rect 371970 272116 371976 272128
rect 340748 272088 371976 272116
rect 340748 272076 340754 272088
rect 371970 272076 371976 272088
rect 372028 272076 372034 272128
rect 380894 272116 380900 272128
rect 372448 272088 380900 272116
rect 355870 271940 355876 271992
rect 355928 271980 355934 271992
rect 372448 271980 372476 272088
rect 380894 272076 380900 272088
rect 380952 272076 380958 272128
rect 382182 272076 382188 272128
rect 382240 272116 382246 272128
rect 405568 272116 405596 272224
rect 427078 272212 427084 272264
rect 427136 272252 427142 272264
rect 437382 272252 437388 272264
rect 427136 272224 437388 272252
rect 427136 272212 427142 272224
rect 437382 272212 437388 272224
rect 437440 272212 437446 272264
rect 437566 272212 437572 272264
rect 437624 272252 437630 272264
rect 447686 272252 447692 272264
rect 437624 272224 447692 272252
rect 437624 272212 437630 272224
rect 447686 272212 447692 272224
rect 447744 272212 447750 272264
rect 447870 272212 447876 272264
rect 447928 272252 447934 272264
rect 489730 272252 489736 272264
rect 447928 272224 489736 272252
rect 447928 272212 447934 272224
rect 489730 272212 489736 272224
rect 489788 272212 489794 272264
rect 490190 272212 490196 272264
rect 490248 272252 490254 272264
rect 561214 272252 561220 272264
rect 490248 272224 561220 272252
rect 490248 272212 490254 272224
rect 561214 272212 561220 272224
rect 561272 272212 561278 272264
rect 382240 272088 405596 272116
rect 382240 272076 382246 272088
rect 411898 272076 411904 272128
rect 411956 272116 411962 272128
rect 487798 272116 487804 272128
rect 411956 272088 487804 272116
rect 411956 272076 411962 272088
rect 487798 272076 487804 272088
rect 487856 272076 487862 272128
rect 499022 272076 499028 272128
rect 499080 272116 499086 272128
rect 499666 272116 499672 272128
rect 499080 272088 499672 272116
rect 499080 272076 499086 272088
rect 499666 272076 499672 272088
rect 499724 272076 499730 272128
rect 500218 272076 500224 272128
rect 500276 272116 500282 272128
rect 552658 272116 552664 272128
rect 500276 272088 552664 272116
rect 500276 272076 500282 272088
rect 552658 272076 552664 272088
rect 552716 272076 552722 272128
rect 490006 272008 490012 272060
rect 490064 272048 490070 272060
rect 498838 272048 498844 272060
rect 490064 272020 498844 272048
rect 490064 272008 490070 272020
rect 498838 272008 498844 272020
rect 498896 272008 498902 272060
rect 355928 271952 372476 271980
rect 355928 271940 355934 271952
rect 378778 271940 378784 271992
rect 378836 271980 378842 271992
rect 388438 271980 388444 271992
rect 378836 271952 388444 271980
rect 378836 271940 378842 271952
rect 388438 271940 388444 271952
rect 388496 271940 388502 271992
rect 388622 271940 388628 271992
rect 388680 271980 388686 271992
rect 394970 271980 394976 271992
rect 388680 271952 394976 271980
rect 388680 271940 388686 271952
rect 394970 271940 394976 271952
rect 395028 271940 395034 271992
rect 405366 271940 405372 271992
rect 405424 271980 405430 271992
rect 415210 271980 415216 271992
rect 405424 271952 415216 271980
rect 405424 271940 405430 271952
rect 415210 271940 415216 271952
rect 415268 271940 415274 271992
rect 415670 271940 415676 271992
rect 415728 271980 415734 271992
rect 427078 271980 427084 271992
rect 415728 271952 427084 271980
rect 415728 271940 415734 271952
rect 427078 271940 427084 271952
rect 427136 271940 427142 271992
rect 427722 271940 427728 271992
rect 427780 271980 427786 271992
rect 489868 271980 489874 271992
rect 427780 271952 489874 271980
rect 427780 271940 427786 271952
rect 489868 271940 489874 271952
rect 489926 271940 489932 271992
rect 499528 271940 499534 271992
rect 499586 271980 499592 271992
rect 532786 271980 532792 271992
rect 499586 271952 532792 271980
rect 499586 271940 499592 271952
rect 532786 271940 532792 271952
rect 532844 271940 532850 271992
rect 551554 271940 551560 271992
rect 551612 271980 551618 271992
rect 555234 271980 555240 271992
rect 551612 271952 555240 271980
rect 551612 271940 551618 271952
rect 555234 271940 555240 271952
rect 555292 271940 555298 271992
rect 101306 271804 101312 271856
rect 101364 271844 101370 271856
rect 157610 271844 157616 271856
rect 101364 271816 157616 271844
rect 101364 271804 101370 271816
rect 157610 271804 157616 271816
rect 157668 271804 157674 271856
rect 179138 271804 179144 271856
rect 179196 271844 179202 271856
rect 204898 271844 204904 271856
rect 179196 271816 204904 271844
rect 179196 271804 179202 271816
rect 204898 271804 204904 271816
rect 204956 271804 204962 271856
rect 232498 271804 232504 271856
rect 232556 271844 232562 271856
rect 233878 271844 233884 271856
rect 232556 271816 233884 271844
rect 232556 271804 232562 271816
rect 233878 271804 233884 271816
rect 233936 271804 233942 271856
rect 304902 271804 304908 271856
rect 304960 271844 304966 271856
rect 334158 271844 334164 271856
rect 304960 271816 334164 271844
rect 304960 271804 304966 271816
rect 334158 271804 334164 271816
rect 334216 271804 334222 271856
rect 334618 271804 334624 271856
rect 334676 271844 334682 271856
rect 349614 271844 349620 271856
rect 334676 271816 349620 271844
rect 334676 271804 334682 271816
rect 349614 271804 349620 271816
rect 349672 271804 349678 271856
rect 361298 271804 361304 271856
rect 361356 271844 361362 271856
rect 426434 271844 426440 271856
rect 361356 271816 426440 271844
rect 361356 271804 361362 271816
rect 426434 271804 426440 271816
rect 426492 271804 426498 271856
rect 427538 271804 427544 271856
rect 427596 271844 427602 271856
rect 531590 271844 531596 271856
rect 427596 271816 531596 271844
rect 427596 271804 427602 271816
rect 531590 271804 531596 271816
rect 531648 271804 531654 271856
rect 538766 271844 538772 271856
rect 533356 271816 538772 271844
rect 263410 271736 263416 271788
rect 263468 271776 263474 271788
rect 269206 271776 269212 271788
rect 263468 271748 269212 271776
rect 263468 271736 263474 271748
rect 269206 271736 269212 271748
rect 269264 271736 269270 271788
rect 349816 271748 354674 271776
rect 88610 271668 88616 271720
rect 88668 271708 88674 271720
rect 145650 271708 145656 271720
rect 88668 271680 145656 271708
rect 88668 271668 88674 271680
rect 145650 271668 145656 271680
rect 145708 271668 145714 271720
rect 170122 271668 170128 271720
rect 170180 271708 170186 271720
rect 201034 271708 201040 271720
rect 170180 271680 201040 271708
rect 170180 271668 170186 271680
rect 201034 271668 201040 271680
rect 201092 271668 201098 271720
rect 296622 271668 296628 271720
rect 296680 271708 296686 271720
rect 301130 271708 301136 271720
rect 296680 271680 301136 271708
rect 296680 271668 296686 271680
rect 301130 271668 301136 271680
rect 301188 271668 301194 271720
rect 309042 271668 309048 271720
rect 309100 271708 309106 271720
rect 342438 271708 342444 271720
rect 309100 271680 342444 271708
rect 309100 271668 309106 271680
rect 342438 271668 342444 271680
rect 342496 271668 342502 271720
rect 347774 271668 347780 271720
rect 347832 271708 347838 271720
rect 349816 271708 349844 271748
rect 347832 271680 349844 271708
rect 354646 271708 354674 271748
rect 363598 271708 363604 271720
rect 354646 271680 363604 271708
rect 347832 271668 347838 271680
rect 363598 271668 363604 271680
rect 363656 271668 363662 271720
rect 363782 271668 363788 271720
rect 363840 271708 363846 271720
rect 429746 271708 429752 271720
rect 363840 271680 429752 271708
rect 363840 271668 363846 271680
rect 429746 271668 429752 271680
rect 429804 271668 429810 271720
rect 435174 271708 435180 271720
rect 430040 271680 435180 271708
rect 352190 271640 352196 271652
rect 350506 271612 352196 271640
rect 98914 271532 98920 271584
rect 98972 271572 98978 271584
rect 156506 271572 156512 271584
rect 98972 271544 156512 271572
rect 98972 271532 98978 271544
rect 156506 271532 156512 271544
rect 156564 271532 156570 271584
rect 165154 271532 165160 271584
rect 165212 271572 165218 271584
rect 197354 271572 197360 271584
rect 165212 271544 197360 271572
rect 165212 271532 165218 271544
rect 197354 271532 197360 271544
rect 197412 271532 197418 271584
rect 213638 271532 213644 271584
rect 213696 271572 213702 271584
rect 228266 271572 228272 271584
rect 213696 271544 228272 271572
rect 213696 271532 213702 271544
rect 228266 271532 228272 271544
rect 228324 271532 228330 271584
rect 289630 271532 289636 271584
rect 289688 271572 289694 271584
rect 297266 271572 297272 271584
rect 289688 271544 297272 271572
rect 289688 271532 289694 271544
rect 297266 271532 297272 271544
rect 297324 271532 297330 271584
rect 301498 271532 301504 271584
rect 301556 271572 301562 271584
rect 314102 271572 314108 271584
rect 301556 271544 314108 271572
rect 301556 271532 301562 271544
rect 314102 271532 314108 271544
rect 314160 271532 314166 271584
rect 315942 271532 315948 271584
rect 316000 271572 316006 271584
rect 345658 271572 345664 271584
rect 316000 271544 345664 271572
rect 316000 271532 316006 271544
rect 345658 271532 345664 271544
rect 345716 271532 345722 271584
rect 346578 271532 346584 271584
rect 346636 271572 346642 271584
rect 350506 271572 350534 271612
rect 352190 271600 352196 271612
rect 352248 271600 352254 271652
rect 346636 271544 350534 271572
rect 346636 271532 346642 271544
rect 359458 271532 359464 271584
rect 359516 271572 359522 271584
rect 365438 271572 365444 271584
rect 359516 271544 365444 271572
rect 359516 271532 359522 271544
rect 365438 271532 365444 271544
rect 365496 271532 365502 271584
rect 383194 271532 383200 271584
rect 383252 271572 383258 271584
rect 388622 271572 388628 271584
rect 383252 271544 388628 271572
rect 383252 271532 383258 271544
rect 388622 271532 388628 271544
rect 388680 271532 388686 271584
rect 388806 271532 388812 271584
rect 388864 271572 388870 271584
rect 391750 271572 391756 271584
rect 388864 271544 391756 271572
rect 388864 271532 388870 271544
rect 391750 271532 391756 271544
rect 391808 271532 391814 271584
rect 391934 271532 391940 271584
rect 391992 271572 391998 271584
rect 430040 271572 430068 271680
rect 435174 271668 435180 271680
rect 435232 271668 435238 271720
rect 435358 271668 435364 271720
rect 435416 271708 435422 271720
rect 533356 271708 533384 271816
rect 538766 271804 538772 271816
rect 538824 271804 538830 271856
rect 435416 271680 533384 271708
rect 435416 271668 435422 271680
rect 533522 271668 533528 271720
rect 533580 271708 533586 271720
rect 551738 271708 551744 271720
rect 533580 271680 551744 271708
rect 533580 271668 533586 271680
rect 551738 271668 551744 271680
rect 551796 271668 551802 271720
rect 554038 271668 554044 271720
rect 554096 271708 554102 271720
rect 615678 271708 615684 271720
rect 554096 271680 615684 271708
rect 554096 271668 554102 271680
rect 615678 271668 615684 271680
rect 615736 271668 615742 271720
rect 391992 271544 430068 271572
rect 391992 271532 391998 271544
rect 430206 271532 430212 271584
rect 430264 271572 430270 271584
rect 440602 271572 440608 271584
rect 430264 271544 440608 271572
rect 430264 271532 430270 271544
rect 440602 271532 440608 271544
rect 440660 271532 440666 271584
rect 440970 271532 440976 271584
rect 441028 271572 441034 271584
rect 441028 271544 446904 271572
rect 441028 271532 441034 271544
rect 446876 271504 446904 271544
rect 447088 271532 447094 271584
rect 447146 271572 447152 271584
rect 451228 271572 451234 271584
rect 447146 271544 451234 271572
rect 447146 271532 447152 271544
rect 451228 271532 451234 271544
rect 451286 271532 451292 271584
rect 451366 271532 451372 271584
rect 451424 271572 451430 271584
rect 480254 271572 480260 271584
rect 451424 271544 480260 271572
rect 451424 271532 451430 271544
rect 480254 271532 480260 271544
rect 480312 271532 480318 271584
rect 480530 271532 480536 271584
rect 480588 271572 480594 271584
rect 489270 271572 489276 271584
rect 480588 271544 489276 271572
rect 480588 271532 480594 271544
rect 489270 271532 489276 271544
rect 489328 271532 489334 271584
rect 489638 271532 489644 271584
rect 489696 271572 489702 271584
rect 562410 271572 562416 271584
rect 489696 271544 562416 271572
rect 489696 271532 489702 271544
rect 562410 271532 562416 271544
rect 562468 271532 562474 271584
rect 625798 271532 625804 271584
rect 625856 271572 625862 271584
rect 629754 271572 629760 271584
rect 625856 271544 629760 271572
rect 625856 271532 625862 271544
rect 629754 271532 629760 271544
rect 629812 271532 629818 271584
rect 446876 271476 446996 271504
rect 92474 271396 92480 271448
rect 92532 271436 92538 271448
rect 150434 271436 150440 271448
rect 92532 271408 150440 271436
rect 92532 271396 92538 271408
rect 150434 271396 150440 271408
rect 150492 271396 150498 271448
rect 150986 271396 150992 271448
rect 151044 271436 151050 271448
rect 188246 271436 188252 271448
rect 151044 271408 188252 271436
rect 151044 271396 151050 271408
rect 188246 271396 188252 271408
rect 188304 271396 188310 271448
rect 201770 271396 201776 271448
rect 201828 271436 201834 271448
rect 220998 271436 221004 271448
rect 201828 271408 221004 271436
rect 201828 271396 201834 271408
rect 220998 271396 221004 271408
rect 221056 271396 221062 271448
rect 229002 271396 229008 271448
rect 229060 271436 229066 271448
rect 237834 271436 237840 271448
rect 229060 271408 237840 271436
rect 229060 271396 229066 271408
rect 237834 271396 237840 271408
rect 237892 271396 237898 271448
rect 268838 271396 268844 271448
rect 268896 271436 268902 271448
rect 277486 271436 277492 271448
rect 268896 271408 277492 271436
rect 268896 271396 268902 271408
rect 277486 271396 277492 271408
rect 277544 271396 277550 271448
rect 286318 271396 286324 271448
rect 286376 271436 286382 271448
rect 296346 271436 296352 271448
rect 286376 271408 296352 271436
rect 286376 271396 286382 271408
rect 296346 271396 296352 271408
rect 296404 271396 296410 271448
rect 300670 271396 300676 271448
rect 300728 271436 300734 271448
rect 311066 271436 311072 271448
rect 300728 271408 311072 271436
rect 300728 271396 300734 271408
rect 311066 271396 311072 271408
rect 311124 271396 311130 271448
rect 311710 271396 311716 271448
rect 311768 271436 311774 271448
rect 346762 271436 346768 271448
rect 311768 271408 346768 271436
rect 311768 271396 311774 271408
rect 346762 271396 346768 271408
rect 346820 271396 346826 271448
rect 350074 271396 350080 271448
rect 350132 271436 350138 271448
rect 388070 271436 388076 271448
rect 350132 271408 388076 271436
rect 350132 271396 350138 271408
rect 388070 271396 388076 271408
rect 388128 271396 388134 271448
rect 413462 271436 413468 271448
rect 388456 271408 413468 271436
rect 84746 271260 84752 271312
rect 84804 271300 84810 271312
rect 147674 271300 147680 271312
rect 84804 271272 147680 271300
rect 84804 271260 84810 271272
rect 147674 271260 147680 271272
rect 147732 271260 147738 271312
rect 155678 271260 155684 271312
rect 155736 271300 155742 271312
rect 192202 271300 192208 271312
rect 155736 271272 192208 271300
rect 155736 271260 155742 271272
rect 192202 271260 192208 271272
rect 192260 271260 192266 271312
rect 193490 271260 193496 271312
rect 193548 271300 193554 271312
rect 215754 271300 215760 271312
rect 193548 271272 215760 271300
rect 193548 271260 193554 271272
rect 215754 271260 215760 271272
rect 215812 271260 215818 271312
rect 221918 271260 221924 271312
rect 221976 271300 221982 271312
rect 232498 271300 232504 271312
rect 221976 271272 232504 271300
rect 221976 271260 221982 271272
rect 232498 271260 232504 271272
rect 232556 271260 232562 271312
rect 273070 271260 273076 271312
rect 273128 271300 273134 271312
rect 284570 271300 284576 271312
rect 273128 271272 284576 271300
rect 273128 271260 273134 271272
rect 284570 271260 284576 271272
rect 284628 271260 284634 271312
rect 285306 271260 285312 271312
rect 285364 271300 285370 271312
rect 304626 271300 304632 271312
rect 285364 271272 304632 271300
rect 285364 271260 285370 271272
rect 304626 271260 304632 271272
rect 304684 271260 304690 271312
rect 319990 271260 319996 271312
rect 320048 271300 320054 271312
rect 360194 271300 360200 271312
rect 320048 271272 360200 271300
rect 320048 271260 320054 271272
rect 360194 271260 360200 271272
rect 360252 271260 360258 271312
rect 370314 271260 370320 271312
rect 370372 271300 370378 271312
rect 388456 271300 388484 271408
rect 413462 271396 413468 271408
rect 413520 271396 413526 271448
rect 413922 271396 413928 271448
rect 413980 271436 413986 271448
rect 427078 271436 427084 271448
rect 413980 271408 427084 271436
rect 413980 271396 413986 271408
rect 427078 271396 427084 271408
rect 427136 271396 427142 271448
rect 430022 271396 430028 271448
rect 430080 271436 430086 271448
rect 433426 271436 433432 271448
rect 430080 271408 433432 271436
rect 430080 271396 430086 271408
rect 433426 271396 433432 271408
rect 433484 271396 433490 271448
rect 433610 271396 433616 271448
rect 433668 271436 433674 271448
rect 435358 271436 435364 271448
rect 433668 271408 435364 271436
rect 433668 271396 433674 271408
rect 435358 271396 435364 271408
rect 435416 271396 435422 271448
rect 439130 271396 439136 271448
rect 439188 271436 439194 271448
rect 446674 271436 446680 271448
rect 439188 271408 446680 271436
rect 439188 271396 439194 271408
rect 446674 271396 446680 271408
rect 446732 271396 446738 271448
rect 446968 271436 446996 271476
rect 553854 271436 553860 271448
rect 446968 271408 489408 271436
rect 489380 271368 489408 271408
rect 489656 271408 553860 271436
rect 489656 271368 489684 271408
rect 553854 271396 553860 271408
rect 553912 271396 553918 271448
rect 489380 271340 489684 271368
rect 370372 271272 388484 271300
rect 370372 271260 370378 271272
rect 388622 271260 388628 271312
rect 388680 271300 388686 271312
rect 461578 271300 461584 271312
rect 388680 271272 461584 271300
rect 388680 271260 388686 271272
rect 461578 271260 461584 271272
rect 461636 271260 461642 271312
rect 461762 271260 461768 271312
rect 461820 271300 461826 271312
rect 465166 271300 465172 271312
rect 461820 271272 465172 271300
rect 461820 271260 461826 271272
rect 465166 271260 465172 271272
rect 465224 271260 465230 271312
rect 465350 271260 465356 271312
rect 465408 271300 465414 271312
rect 465408 271272 480484 271300
rect 465408 271260 465414 271272
rect 480456 271232 480484 271272
rect 480714 271260 480720 271312
rect 480772 271300 480778 271312
rect 487614 271300 487620 271312
rect 480772 271272 487620 271300
rect 480772 271260 480778 271272
rect 487614 271260 487620 271272
rect 487672 271260 487678 271312
rect 580074 271300 580080 271312
rect 489748 271272 580080 271300
rect 489748 271232 489776 271272
rect 580074 271260 580080 271272
rect 580132 271260 580138 271312
rect 480456 271204 480576 271232
rect 65886 271124 65892 271176
rect 65944 271164 65950 271176
rect 136634 271164 136640 271176
rect 65944 271136 136640 271164
rect 65944 271124 65950 271136
rect 136634 271124 136640 271136
rect 136692 271124 136698 271176
rect 139118 271124 139124 271176
rect 139176 271164 139182 271176
rect 140498 271164 140504 271176
rect 139176 271136 140504 271164
rect 139176 271124 139182 271136
rect 140498 271124 140504 271136
rect 140556 271124 140562 271176
rect 145006 271124 145012 271176
rect 145064 271164 145070 271176
rect 184934 271164 184940 271176
rect 145064 271136 184940 271164
rect 145064 271124 145070 271136
rect 184934 271124 184940 271136
rect 184992 271124 184998 271176
rect 185578 271124 185584 271176
rect 185636 271164 185642 271176
rect 191834 271164 191840 271176
rect 185636 271136 191840 271164
rect 185636 271124 185642 271136
rect 191834 271124 191840 271136
rect 191892 271124 191898 271176
rect 192386 271124 192392 271176
rect 192444 271164 192450 271176
rect 215294 271164 215300 271176
rect 192444 271136 215300 271164
rect 192444 271124 192450 271136
rect 215294 271124 215300 271136
rect 215352 271124 215358 271176
rect 215938 271124 215944 271176
rect 215996 271164 216002 271176
rect 229738 271164 229744 271176
rect 215996 271136 229744 271164
rect 215996 271124 216002 271136
rect 229738 271124 229744 271136
rect 229796 271124 229802 271176
rect 233694 271124 233700 271176
rect 233752 271164 233758 271176
rect 240778 271164 240784 271176
rect 233752 271136 240784 271164
rect 233752 271124 233758 271136
rect 240778 271124 240784 271136
rect 240836 271124 240842 271176
rect 277302 271124 277308 271176
rect 277360 271164 277366 271176
rect 291654 271164 291660 271176
rect 277360 271136 291660 271164
rect 277360 271124 277366 271136
rect 291654 271124 291660 271136
rect 291712 271124 291718 271176
rect 292390 271124 292396 271176
rect 292448 271164 292454 271176
rect 315298 271164 315304 271176
rect 292448 271136 315304 271164
rect 292448 271124 292454 271136
rect 315298 271124 315304 271136
rect 315356 271124 315362 271176
rect 321278 271124 321284 271176
rect 321336 271164 321342 271176
rect 362586 271164 362592 271176
rect 321336 271136 362592 271164
rect 321336 271124 321342 271136
rect 362586 271124 362592 271136
rect 362644 271124 362650 271176
rect 365622 271124 365628 271176
rect 365680 271164 365686 271176
rect 424502 271164 424508 271176
rect 365680 271136 424508 271164
rect 365680 271124 365686 271136
rect 424502 271124 424508 271136
rect 424560 271124 424566 271176
rect 430206 271164 430212 271176
rect 424888 271136 430212 271164
rect 114278 270988 114284 271040
rect 114336 271028 114342 271040
rect 167178 271028 167184 271040
rect 114336 271000 167184 271028
rect 114336 270988 114342 271000
rect 167178 270988 167184 271000
rect 167236 270988 167242 271040
rect 337746 270988 337752 271040
rect 337804 271028 337810 271040
rect 359458 271028 359464 271040
rect 337804 271000 359464 271028
rect 337804 270988 337810 271000
rect 359458 270988 359464 271000
rect 359516 270988 359522 271040
rect 360102 270988 360108 271040
rect 360160 271028 360166 271040
rect 413278 271028 413284 271040
rect 360160 271000 413284 271028
rect 360160 270988 360166 271000
rect 413278 270988 413284 271000
rect 413336 270988 413342 271040
rect 413462 270988 413468 271040
rect 413520 271028 413526 271040
rect 424888 271028 424916 271136
rect 430206 271124 430212 271136
rect 430264 271124 430270 271176
rect 456748 271164 456754 271176
rect 430408 271136 456754 271164
rect 413520 271000 424916 271028
rect 413520 270988 413526 271000
rect 427078 270988 427084 271040
rect 427136 271028 427142 271040
rect 430408 271028 430436 271136
rect 456748 271124 456754 271136
rect 456806 271124 456812 271176
rect 456886 271124 456892 271176
rect 456944 271164 456950 271176
rect 466408 271164 466414 271176
rect 456944 271136 466414 271164
rect 456944 271124 456950 271136
rect 466408 271124 466414 271136
rect 466466 271124 466472 271176
rect 466546 271124 466552 271176
rect 466604 271164 466610 271176
rect 480254 271164 480260 271176
rect 466604 271136 480260 271164
rect 466604 271124 466610 271136
rect 480254 271124 480260 271136
rect 480312 271124 480318 271176
rect 480548 271164 480576 271204
rect 489564 271204 489776 271232
rect 489564 271164 489592 271204
rect 480548 271136 489592 271164
rect 489914 271124 489920 271176
rect 489972 271164 489978 271176
rect 594334 271164 594340 271176
rect 489972 271136 594340 271164
rect 489972 271124 489978 271136
rect 594334 271124 594340 271136
rect 594392 271124 594398 271176
rect 427136 271000 430436 271028
rect 427136 270988 427142 271000
rect 431770 270988 431776 271040
rect 431828 271028 431834 271040
rect 539870 271028 539876 271040
rect 431828 271000 539876 271028
rect 431828 270988 431834 271000
rect 539870 270988 539876 271000
rect 539928 270988 539934 271040
rect 123754 270852 123760 270904
rect 123812 270892 123818 270904
rect 172698 270892 172704 270904
rect 123812 270864 172704 270892
rect 123812 270852 123818 270864
rect 172698 270852 172704 270864
rect 172756 270852 172762 270904
rect 344186 270852 344192 270904
rect 344244 270892 344250 270904
rect 356882 270892 356888 270904
rect 344244 270864 356888 270892
rect 344244 270852 344250 270864
rect 356882 270852 356888 270864
rect 356940 270852 356946 270904
rect 357158 270852 357164 270904
rect 357216 270892 357222 270904
rect 417694 270892 417700 270904
rect 357216 270864 417700 270892
rect 357216 270852 357222 270864
rect 417694 270852 417700 270864
rect 417752 270852 417758 270904
rect 418154 270852 418160 270904
rect 418212 270892 418218 270904
rect 418982 270892 418988 270904
rect 418212 270864 418988 270892
rect 418212 270852 418218 270864
rect 418982 270852 418988 270864
rect 419040 270852 419046 270904
rect 419442 270852 419448 270904
rect 419500 270892 419506 270904
rect 509188 270892 509194 270904
rect 419500 270864 509194 270892
rect 419500 270852 419506 270864
rect 509188 270852 509194 270864
rect 509246 270852 509252 270904
rect 509418 270852 509424 270904
rect 509476 270892 509482 270904
rect 533522 270892 533528 270904
rect 509476 270864 533528 270892
rect 509476 270852 509482 270864
rect 533522 270852 533528 270864
rect 533580 270852 533586 270904
rect 538858 270852 538864 270904
rect 538916 270892 538922 270904
rect 597830 270892 597836 270904
rect 538916 270864 597836 270892
rect 538916 270852 538922 270864
rect 597830 270852 597836 270864
rect 597888 270852 597894 270904
rect 134426 270716 134432 270768
rect 134484 270756 134490 270768
rect 178954 270756 178960 270768
rect 134484 270728 178960 270756
rect 134484 270716 134490 270728
rect 178954 270716 178960 270728
rect 179012 270716 179018 270768
rect 345658 270716 345664 270768
rect 345716 270756 345722 270768
rect 353110 270756 353116 270768
rect 345716 270728 353116 270756
rect 345716 270716 345722 270728
rect 353110 270716 353116 270728
rect 353168 270716 353174 270768
rect 354582 270716 354588 270768
rect 354640 270756 354646 270768
rect 402882 270756 402888 270768
rect 354640 270728 402888 270756
rect 354640 270716 354646 270728
rect 402882 270716 402888 270728
rect 402940 270716 402946 270768
rect 403066 270716 403072 270768
rect 403124 270756 403130 270768
rect 403986 270756 403992 270768
rect 403124 270728 403992 270756
rect 403124 270716 403130 270728
rect 403986 270716 403992 270728
rect 404044 270716 404050 270768
rect 412910 270756 412916 270768
rect 405476 270728 412916 270756
rect 405476 270688 405504 270728
rect 412910 270716 412916 270728
rect 412968 270716 412974 270768
rect 413278 270716 413284 270768
rect 413336 270756 413342 270768
rect 422478 270756 422484 270768
rect 413336 270728 422484 270756
rect 413336 270716 413342 270728
rect 422478 270716 422484 270728
rect 422536 270716 422542 270768
rect 424502 270716 424508 270768
rect 424560 270756 424566 270768
rect 430022 270756 430028 270768
rect 424560 270728 430028 270756
rect 424560 270716 424566 270728
rect 430022 270716 430028 270728
rect 430080 270716 430086 270768
rect 430298 270716 430304 270768
rect 430356 270756 430362 270768
rect 431310 270756 431316 270768
rect 430356 270728 431316 270756
rect 430356 270716 430362 270728
rect 431310 270716 431316 270728
rect 431368 270716 431374 270768
rect 432414 270716 432420 270768
rect 432472 270756 432478 270768
rect 436094 270756 436100 270768
rect 432472 270728 436100 270756
rect 432472 270716 432478 270728
rect 436094 270716 436100 270728
rect 436152 270716 436158 270768
rect 436278 270716 436284 270768
rect 436336 270756 436342 270768
rect 535178 270756 535184 270768
rect 436336 270728 535184 270756
rect 436336 270716 436342 270728
rect 535178 270716 535184 270728
rect 535236 270716 535242 270768
rect 405384 270660 405504 270688
rect 142982 270580 142988 270632
rect 143040 270620 143046 270632
rect 165706 270620 165712 270632
rect 143040 270592 165712 270620
rect 143040 270580 143046 270592
rect 165706 270580 165712 270592
rect 165764 270580 165770 270632
rect 343358 270580 343364 270632
rect 343416 270620 343422 270632
rect 348142 270620 348148 270632
rect 343416 270592 348148 270620
rect 343416 270580 343422 270592
rect 348142 270580 348148 270592
rect 348200 270580 348206 270632
rect 353202 270580 353208 270632
rect 353260 270620 353266 270632
rect 402790 270620 402796 270632
rect 353260 270592 402796 270620
rect 353260 270580 353266 270592
rect 402790 270580 402796 270592
rect 402848 270580 402854 270632
rect 402928 270580 402934 270632
rect 402986 270620 402992 270632
rect 405384 270620 405412 270660
rect 402986 270592 405412 270620
rect 402986 270580 402992 270592
rect 405918 270580 405924 270632
rect 405976 270620 405982 270632
rect 489914 270620 489920 270632
rect 405976 270592 489920 270620
rect 405976 270580 405982 270592
rect 489914 270580 489920 270592
rect 489972 270580 489978 270632
rect 490098 270580 490104 270632
rect 490156 270620 490162 270632
rect 499482 270620 499488 270632
rect 490156 270592 499488 270620
rect 490156 270580 490162 270592
rect 499482 270580 499488 270592
rect 499540 270580 499546 270632
rect 499666 270580 499672 270632
rect 499724 270620 499730 270632
rect 639230 270620 639236 270632
rect 499724 270592 639236 270620
rect 499724 270580 499730 270592
rect 639230 270580 639236 270592
rect 639288 270580 639294 270632
rect 108942 270444 108948 270496
rect 109000 270484 109006 270496
rect 162394 270484 162400 270496
rect 109000 270456 162400 270484
rect 109000 270444 109006 270456
rect 162394 270444 162400 270456
rect 162452 270444 162458 270496
rect 176930 270444 176936 270496
rect 176988 270484 176994 270496
rect 176988 270456 178724 270484
rect 176988 270444 176994 270456
rect 78858 270308 78864 270360
rect 78916 270348 78922 270360
rect 132586 270348 132592 270360
rect 78916 270320 132592 270348
rect 78916 270308 78922 270320
rect 132586 270308 132592 270320
rect 132644 270308 132650 270360
rect 133782 270308 133788 270360
rect 133840 270348 133846 270360
rect 177574 270348 177580 270360
rect 133840 270320 177580 270348
rect 133840 270308 133846 270320
rect 177574 270308 177580 270320
rect 177632 270308 177638 270360
rect 178696 270348 178724 270456
rect 179138 270444 179144 270496
rect 179196 270484 179202 270496
rect 202138 270484 202144 270496
rect 179196 270456 202144 270484
rect 179196 270444 179202 270456
rect 202138 270444 202144 270456
rect 202196 270444 202202 270496
rect 207014 270444 207020 270496
rect 207072 270484 207078 270496
rect 209498 270484 209504 270496
rect 207072 270456 209504 270484
rect 207072 270444 207078 270456
rect 209498 270444 209504 270456
rect 209556 270444 209562 270496
rect 221734 270444 221740 270496
rect 221792 270484 221798 270496
rect 229370 270484 229376 270496
rect 221792 270456 229376 270484
rect 221792 270444 221798 270456
rect 229370 270444 229376 270456
rect 229428 270444 229434 270496
rect 244366 270444 244372 270496
rect 244424 270484 244430 270496
rect 247770 270484 247776 270496
rect 244424 270456 247776 270484
rect 244424 270444 244430 270456
rect 247770 270444 247776 270456
rect 247828 270444 247834 270496
rect 250162 270444 250168 270496
rect 250220 270484 250226 270496
rect 251450 270484 251456 270496
rect 250220 270456 251456 270484
rect 250220 270444 250226 270456
rect 251450 270444 251456 270456
rect 251508 270444 251514 270496
rect 258810 270444 258816 270496
rect 258868 270484 258874 270496
rect 261294 270484 261300 270496
rect 258868 270456 261300 270484
rect 258868 270444 258874 270456
rect 261294 270444 261300 270456
rect 261352 270444 261358 270496
rect 292666 270444 292672 270496
rect 292724 270484 292730 270496
rect 305086 270484 305092 270496
rect 292724 270456 305092 270484
rect 292724 270444 292730 270456
rect 305086 270444 305092 270456
rect 305144 270444 305150 270496
rect 325786 270444 325792 270496
rect 325844 270484 325850 270496
rect 355318 270484 355324 270496
rect 325844 270456 355324 270484
rect 325844 270444 325850 270456
rect 355318 270444 355324 270456
rect 355376 270444 355382 270496
rect 367738 270444 367744 270496
rect 367796 270484 367802 270496
rect 432414 270484 432420 270496
rect 367796 270456 432420 270484
rect 367796 270444 367802 270456
rect 432414 270444 432420 270456
rect 432472 270444 432478 270496
rect 432598 270444 432604 270496
rect 432656 270484 432662 270496
rect 442258 270484 442264 270496
rect 432656 270456 442264 270484
rect 432656 270444 432662 270456
rect 442258 270444 442264 270456
rect 442316 270444 442322 270496
rect 442442 270444 442448 270496
rect 442500 270484 442506 270496
rect 444926 270484 444932 270496
rect 442500 270456 444932 270484
rect 442500 270444 442506 270456
rect 444926 270444 444932 270456
rect 444984 270444 444990 270496
rect 445110 270444 445116 270496
rect 445168 270484 445174 270496
rect 549530 270484 549536 270496
rect 445168 270456 549536 270484
rect 445168 270444 445174 270456
rect 549530 270444 549536 270456
rect 549588 270444 549594 270496
rect 205818 270348 205824 270360
rect 178696 270320 205824 270348
rect 205818 270308 205824 270320
rect 205876 270308 205882 270360
rect 208394 270308 208400 270360
rect 208452 270348 208458 270360
rect 224954 270348 224960 270360
rect 208452 270320 224960 270348
rect 208452 270308 208458 270320
rect 224954 270308 224960 270320
rect 225012 270308 225018 270360
rect 243170 270308 243176 270360
rect 243228 270348 243234 270360
rect 247034 270348 247040 270360
rect 243228 270320 247040 270348
rect 243228 270308 243234 270320
rect 247034 270308 247040 270320
rect 247092 270308 247098 270360
rect 261018 270308 261024 270360
rect 261076 270348 261082 270360
rect 264974 270348 264980 270360
rect 261076 270320 264980 270348
rect 261076 270308 261082 270320
rect 264974 270308 264980 270320
rect 265032 270308 265038 270360
rect 274818 270308 274824 270360
rect 274876 270348 274882 270360
rect 278958 270348 278964 270360
rect 274876 270320 278964 270348
rect 274876 270308 274882 270320
rect 278958 270308 278964 270320
rect 279016 270308 279022 270360
rect 301958 270308 301964 270360
rect 302016 270348 302022 270360
rect 320174 270348 320180 270360
rect 302016 270320 320180 270348
rect 302016 270308 302022 270320
rect 320174 270308 320180 270320
rect 320232 270308 320238 270360
rect 332318 270308 332324 270360
rect 332376 270348 332382 270360
rect 379146 270348 379152 270360
rect 332376 270320 379152 270348
rect 332376 270308 332382 270320
rect 379146 270308 379152 270320
rect 379204 270308 379210 270360
rect 379330 270308 379336 270360
rect 379388 270348 379394 270360
rect 383378 270348 383384 270360
rect 379388 270320 383384 270348
rect 379388 270308 379394 270320
rect 383378 270308 383384 270320
rect 383436 270308 383442 270360
rect 383562 270308 383568 270360
rect 383620 270348 383626 270360
rect 388438 270348 388444 270360
rect 383620 270320 388444 270348
rect 383620 270308 383626 270320
rect 388438 270308 388444 270320
rect 388496 270308 388502 270360
rect 388622 270308 388628 270360
rect 388680 270348 388686 270360
rect 459830 270348 459836 270360
rect 388680 270320 459836 270348
rect 388680 270308 388686 270320
rect 459830 270308 459836 270320
rect 459888 270308 459894 270360
rect 469766 270348 469772 270360
rect 461596 270320 469772 270348
rect 94222 270172 94228 270224
rect 94280 270212 94286 270224
rect 153562 270212 153568 270224
rect 94280 270184 153568 270212
rect 94280 270172 94286 270184
rect 153562 270172 153568 270184
rect 153620 270172 153626 270224
rect 163682 270172 163688 270224
rect 163740 270212 163746 270224
rect 166442 270212 166448 270224
rect 163740 270184 166448 270212
rect 163740 270172 163746 270184
rect 166442 270172 166448 270184
rect 166500 270172 166506 270224
rect 172422 270172 172428 270224
rect 172480 270212 172486 270224
rect 179138 270212 179144 270224
rect 172480 270184 179144 270212
rect 172480 270172 172486 270184
rect 179138 270172 179144 270184
rect 179196 270172 179202 270224
rect 179506 270172 179512 270224
rect 179564 270212 179570 270224
rect 203610 270212 203616 270224
rect 179564 270184 203616 270212
rect 179564 270172 179570 270184
rect 203610 270172 203616 270184
rect 203668 270172 203674 270224
rect 205542 270172 205548 270224
rect 205600 270212 205606 270224
rect 223482 270212 223488 270224
rect 205600 270184 223488 270212
rect 205600 270172 205606 270184
rect 223482 270172 223488 270184
rect 223540 270172 223546 270224
rect 278866 270172 278872 270224
rect 278924 270212 278930 270224
rect 288434 270212 288440 270224
rect 278924 270184 288440 270212
rect 278924 270172 278930 270184
rect 288434 270172 288440 270184
rect 288492 270172 288498 270224
rect 290458 270172 290464 270224
rect 290516 270212 290522 270224
rect 311894 270212 311900 270224
rect 290516 270184 311900 270212
rect 290516 270172 290522 270184
rect 311894 270172 311900 270184
rect 311952 270172 311958 270224
rect 312814 270172 312820 270224
rect 312872 270212 312878 270224
rect 331398 270212 331404 270224
rect 312872 270184 331404 270212
rect 312872 270172 312878 270184
rect 331398 270172 331404 270184
rect 331456 270172 331462 270224
rect 351638 270172 351644 270224
rect 351696 270212 351702 270224
rect 359642 270212 359648 270224
rect 351696 270184 359648 270212
rect 351696 270172 351702 270184
rect 359642 270172 359648 270184
rect 359700 270172 359706 270224
rect 359826 270172 359832 270224
rect 359884 270212 359890 270224
rect 359884 270184 374684 270212
rect 359884 270172 359890 270184
rect 67542 270036 67548 270088
rect 67600 270076 67606 270088
rect 78582 270076 78588 270088
rect 67600 270048 78588 270076
rect 67600 270036 67606 270048
rect 78582 270036 78588 270048
rect 78640 270036 78646 270088
rect 80054 270036 80060 270088
rect 80112 270076 80118 270088
rect 144454 270076 144460 270088
rect 80112 270048 144460 270076
rect 80112 270036 80118 270048
rect 144454 270036 144460 270048
rect 144512 270036 144518 270088
rect 152734 270036 152740 270088
rect 152792 270076 152798 270088
rect 179782 270076 179788 270088
rect 152792 270048 179788 270076
rect 152792 270036 152798 270048
rect 179782 270036 179788 270048
rect 179840 270036 179846 270088
rect 183462 270036 183468 270088
rect 183520 270076 183526 270088
rect 194502 270076 194508 270088
rect 183520 270048 194508 270076
rect 183520 270036 183526 270048
rect 194502 270036 194508 270048
rect 194560 270036 194566 270088
rect 202966 270036 202972 270088
rect 203024 270076 203030 270088
rect 222010 270076 222016 270088
rect 203024 270048 222016 270076
rect 203024 270036 203030 270048
rect 222010 270036 222016 270048
rect 222068 270036 222074 270088
rect 226610 270036 226616 270088
rect 226668 270076 226674 270088
rect 236730 270076 236736 270088
rect 226668 270048 236736 270076
rect 226668 270036 226674 270048
rect 236730 270036 236736 270048
rect 236788 270036 236794 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 273254 270076 273260 270088
rect 266228 270048 273260 270076
rect 266228 270036 266234 270048
rect 273254 270036 273260 270048
rect 273312 270036 273318 270088
rect 276474 270036 276480 270088
rect 276532 270076 276538 270088
rect 289814 270076 289820 270088
rect 276532 270048 289820 270076
rect 276532 270036 276538 270048
rect 289814 270036 289820 270048
rect 289872 270036 289878 270088
rect 297818 270036 297824 270088
rect 297876 270076 297882 270088
rect 324314 270076 324320 270088
rect 297876 270048 324320 270076
rect 297876 270036 297882 270048
rect 324314 270036 324320 270048
rect 324372 270036 324378 270088
rect 334986 270036 334992 270088
rect 335044 270076 335050 270088
rect 374454 270076 374460 270088
rect 335044 270048 374460 270076
rect 335044 270036 335050 270048
rect 374454 270036 374460 270048
rect 374512 270036 374518 270088
rect 374656 270076 374684 270184
rect 374822 270172 374828 270224
rect 374880 270212 374886 270224
rect 376754 270212 376760 270224
rect 374880 270184 376760 270212
rect 374880 270172 374886 270184
rect 376754 270172 376760 270184
rect 376812 270172 376818 270224
rect 376938 270172 376944 270224
rect 376996 270212 377002 270224
rect 405734 270212 405740 270224
rect 376996 270184 405740 270212
rect 376996 270172 377002 270184
rect 405734 270172 405740 270184
rect 405792 270172 405798 270224
rect 405918 270172 405924 270224
rect 405976 270212 405982 270224
rect 406746 270212 406752 270224
rect 405976 270184 406752 270212
rect 405976 270172 405982 270184
rect 406746 270172 406752 270184
rect 406804 270172 406810 270224
rect 407390 270172 407396 270224
rect 407448 270212 407454 270224
rect 407448 270184 407896 270212
rect 407448 270172 407454 270184
rect 393682 270076 393688 270088
rect 374656 270048 393688 270076
rect 393682 270036 393688 270048
rect 393740 270036 393746 270088
rect 397638 270076 397644 270088
rect 395356 270048 397644 270076
rect 75822 269900 75828 269952
rect 75880 269940 75886 269952
rect 141786 269940 141792 269952
rect 75880 269912 141792 269940
rect 75880 269900 75886 269912
rect 141786 269900 141792 269912
rect 141844 269900 141850 269952
rect 143902 269900 143908 269952
rect 143960 269940 143966 269952
rect 184474 269940 184480 269952
rect 143960 269912 184480 269940
rect 143960 269900 143966 269912
rect 184474 269900 184480 269912
rect 184532 269900 184538 269952
rect 191650 269900 191656 269952
rect 191708 269940 191714 269952
rect 211154 269940 211160 269952
rect 191708 269912 211160 269940
rect 191708 269900 191714 269912
rect 211154 269900 211160 269912
rect 211212 269900 211218 269952
rect 212258 269900 212264 269952
rect 212316 269940 212322 269952
rect 219434 269940 219440 269952
rect 212316 269912 219440 269940
rect 212316 269900 212322 269912
rect 219434 269900 219440 269912
rect 219492 269900 219498 269952
rect 219618 269900 219624 269952
rect 219676 269940 219682 269952
rect 227714 269940 227720 269952
rect 219676 269912 227720 269940
rect 219676 269900 219682 269912
rect 227714 269900 227720 269912
rect 227772 269900 227778 269952
rect 230382 269900 230388 269952
rect 230440 269940 230446 269952
rect 238938 269940 238944 269952
rect 230440 269912 238944 269940
rect 230440 269900 230446 269912
rect 238938 269900 238944 269912
rect 238996 269900 239002 269952
rect 266906 269900 266912 269952
rect 266964 269940 266970 269952
rect 274634 269940 274640 269952
rect 266964 269912 274640 269940
rect 266964 269900 266970 269912
rect 274634 269900 274640 269912
rect 274692 269900 274698 269952
rect 275002 269900 275008 269952
rect 275060 269940 275066 269952
rect 287054 269940 287060 269952
rect 275060 269912 287060 269940
rect 275060 269900 275066 269912
rect 287054 269900 287060 269912
rect 287112 269900 287118 269952
rect 287514 269900 287520 269952
rect 287572 269940 287578 269952
rect 307754 269940 307760 269952
rect 287572 269912 307760 269940
rect 287572 269900 287578 269912
rect 307754 269900 307760 269912
rect 307812 269900 307818 269952
rect 310330 269900 310336 269952
rect 310388 269940 310394 269952
rect 338850 269940 338856 269952
rect 310388 269912 338856 269940
rect 310388 269900 310394 269912
rect 338850 269900 338856 269912
rect 338908 269900 338914 269952
rect 339034 269900 339040 269952
rect 339092 269940 339098 269952
rect 359458 269940 359464 269952
rect 339092 269912 359464 269940
rect 339092 269900 339098 269912
rect 359458 269900 359464 269912
rect 359516 269900 359522 269952
rect 359642 269900 359648 269952
rect 359700 269940 359706 269952
rect 395356 269940 395384 270048
rect 397638 270036 397644 270048
rect 397696 270036 397702 270088
rect 398282 270036 398288 270088
rect 398340 270076 398346 270088
rect 407868 270076 407896 270184
rect 408034 270172 408040 270224
rect 408092 270212 408098 270224
rect 408494 270212 408500 270224
rect 408092 270184 408500 270212
rect 408092 270172 408098 270184
rect 408494 270172 408500 270184
rect 408552 270172 408558 270224
rect 408770 270172 408776 270224
rect 408828 270212 408834 270224
rect 442074 270212 442080 270224
rect 408828 270184 442080 270212
rect 408828 270172 408834 270184
rect 442074 270172 442080 270184
rect 442132 270172 442138 270224
rect 442258 270172 442264 270224
rect 442316 270212 442322 270224
rect 461596 270212 461624 270320
rect 469766 270308 469772 270320
rect 469824 270308 469830 270360
rect 469950 270308 469956 270360
rect 470008 270348 470014 270360
rect 474734 270348 474740 270360
rect 470008 270320 474740 270348
rect 470008 270308 470014 270320
rect 474734 270308 474740 270320
rect 474792 270308 474798 270360
rect 474918 270308 474924 270360
rect 474976 270348 474982 270360
rect 599302 270348 599308 270360
rect 474976 270320 599308 270348
rect 474976 270308 474982 270320
rect 599302 270308 599308 270320
rect 599360 270308 599366 270360
rect 442316 270184 461624 270212
rect 442316 270172 442322 270184
rect 461762 270172 461768 270224
rect 461820 270212 461826 270224
rect 582742 270212 582748 270224
rect 461820 270184 582748 270212
rect 461820 270172 461826 270184
rect 582742 270172 582748 270184
rect 582800 270172 582806 270224
rect 620278 270212 620284 270224
rect 605806 270184 620284 270212
rect 408586 270076 408592 270088
rect 398340 270048 407804 270076
rect 407868 270048 408592 270076
rect 398340 270036 398346 270048
rect 359700 269912 395384 269940
rect 359700 269900 359706 269912
rect 395890 269900 395896 269952
rect 395948 269940 395954 269952
rect 407574 269940 407580 269952
rect 395948 269912 407580 269940
rect 395948 269900 395954 269912
rect 407574 269900 407580 269912
rect 407632 269900 407638 269952
rect 407776 269940 407804 270048
rect 408586 270036 408592 270048
rect 408644 270036 408650 270088
rect 408954 270036 408960 270088
rect 409012 270076 409018 270088
rect 499390 270076 499396 270088
rect 409012 270048 499396 270076
rect 409012 270036 409018 270048
rect 499390 270036 499396 270048
rect 499448 270036 499454 270088
rect 499528 270036 499534 270088
rect 499586 270076 499592 270088
rect 605806 270076 605834 270184
rect 620278 270172 620284 270184
rect 620336 270172 620342 270224
rect 626534 270076 626540 270088
rect 499586 270048 605834 270076
rect 619192 270048 626540 270076
rect 499586 270036 499592 270048
rect 407776 269912 480254 269940
rect 69382 269764 69388 269816
rect 69440 269804 69446 269816
rect 138842 269804 138848 269816
rect 69440 269776 138848 269804
rect 69440 269764 69446 269776
rect 138842 269764 138848 269776
rect 138900 269764 138906 269816
rect 140682 269764 140688 269816
rect 140740 269804 140746 269816
rect 173526 269804 173532 269816
rect 140740 269776 173532 269804
rect 140740 269764 140746 269776
rect 173526 269764 173532 269776
rect 173584 269764 173590 269816
rect 195514 269804 195520 269816
rect 173728 269776 195520 269804
rect 122742 269628 122748 269680
rect 122800 269668 122806 269680
rect 122800 269640 166304 269668
rect 122800 269628 122806 269640
rect 84102 269492 84108 269544
rect 84160 269532 84166 269544
rect 126698 269532 126704 269544
rect 84160 269504 126704 269532
rect 84160 269492 84166 269504
rect 126698 269492 126704 269504
rect 126756 269492 126762 269544
rect 126882 269492 126888 269544
rect 126940 269532 126946 269544
rect 166074 269532 166080 269544
rect 126940 269504 166080 269532
rect 126940 269492 126946 269504
rect 166074 269492 166080 269504
rect 166132 269492 166138 269544
rect 166276 269532 166304 269640
rect 166442 269628 166448 269680
rect 166500 269668 166506 269680
rect 173728 269668 173756 269776
rect 195514 269764 195520 269776
rect 195572 269764 195578 269816
rect 195882 269764 195888 269816
rect 195940 269804 195946 269816
rect 216858 269804 216864 269816
rect 195940 269776 216864 269804
rect 195940 269764 195946 269776
rect 216858 269764 216864 269776
rect 216916 269764 216922 269816
rect 223298 269764 223304 269816
rect 223356 269804 223362 269816
rect 234522 269804 234528 269816
rect 223356 269776 234528 269804
rect 223356 269764 223362 269776
rect 234522 269764 234528 269776
rect 234580 269764 234586 269816
rect 237190 269764 237196 269816
rect 237248 269804 237254 269816
rect 243354 269804 243360 269816
rect 237248 269776 243360 269804
rect 237248 269764 237254 269776
rect 243354 269764 243360 269776
rect 243412 269764 243418 269816
rect 261754 269764 261760 269816
rect 261812 269804 261818 269816
rect 263594 269804 263600 269816
rect 261812 269776 263600 269804
rect 261812 269764 261818 269776
rect 263594 269764 263600 269776
rect 263652 269764 263658 269816
rect 265434 269764 265440 269816
rect 265492 269804 265498 269816
rect 271874 269804 271880 269816
rect 265492 269776 271880 269804
rect 265492 269764 265498 269776
rect 271874 269764 271880 269776
rect 271932 269764 271938 269816
rect 283098 269764 283104 269816
rect 283156 269804 283162 269816
rect 300854 269804 300860 269816
rect 283156 269776 300860 269804
rect 283156 269764 283162 269776
rect 300854 269764 300860 269776
rect 300912 269764 300918 269816
rect 306098 269764 306104 269816
rect 306156 269804 306162 269816
rect 335354 269804 335360 269816
rect 306156 269776 335360 269804
rect 306156 269764 306162 269776
rect 335354 269764 335360 269776
rect 335412 269764 335418 269816
rect 337194 269764 337200 269816
rect 337252 269804 337258 269816
rect 383562 269804 383568 269816
rect 337252 269776 383568 269804
rect 337252 269764 337258 269776
rect 383562 269764 383568 269776
rect 383620 269764 383626 269816
rect 383746 269764 383752 269816
rect 383804 269804 383810 269816
rect 383804 269776 398144 269804
rect 383804 269764 383810 269776
rect 166500 269640 173756 269668
rect 166500 269628 166506 269640
rect 173894 269628 173900 269680
rect 173952 269668 173958 269680
rect 179506 269668 179512 269680
rect 173952 269640 179512 269668
rect 173952 269628 173958 269640
rect 179506 269628 179512 269640
rect 179564 269628 179570 269680
rect 179966 269628 179972 269680
rect 180024 269668 180030 269680
rect 189626 269668 189632 269680
rect 180024 269640 189632 269668
rect 180024 269628 180030 269640
rect 189626 269628 189632 269640
rect 189684 269628 189690 269680
rect 197538 269628 197544 269680
rect 197596 269668 197602 269680
rect 205082 269668 205088 269680
rect 197596 269640 205088 269668
rect 197596 269628 197602 269640
rect 205082 269628 205088 269640
rect 205140 269628 205146 269680
rect 271874 269628 271880 269680
rect 271932 269668 271938 269680
rect 281534 269668 281540 269680
rect 271932 269640 281540 269668
rect 271932 269628 271938 269640
rect 281534 269628 281540 269640
rect 281592 269628 281598 269680
rect 313918 269628 313924 269680
rect 313976 269668 313982 269680
rect 338114 269668 338120 269680
rect 313976 269640 338120 269668
rect 313976 269628 313982 269640
rect 338114 269628 338120 269640
rect 338172 269628 338178 269680
rect 341242 269628 341248 269680
rect 341300 269668 341306 269680
rect 359274 269668 359280 269680
rect 341300 269640 359280 269668
rect 341300 269628 341306 269640
rect 359274 269628 359280 269640
rect 359332 269628 359338 269680
rect 359458 269628 359464 269680
rect 359516 269668 359522 269680
rect 373718 269668 373724 269680
rect 359516 269640 373724 269668
rect 359516 269628 359522 269640
rect 373718 269628 373724 269640
rect 373776 269628 373782 269680
rect 397914 269668 397920 269680
rect 373920 269640 397920 269668
rect 171226 269532 171232 269544
rect 166276 269504 171232 269532
rect 171226 269492 171232 269504
rect 171284 269492 171290 269544
rect 173526 269492 173532 269544
rect 173584 269532 173590 269544
rect 182266 269532 182272 269544
rect 173584 269504 182272 269532
rect 173584 269492 173590 269504
rect 182266 269492 182272 269504
rect 182324 269492 182330 269544
rect 310790 269492 310796 269544
rect 310848 269532 310854 269544
rect 327534 269532 327540 269544
rect 310848 269504 327540 269532
rect 310848 269492 310854 269504
rect 327534 269492 327540 269504
rect 327592 269492 327598 269544
rect 330202 269492 330208 269544
rect 330260 269532 330266 269544
rect 372982 269532 372988 269544
rect 330260 269504 372988 269532
rect 330260 269492 330266 269504
rect 372982 269492 372988 269504
rect 373040 269492 373046 269544
rect 373442 269492 373448 269544
rect 373500 269532 373506 269544
rect 373920 269532 373948 269640
rect 397914 269628 397920 269640
rect 397972 269628 397978 269680
rect 398116 269668 398144 269776
rect 398466 269764 398472 269816
rect 398524 269804 398530 269816
rect 476022 269804 476028 269816
rect 398524 269776 476028 269804
rect 398524 269764 398530 269776
rect 476022 269764 476028 269776
rect 476080 269764 476086 269816
rect 477034 269764 477040 269816
rect 477092 269804 477098 269816
rect 480070 269804 480076 269816
rect 477092 269776 480076 269804
rect 477092 269764 477098 269776
rect 480070 269764 480076 269776
rect 480128 269764 480134 269816
rect 480226 269804 480254 269912
rect 480530 269900 480536 269952
rect 480588 269940 480594 269952
rect 488166 269940 488172 269952
rect 480588 269912 488172 269940
rect 480588 269900 480594 269912
rect 488166 269900 488172 269912
rect 488224 269900 488230 269952
rect 488350 269900 488356 269952
rect 488408 269940 488414 269952
rect 494514 269940 494520 269952
rect 488408 269912 494520 269940
rect 488408 269900 488414 269912
rect 494514 269900 494520 269912
rect 494572 269900 494578 269952
rect 619192 269940 619220 270048
rect 626534 270036 626540 270048
rect 626592 270036 626598 270088
rect 494716 269912 619220 269940
rect 484486 269804 484492 269816
rect 480226 269776 484492 269804
rect 484486 269764 484492 269776
rect 484544 269764 484550 269816
rect 486234 269764 486240 269816
rect 486292 269804 486298 269816
rect 494716 269804 494744 269912
rect 620278 269900 620284 269952
rect 620336 269940 620342 269952
rect 630674 269940 630680 269952
rect 620336 269912 630680 269940
rect 620336 269900 620342 269912
rect 630674 269900 630680 269912
rect 630732 269900 630738 269952
rect 486292 269776 494744 269804
rect 486292 269764 486298 269776
rect 494882 269764 494888 269816
rect 494940 269804 494946 269816
rect 499298 269804 499304 269816
rect 494940 269776 499304 269804
rect 494940 269764 494946 269776
rect 499298 269764 499304 269776
rect 499356 269764 499362 269816
rect 499574 269764 499580 269816
rect 499632 269804 499638 269816
rect 619634 269804 619640 269816
rect 499632 269776 619640 269804
rect 499632 269764 499638 269776
rect 619634 269764 619640 269776
rect 619692 269764 619698 269816
rect 636194 269764 636200 269816
rect 636252 269804 636258 269816
rect 647234 269804 647240 269816
rect 636252 269776 647240 269804
rect 636252 269764 636258 269776
rect 647234 269764 647240 269776
rect 647292 269764 647298 269816
rect 407390 269668 407396 269680
rect 398116 269640 407396 269668
rect 407390 269628 407396 269640
rect 407448 269628 407454 269680
rect 407574 269628 407580 269680
rect 407632 269668 407638 269680
rect 413462 269668 413468 269680
rect 407632 269640 413468 269668
rect 407632 269628 407638 269640
rect 413462 269628 413468 269640
rect 413520 269628 413526 269680
rect 414106 269628 414112 269680
rect 414164 269668 414170 269680
rect 509050 269668 509056 269680
rect 414164 269640 509056 269668
rect 414164 269628 414170 269640
rect 509050 269628 509056 269640
rect 509108 269628 509114 269680
rect 509234 269628 509240 269680
rect 509292 269668 509298 269680
rect 633618 269668 633624 269680
rect 509292 269640 633624 269668
rect 509292 269628 509298 269640
rect 633618 269628 633624 269640
rect 633676 269628 633682 269680
rect 373500 269504 373948 269532
rect 373500 269492 373506 269504
rect 375190 269492 375196 269544
rect 375248 269532 375254 269544
rect 384114 269532 384120 269544
rect 375248 269504 384120 269532
rect 375248 269492 375254 269504
rect 384114 269492 384120 269504
rect 384172 269492 384178 269544
rect 384482 269492 384488 269544
rect 384540 269532 384546 269544
rect 388622 269532 388628 269544
rect 384540 269504 388628 269532
rect 384540 269492 384546 269504
rect 388622 269492 388628 269504
rect 388680 269492 388686 269544
rect 388990 269492 388996 269544
rect 389048 269532 389054 269544
rect 390554 269532 390560 269544
rect 389048 269504 390560 269532
rect 389048 269492 389054 269504
rect 390554 269492 390560 269504
rect 390612 269492 390618 269544
rect 391290 269492 391296 269544
rect 391348 269532 391354 269544
rect 469582 269532 469588 269544
rect 391348 269504 469588 269532
rect 391348 269492 391354 269504
rect 469582 269492 469588 269504
rect 469640 269492 469646 269544
rect 469766 269492 469772 269544
rect 469824 269532 469830 269544
rect 481634 269532 481640 269544
rect 469824 269504 481640 269532
rect 469824 269492 469830 269504
rect 481634 269492 481640 269504
rect 481692 269492 481698 269544
rect 484302 269492 484308 269544
rect 484360 269532 484366 269544
rect 489730 269532 489736 269544
rect 484360 269504 489736 269532
rect 484360 269492 484366 269504
rect 489730 269492 489736 269504
rect 489788 269492 489794 269544
rect 489914 269492 489920 269544
rect 489972 269532 489978 269544
rect 590654 269532 590660 269544
rect 489972 269504 590660 269532
rect 489972 269492 489978 269504
rect 590654 269492 590660 269504
rect 590712 269492 590718 269544
rect 259730 269424 259736 269476
rect 259788 269464 259794 269476
rect 260834 269464 260840 269476
rect 259788 269436 260840 269464
rect 259788 269424 259794 269436
rect 260834 269424 260840 269436
rect 260892 269424 260898 269476
rect 129366 269356 129372 269408
rect 129424 269396 129430 269408
rect 175642 269396 175648 269408
rect 129424 269368 175648 269396
rect 129424 269356 129430 269368
rect 175642 269356 175648 269368
rect 175700 269356 175706 269408
rect 354766 269356 354772 269408
rect 354824 269396 354830 269408
rect 393682 269396 393688 269408
rect 354824 269368 393688 269396
rect 354824 269356 354830 269368
rect 393682 269356 393688 269368
rect 393740 269356 393746 269408
rect 393866 269356 393872 269408
rect 393924 269396 393930 269408
rect 398466 269396 398472 269408
rect 393924 269368 398472 269396
rect 393924 269356 393930 269368
rect 398466 269356 398472 269368
rect 398524 269356 398530 269408
rect 398926 269356 398932 269408
rect 398984 269396 398990 269408
rect 401778 269396 401784 269408
rect 398984 269368 401784 269396
rect 398984 269356 398990 269368
rect 401778 269356 401784 269368
rect 401836 269356 401842 269408
rect 401962 269356 401968 269408
rect 402020 269396 402026 269408
rect 402020 269368 413324 269396
rect 402020 269356 402026 269368
rect 264698 269288 264704 269340
rect 264756 269328 264762 269340
rect 265894 269328 265900 269340
rect 264756 269300 265900 269328
rect 264756 269288 264762 269300
rect 265894 269288 265900 269300
rect 265952 269288 265958 269340
rect 128538 269220 128544 269272
rect 128596 269260 128602 269272
rect 163590 269260 163596 269272
rect 128596 269232 163596 269260
rect 128596 269220 128602 269232
rect 163590 269220 163596 269232
rect 163648 269220 163654 269272
rect 166074 269220 166080 269272
rect 166132 269260 166138 269272
rect 173434 269260 173440 269272
rect 166132 269232 173440 269260
rect 166132 269220 166138 269232
rect 173434 269220 173440 269232
rect 173492 269220 173498 269272
rect 327994 269220 328000 269272
rect 328052 269260 328058 269272
rect 372614 269260 372620 269272
rect 328052 269232 372620 269260
rect 328052 269220 328058 269232
rect 372614 269220 372620 269232
rect 372672 269220 372678 269272
rect 372982 269220 372988 269272
rect 373040 269260 373046 269272
rect 374270 269260 374276 269272
rect 373040 269232 374276 269260
rect 373040 269220 373046 269232
rect 374270 269220 374276 269232
rect 374328 269220 374334 269272
rect 383930 269260 383936 269272
rect 383626 269232 383936 269260
rect 374454 269152 374460 269204
rect 374512 269192 374518 269204
rect 383626 269192 383654 269232
rect 383930 269220 383936 269232
rect 383988 269220 383994 269272
rect 388438 269220 388444 269272
rect 388496 269260 388502 269272
rect 408448 269260 408454 269272
rect 388496 269232 408454 269260
rect 388496 269220 388502 269232
rect 408448 269220 408454 269232
rect 408506 269220 408512 269272
rect 408678 269220 408684 269272
rect 408736 269260 408742 269272
rect 412634 269260 412640 269272
rect 408736 269232 412640 269260
rect 408736 269220 408742 269232
rect 412634 269220 412640 269232
rect 412692 269220 412698 269272
rect 413296 269260 413324 269368
rect 413462 269356 413468 269408
rect 413520 269396 413526 269408
rect 432598 269396 432604 269408
rect 413520 269368 432604 269396
rect 413520 269356 413526 269368
rect 432598 269356 432604 269368
rect 432656 269356 432662 269408
rect 432782 269356 432788 269408
rect 432840 269396 432846 269408
rect 535454 269396 535460 269408
rect 432840 269368 535460 269396
rect 432840 269356 432846 269368
rect 535454 269356 535460 269368
rect 535512 269356 535518 269408
rect 423674 269260 423680 269272
rect 413296 269232 423680 269260
rect 423674 269220 423680 269232
rect 423732 269220 423738 269272
rect 423858 269220 423864 269272
rect 423916 269260 423922 269272
rect 521654 269260 521660 269272
rect 423916 269232 521660 269260
rect 423916 269220 423922 269232
rect 521654 269220 521660 269232
rect 521712 269220 521718 269272
rect 374512 269164 383654 269192
rect 374512 269152 374518 269164
rect 384114 269152 384120 269204
rect 384172 269192 384178 269204
rect 384482 269192 384488 269204
rect 384172 269164 384488 269192
rect 384172 269152 384178 269164
rect 384482 269152 384488 269164
rect 384540 269152 384546 269204
rect 248322 269084 248328 269136
rect 248380 269124 248386 269136
rect 249978 269124 249984 269136
rect 248380 269096 249984 269124
rect 248380 269084 248386 269096
rect 249978 269084 249984 269096
rect 250036 269084 250042 269136
rect 42426 269016 42432 269068
rect 42484 269056 42490 269068
rect 45554 269056 45560 269068
rect 42484 269028 45560 269056
rect 42484 269016 42490 269028
rect 45554 269016 45560 269028
rect 45612 269016 45618 269068
rect 118602 269016 118608 269068
rect 118660 269056 118666 269068
rect 169754 269056 169760 269068
rect 118660 269028 169760 269056
rect 118660 269016 118666 269028
rect 169754 269016 169760 269028
rect 169812 269016 169818 269068
rect 225414 269016 225420 269068
rect 225472 269056 225478 269068
rect 226334 269056 226340 269068
rect 225472 269028 226340 269056
rect 225472 269016 225478 269028
rect 226334 269016 226340 269028
rect 226392 269016 226398 269068
rect 324314 269016 324320 269068
rect 324372 269056 324378 269068
rect 336734 269056 336740 269068
rect 324372 269028 336740 269056
rect 324372 269016 324378 269028
rect 336734 269016 336740 269028
rect 336792 269016 336798 269068
rect 339402 269016 339408 269068
rect 339460 269056 339466 269068
rect 358906 269056 358912 269068
rect 339460 269028 358912 269056
rect 339460 269016 339466 269028
rect 358906 269016 358912 269028
rect 358964 269016 358970 269068
rect 375834 269016 375840 269068
rect 375892 269056 375898 269068
rect 407758 269056 407764 269068
rect 375892 269028 407764 269056
rect 375892 269016 375898 269028
rect 407758 269016 407764 269028
rect 407816 269016 407822 269068
rect 407942 269016 407948 269068
rect 408000 269056 408006 269068
rect 408000 269028 432644 269056
rect 408000 269016 408006 269028
rect 104894 268880 104900 268932
rect 104952 268920 104958 268932
rect 160186 268920 160192 268932
rect 104952 268892 160192 268920
rect 104952 268880 104958 268892
rect 160186 268880 160192 268892
rect 160244 268880 160250 268932
rect 203886 268880 203892 268932
rect 203944 268920 203950 268932
rect 203944 268892 209774 268920
rect 203944 268880 203950 268892
rect 209746 268852 209774 268892
rect 269114 268880 269120 268932
rect 269172 268920 269178 268932
rect 276658 268920 276664 268932
rect 269172 268892 276664 268920
rect 269172 268880 269178 268892
rect 276658 268880 276664 268892
rect 276716 268880 276722 268932
rect 299290 268880 299296 268932
rect 299348 268920 299354 268932
rect 319622 268920 319628 268932
rect 299348 268892 319628 268920
rect 299348 268880 299354 268892
rect 319622 268880 319628 268892
rect 319680 268880 319686 268932
rect 319806 268880 319812 268932
rect 319864 268920 319870 268932
rect 345198 268920 345204 268932
rect 319864 268892 345204 268920
rect 319864 268880 319870 268892
rect 345198 268880 345204 268892
rect 345256 268880 345262 268932
rect 349338 268880 349344 268932
rect 349396 268920 349402 268932
rect 349396 268892 354674 268920
rect 349396 268880 349402 268892
rect 209866 268852 209872 268864
rect 209746 268824 209872 268852
rect 209866 268812 209872 268824
rect 209924 268812 209930 268864
rect 77202 268744 77208 268796
rect 77260 268784 77266 268796
rect 104894 268784 104900 268796
rect 77260 268756 104900 268784
rect 77260 268744 77266 268756
rect 104894 268744 104900 268756
rect 104952 268744 104958 268796
rect 106274 268744 106280 268796
rect 106332 268784 106338 268796
rect 161658 268784 161664 268796
rect 106332 268756 161664 268784
rect 106332 268744 106338 268756
rect 161658 268744 161664 268756
rect 161716 268744 161722 268796
rect 187602 268744 187608 268796
rect 187660 268784 187666 268796
rect 208486 268784 208492 268796
rect 187660 268756 208492 268784
rect 187660 268744 187666 268756
rect 208486 268744 208492 268756
rect 208544 268744 208550 268796
rect 316954 268744 316960 268796
rect 317012 268784 317018 268796
rect 353386 268784 353392 268796
rect 317012 268756 353392 268784
rect 317012 268744 317018 268756
rect 353386 268744 353392 268756
rect 353444 268744 353450 268796
rect 354646 268784 354674 268892
rect 358538 268880 358544 268932
rect 358596 268920 358602 268932
rect 369302 268920 369308 268932
rect 358596 268892 369308 268920
rect 358596 268880 358602 268892
rect 369302 268880 369308 268892
rect 369360 268880 369366 268932
rect 369486 268880 369492 268932
rect 369544 268920 369550 268932
rect 432616 268920 432644 269028
rect 432782 269016 432788 269068
rect 432840 269056 432846 269068
rect 449894 269056 449900 269068
rect 432840 269028 449900 269056
rect 432840 269016 432846 269028
rect 449894 269016 449900 269028
rect 449952 269016 449958 269068
rect 453114 269016 453120 269068
rect 453172 269056 453178 269068
rect 453172 269028 461624 269056
rect 453172 269016 453178 269028
rect 441338 268920 441344 268932
rect 369544 268892 432552 268920
rect 432616 268892 441344 268920
rect 369544 268880 369550 268892
rect 354646 268756 364334 268784
rect 95418 268608 95424 268660
rect 95476 268648 95482 268660
rect 155034 268648 155040 268660
rect 95476 268620 155040 268648
rect 95476 268608 95482 268620
rect 155034 268608 155040 268620
rect 155092 268608 155098 268660
rect 162578 268608 162584 268660
rect 162636 268648 162642 268660
rect 190086 268648 190092 268660
rect 162636 268620 190092 268648
rect 162636 268608 162642 268620
rect 190086 268608 190092 268620
rect 190144 268608 190150 268660
rect 190362 268608 190368 268660
rect 190420 268648 190426 268660
rect 203334 268648 203340 268660
rect 190420 268620 203340 268648
rect 190420 268608 190426 268620
rect 203334 268608 203340 268620
rect 203392 268608 203398 268660
rect 273530 268608 273536 268660
rect 273588 268648 273594 268660
rect 282914 268648 282920 268660
rect 273588 268620 282920 268648
rect 273588 268608 273594 268620
rect 282914 268608 282920 268620
rect 282972 268608 282978 268660
rect 294874 268608 294880 268660
rect 294932 268648 294938 268660
rect 317138 268648 317144 268660
rect 294932 268620 317144 268648
rect 294932 268608 294938 268620
rect 317138 268608 317144 268620
rect 317196 268608 317202 268660
rect 329466 268608 329472 268660
rect 329524 268648 329530 268660
rect 340874 268648 340880 268660
rect 329524 268620 340880 268648
rect 329524 268608 329530 268620
rect 340874 268608 340880 268620
rect 340932 268608 340938 268660
rect 353754 268608 353760 268660
rect 353812 268648 353818 268660
rect 364306 268648 364334 268756
rect 364794 268744 364800 268796
rect 364852 268784 364858 268796
rect 432230 268784 432236 268796
rect 364852 268756 432236 268784
rect 364852 268744 364858 268756
rect 432230 268744 432236 268756
rect 432288 268744 432294 268796
rect 432524 268784 432552 268892
rect 441338 268880 441344 268892
rect 441396 268880 441402 268932
rect 447042 268920 447048 268932
rect 441540 268892 447048 268920
rect 437014 268784 437020 268796
rect 432524 268756 437020 268784
rect 437014 268744 437020 268756
rect 437072 268744 437078 268796
rect 437382 268744 437388 268796
rect 437440 268784 437446 268796
rect 441540 268784 441568 268892
rect 447042 268880 447048 268892
rect 447100 268880 447106 268932
rect 452378 268880 452384 268932
rect 452436 268920 452442 268932
rect 455598 268920 455604 268932
rect 452436 268892 455604 268920
rect 452436 268880 452442 268892
rect 455598 268880 455604 268892
rect 455656 268880 455662 268932
rect 456794 268880 456800 268932
rect 456852 268920 456858 268932
rect 460014 268920 460020 268932
rect 456852 268892 460020 268920
rect 456852 268880 456858 268892
rect 460014 268880 460020 268892
rect 460072 268880 460078 268932
rect 461394 268880 461400 268932
rect 461452 268880 461458 268932
rect 452654 268784 452660 268796
rect 437440 268756 441568 268784
rect 441632 268756 452660 268784
rect 437440 268744 437446 268756
rect 369946 268648 369952 268660
rect 353812 268620 359504 268648
rect 364306 268620 369952 268648
rect 353812 268608 353818 268620
rect 87138 268472 87144 268524
rect 87196 268512 87202 268524
rect 149882 268512 149888 268524
rect 87196 268484 149888 268512
rect 87196 268472 87202 268484
rect 149882 268472 149888 268484
rect 149940 268472 149946 268524
rect 162762 268472 162768 268524
rect 162820 268512 162826 268524
rect 196986 268512 196992 268524
rect 162820 268484 196992 268512
rect 162820 268472 162826 268484
rect 196986 268472 196992 268484
rect 197044 268472 197050 268524
rect 208854 268472 208860 268524
rect 208912 268512 208918 268524
rect 225690 268512 225696 268524
rect 208912 268484 225696 268512
rect 208912 268472 208918 268484
rect 225690 268472 225696 268484
rect 225748 268472 225754 268524
rect 282362 268472 282368 268524
rect 282420 268512 282426 268524
rect 295334 268512 295340 268524
rect 282420 268484 295340 268512
rect 282420 268472 282426 268484
rect 295334 268472 295340 268484
rect 295392 268472 295398 268524
rect 297082 268472 297088 268524
rect 297140 268512 297146 268524
rect 322934 268512 322940 268524
rect 297140 268484 322940 268512
rect 297140 268472 297146 268484
rect 322934 268472 322940 268484
rect 322992 268472 322998 268524
rect 324682 268472 324688 268524
rect 324740 268512 324746 268524
rect 359274 268512 359280 268524
rect 324740 268484 359280 268512
rect 324740 268472 324746 268484
rect 359274 268472 359280 268484
rect 359332 268472 359338 268524
rect 359476 268512 359504 268620
rect 369946 268608 369952 268620
rect 370004 268608 370010 268660
rect 374638 268608 374644 268660
rect 374696 268648 374702 268660
rect 385034 268648 385040 268660
rect 374696 268620 385040 268648
rect 374696 268608 374702 268620
rect 385034 268608 385040 268620
rect 385092 268608 385098 268660
rect 388346 268608 388352 268660
rect 388404 268648 388410 268660
rect 441632 268648 441660 268756
rect 452654 268744 452660 268756
rect 452712 268744 452718 268796
rect 461412 268784 461440 268880
rect 461596 268852 461624 269028
rect 461762 269016 461768 269068
rect 461820 269056 461826 269068
rect 572714 269056 572720 269068
rect 461820 269028 572720 269056
rect 461820 269016 461826 269028
rect 572714 269016 572720 269028
rect 572772 269016 572778 269068
rect 461854 268880 461860 268932
rect 461912 268920 461918 268932
rect 576854 268920 576860 268932
rect 461912 268892 576860 268920
rect 461912 268880 461918 268892
rect 576854 268880 576860 268892
rect 576912 268880 576918 268932
rect 461596 268824 461716 268852
rect 455432 268756 461440 268784
rect 388404 268620 441660 268648
rect 388404 268608 388410 268620
rect 442074 268608 442080 268660
rect 442132 268648 442138 268660
rect 455432 268648 455460 268756
rect 442132 268620 455460 268648
rect 442132 268608 442138 268620
rect 455598 268608 455604 268660
rect 455656 268648 455662 268660
rect 461394 268648 461400 268660
rect 455656 268620 461400 268648
rect 455656 268608 455662 268620
rect 461394 268608 461400 268620
rect 461452 268608 461458 268660
rect 461688 268648 461716 268824
rect 462130 268744 462136 268796
rect 462188 268784 462194 268796
rect 466408 268784 466414 268796
rect 462188 268756 466414 268784
rect 462188 268744 462194 268756
rect 466408 268744 466414 268756
rect 466466 268744 466472 268796
rect 467006 268744 467012 268796
rect 467064 268784 467070 268796
rect 583846 268784 583852 268796
rect 467064 268756 583852 268784
rect 467064 268744 467070 268756
rect 583846 268744 583852 268756
rect 583904 268744 583910 268796
rect 466270 268648 466276 268660
rect 461688 268620 466276 268648
rect 466270 268608 466276 268620
rect 466328 268608 466334 268660
rect 466822 268608 466828 268660
rect 466880 268648 466886 268660
rect 499390 268648 499396 268660
rect 466880 268620 499396 268648
rect 466880 268608 466886 268620
rect 499390 268608 499396 268620
rect 499448 268608 499454 268660
rect 499528 268608 499534 268660
rect 499586 268648 499592 268660
rect 580994 268648 581000 268660
rect 499586 268620 581000 268648
rect 499586 268608 499592 268620
rect 580994 268608 581000 268620
rect 581052 268608 581058 268660
rect 359476 268484 379514 268512
rect 82722 268336 82728 268388
rect 82780 268376 82786 268388
rect 146938 268376 146944 268388
rect 82780 268348 146944 268376
rect 82780 268336 82786 268348
rect 146938 268336 146944 268348
rect 146996 268336 147002 268388
rect 148870 268336 148876 268388
rect 148928 268376 148934 268388
rect 187878 268376 187884 268388
rect 148928 268348 187884 268376
rect 148928 268336 148934 268348
rect 187878 268336 187884 268348
rect 187936 268336 187942 268388
rect 188062 268336 188068 268388
rect 188120 268376 188126 268388
rect 188120 268348 200114 268376
rect 188120 268336 188126 268348
rect 115842 268200 115848 268252
rect 115900 268240 115906 268252
rect 166810 268240 166816 268252
rect 115900 268212 166816 268240
rect 115900 268200 115906 268212
rect 166810 268200 166816 268212
rect 166868 268200 166874 268252
rect 200086 268240 200114 268348
rect 210878 268336 210884 268388
rect 210936 268376 210942 268388
rect 219802 268376 219808 268388
rect 210936 268348 219808 268376
rect 210936 268336 210942 268348
rect 219802 268336 219808 268348
rect 219860 268336 219866 268388
rect 220722 268336 220728 268388
rect 220780 268376 220786 268388
rect 233050 268376 233056 268388
rect 220780 268348 233056 268376
rect 220780 268336 220786 268348
rect 233050 268336 233056 268348
rect 233108 268336 233114 268388
rect 281626 268336 281632 268388
rect 281684 268376 281690 268388
rect 298094 268376 298100 268388
rect 281684 268348 298100 268376
rect 281684 268336 281690 268348
rect 298094 268336 298100 268348
rect 298152 268336 298158 268388
rect 304166 268336 304172 268388
rect 304224 268376 304230 268388
rect 329834 268376 329840 268388
rect 304224 268348 329840 268376
rect 304224 268336 304230 268348
rect 329834 268336 329840 268348
rect 329892 268336 329898 268388
rect 342162 268336 342168 268388
rect 342220 268376 342226 268388
rect 374638 268376 374644 268388
rect 342220 268348 374644 268376
rect 342220 268336 342226 268348
rect 374638 268336 374644 268348
rect 374696 268336 374702 268388
rect 379486 268376 379514 268484
rect 382458 268472 382464 268524
rect 382516 268512 382522 268524
rect 455138 268512 455144 268524
rect 382516 268484 455144 268512
rect 382516 268472 382522 268484
rect 455138 268472 455144 268484
rect 455196 268472 455202 268524
rect 455322 268472 455328 268524
rect 455380 268512 455386 268524
rect 461762 268512 461768 268524
rect 455380 268484 461768 268512
rect 455380 268472 455386 268484
rect 461762 268472 461768 268484
rect 461820 268472 461826 268524
rect 461946 268472 461952 268524
rect 462004 268512 462010 268524
rect 480070 268512 480076 268524
rect 462004 268484 480076 268512
rect 462004 268472 462010 268484
rect 480070 268472 480076 268484
rect 480128 268472 480134 268524
rect 594794 268512 594800 268524
rect 480226 268484 594800 268512
rect 382826 268376 382832 268388
rect 379486 268348 382832 268376
rect 382826 268336 382832 268348
rect 382884 268336 382890 268388
rect 387610 268336 387616 268388
rect 387668 268376 387674 268388
rect 462130 268376 462136 268388
rect 387668 268348 462136 268376
rect 387668 268336 387674 268348
rect 462130 268336 462136 268348
rect 462188 268336 462194 268388
rect 462314 268336 462320 268388
rect 462372 268376 462378 268388
rect 466546 268376 466552 268388
rect 462372 268348 466552 268376
rect 462372 268336 462378 268348
rect 466546 268336 466552 268348
rect 466604 268336 466610 268388
rect 466730 268336 466736 268388
rect 466788 268376 466794 268388
rect 480226 268376 480254 268484
rect 594794 268472 594800 268484
rect 594852 268472 594858 268524
rect 601602 268472 601608 268524
rect 601660 268512 601666 268524
rect 645854 268512 645860 268524
rect 601660 268484 645860 268512
rect 601660 268472 601666 268484
rect 645854 268472 645860 268484
rect 645912 268472 645918 268524
rect 466788 268348 480254 268376
rect 466788 268336 466794 268348
rect 480346 268336 480352 268388
rect 480404 268376 480410 268388
rect 608870 268376 608876 268388
rect 480404 268348 608876 268376
rect 480404 268336 480410 268348
rect 608870 268336 608876 268348
rect 608928 268336 608934 268388
rect 210970 268240 210976 268252
rect 200086 268212 210976 268240
rect 210970 268200 210976 268212
rect 211028 268200 211034 268252
rect 317690 268200 317696 268252
rect 317748 268240 317754 268252
rect 356054 268240 356060 268252
rect 317748 268212 356060 268240
rect 317748 268200 317754 268212
rect 356054 268200 356060 268212
rect 356112 268200 356118 268252
rect 359274 268200 359280 268252
rect 359332 268240 359338 268252
rect 367186 268240 367192 268252
rect 359332 268212 367192 268240
rect 359332 268200 359338 268212
rect 367186 268200 367192 268212
rect 367244 268200 367250 268252
rect 413094 268240 413100 268252
rect 369136 268212 413100 268240
rect 135254 268064 135260 268116
rect 135312 268104 135318 268116
rect 138106 268104 138112 268116
rect 135312 268076 138112 268104
rect 135312 268064 135318 268076
rect 138106 268064 138112 268076
rect 138164 268064 138170 268116
rect 147490 268064 147496 268116
rect 147548 268104 147554 268116
rect 186682 268104 186688 268116
rect 147548 268076 186688 268104
rect 147548 268064 147554 268076
rect 186682 268064 186688 268076
rect 186740 268064 186746 268116
rect 360378 268064 360384 268116
rect 360436 268104 360442 268116
rect 369136 268104 369164 268212
rect 413094 268200 413100 268212
rect 413152 268200 413158 268252
rect 432414 268240 432420 268252
rect 413296 268212 432420 268240
rect 360436 268076 369164 268104
rect 360436 268064 360442 268076
rect 369302 268064 369308 268116
rect 369360 268104 369366 268116
rect 407298 268104 407304 268116
rect 369360 268076 407304 268104
rect 369360 268064 369366 268076
rect 407298 268064 407304 268076
rect 407356 268064 407362 268116
rect 407758 268064 407764 268116
rect 407816 268104 407822 268116
rect 413296 268104 413324 268212
rect 432414 268200 432420 268212
rect 432472 268200 432478 268252
rect 432598 268200 432604 268252
rect 432656 268240 432662 268252
rect 442074 268240 442080 268252
rect 432656 268212 442080 268240
rect 432656 268200 432662 268212
rect 442074 268200 442080 268212
rect 442132 268200 442138 268252
rect 547874 268240 547880 268252
rect 442276 268212 547880 268240
rect 407816 268076 413324 268104
rect 407816 268064 407822 268076
rect 413462 268064 413468 268116
rect 413520 268104 413526 268116
rect 416682 268104 416688 268116
rect 413520 268076 416688 268104
rect 413520 268064 413526 268076
rect 416682 268064 416688 268076
rect 416740 268064 416746 268116
rect 416866 268064 416872 268116
rect 416924 268104 416930 268116
rect 437014 268104 437020 268116
rect 416924 268076 437020 268104
rect 416924 268064 416930 268076
rect 437014 268064 437020 268076
rect 437072 268064 437078 268116
rect 437198 268064 437204 268116
rect 437256 268104 437262 268116
rect 442276 268104 442304 268212
rect 547874 268200 547880 268212
rect 547932 268200 547938 268252
rect 664438 268132 664444 268184
rect 664496 268172 664502 268184
rect 675294 268172 675300 268184
rect 664496 268144 675300 268172
rect 664496 268132 664502 268144
rect 675294 268132 675300 268144
rect 675352 268132 675358 268184
rect 437256 268076 442304 268104
rect 437256 268064 437262 268076
rect 442442 268064 442448 268116
rect 442500 268104 442506 268116
rect 541250 268104 541256 268116
rect 442500 268076 541256 268104
rect 442500 268064 442506 268076
rect 541250 268064 541256 268076
rect 541308 268064 541314 268116
rect 659286 267996 659292 268048
rect 659344 268036 659350 268048
rect 668946 268036 668952 268048
rect 659344 268008 668952 268036
rect 659344 267996 659350 268008
rect 668946 267996 668952 268008
rect 669004 267996 669010 268048
rect 675478 268036 675484 268048
rect 669286 268008 675484 268036
rect 158714 267928 158720 267980
rect 158772 267968 158778 267980
rect 180794 267968 180800 267980
rect 158772 267940 180800 267968
rect 158772 267928 158778 267940
rect 180794 267928 180800 267940
rect 180852 267928 180858 267980
rect 365806 267928 365812 267980
rect 365864 267968 365870 267980
rect 365864 267940 393314 267968
rect 365864 267928 365870 267940
rect 347130 267792 347136 267844
rect 347188 267832 347194 267844
rect 376110 267832 376116 267844
rect 347188 267804 376116 267832
rect 347188 267792 347194 267804
rect 376110 267792 376116 267804
rect 376168 267792 376174 267844
rect 378042 267792 378048 267844
rect 378100 267832 378106 267844
rect 388346 267832 388352 267844
rect 378100 267804 388352 267832
rect 378100 267792 378106 267804
rect 388346 267792 388352 267804
rect 388404 267792 388410 267844
rect 390094 267792 390100 267844
rect 390152 267832 390158 267844
rect 391934 267832 391940 267844
rect 390152 267804 391940 267832
rect 390152 267792 390158 267804
rect 391934 267792 391940 267804
rect 391992 267792 391998 267844
rect 393286 267832 393314 267940
rect 396166 267928 396172 267980
rect 396224 267968 396230 267980
rect 407942 267968 407948 267980
rect 396224 267940 407948 267968
rect 396224 267928 396230 267940
rect 407942 267928 407948 267940
rect 408000 267928 408006 267980
rect 411162 267928 411168 267980
rect 411220 267968 411226 267980
rect 412910 267968 412916 267980
rect 411220 267940 412916 267968
rect 411220 267928 411226 267940
rect 412910 267928 412916 267940
rect 412968 267928 412974 267980
rect 413094 267928 413100 267980
rect 413152 267968 413158 267980
rect 418522 267968 418528 267980
rect 413152 267940 418528 267968
rect 413152 267928 413158 267940
rect 418522 267928 418528 267940
rect 418580 267928 418586 267980
rect 422938 267928 422944 267980
rect 422996 267968 423002 267980
rect 424870 267968 424876 267980
rect 422996 267940 424876 267968
rect 422996 267928 423002 267940
rect 424870 267928 424876 267940
rect 424928 267928 424934 267980
rect 428458 267928 428464 267980
rect 428516 267968 428522 267980
rect 524690 267968 524696 267980
rect 428516 267940 524696 267968
rect 428516 267928 428522 267940
rect 524690 267928 524696 267940
rect 524748 267928 524754 267980
rect 427740 267872 427860 267900
rect 404354 267832 404360 267844
rect 393286 267804 404360 267832
rect 404354 267792 404360 267804
rect 404412 267792 404418 267844
rect 407298 267792 407304 267844
rect 407356 267832 407362 267844
rect 410886 267832 410892 267844
rect 407356 267804 410892 267832
rect 407356 267792 407362 267804
rect 410886 267792 410892 267804
rect 410944 267792 410950 267844
rect 412634 267792 412640 267844
rect 412692 267832 412698 267844
rect 415486 267832 415492 267844
rect 412692 267804 415492 267832
rect 412692 267792 412698 267804
rect 415486 267792 415492 267804
rect 415544 267792 415550 267844
rect 415670 267792 415676 267844
rect 415728 267832 415734 267844
rect 415728 267804 417924 267832
rect 415728 267792 415734 267804
rect 263962 267724 263968 267776
rect 264020 267764 264026 267776
rect 269574 267764 269580 267776
rect 264020 267736 269580 267764
rect 264020 267724 264026 267736
rect 269574 267724 269580 267736
rect 269632 267724 269638 267776
rect 42610 267656 42616 267708
rect 42668 267696 42674 267708
rect 47210 267696 47216 267708
rect 42668 267668 47216 267696
rect 42668 267656 42674 267668
rect 47210 267656 47216 267668
rect 47268 267656 47274 267708
rect 132402 267656 132408 267708
rect 132460 267696 132466 267708
rect 178586 267696 178592 267708
rect 132460 267668 178592 267696
rect 132460 267656 132466 267668
rect 178586 267656 178592 267668
rect 178644 267656 178650 267708
rect 213178 267656 213184 267708
rect 213236 267696 213242 267708
rect 220538 267696 220544 267708
rect 213236 267668 220544 267696
rect 213236 267656 213242 267668
rect 220538 267656 220544 267668
rect 220596 267656 220602 267708
rect 305914 267656 305920 267708
rect 305972 267696 305978 267708
rect 324314 267696 324320 267708
rect 305972 267668 324320 267696
rect 305972 267656 305978 267668
rect 324314 267656 324320 267668
rect 324372 267656 324378 267708
rect 333882 267656 333888 267708
rect 333940 267696 333946 267708
rect 353938 267696 353944 267708
rect 333940 267668 353944 267696
rect 333940 267656 333946 267668
rect 353938 267656 353944 267668
rect 353996 267656 354002 267708
rect 357434 267656 357440 267708
rect 357492 267696 357498 267708
rect 365990 267696 365996 267708
rect 357492 267668 365996 267696
rect 357492 267656 357498 267668
rect 365990 267656 365996 267668
rect 366048 267656 366054 267708
rect 373442 267696 373448 267708
rect 368032 267668 373448 267696
rect 100662 267520 100668 267572
rect 100720 267560 100726 267572
rect 158714 267560 158720 267572
rect 100720 267532 158720 267560
rect 100720 267520 100726 267532
rect 158714 267520 158720 267532
rect 158772 267520 158778 267572
rect 166258 267520 166264 267572
rect 166316 267560 166322 267572
rect 194042 267560 194048 267572
rect 166316 267532 194048 267560
rect 166316 267520 166322 267532
rect 194042 267520 194048 267532
rect 194100 267520 194106 267572
rect 203334 267520 203340 267572
rect 203392 267560 203398 267572
rect 213178 267560 213184 267572
rect 203392 267532 213184 267560
rect 203392 267520 203398 267532
rect 213178 267520 213184 267532
rect 213236 267520 213242 267572
rect 286686 267520 286692 267572
rect 286744 267560 286750 267572
rect 294598 267560 294604 267572
rect 286744 267532 294604 267560
rect 286744 267520 286750 267532
rect 294598 267520 294604 267532
rect 294656 267520 294662 267572
rect 295610 267520 295616 267572
rect 295668 267560 295674 267572
rect 301958 267560 301964 267572
rect 295668 267532 301964 267560
rect 295668 267520 295674 267532
rect 301958 267520 301964 267532
rect 302016 267520 302022 267572
rect 308122 267520 308128 267572
rect 308180 267560 308186 267572
rect 329466 267560 329472 267572
rect 308180 267532 329472 267560
rect 308180 267520 308186 267532
rect 329466 267520 329472 267532
rect 329524 267520 329530 267572
rect 342714 267520 342720 267572
rect 342772 267560 342778 267572
rect 343542 267560 343548 267572
rect 342772 267532 343548 267560
rect 342772 267520 342778 267532
rect 343542 267520 343548 267532
rect 343600 267520 343606 267572
rect 346394 267520 346400 267572
rect 346452 267560 346458 267572
rect 368032 267560 368060 267668
rect 373442 267656 373448 267668
rect 373500 267656 373506 267708
rect 373626 267656 373632 267708
rect 373684 267696 373690 267708
rect 417694 267696 417700 267708
rect 373684 267668 417700 267696
rect 373684 267656 373690 267668
rect 417694 267656 417700 267668
rect 417752 267656 417758 267708
rect 417896 267696 417924 267804
rect 418062 267792 418068 267844
rect 418120 267832 418126 267844
rect 427740 267832 427768 267872
rect 418120 267804 427768 267832
rect 427832 267832 427860 267872
rect 660298 267860 660304 267912
rect 660356 267900 660362 267912
rect 669286 267900 669314 268008
rect 675478 267996 675484 268008
rect 675536 267996 675542 268048
rect 660356 267872 669314 267900
rect 660356 267860 660362 267872
rect 506474 267832 506480 267844
rect 427832 267804 428136 267832
rect 418120 267792 418126 267804
rect 428108 267764 428136 267804
rect 428292 267804 506480 267832
rect 428292 267764 428320 267804
rect 506474 267792 506480 267804
rect 506532 267792 506538 267844
rect 675478 267832 675484 267844
rect 669424 267804 675484 267832
rect 428108 267736 428320 267764
rect 668946 267724 668952 267776
rect 669004 267764 669010 267776
rect 669004 267736 669360 267764
rect 669004 267724 669010 267736
rect 427078 267696 427084 267708
rect 417896 267668 427084 267696
rect 427078 267656 427084 267668
rect 427136 267656 427142 267708
rect 432782 267656 432788 267708
rect 432840 267696 432846 267708
rect 436002 267696 436008 267708
rect 432840 267668 436008 267696
rect 432840 267656 432846 267668
rect 436002 267656 436008 267668
rect 436060 267656 436066 267708
rect 437382 267656 437388 267708
rect 437440 267696 437446 267708
rect 437440 267668 471284 267696
rect 437440 267656 437446 267668
rect 371602 267560 371608 267572
rect 346452 267532 368060 267560
rect 368124 267532 371608 267560
rect 346452 267520 346458 267532
rect 132586 267384 132592 267436
rect 132644 267424 132650 267436
rect 145466 267424 145472 267436
rect 132644 267396 145472 267424
rect 132644 267384 132650 267396
rect 145466 267384 145472 267396
rect 145524 267384 145530 267436
rect 145650 267384 145656 267436
rect 145708 267424 145714 267436
rect 149514 267424 149520 267436
rect 145708 267396 149520 267424
rect 145708 267384 145714 267396
rect 149514 267384 149520 267396
rect 149572 267384 149578 267436
rect 149698 267384 149704 267436
rect 149756 267424 149762 267436
rect 174170 267424 174176 267436
rect 149756 267396 174176 267424
rect 149756 267384 149762 267396
rect 174170 267384 174176 267396
rect 174228 267384 174234 267436
rect 179322 267384 179328 267436
rect 179380 267424 179386 267436
rect 207290 267424 207296 267436
rect 179380 267396 207296 267424
rect 179380 267384 179386 267396
rect 207290 267384 207296 267396
rect 207348 267384 207354 267436
rect 233878 267384 233884 267436
rect 233936 267424 233942 267436
rect 240410 267424 240416 267436
rect 233936 267396 240416 267424
rect 233936 267384 233942 267396
rect 240410 267384 240416 267396
rect 240468 267384 240474 267436
rect 293402 267384 293408 267436
rect 293460 267424 293466 267436
rect 302878 267424 302884 267436
rect 293460 267396 302884 267424
rect 293460 267384 293466 267396
rect 302878 267384 302884 267396
rect 302936 267384 302942 267436
rect 313274 267384 313280 267436
rect 313332 267424 313338 267436
rect 334618 267424 334624 267436
rect 313332 267396 334624 267424
rect 313332 267384 313338 267396
rect 334618 267384 334624 267396
rect 334676 267384 334682 267436
rect 335354 267384 335360 267436
rect 335412 267424 335418 267436
rect 342162 267424 342168 267436
rect 335412 267396 342168 267424
rect 335412 267384 335418 267396
rect 342162 267384 342168 267396
rect 342220 267384 342226 267436
rect 368124 267424 368152 267532
rect 371602 267520 371608 267532
rect 371660 267520 371666 267572
rect 371786 267520 371792 267572
rect 371844 267560 371850 267572
rect 377122 267560 377128 267572
rect 371844 267532 377128 267560
rect 371844 267520 371850 267532
rect 377122 267520 377128 267532
rect 377180 267520 377186 267572
rect 377306 267520 377312 267572
rect 377364 267560 377370 267572
rect 379330 267560 379336 267572
rect 377364 267532 379336 267560
rect 377364 267520 377370 267532
rect 379330 267520 379336 267532
rect 379388 267520 379394 267572
rect 379514 267520 379520 267572
rect 379572 267560 379578 267572
rect 379572 267532 381216 267560
rect 379572 267520 379578 267532
rect 380526 267424 380532 267436
rect 350506 267396 368152 267424
rect 369136 267396 380532 267424
rect 86218 267248 86224 267300
rect 86276 267288 86282 267300
rect 145926 267288 145932 267300
rect 86276 267260 145932 267288
rect 86276 267248 86282 267260
rect 145926 267248 145932 267260
rect 145984 267248 145990 267300
rect 146202 267248 146208 267300
rect 146260 267288 146266 267300
rect 187418 267288 187424 267300
rect 146260 267260 187424 267288
rect 146260 267248 146266 267260
rect 187418 267248 187424 267260
rect 187476 267248 187482 267300
rect 194502 267248 194508 267300
rect 194560 267288 194566 267300
rect 208762 267288 208768 267300
rect 194560 267260 208768 267288
rect 194560 267248 194566 267260
rect 208762 267248 208768 267260
rect 208820 267248 208826 267300
rect 257338 267248 257344 267300
rect 257396 267288 257402 267300
rect 259454 267288 259460 267300
rect 257396 267260 259460 267288
rect 257396 267248 257402 267260
rect 259454 267248 259460 267260
rect 259512 267248 259518 267300
rect 322106 267248 322112 267300
rect 322164 267288 322170 267300
rect 341794 267288 341800 267300
rect 322164 267260 341800 267288
rect 322164 267248 322170 267260
rect 341794 267248 341800 267260
rect 341852 267248 341858 267300
rect 341978 267248 341984 267300
rect 342036 267288 342042 267300
rect 350506 267288 350534 267396
rect 342036 267260 350534 267288
rect 342036 267248 342042 267260
rect 355226 267248 355232 267300
rect 355284 267288 355290 267300
rect 369136 267288 369164 267396
rect 380526 267384 380532 267396
rect 380584 267384 380590 267436
rect 381188 267424 381216 267532
rect 381354 267520 381360 267572
rect 381412 267560 381418 267572
rect 384298 267560 384304 267572
rect 381412 267532 384304 267560
rect 381412 267520 381418 267532
rect 384298 267520 384304 267532
rect 384356 267520 384362 267572
rect 384482 267520 384488 267572
rect 384540 267560 384546 267572
rect 388162 267560 388168 267572
rect 384540 267532 388168 267560
rect 384540 267520 384546 267532
rect 388162 267520 388168 267532
rect 388220 267520 388226 267572
rect 388346 267520 388352 267572
rect 388404 267560 388410 267572
rect 392578 267560 392584 267572
rect 388404 267532 392584 267560
rect 388404 267520 388410 267532
rect 392578 267520 392584 267532
rect 392636 267520 392642 267572
rect 392762 267520 392768 267572
rect 392820 267560 392826 267572
rect 427354 267560 427360 267572
rect 392820 267532 427360 267560
rect 392820 267520 392826 267532
rect 427354 267520 427360 267532
rect 427412 267520 427418 267572
rect 427998 267520 428004 267572
rect 428056 267560 428062 267572
rect 471054 267560 471060 267572
rect 428056 267532 471060 267560
rect 428056 267520 428062 267532
rect 471054 267520 471060 267532
rect 471112 267520 471118 267572
rect 471256 267560 471284 267668
rect 471422 267656 471428 267708
rect 471480 267696 471486 267708
rect 538858 267696 538864 267708
rect 471480 267668 538864 267696
rect 471480 267656 471486 267668
rect 538858 267656 538864 267668
rect 538916 267656 538922 267708
rect 669332 267696 669360 267736
rect 669424 267696 669452 267804
rect 675478 267792 675484 267804
rect 675536 267792 675542 267844
rect 669332 267668 669452 267696
rect 490466 267560 490472 267572
rect 471256 267532 490472 267560
rect 490466 267520 490472 267532
rect 490524 267520 490530 267572
rect 490650 267520 490656 267572
rect 490708 267560 490714 267572
rect 494146 267560 494152 267572
rect 490708 267532 494152 267560
rect 490708 267520 490714 267532
rect 494146 267520 494152 267532
rect 494204 267520 494210 267572
rect 494514 267520 494520 267572
rect 494572 267560 494578 267572
rect 585778 267560 585784 267572
rect 494572 267532 585784 267560
rect 494572 267520 494578 267532
rect 585778 267520 585784 267532
rect 585836 267520 585842 267572
rect 391750 267424 391756 267436
rect 381188 267396 391756 267424
rect 391750 267384 391756 267396
rect 391808 267384 391814 267436
rect 392026 267384 392032 267436
rect 392084 267424 392090 267436
rect 393222 267424 393228 267436
rect 392084 267396 393228 267424
rect 392084 267384 392090 267396
rect 393222 267384 393228 267396
rect 393280 267384 393286 267436
rect 393406 267384 393412 267436
rect 393464 267424 393470 267436
rect 464706 267424 464712 267436
rect 393464 267396 464712 267424
rect 393464 267384 393470 267396
rect 464706 267384 464712 267396
rect 464764 267384 464770 267436
rect 466822 267384 466828 267436
rect 466880 267424 466886 267436
rect 480162 267424 480168 267436
rect 466880 267396 480168 267424
rect 466880 267384 466886 267396
rect 480162 267384 480168 267396
rect 480220 267384 480226 267436
rect 480346 267384 480352 267436
rect 480404 267424 480410 267436
rect 483106 267424 483112 267436
rect 480404 267396 483112 267424
rect 480404 267384 480410 267396
rect 483106 267384 483112 267396
rect 483164 267384 483170 267436
rect 483290 267384 483296 267436
rect 483348 267424 483354 267436
rect 489730 267424 489736 267436
rect 483348 267396 489736 267424
rect 483348 267384 483354 267396
rect 489730 267384 489736 267396
rect 489788 267384 489794 267436
rect 490190 267384 490196 267436
rect 490248 267424 490254 267436
rect 625798 267424 625804 267436
rect 490248 267396 625804 267424
rect 490248 267384 490254 267396
rect 625798 267384 625804 267396
rect 625856 267384 625862 267436
rect 466380 267328 466500 267356
rect 355284 267260 369164 267288
rect 355284 267248 355290 267260
rect 370498 267248 370504 267300
rect 370556 267288 370562 267300
rect 390094 267288 390100 267300
rect 370556 267260 390100 267288
rect 370556 267248 370562 267260
rect 390094 267248 390100 267260
rect 390152 267248 390158 267300
rect 390462 267248 390468 267300
rect 390520 267288 390526 267300
rect 390520 267260 397960 267288
rect 390520 267248 390526 267260
rect 397932 267220 397960 267260
rect 398466 267248 398472 267300
rect 398524 267288 398530 267300
rect 401962 267288 401968 267300
rect 398524 267260 401968 267288
rect 398524 267248 398530 267260
rect 401962 267248 401968 267260
rect 402020 267248 402026 267300
rect 402974 267248 402980 267300
rect 403032 267288 403038 267300
rect 403032 267260 413324 267288
rect 403032 267248 403038 267260
rect 397932 267192 398052 267220
rect 91002 267112 91008 267164
rect 91060 267152 91066 267164
rect 146754 267152 146760 267164
rect 91060 267124 146760 267152
rect 91060 267112 91066 267124
rect 146754 267112 146760 267124
rect 146812 267112 146818 267164
rect 149514 267112 149520 267164
rect 149572 267152 149578 267164
rect 151354 267152 151360 267164
rect 149572 267124 151360 267152
rect 149572 267112 149578 267124
rect 151354 267112 151360 267124
rect 151412 267112 151418 267164
rect 167638 267112 167644 267164
rect 167696 267152 167702 267164
rect 198458 267152 198464 267164
rect 167696 267124 198464 267152
rect 167696 267112 167702 267124
rect 198458 267112 198464 267124
rect 198516 267112 198522 267164
rect 209866 267112 209872 267164
rect 209924 267152 209930 267164
rect 222746 267152 222752 267164
rect 209924 267124 222752 267152
rect 209924 267112 209930 267124
rect 222746 267112 222752 267124
rect 222804 267112 222810 267164
rect 227714 267112 227720 267164
rect 227772 267152 227778 267164
rect 232314 267152 232320 267164
rect 227772 267124 232320 267152
rect 227772 267112 227778 267124
rect 232314 267112 232320 267124
rect 232372 267112 232378 267164
rect 267642 267112 267648 267164
rect 267700 267152 267706 267164
rect 271138 267152 271144 267164
rect 267700 267124 271144 267152
rect 267700 267112 267706 267124
rect 271138 267112 271144 267124
rect 271196 267112 271202 267164
rect 272058 267112 272064 267164
rect 272116 267152 272122 267164
rect 280706 267152 280712 267164
rect 272116 267124 280712 267152
rect 272116 267112 272122 267124
rect 280706 267112 280712 267124
rect 280764 267112 280770 267164
rect 291194 267112 291200 267164
rect 291252 267152 291258 267164
rect 301498 267152 301504 267164
rect 291252 267124 301504 267152
rect 291252 267112 291258 267124
rect 301498 267112 301504 267124
rect 301556 267112 301562 267164
rect 302234 267112 302240 267164
rect 302292 267152 302298 267164
rect 312814 267152 312820 267164
rect 302292 267124 312820 267152
rect 302292 267112 302298 267124
rect 312814 267112 312820 267124
rect 312872 267112 312878 267164
rect 312998 267112 313004 267164
rect 313056 267152 313062 267164
rect 343358 267152 343364 267164
rect 313056 267124 343364 267152
rect 313056 267112 313062 267124
rect 343358 267112 343364 267124
rect 343416 267112 343422 267164
rect 350810 267112 350816 267164
rect 350868 267152 350874 267164
rect 350868 267124 369992 267152
rect 350868 267112 350874 267124
rect 73798 266976 73804 267028
rect 73856 267016 73862 267028
rect 140314 267016 140320 267028
rect 73856 266988 140320 267016
rect 73856 266976 73862 266988
rect 140314 266976 140320 266988
rect 140372 266976 140378 267028
rect 140498 266976 140504 267028
rect 140556 267016 140562 267028
rect 183002 267016 183008 267028
rect 140556 266988 183008 267016
rect 140556 266976 140562 266988
rect 183002 266976 183008 266988
rect 183060 266976 183066 267028
rect 186958 266976 186964 267028
rect 187016 267016 187022 267028
rect 211706 267016 211712 267028
rect 187016 266988 211712 267016
rect 187016 266976 187022 266988
rect 211706 266976 211712 266988
rect 211764 266976 211770 267028
rect 212442 266976 212448 267028
rect 212500 267016 212506 267028
rect 212500 266988 219434 267016
rect 212500 266976 212506 266988
rect 104894 266840 104900 266892
rect 104952 266880 104958 266892
rect 143258 266880 143264 266892
rect 104952 266852 143264 266880
rect 104952 266840 104958 266852
rect 143258 266840 143264 266852
rect 143316 266840 143322 266892
rect 146754 266840 146760 266892
rect 146812 266880 146818 266892
rect 152090 266880 152096 266892
rect 146812 266852 152096 266880
rect 146812 266840 146818 266852
rect 152090 266840 152096 266852
rect 152148 266840 152154 266892
rect 153838 266840 153844 266892
rect 153896 266880 153902 266892
rect 163130 266880 163136 266892
rect 153896 266852 163136 266880
rect 153896 266840 153902 266852
rect 163130 266840 163136 266852
rect 163188 266840 163194 266892
rect 163682 266840 163688 266892
rect 163740 266880 163746 266892
rect 176378 266880 176384 266892
rect 163740 266852 176384 266880
rect 163740 266840 163746 266852
rect 176378 266840 176384 266852
rect 176436 266840 176442 266892
rect 202874 266880 202880 266892
rect 180766 266852 202880 266880
rect 119338 266704 119344 266756
rect 119396 266744 119402 266756
rect 156230 266744 156236 266756
rect 119396 266716 156236 266744
rect 119396 266704 119402 266716
rect 156230 266704 156236 266716
rect 156288 266704 156294 266756
rect 156782 266704 156788 266756
rect 156840 266744 156846 266756
rect 165338 266744 165344 266756
rect 156840 266716 165344 266744
rect 156840 266704 156846 266716
rect 165338 266704 165344 266716
rect 165396 266704 165402 266756
rect 175918 266704 175924 266756
rect 175976 266744 175982 266756
rect 180766 266744 180794 266852
rect 202874 266840 202880 266852
rect 202932 266840 202938 266892
rect 219406 266880 219434 266988
rect 226334 266976 226340 267028
rect 226392 267016 226398 267028
rect 235994 267016 236000 267028
rect 226392 266988 236000 267016
rect 226392 266976 226398 266988
rect 235994 266976 236000 266988
rect 236052 266976 236058 267028
rect 278682 266976 278688 267028
rect 278740 267016 278746 267028
rect 293218 267016 293224 267028
rect 278740 266988 293224 267016
rect 278740 266976 278746 266988
rect 293218 266976 293224 266988
rect 293276 266976 293282 267028
rect 300394 266976 300400 267028
rect 300452 267016 300458 267028
rect 310790 267016 310796 267028
rect 300452 266988 310796 267016
rect 300452 266976 300458 266988
rect 310790 266976 310796 266988
rect 310848 266976 310854 267028
rect 314746 266976 314752 267028
rect 314804 267016 314810 267028
rect 340046 267016 340052 267028
rect 314804 266988 340052 267016
rect 314804 266976 314810 266988
rect 340046 266976 340052 266988
rect 340104 266976 340110 267028
rect 340248 266988 340874 267016
rect 227162 266880 227168 266892
rect 219406 266852 227168 266880
rect 227162 266840 227168 266852
rect 227220 266840 227226 266892
rect 256510 266840 256516 266892
rect 256568 266880 256574 266892
rect 258074 266880 258080 266892
rect 256568 266852 258080 266880
rect 256568 266840 256574 266852
rect 258074 266840 258080 266852
rect 258132 266840 258138 266892
rect 262858 266840 262864 266892
rect 262916 266880 262922 266892
rect 267918 266880 267924 266892
rect 262916 266852 267924 266880
rect 262916 266840 262922 266852
rect 267918 266840 267924 266852
rect 267976 266840 267982 266892
rect 275738 266840 275744 266892
rect 275796 266880 275802 266892
rect 278866 266880 278872 266892
rect 275796 266852 278872 266880
rect 275796 266840 275802 266852
rect 278866 266840 278872 266852
rect 278924 266840 278930 266892
rect 288986 266840 288992 266892
rect 289044 266880 289050 266892
rect 298738 266880 298744 266892
rect 289044 266852 298744 266880
rect 289044 266840 289050 266852
rect 298738 266840 298744 266852
rect 298796 266840 298802 266892
rect 311066 266840 311072 266892
rect 311124 266880 311130 266892
rect 319806 266880 319812 266892
rect 311124 266852 319812 266880
rect 311124 266840 311130 266852
rect 319806 266840 319812 266852
rect 319864 266840 319870 266892
rect 327258 266840 327264 266892
rect 327316 266880 327322 266892
rect 333422 266880 333428 266892
rect 327316 266852 333428 266880
rect 327316 266840 327322 266852
rect 333422 266840 333428 266852
rect 333480 266840 333486 266892
rect 338298 266840 338304 266892
rect 338356 266880 338362 266892
rect 340248 266880 340276 266988
rect 338356 266852 340276 266880
rect 340846 266880 340874 266988
rect 341794 266976 341800 267028
rect 341852 267016 341858 267028
rect 347774 267016 347780 267028
rect 341852 266988 347780 267016
rect 341852 266976 341858 266988
rect 347774 266976 347780 266988
rect 347832 266976 347838 267028
rect 348602 266976 348608 267028
rect 348660 267016 348666 267028
rect 348660 266988 364334 267016
rect 348660 266976 348666 266988
rect 358078 266880 358084 266892
rect 340846 266852 358084 266880
rect 338356 266840 338362 266852
rect 358078 266840 358084 266852
rect 358136 266840 358142 266892
rect 359642 266840 359648 266892
rect 359700 266880 359706 266892
rect 362954 266880 362960 266892
rect 359700 266852 362960 266880
rect 359700 266840 359706 266852
rect 362954 266840 362960 266852
rect 363012 266840 363018 266892
rect 364306 266880 364334 266988
rect 365990 266976 365996 267028
rect 366048 267016 366054 267028
rect 369964 267016 369992 267124
rect 371418 267112 371424 267164
rect 371476 267152 371482 267164
rect 396166 267152 396172 267164
rect 371476 267124 396172 267152
rect 371476 267112 371482 267124
rect 396166 267112 396172 267124
rect 396224 267112 396230 267164
rect 398024 267152 398052 267192
rect 398024 267124 413232 267152
rect 378962 267016 378968 267028
rect 366048 266988 369854 267016
rect 369964 266988 378968 267016
rect 366048 266976 366054 266988
rect 369118 266880 369124 266892
rect 364306 266852 369124 266880
rect 369118 266840 369124 266852
rect 369176 266840 369182 266892
rect 369826 266880 369854 266988
rect 378962 266976 378968 266988
rect 379020 266976 379026 267028
rect 379698 266976 379704 267028
rect 379756 267016 379762 267028
rect 413002 267016 413008 267028
rect 379756 266988 413008 267016
rect 379756 266976 379762 266988
rect 413002 266976 413008 266988
rect 413060 266976 413066 267028
rect 369826 266852 370176 266880
rect 175976 266716 180794 266744
rect 175976 266704 175982 266716
rect 319162 266704 319168 266756
rect 319220 266744 319226 266756
rect 339402 266744 339408 266756
rect 319220 266716 339408 266744
rect 319220 266704 319226 266716
rect 339402 266704 339408 266716
rect 339460 266704 339466 266756
rect 340046 266704 340052 266756
rect 340104 266744 340110 266756
rect 340104 266716 340874 266744
rect 340104 266704 340110 266716
rect 206278 266636 206284 266688
rect 206336 266676 206342 266688
rect 210234 266676 210240 266688
rect 206336 266648 210240 266676
rect 206336 266636 206342 266648
rect 210234 266636 210240 266648
rect 210292 266636 210298 266688
rect 126698 266568 126704 266620
rect 126756 266608 126762 266620
rect 148410 266608 148416 266620
rect 126756 266580 148416 266608
rect 126756 266568 126762 266580
rect 148410 266568 148416 266580
rect 148468 266568 148474 266620
rect 159634 266568 159640 266620
rect 159692 266608 159698 266620
rect 168282 266608 168288 266620
rect 159692 266580 168288 266608
rect 159692 266568 159698 266580
rect 168282 266568 168288 266580
rect 168340 266568 168346 266620
rect 246298 266568 246304 266620
rect 246356 266608 246362 266620
rect 248506 266608 248512 266620
rect 246356 266580 248512 266608
rect 246356 266568 246362 266580
rect 248506 266568 248512 266580
rect 248564 266568 248570 266620
rect 333422 266568 333428 266620
rect 333480 266608 333486 266620
rect 340846 266608 340874 266716
rect 343450 266704 343456 266756
rect 343508 266744 343514 266756
rect 351638 266744 351644 266756
rect 343508 266716 351644 266744
rect 343508 266704 343514 266716
rect 351638 266704 351644 266716
rect 351696 266704 351702 266756
rect 353018 266704 353024 266756
rect 353076 266744 353082 266756
rect 369302 266744 369308 266756
rect 353076 266716 369308 266744
rect 353076 266704 353082 266716
rect 369302 266704 369308 266716
rect 369360 266704 369366 266756
rect 370148 266744 370176 266852
rect 370682 266840 370688 266892
rect 370740 266880 370746 266892
rect 412818 266880 412824 266892
rect 370740 266852 412824 266880
rect 370740 266840 370746 266852
rect 412818 266840 412824 266852
rect 412876 266840 412882 266892
rect 413204 266880 413232 267124
rect 413296 267084 413324 267260
rect 417050 267248 417056 267300
rect 417108 267288 417114 267300
rect 417878 267288 417884 267300
rect 417108 267260 417884 267288
rect 417108 267248 417114 267260
rect 417878 267248 417884 267260
rect 417936 267248 417942 267300
rect 418062 267248 418068 267300
rect 418120 267288 418126 267300
rect 466380 267288 466408 267328
rect 418120 267260 466408 267288
rect 466472 267288 466500 267328
rect 466472 267260 466868 267288
rect 418120 267248 418126 267260
rect 413462 267180 413468 267232
rect 413520 267220 413526 267232
rect 416866 267220 416872 267232
rect 413520 267192 416872 267220
rect 413520 267180 413526 267192
rect 416866 267180 416872 267192
rect 416924 267180 416930 267232
rect 466178 267152 466184 267164
rect 417068 267124 466184 267152
rect 417068 267084 417096 267124
rect 466178 267112 466184 267124
rect 466236 267112 466242 267164
rect 413296 267056 417096 267084
rect 417234 266976 417240 267028
rect 417292 267016 417298 267028
rect 421742 267016 421748 267028
rect 417292 266988 421748 267016
rect 417292 266976 417298 266988
rect 421742 266976 421748 266988
rect 421800 266976 421806 267028
rect 426894 267016 426900 267028
rect 421944 266988 426900 267016
rect 421944 266880 421972 266988
rect 426894 266976 426900 266988
rect 426952 266976 426958 267028
rect 427078 266976 427084 267028
rect 427136 267016 427142 267028
rect 466178 267016 466184 267028
rect 427136 266988 466184 267016
rect 427136 266976 427142 266988
rect 466178 266976 466184 266988
rect 466236 266976 466242 267028
rect 466840 267016 466868 267260
rect 469674 267248 469680 267300
rect 469732 267288 469738 267300
rect 470502 267288 470508 267300
rect 469732 267260 470508 267288
rect 469732 267248 469738 267260
rect 470502 267248 470508 267260
rect 470560 267248 470566 267300
rect 471054 267248 471060 267300
rect 471112 267288 471118 267300
rect 476298 267288 476304 267300
rect 471112 267260 476304 267288
rect 471112 267248 471118 267260
rect 476298 267248 476304 267260
rect 476356 267248 476362 267300
rect 476482 267248 476488 267300
rect 476540 267288 476546 267300
rect 543734 267288 543740 267300
rect 476540 267260 543740 267288
rect 476540 267248 476546 267260
rect 543734 267248 543740 267260
rect 543792 267248 543798 267300
rect 467006 267112 467012 267164
rect 467064 267152 467070 267164
rect 487798 267152 487804 267164
rect 467064 267124 487804 267152
rect 467064 267112 467070 267124
rect 487798 267112 487804 267124
rect 487856 267112 487862 267164
rect 489914 267112 489920 267164
rect 489972 267152 489978 267164
rect 491202 267152 491208 267164
rect 489972 267124 491208 267152
rect 489972 267112 489978 267124
rect 491202 267112 491208 267124
rect 491260 267112 491266 267164
rect 491386 267112 491392 267164
rect 491444 267152 491450 267164
rect 494698 267152 494704 267164
rect 491444 267124 494704 267152
rect 491444 267112 491450 267124
rect 494698 267112 494704 267124
rect 494756 267112 494762 267164
rect 494882 267112 494888 267164
rect 494940 267152 494946 267164
rect 497642 267152 497648 267164
rect 494940 267124 497648 267152
rect 494940 267112 494946 267124
rect 497642 267112 497648 267124
rect 497700 267112 497706 267164
rect 499528 267112 499534 267164
rect 499586 267152 499592 267164
rect 632698 267152 632704 267164
rect 499586 267124 632704 267152
rect 499586 267112 499592 267124
rect 632698 267112 632704 267124
rect 632756 267112 632762 267164
rect 479518 267016 479524 267028
rect 466840 266988 479524 267016
rect 479518 266976 479524 266988
rect 479576 266976 479582 267028
rect 479702 266976 479708 267028
rect 479760 267016 479766 267028
rect 554038 267016 554044 267028
rect 479760 266988 554044 267016
rect 479760 266976 479766 266988
rect 554038 266976 554044 266988
rect 554096 266976 554102 267028
rect 413204 266852 421972 266880
rect 422386 266840 422392 266892
rect 422444 266880 422450 266892
rect 514018 266880 514024 266892
rect 422444 266852 514024 266880
rect 422444 266840 422450 266852
rect 514018 266840 514024 266852
rect 514076 266840 514082 266892
rect 514202 266840 514208 266892
rect 514260 266880 514266 266892
rect 525886 266880 525892 266892
rect 514260 266852 525892 266880
rect 514260 266840 514266 266852
rect 525886 266840 525892 266852
rect 525944 266840 525950 266892
rect 374086 266744 374092 266756
rect 370148 266716 374092 266744
rect 374086 266704 374092 266716
rect 374144 266704 374150 266756
rect 375098 266704 375104 266756
rect 375156 266744 375162 266756
rect 379698 266744 379704 266756
rect 375156 266716 379704 266744
rect 375156 266704 375162 266716
rect 379698 266704 379704 266716
rect 379756 266704 379762 266756
rect 380986 266704 380992 266756
rect 381044 266744 381050 266756
rect 382182 266744 382188 266756
rect 381044 266716 382188 266744
rect 381044 266704 381050 266716
rect 382182 266704 382188 266716
rect 382240 266704 382246 266756
rect 385402 266704 385408 266756
rect 385460 266744 385466 266756
rect 388806 266744 388812 266756
rect 385460 266716 388812 266744
rect 385460 266704 385466 266716
rect 388806 266704 388812 266716
rect 388864 266704 388870 266756
rect 390554 266704 390560 266756
rect 390612 266744 390618 266756
rect 391566 266744 391572 266756
rect 390612 266716 391572 266744
rect 390612 266704 390618 266716
rect 391566 266704 391572 266716
rect 391624 266704 391630 266756
rect 391750 266704 391756 266756
rect 391808 266744 391814 266756
rect 424962 266744 424968 266756
rect 391808 266716 424968 266744
rect 391808 266704 391814 266716
rect 424962 266704 424968 266716
rect 425020 266704 425026 266756
rect 425146 266704 425152 266756
rect 425204 266744 425210 266756
rect 426250 266744 426256 266756
rect 425204 266716 426256 266744
rect 425204 266704 425210 266716
rect 426250 266704 426256 266716
rect 426308 266704 426314 266756
rect 426618 266704 426624 266756
rect 426676 266744 426682 266756
rect 427538 266744 427544 266756
rect 426676 266716 427544 266744
rect 426676 266704 426682 266716
rect 427538 266704 427544 266716
rect 427596 266704 427602 266756
rect 427906 266704 427912 266756
rect 427964 266744 427970 266756
rect 432782 266744 432788 266756
rect 427964 266716 432788 266744
rect 427964 266704 427970 266716
rect 432782 266704 432788 266716
rect 432840 266704 432846 266756
rect 433242 266704 433248 266756
rect 433300 266744 433306 266756
rect 437382 266744 437388 266756
rect 433300 266716 437388 266744
rect 433300 266704 433306 266716
rect 437382 266704 437388 266716
rect 437440 266704 437446 266756
rect 437658 266704 437664 266756
rect 437716 266744 437722 266756
rect 476482 266744 476488 266756
rect 437716 266716 476488 266744
rect 437716 266704 437722 266716
rect 476482 266704 476488 266716
rect 476540 266704 476546 266756
rect 478874 266704 478880 266756
rect 478932 266744 478938 266756
rect 479702 266744 479708 266756
rect 478932 266716 479708 266744
rect 478932 266704 478938 266716
rect 479702 266704 479708 266716
rect 479760 266704 479766 266756
rect 479886 266704 479892 266756
rect 479944 266744 479950 266756
rect 571978 266744 571984 266756
rect 479944 266716 571984 266744
rect 479944 266704 479950 266716
rect 571978 266704 571984 266716
rect 572036 266704 572042 266756
rect 666370 266636 666376 266688
rect 666428 266676 666434 266688
rect 675478 266676 675484 266688
rect 666428 266648 675484 266676
rect 666428 266636 666434 266648
rect 675478 266636 675484 266648
rect 675536 266636 675542 266688
rect 346578 266608 346584 266620
rect 333480 266580 335354 266608
rect 340846 266580 346584 266608
rect 333480 266568 333486 266580
rect 211154 266500 211160 266552
rect 211212 266540 211218 266552
rect 214650 266540 214656 266552
rect 211212 266512 214656 266540
rect 211212 266500 211218 266512
rect 214650 266500 214656 266512
rect 214708 266500 214714 266552
rect 241330 266500 241336 266552
rect 241388 266540 241394 266552
rect 245562 266540 245568 266552
rect 241388 266512 245568 266540
rect 241388 266500 241394 266512
rect 245562 266500 245568 266512
rect 245620 266500 245626 266552
rect 259546 266500 259552 266552
rect 259604 266540 259610 266552
rect 262582 266540 262588 266552
rect 259604 266512 262588 266540
rect 259604 266500 259610 266512
rect 262582 266500 262588 266512
rect 262640 266500 262646 266552
rect 269850 266500 269856 266552
rect 269908 266540 269914 266552
rect 274818 266540 274824 266552
rect 269908 266512 274824 266540
rect 269908 266500 269914 266512
rect 274818 266500 274824 266512
rect 274876 266500 274882 266552
rect 280154 266500 280160 266552
rect 280212 266540 280218 266552
rect 286318 266540 286324 266552
rect 280212 266512 286324 266540
rect 280212 266500 280218 266512
rect 286318 266500 286324 266512
rect 286376 266500 286382 266552
rect 301498 266500 301504 266552
rect 301556 266540 301562 266552
rect 304166 266540 304172 266552
rect 301556 266512 304172 266540
rect 301556 266500 301562 266512
rect 304166 266500 304172 266512
rect 304224 266500 304230 266552
rect 304442 266500 304448 266552
rect 304500 266540 304506 266552
rect 306098 266540 306104 266552
rect 304500 266512 306104 266540
rect 304500 266500 304506 266512
rect 306098 266500 306104 266512
rect 306156 266500 306162 266552
rect 330938 266500 330944 266552
rect 330996 266540 331002 266552
rect 333238 266540 333244 266552
rect 330996 266512 333244 266540
rect 330996 266500 331002 266512
rect 333238 266500 333244 266512
rect 333296 266500 333302 266552
rect 78582 266432 78588 266484
rect 78640 266472 78646 266484
rect 137370 266472 137376 266484
rect 78640 266444 137376 266472
rect 78640 266432 78646 266444
rect 137370 266432 137376 266444
rect 137428 266432 137434 266484
rect 137554 266432 137560 266484
rect 137612 266472 137618 266484
rect 154298 266472 154304 266484
rect 137612 266444 154304 266472
rect 137612 266432 137618 266444
rect 154298 266432 154304 266444
rect 154356 266432 154362 266484
rect 335326 266472 335354 266580
rect 346578 266568 346584 266580
rect 346636 266568 346642 266620
rect 347866 266568 347872 266620
rect 347924 266608 347930 266620
rect 365806 266608 365812 266620
rect 347924 266580 365812 266608
rect 347924 266568 347930 266580
rect 365806 266568 365812 266580
rect 365864 266568 365870 266620
rect 372890 266568 372896 266620
rect 372948 266608 372954 266620
rect 405918 266608 405924 266620
rect 372948 266580 405924 266608
rect 372948 266568 372954 266580
rect 405918 266568 405924 266580
rect 405976 266568 405982 266620
rect 490098 266608 490104 266620
rect 417804 266580 466316 266608
rect 406378 266500 406384 266552
rect 406436 266540 406442 266552
rect 417602 266540 417608 266552
rect 406436 266512 417608 266540
rect 406436 266500 406442 266512
rect 417602 266500 417608 266512
rect 417660 266500 417666 266552
rect 345474 266472 345480 266484
rect 335326 266444 345480 266472
rect 345474 266432 345480 266444
rect 345532 266432 345538 266484
rect 362954 266432 362960 266484
rect 363012 266472 363018 266484
rect 396258 266472 396264 266484
rect 363012 266444 396264 266472
rect 363012 266432 363018 266444
rect 396258 266432 396264 266444
rect 396316 266432 396322 266484
rect 157886 266364 157892 266416
rect 157944 266404 157950 266416
rect 159450 266404 159456 266416
rect 157944 266376 159456 266404
rect 157944 266364 157950 266376
rect 159450 266364 159456 266376
rect 159508 266364 159514 266416
rect 204898 266364 204904 266416
rect 204956 266404 204962 266416
rect 206554 266404 206560 266416
rect 204956 266376 206560 266404
rect 204956 266364 204962 266376
rect 206554 266364 206560 266376
rect 206612 266364 206618 266416
rect 208486 266364 208492 266416
rect 208544 266404 208550 266416
rect 212442 266404 212448 266416
rect 208544 266376 212448 266404
rect 208544 266364 208550 266376
rect 212442 266364 212448 266376
rect 212500 266364 212506 266416
rect 219434 266364 219440 266416
rect 219492 266404 219498 266416
rect 227898 266404 227904 266416
rect 219492 266376 227904 266404
rect 219492 266364 219498 266376
rect 227898 266364 227904 266376
rect 227956 266364 227962 266416
rect 232498 266364 232504 266416
rect 232556 266404 232562 266416
rect 233786 266404 233792 266416
rect 232556 266376 233792 266404
rect 232556 266364 232562 266376
rect 233786 266364 233792 266376
rect 233844 266364 233850 266416
rect 239490 266364 239496 266416
rect 239548 266404 239554 266416
rect 241882 266404 241888 266416
rect 239548 266376 241888 266404
rect 239548 266364 239554 266376
rect 241882 266364 241888 266376
rect 241940 266364 241946 266416
rect 251174 266364 251180 266416
rect 251232 266404 251238 266416
rect 252186 266404 252192 266416
rect 251232 266376 252192 266404
rect 251232 266364 251238 266376
rect 252186 266364 252192 266376
rect 252244 266364 252250 266416
rect 255866 266364 255872 266416
rect 255924 266404 255930 266416
rect 256694 266404 256700 266416
rect 255924 266376 256700 266404
rect 255924 266364 255930 266376
rect 256694 266364 256700 266376
rect 256752 266364 256758 266416
rect 258074 266364 258080 266416
rect 258132 266404 258138 266416
rect 259730 266404 259736 266416
rect 258132 266376 259736 266404
rect 258132 266364 258138 266376
rect 259730 266364 259736 266376
rect 259788 266364 259794 266416
rect 260282 266364 260288 266416
rect 260340 266404 260346 266416
rect 261754 266404 261760 266416
rect 260340 266376 261760 266404
rect 260340 266364 260346 266376
rect 261754 266364 261760 266376
rect 261812 266364 261818 266416
rect 262122 266364 262128 266416
rect 262180 266404 262186 266416
rect 266354 266404 266360 266416
rect 262180 266376 266360 266404
rect 262180 266364 262186 266376
rect 266354 266364 266360 266376
rect 266412 266364 266418 266416
rect 270586 266364 270592 266416
rect 270644 266404 270650 266416
rect 271598 266404 271604 266416
rect 270644 266376 271604 266404
rect 270644 266364 270650 266376
rect 271598 266364 271604 266376
rect 271656 266364 271662 266416
rect 280890 266364 280896 266416
rect 280948 266404 280954 266416
rect 282178 266404 282184 266416
rect 280948 266376 282184 266404
rect 280948 266364 280954 266376
rect 282178 266364 282184 266376
rect 282236 266364 282242 266416
rect 284570 266364 284576 266416
rect 284628 266404 284634 266416
rect 285490 266404 285496 266416
rect 284628 266376 285496 266404
rect 284628 266364 284634 266376
rect 285490 266364 285496 266376
rect 285548 266364 285554 266416
rect 286042 266364 286048 266416
rect 286100 266404 286106 266416
rect 286870 266404 286876 266416
rect 286100 266376 286876 266404
rect 286100 266364 286106 266376
rect 286870 266364 286876 266376
rect 286928 266364 286934 266416
rect 294138 266364 294144 266416
rect 294196 266404 294202 266416
rect 295058 266404 295064 266416
rect 294196 266376 295064 266404
rect 294196 266364 294202 266376
rect 295058 266364 295064 266376
rect 295116 266364 295122 266416
rect 298554 266364 298560 266416
rect 298612 266404 298618 266416
rect 300118 266404 300124 266416
rect 298612 266376 300124 266404
rect 298612 266364 298618 266376
rect 300118 266364 300124 266376
rect 300176 266364 300182 266416
rect 303706 266364 303712 266416
rect 303764 266404 303770 266416
rect 304902 266404 304908 266416
rect 303764 266376 304908 266404
rect 303764 266364 303770 266376
rect 304902 266364 304908 266376
rect 304960 266364 304966 266416
rect 305178 266364 305184 266416
rect 305236 266404 305242 266416
rect 306282 266404 306288 266416
rect 305236 266376 306288 266404
rect 305236 266364 305242 266376
rect 306282 266364 306288 266376
rect 306340 266364 306346 266416
rect 306650 266364 306656 266416
rect 306708 266404 306714 266416
rect 313918 266404 313924 266416
rect 306708 266376 313924 266404
rect 306708 266364 306714 266376
rect 313918 266364 313924 266376
rect 313976 266364 313982 266416
rect 316218 266364 316224 266416
rect 316276 266404 316282 266416
rect 317322 266404 317328 266416
rect 316276 266376 317328 266404
rect 316276 266364 316282 266376
rect 317322 266364 317328 266376
rect 317380 266364 317386 266416
rect 320634 266364 320640 266416
rect 320692 266404 320698 266416
rect 321462 266404 321468 266416
rect 320692 266376 321468 266404
rect 320692 266364 320698 266376
rect 321462 266364 321468 266376
rect 321520 266364 321526 266416
rect 331674 266364 331680 266416
rect 331732 266404 331738 266416
rect 332502 266404 332508 266416
rect 331732 266376 332508 266404
rect 331732 266364 331738 266376
rect 332502 266364 332508 266376
rect 332560 266364 332566 266416
rect 345658 266364 345664 266416
rect 345716 266404 345722 266416
rect 345716 266376 352144 266404
rect 345716 266364 345722 266376
rect 352116 266268 352144 266376
rect 352282 266364 352288 266416
rect 352340 266404 352346 266416
rect 353202 266404 353208 266416
rect 352340 266376 353208 266404
rect 352340 266364 352346 266376
rect 353202 266364 353208 266376
rect 353260 266364 353266 266416
rect 354766 266404 354772 266416
rect 353404 266376 354772 266404
rect 353404 266268 353432 266376
rect 354766 266364 354772 266376
rect 354824 266364 354830 266416
rect 358906 266364 358912 266416
rect 358964 266404 358970 266416
rect 360102 266404 360108 266416
rect 358964 266376 360108 266404
rect 358964 266364 358970 266376
rect 360102 266364 360108 266376
rect 360160 266364 360166 266416
rect 361850 266364 361856 266416
rect 361908 266404 361914 266416
rect 362770 266404 362776 266416
rect 361908 266376 362776 266404
rect 361908 266364 361914 266376
rect 362770 266364 362776 266376
rect 362828 266364 362834 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 397472 266376 401456 266404
rect 352116 266240 353432 266268
rect 397178 266228 397184 266280
rect 397236 266268 397242 266280
rect 397472 266268 397500 266376
rect 397236 266240 397500 266268
rect 401428 266268 401456 266376
rect 401594 266364 401600 266416
rect 401652 266404 401658 266416
rect 402882 266404 402888 266416
rect 401652 266376 402888 266404
rect 401652 266364 401658 266376
rect 402882 266364 402888 266376
rect 402940 266364 402946 266416
rect 403066 266364 403072 266416
rect 403124 266404 403130 266416
rect 404170 266404 404176 266416
rect 403124 266376 404176 266404
rect 403124 266364 403130 266376
rect 404170 266364 404176 266376
rect 404228 266364 404234 266416
rect 404372 266376 414704 266404
rect 404372 266268 404400 266376
rect 401428 266240 404400 266268
rect 414676 266268 414704 266376
rect 414842 266364 414848 266416
rect 414900 266404 414906 266416
rect 417234 266404 417240 266416
rect 414900 266376 417240 266404
rect 414900 266364 414906 266376
rect 417234 266364 417240 266376
rect 417292 266364 417298 266416
rect 417418 266364 417424 266416
rect 417476 266404 417482 266416
rect 417804 266404 417832 266580
rect 466288 266540 466316 266580
rect 466748 266580 490104 266608
rect 466748 266540 466776 266580
rect 490098 266568 490104 266580
rect 490156 266568 490162 266620
rect 493318 266608 493324 266620
rect 491588 266580 493324 266608
rect 466288 266512 466776 266540
rect 421926 266432 421932 266484
rect 421984 266472 421990 266484
rect 465810 266472 465816 266484
rect 421984 266444 465816 266472
rect 421984 266432 421990 266444
rect 465810 266432 465816 266444
rect 465868 266432 465874 266484
rect 466914 266432 466920 266484
rect 466972 266472 466978 266484
rect 491588 266472 491616 266580
rect 493318 266568 493324 266580
rect 493376 266568 493382 266620
rect 494698 266568 494704 266620
rect 494756 266608 494762 266620
rect 513834 266608 513840 266620
rect 494756 266580 513840 266608
rect 494756 266568 494762 266580
rect 513834 266568 513840 266580
rect 513892 266568 513898 266620
rect 514018 266568 514024 266620
rect 514076 266608 514082 266620
rect 518894 266608 518900 266620
rect 514076 266580 518900 266608
rect 514076 266568 514082 266580
rect 518894 266568 518900 266580
rect 518952 266568 518958 266620
rect 664254 266500 664260 266552
rect 664312 266540 664318 266552
rect 675110 266540 675116 266552
rect 664312 266512 675116 266540
rect 664312 266500 664318 266512
rect 675110 266500 675116 266512
rect 675168 266500 675174 266552
rect 466972 266444 491616 266472
rect 466972 266432 466978 266444
rect 492858 266432 492864 266484
rect 492916 266472 492922 266484
rect 493686 266472 493692 266484
rect 492916 266444 493692 266472
rect 492916 266432 492922 266444
rect 493686 266432 493692 266444
rect 493744 266432 493750 266484
rect 494330 266432 494336 266484
rect 494388 266472 494394 266484
rect 495342 266472 495348 266484
rect 494388 266444 495348 266472
rect 494388 266432 494394 266444
rect 495342 266432 495348 266444
rect 495400 266432 495406 266484
rect 495802 266432 495808 266484
rect 495860 266472 495866 266484
rect 496722 266472 496728 266484
rect 495860 266444 496728 266472
rect 495860 266432 495866 266444
rect 496722 266432 496728 266444
rect 496780 266432 496786 266484
rect 498654 266432 498660 266484
rect 498712 266472 498718 266484
rect 499206 266472 499212 266484
rect 498712 266444 499212 266472
rect 498712 266432 498718 266444
rect 499206 266432 499212 266444
rect 499264 266432 499270 266484
rect 499390 266432 499396 266484
rect 499448 266472 499454 266484
rect 601602 266472 601608 266484
rect 499448 266444 601608 266472
rect 499448 266432 499454 266444
rect 601602 266432 601608 266444
rect 601660 266432 601666 266484
rect 417476 266376 417832 266404
rect 417476 266364 417482 266376
rect 418522 266364 418528 266416
rect 418580 266404 418586 266416
rect 419442 266404 419448 266416
rect 418580 266376 419448 266404
rect 418580 266364 418586 266376
rect 419442 266364 419448 266376
rect 419500 266364 419506 266416
rect 419644 266376 421788 266404
rect 415670 266268 415676 266280
rect 414676 266240 415676 266268
rect 397236 266228 397242 266240
rect 415670 266228 415676 266240
rect 415728 266228 415734 266280
rect 419442 266228 419448 266280
rect 419500 266268 419506 266280
rect 419644 266268 419672 266376
rect 421760 266336 421788 266376
rect 664438 266364 664444 266416
rect 664496 266404 664502 266416
rect 675294 266404 675300 266416
rect 664496 266376 675300 266404
rect 664496 266364 664502 266376
rect 675294 266364 675300 266376
rect 675352 266364 675358 266416
rect 422386 266336 422392 266348
rect 421760 266308 422392 266336
rect 422386 266296 422392 266308
rect 422444 266296 422450 266348
rect 424042 266296 424048 266348
rect 424100 266336 424106 266348
rect 427906 266336 427912 266348
rect 424100 266308 427912 266336
rect 424100 266296 424106 266308
rect 427906 266296 427912 266308
rect 427964 266296 427970 266348
rect 435082 266296 435088 266348
rect 435140 266336 435146 266348
rect 437658 266336 437664 266348
rect 435140 266308 437664 266336
rect 435140 266296 435146 266308
rect 437658 266296 437664 266308
rect 437716 266296 437722 266348
rect 448698 266296 448704 266348
rect 448756 266336 448762 266348
rect 566090 266336 566096 266348
rect 448756 266308 566096 266336
rect 448756 266296 448762 266308
rect 566090 266296 566096 266308
rect 566148 266296 566154 266348
rect 419500 266240 419672 266268
rect 419500 266228 419506 266240
rect 382090 266160 382096 266212
rect 382148 266200 382154 266212
rect 384114 266200 384120 266212
rect 382148 266172 384120 266200
rect 382148 266160 382154 266172
rect 384114 266160 384120 266172
rect 384172 266160 384178 266212
rect 421834 266160 421840 266212
rect 421892 266200 421898 266212
rect 422202 266200 422208 266212
rect 421892 266172 422208 266200
rect 421892 266160 421898 266172
rect 422202 266160 422208 266172
rect 422260 266160 422266 266212
rect 442074 266160 442080 266212
rect 442132 266200 442138 266212
rect 448882 266200 448888 266212
rect 442132 266172 448888 266200
rect 442132 266160 442138 266172
rect 448882 266160 448888 266172
rect 448940 266160 448946 266212
rect 449066 266160 449072 266212
rect 449124 266200 449130 266212
rect 456748 266200 456754 266212
rect 449124 266172 456754 266200
rect 449124 266160 449130 266172
rect 456748 266160 456754 266172
rect 456806 266160 456812 266212
rect 456886 266160 456892 266212
rect 456944 266200 456950 266212
rect 575658 266200 575664 266212
rect 456944 266172 575664 266200
rect 456944 266160 456950 266172
rect 575658 266160 575664 266172
rect 575716 266160 575722 266212
rect 362586 266024 362592 266076
rect 362644 266064 362650 266076
rect 428274 266064 428280 266076
rect 362644 266036 428280 266064
rect 362644 266024 362650 266036
rect 428274 266024 428280 266036
rect 428332 266024 428338 266076
rect 447594 266024 447600 266076
rect 447652 266064 447658 266076
rect 448330 266064 448336 266076
rect 447652 266036 448336 266064
rect 447652 266024 447658 266036
rect 448330 266024 448336 266036
rect 448388 266024 448394 266076
rect 448514 266024 448520 266076
rect 448572 266064 448578 266076
rect 448572 266036 461256 266064
rect 448572 266024 448578 266036
rect 184934 265888 184940 265940
rect 184992 265928 184998 265940
rect 185670 265928 185676 265940
rect 184992 265900 185676 265928
rect 184992 265888 184998 265900
rect 185670 265888 185676 265900
rect 185728 265888 185734 265940
rect 198734 265888 198740 265940
rect 198792 265928 198798 265940
rect 199654 265928 199660 265940
rect 198792 265900 199660 265928
rect 198792 265888 198798 265900
rect 199654 265888 199660 265900
rect 199712 265888 199718 265940
rect 384666 265888 384672 265940
rect 384724 265928 384730 265940
rect 461026 265928 461032 265940
rect 384724 265900 461032 265928
rect 384724 265888 384730 265900
rect 461026 265888 461032 265900
rect 461084 265888 461090 265940
rect 461228 265928 461256 266036
rect 461762 266024 461768 266076
rect 461820 266064 461826 266076
rect 463970 266064 463976 266076
rect 461820 266036 463976 266064
rect 461820 266024 461826 266036
rect 463970 266024 463976 266036
rect 464028 266024 464034 266076
rect 464154 266024 464160 266076
rect 464212 266064 464218 266076
rect 591022 266064 591028 266076
rect 464212 266036 591028 266064
rect 464212 266024 464218 266036
rect 591022 266024 591028 266036
rect 591080 266024 591086 266076
rect 467374 265928 467380 265940
rect 461228 265900 467380 265928
rect 467374 265888 467380 265900
rect 467432 265888 467438 265940
rect 470778 265888 470784 265940
rect 470836 265928 470842 265940
rect 601786 265928 601792 265940
rect 470836 265900 601792 265928
rect 470836 265888 470842 265900
rect 601786 265888 601792 265900
rect 601844 265888 601850 265940
rect 670418 265820 670424 265872
rect 670476 265860 670482 265872
rect 675294 265860 675300 265872
rect 670476 265832 675300 265860
rect 670476 265820 670482 265832
rect 675294 265820 675300 265832
rect 675352 265820 675358 265872
rect 368474 265752 368480 265804
rect 368532 265792 368538 265804
rect 369762 265792 369768 265804
rect 368532 265764 369768 265792
rect 368532 265752 368538 265764
rect 369762 265752 369768 265764
rect 369820 265752 369826 265804
rect 389082 265752 389088 265804
rect 389140 265792 389146 265804
rect 470594 265792 470600 265804
rect 389140 265764 470600 265792
rect 389140 265752 389146 265764
rect 470594 265752 470600 265764
rect 470652 265752 470658 265804
rect 477402 265752 477408 265804
rect 477460 265792 477466 265804
rect 612734 265792 612740 265804
rect 477460 265764 612740 265792
rect 477460 265752 477466 265764
rect 612734 265752 612740 265764
rect 612792 265752 612798 265804
rect 404538 265616 404544 265668
rect 404596 265656 404602 265668
rect 495618 265656 495624 265668
rect 404596 265628 495624 265656
rect 404596 265616 404602 265628
rect 495618 265616 495624 265628
rect 495676 265616 495682 265668
rect 497274 265616 497280 265668
rect 497332 265656 497338 265668
rect 643738 265656 643744 265668
rect 497332 265628 643744 265656
rect 497332 265616 497338 265628
rect 643738 265616 643744 265628
rect 643796 265616 643802 265668
rect 669314 265548 669320 265600
rect 669372 265588 669378 265600
rect 675478 265588 675484 265600
rect 669372 265560 675484 265588
rect 669372 265548 669378 265560
rect 675478 265548 675484 265560
rect 675536 265548 675542 265600
rect 403802 265480 403808 265532
rect 403860 265520 403866 265532
rect 448514 265520 448520 265532
rect 403860 265492 448520 265520
rect 403860 265480 403866 265492
rect 448514 265480 448520 265492
rect 448572 265480 448578 265532
rect 559282 265520 559288 265532
rect 448716 265492 559288 265520
rect 444282 265344 444288 265396
rect 444340 265384 444346 265396
rect 448716 265384 448744 265492
rect 559282 265480 559288 265492
rect 559340 265480 559346 265532
rect 444340 265356 448744 265384
rect 444340 265344 444346 265356
rect 448882 265344 448888 265396
rect 448940 265384 448946 265396
rect 552842 265384 552848 265396
rect 448940 265356 552848 265384
rect 448940 265344 448946 265356
rect 552842 265344 552848 265356
rect 552900 265344 552906 265396
rect 417786 265208 417792 265260
rect 417844 265248 417850 265260
rect 516410 265248 516416 265260
rect 417844 265220 516416 265248
rect 417844 265208 417850 265220
rect 516410 265208 516416 265220
rect 516468 265208 516474 265260
rect 666002 265208 666008 265260
rect 666060 265248 666066 265260
rect 675478 265248 675484 265260
rect 666060 265220 675484 265248
rect 666060 265208 666066 265220
rect 675478 265208 675484 265220
rect 675536 265208 675542 265260
rect 439866 265072 439872 265124
rect 439924 265112 439930 265124
rect 537754 265112 537760 265124
rect 439924 265084 537760 265112
rect 439924 265072 439930 265084
rect 537754 265072 537760 265084
rect 537812 265072 537818 265124
rect 664990 265072 664996 265124
rect 665048 265112 665054 265124
rect 665048 265084 669452 265112
rect 665048 265072 665054 265084
rect 669424 265044 669452 265084
rect 675478 265044 675484 265056
rect 669424 265016 675484 265044
rect 675478 265004 675484 265016
rect 675536 265004 675542 265056
rect 437658 264936 437664 264988
rect 437716 264976 437722 264988
rect 523678 264976 523684 264988
rect 437716 264948 523684 264976
rect 437716 264936 437722 264948
rect 523678 264936 523684 264948
rect 523736 264936 523742 264988
rect 664254 264936 664260 264988
rect 664312 264976 664318 264988
rect 664312 264948 669314 264976
rect 664312 264936 664318 264948
rect 669286 264920 669314 264948
rect 669286 264880 669320 264920
rect 669314 264868 669320 264880
rect 669372 264868 669378 264920
rect 435450 264732 435456 264784
rect 435508 264772 435514 264784
rect 545114 264772 545120 264784
rect 435508 264744 545120 264772
rect 435508 264732 435514 264744
rect 545114 264732 545120 264744
rect 545172 264732 545178 264784
rect 461210 264596 461216 264648
rect 461268 264636 461274 264648
rect 586514 264636 586520 264648
rect 461268 264608 586520 264636
rect 461268 264596 461274 264608
rect 586514 264596 586520 264608
rect 586572 264596 586578 264648
rect 471882 264460 471888 264512
rect 471940 264500 471946 264512
rect 603074 264500 603080 264512
rect 471940 264472 603080 264500
rect 471940 264460 471946 264472
rect 603074 264460 603080 264472
rect 603132 264460 603138 264512
rect 482186 264324 482192 264376
rect 482244 264364 482250 264376
rect 618898 264364 618904 264376
rect 482244 264336 618904 264364
rect 482244 264324 482250 264336
rect 618898 264324 618904 264336
rect 618956 264324 618962 264376
rect 51902 264188 51908 264240
rect 51960 264228 51966 264240
rect 655698 264228 655704 264240
rect 51960 264200 655704 264228
rect 51960 264188 51966 264200
rect 655698 264188 655704 264200
rect 655756 264188 655762 264240
rect 665082 263576 665088 263628
rect 665140 263616 665146 263628
rect 675478 263616 675484 263628
rect 665140 263588 675484 263616
rect 665140 263576 665146 263588
rect 675478 263576 675484 263588
rect 675536 263576 675542 263628
rect 673270 262896 673276 262948
rect 673328 262936 673334 262948
rect 675478 262936 675484 262948
rect 673328 262908 675484 262936
rect 673328 262896 673334 262908
rect 675478 262896 675484 262908
rect 675536 262896 675542 262948
rect 511534 261468 511540 261520
rect 511592 261508 511598 261520
rect 568574 261508 568580 261520
rect 511592 261480 568580 261508
rect 511592 261468 511598 261480
rect 568574 261468 568580 261480
rect 568632 261468 568638 261520
rect 671798 261264 671804 261316
rect 671856 261304 671862 261316
rect 675478 261304 675484 261316
rect 671856 261276 675484 261304
rect 671856 261264 671862 261276
rect 675478 261264 675484 261276
rect 675536 261264 675542 261316
rect 511350 259972 511356 260024
rect 511408 260012 511414 260024
rect 514018 260012 514024 260024
rect 511408 259984 514024 260012
rect 511408 259972 511414 259984
rect 514018 259972 514024 259984
rect 514076 259972 514082 260024
rect 669222 259700 669228 259752
rect 669280 259740 669286 259752
rect 675478 259740 675484 259752
rect 669280 259712 675484 259740
rect 669280 259700 669286 259712
rect 675478 259700 675484 259712
rect 675536 259700 675542 259752
rect 666370 259564 666376 259616
rect 666428 259604 666434 259616
rect 675478 259604 675484 259616
rect 666428 259576 675484 259604
rect 666428 259564 666434 259576
rect 675478 259564 675484 259576
rect 675536 259564 675542 259616
rect 666186 259428 666192 259480
rect 666244 259468 666250 259480
rect 675294 259468 675300 259480
rect 666244 259440 675300 259468
rect 666244 259428 666250 259440
rect 675294 259428 675300 259440
rect 675352 259428 675358 259480
rect 670418 259224 670424 259276
rect 670476 259264 670482 259276
rect 675478 259264 675484 259276
rect 670476 259236 675484 259264
rect 670476 259224 670482 259236
rect 675478 259224 675484 259236
rect 675536 259224 675542 259276
rect 672350 258408 672356 258460
rect 672408 258448 672414 258460
rect 675478 258448 675484 258460
rect 672408 258420 675484 258448
rect 672408 258408 672414 258420
rect 675478 258408 675484 258420
rect 675536 258408 675542 258460
rect 35802 258204 35808 258256
rect 35860 258244 35866 258256
rect 39942 258244 39948 258256
rect 35860 258216 39948 258244
rect 35860 258204 35866 258216
rect 39942 258204 39948 258216
rect 40000 258204 40006 258256
rect 35802 257116 35808 257168
rect 35860 257156 35866 257168
rect 39574 257156 39580 257168
rect 35860 257128 39580 257156
rect 35860 257116 35866 257128
rect 39574 257116 39580 257128
rect 39632 257116 39638 257168
rect 42058 256980 42064 257032
rect 42116 257020 42122 257032
rect 43806 257020 43812 257032
rect 42116 256992 43812 257020
rect 42116 256980 42122 256992
rect 43806 256980 43812 256992
rect 43864 256980 43870 257032
rect 41690 256952 41696 256964
rect 36004 256924 41696 256952
rect 35618 256844 35624 256896
rect 35676 256884 35682 256896
rect 36004 256884 36032 256924
rect 41690 256912 41696 256924
rect 41748 256912 41754 256964
rect 35676 256856 36032 256884
rect 35676 256844 35682 256856
rect 35434 256708 35440 256760
rect 35492 256748 35498 256760
rect 41690 256748 41696 256760
rect 35492 256720 41696 256748
rect 35492 256708 35498 256720
rect 41690 256708 41696 256720
rect 41748 256708 41754 256760
rect 42058 256708 42064 256760
rect 42116 256748 42122 256760
rect 45186 256748 45192 256760
rect 42116 256720 45192 256748
rect 42116 256708 42122 256720
rect 45186 256708 45192 256720
rect 45244 256708 45250 256760
rect 511442 256708 511448 256760
rect 511500 256748 511506 256760
rect 519538 256748 519544 256760
rect 511500 256720 519544 256748
rect 511500 256708 511506 256720
rect 519538 256708 519544 256720
rect 519596 256708 519602 256760
rect 675938 256708 675944 256760
rect 675996 256748 676002 256760
rect 683114 256748 683120 256760
rect 675996 256720 683120 256748
rect 675996 256708 676002 256720
rect 683114 256708 683120 256720
rect 683172 256708 683178 256760
rect 669774 256572 669780 256624
rect 669832 256612 669838 256624
rect 675478 256612 675484 256624
rect 669832 256584 675484 256612
rect 669832 256572 669838 256584
rect 675478 256572 675484 256584
rect 675536 256572 675542 256624
rect 35802 255688 35808 255740
rect 35860 255728 35866 255740
rect 40402 255728 40408 255740
rect 35860 255700 40408 255728
rect 35860 255688 35866 255700
rect 40402 255688 40408 255700
rect 40460 255688 40466 255740
rect 41690 255524 41696 255536
rect 41386 255496 41696 255524
rect 35618 255416 35624 255468
rect 35676 255456 35682 255468
rect 41386 255456 41414 255496
rect 41690 255484 41696 255496
rect 41748 255484 41754 255536
rect 42058 255484 42064 255536
rect 42116 255524 42122 255536
rect 42794 255524 42800 255536
rect 42116 255496 42800 255524
rect 42116 255484 42122 255496
rect 42794 255484 42800 255496
rect 42852 255484 42858 255536
rect 35676 255428 41414 255456
rect 35676 255416 35682 255428
rect 35434 255280 35440 255332
rect 35492 255320 35498 255332
rect 41690 255320 41696 255332
rect 35492 255292 41696 255320
rect 35492 255280 35498 255292
rect 41690 255280 41696 255292
rect 41748 255280 41754 255332
rect 42058 255280 42064 255332
rect 42116 255320 42122 255332
rect 45002 255320 45008 255332
rect 42116 255292 45008 255320
rect 42116 255280 42122 255292
rect 45002 255280 45008 255292
rect 45060 255280 45066 255332
rect 35802 254532 35808 254584
rect 35860 254572 35866 254584
rect 39758 254572 39764 254584
rect 35860 254544 39764 254572
rect 35860 254532 35866 254544
rect 39758 254532 39764 254544
rect 39816 254532 39822 254584
rect 35802 254260 35808 254312
rect 35860 254300 35866 254312
rect 40034 254300 40040 254312
rect 35860 254272 40040 254300
rect 35860 254260 35866 254272
rect 40034 254260 40040 254272
rect 40092 254260 40098 254312
rect 35618 254124 35624 254176
rect 35676 254164 35682 254176
rect 35676 254136 38654 254164
rect 35676 254124 35682 254136
rect 38626 254096 38654 254136
rect 41230 254096 41236 254108
rect 38626 254068 41236 254096
rect 41230 254056 41236 254068
rect 41288 254056 41294 254108
rect 35434 253920 35440 253972
rect 35492 253960 35498 253972
rect 41690 253960 41696 253972
rect 35492 253932 41696 253960
rect 35492 253920 35498 253932
rect 41690 253920 41696 253932
rect 41748 253920 41754 253972
rect 42058 253920 42064 253972
rect 42116 253960 42122 253972
rect 44542 253960 44548 253972
rect 42116 253932 44548 253960
rect 42116 253920 42122 253932
rect 44542 253920 44548 253932
rect 44600 253920 44606 253972
rect 35802 252696 35808 252748
rect 35860 252736 35866 252748
rect 41690 252736 41696 252748
rect 35860 252708 41696 252736
rect 35860 252696 35866 252708
rect 41690 252696 41696 252708
rect 41748 252696 41754 252748
rect 35526 252560 35532 252612
rect 35584 252600 35590 252612
rect 40034 252600 40040 252612
rect 35584 252572 40040 252600
rect 35584 252560 35590 252572
rect 40034 252560 40040 252572
rect 40092 252560 40098 252612
rect 511902 252560 511908 252612
rect 511960 252600 511966 252612
rect 562318 252600 562324 252612
rect 511960 252572 562324 252600
rect 511960 252560 511966 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 35802 251472 35808 251524
rect 35860 251512 35866 251524
rect 41506 251512 41512 251524
rect 35860 251484 41512 251512
rect 35860 251472 35866 251484
rect 41506 251472 41512 251484
rect 41564 251472 41570 251524
rect 35526 251200 35532 251252
rect 35584 251240 35590 251252
rect 41690 251240 41696 251252
rect 35584 251212 41696 251240
rect 35584 251200 35590 251212
rect 41690 251200 41696 251212
rect 41748 251200 41754 251252
rect 35802 250180 35808 250232
rect 35860 250220 35866 250232
rect 39390 250220 39396 250232
rect 35860 250192 39396 250220
rect 35860 250180 35866 250192
rect 39390 250180 39396 250192
rect 39448 250180 39454 250232
rect 35434 249908 35440 249960
rect 35492 249948 35498 249960
rect 39850 249948 39856 249960
rect 35492 249920 39856 249948
rect 35492 249908 35498 249920
rect 39850 249908 39856 249920
rect 39908 249908 39914 249960
rect 35618 249772 35624 249824
rect 35676 249812 35682 249824
rect 41690 249812 41696 249824
rect 35676 249784 41696 249812
rect 35676 249772 35682 249784
rect 41690 249772 41696 249784
rect 41748 249772 41754 249824
rect 42058 249772 42064 249824
rect 42116 249812 42122 249824
rect 47210 249812 47216 249824
rect 42116 249784 47216 249812
rect 42116 249772 42122 249784
rect 47210 249772 47216 249784
rect 47268 249772 47274 249824
rect 510614 249772 510620 249824
rect 510672 249812 510678 249824
rect 513282 249812 513288 249824
rect 510672 249784 513288 249812
rect 510672 249772 510678 249784
rect 513282 249772 513288 249784
rect 513340 249772 513346 249824
rect 40034 249500 40040 249552
rect 40092 249540 40098 249552
rect 41690 249540 41696 249552
rect 40092 249512 41696 249540
rect 40092 249500 40098 249512
rect 41690 249500 41696 249512
rect 41748 249500 41754 249552
rect 42058 249432 42064 249484
rect 42116 249472 42122 249484
rect 42610 249472 42616 249484
rect 42116 249444 42616 249472
rect 42116 249432 42122 249444
rect 42610 249432 42616 249444
rect 42668 249432 42674 249484
rect 511166 249024 511172 249076
rect 511224 249064 511230 249076
rect 571334 249064 571340 249076
rect 511224 249036 571340 249064
rect 511224 249024 511230 249036
rect 571334 249024 571340 249036
rect 571392 249024 571398 249076
rect 35802 248820 35808 248872
rect 35860 248860 35866 248872
rect 40126 248860 40132 248872
rect 35860 248832 40132 248860
rect 35860 248820 35866 248832
rect 40126 248820 40132 248832
rect 40184 248820 40190 248872
rect 35434 248548 35440 248600
rect 35492 248588 35498 248600
rect 39114 248588 39120 248600
rect 35492 248560 39120 248588
rect 35492 248548 35498 248560
rect 39114 248548 39120 248560
rect 39172 248548 39178 248600
rect 35618 248412 35624 248464
rect 35676 248452 35682 248464
rect 41690 248452 41696 248464
rect 35676 248424 41696 248452
rect 35676 248412 35682 248424
rect 41690 248412 41696 248424
rect 41748 248412 41754 248464
rect 42058 248412 42064 248464
rect 42116 248452 42122 248464
rect 44358 248452 44364 248464
rect 42116 248424 44364 248452
rect 42116 248412 42122 248424
rect 44358 248412 44364 248424
rect 44416 248412 44422 248464
rect 35802 247460 35808 247512
rect 35860 247500 35866 247512
rect 40402 247500 40408 247512
rect 35860 247472 40408 247500
rect 35860 247460 35866 247472
rect 40402 247460 40408 247472
rect 40460 247460 40466 247512
rect 35618 247188 35624 247240
rect 35676 247228 35682 247240
rect 41690 247228 41696 247240
rect 35676 247200 41696 247228
rect 35676 247188 35682 247200
rect 41690 247188 41696 247200
rect 41748 247188 41754 247240
rect 42058 247188 42064 247240
rect 42116 247228 42122 247240
rect 128998 247228 129004 247240
rect 42116 247200 129004 247228
rect 42116 247188 42122 247200
rect 128998 247188 129004 247200
rect 129056 247188 129062 247240
rect 35802 247052 35808 247104
rect 35860 247092 35866 247104
rect 41690 247092 41696 247104
rect 35860 247064 41696 247092
rect 35860 247052 35866 247064
rect 41690 247052 41696 247064
rect 41748 247052 41754 247104
rect 42058 247052 42064 247104
rect 42116 247092 42122 247104
rect 128814 247092 128820 247104
rect 42116 247064 128820 247092
rect 42116 247052 42122 247064
rect 128814 247052 128820 247064
rect 128872 247052 128878 247104
rect 674466 246984 674472 247036
rect 674524 247024 674530 247036
rect 674834 247024 674840 247036
rect 674524 246996 674840 247024
rect 674524 246984 674530 246996
rect 674834 246984 674840 246996
rect 674892 246984 674898 247036
rect 513282 246304 513288 246356
rect 513340 246344 513346 246356
rect 569954 246344 569960 246356
rect 513340 246316 569960 246344
rect 513340 246304 513346 246316
rect 569954 246304 569960 246316
rect 570012 246304 570018 246356
rect 669406 245148 669412 245200
rect 669464 245188 669470 245200
rect 675386 245188 675392 245200
rect 669464 245160 675392 245188
rect 669464 245148 669470 245160
rect 675386 245148 675392 245160
rect 675444 245148 675450 245200
rect 666186 242836 666192 242888
rect 666244 242876 666250 242888
rect 669406 242876 669412 242888
rect 666244 242848 669412 242876
rect 666244 242836 666250 242848
rect 669406 242836 669412 242848
rect 669464 242836 669470 242888
rect 670418 242836 670424 242888
rect 670476 242876 670482 242888
rect 675110 242876 675116 242888
rect 670476 242848 675116 242876
rect 670476 242836 670482 242848
rect 675110 242836 675116 242848
rect 675168 242836 675174 242888
rect 511258 242292 511264 242344
rect 511316 242332 511322 242344
rect 628558 242332 628564 242344
rect 511316 242304 628564 242332
rect 511316 242292 511322 242304
rect 628558 242292 628564 242304
rect 628616 242292 628622 242344
rect 31018 242156 31024 242208
rect 31076 242196 31082 242208
rect 41690 242196 41696 242208
rect 31076 242168 41696 242196
rect 31076 242156 31082 242168
rect 41690 242156 41696 242168
rect 41748 242156 41754 242208
rect 511994 242156 512000 242208
rect 512052 242196 512058 242208
rect 633434 242196 633440 242208
rect 512052 242168 633440 242196
rect 512052 242156 512058 242168
rect 633434 242156 633440 242168
rect 633492 242156 633498 242208
rect 669222 241680 669228 241732
rect 669280 241720 669286 241732
rect 675110 241720 675116 241732
rect 669280 241692 675116 241720
rect 669280 241680 669286 241692
rect 675110 241680 675116 241692
rect 675168 241680 675174 241732
rect 674650 241408 674656 241460
rect 674708 241448 674714 241460
rect 675110 241448 675116 241460
rect 674708 241420 675116 241448
rect 674708 241408 674714 241420
rect 675110 241408 675116 241420
rect 675168 241408 675174 241460
rect 519538 240728 519544 240780
rect 519596 240768 519602 240780
rect 567194 240768 567200 240780
rect 519596 240740 567200 240768
rect 519596 240728 519602 240740
rect 567194 240728 567200 240740
rect 567252 240728 567258 240780
rect 44174 239912 44180 239964
rect 44232 239952 44238 239964
rect 44634 239952 44640 239964
rect 44232 239924 44640 239952
rect 44232 239912 44238 239924
rect 44634 239912 44640 239924
rect 44692 239912 44698 239964
rect 514018 238144 514024 238196
rect 514076 238184 514082 238196
rect 568758 238184 568764 238196
rect 514076 238156 568764 238184
rect 514076 238144 514082 238156
rect 568758 238144 568764 238156
rect 568816 238144 568822 238196
rect 511258 238008 511264 238060
rect 511316 238048 511322 238060
rect 632698 238048 632704 238060
rect 511316 238020 632704 238048
rect 511316 238008 511322 238020
rect 632698 238008 632704 238020
rect 632756 238008 632762 238060
rect 666370 237328 666376 237380
rect 666428 237368 666434 237380
rect 675294 237368 675300 237380
rect 666428 237340 675300 237368
rect 666428 237328 666434 237340
rect 675294 237328 675300 237340
rect 675352 237328 675358 237380
rect 42426 235900 42432 235952
rect 42484 235940 42490 235952
rect 44634 235940 44640 235952
rect 42484 235912 44640 235940
rect 42484 235900 42490 235912
rect 44634 235900 44640 235912
rect 44692 235900 44698 235952
rect 42426 234540 42432 234592
rect 42484 234580 42490 234592
rect 43806 234580 43812 234592
rect 42484 234552 43812 234580
rect 42484 234540 42490 234552
rect 43806 234540 43812 234552
rect 43864 234540 43870 234592
rect 42426 234200 42432 234252
rect 42484 234240 42490 234252
rect 42978 234240 42984 234252
rect 42484 234212 42984 234240
rect 42484 234200 42490 234212
rect 42978 234200 42984 234212
rect 43036 234200 43042 234252
rect 510890 233996 510896 234048
rect 510948 234036 510954 234048
rect 577498 234036 577504 234048
rect 510948 234008 577504 234036
rect 510948 233996 510954 234008
rect 577498 233996 577504 234008
rect 577556 233996 577562 234048
rect 510706 233860 510712 233912
rect 510764 233900 510770 233912
rect 629938 233900 629944 233912
rect 510764 233872 629944 233900
rect 510764 233860 510770 233872
rect 629938 233860 629944 233872
rect 629996 233860 630002 233912
rect 42426 231820 42432 231872
rect 42484 231860 42490 231872
rect 47026 231860 47032 231872
rect 42484 231832 47032 231860
rect 42484 231820 42490 231832
rect 47026 231820 47032 231832
rect 47084 231820 47090 231872
rect 55858 231752 55864 231804
rect 55916 231792 55922 231804
rect 646038 231792 646044 231804
rect 55916 231764 646044 231792
rect 55916 231752 55922 231764
rect 646038 231752 646044 231764
rect 646096 231752 646102 231804
rect 42426 231684 42432 231736
rect 42484 231724 42490 231736
rect 44358 231724 44364 231736
rect 42484 231696 44364 231724
rect 42484 231684 42490 231696
rect 44358 231684 44364 231696
rect 44416 231684 44422 231736
rect 46198 231616 46204 231668
rect 46256 231656 46262 231668
rect 643094 231656 643100 231668
rect 46256 231628 643100 231656
rect 46256 231616 46262 231628
rect 643094 231616 643100 231628
rect 643152 231616 643158 231668
rect 51718 231480 51724 231532
rect 51776 231520 51782 231532
rect 650546 231520 650552 231532
rect 51776 231492 650552 231520
rect 51776 231480 51782 231492
rect 650546 231480 650552 231492
rect 650604 231480 650610 231532
rect 47578 231344 47584 231396
rect 47636 231384 47642 231396
rect 645854 231384 645860 231396
rect 47636 231356 645860 231384
rect 47636 231344 47642 231356
rect 645854 231344 645860 231356
rect 645912 231344 645918 231396
rect 44818 231208 44824 231260
rect 44876 231248 44882 231260
rect 644474 231248 644480 231260
rect 44876 231220 644480 231248
rect 44876 231208 44882 231220
rect 644474 231208 644480 231220
rect 644532 231208 644538 231260
rect 50522 231072 50528 231124
rect 50580 231112 50586 231124
rect 652754 231112 652760 231124
rect 50580 231084 652760 231112
rect 50580 231072 50586 231084
rect 652754 231072 652760 231084
rect 652812 231072 652818 231124
rect 53098 230936 53104 230988
rect 53156 230976 53162 230988
rect 641806 230976 641812 230988
rect 53156 230948 641812 230976
rect 53156 230936 53162 230948
rect 641806 230936 641812 230948
rect 641864 230936 641870 230988
rect 132586 230800 132592 230852
rect 132644 230840 132650 230852
rect 661310 230840 661316 230852
rect 132644 230812 661316 230840
rect 132644 230800 132650 230812
rect 661310 230800 661316 230812
rect 661368 230800 661374 230852
rect 108942 230732 108948 230784
rect 109000 230772 109006 230784
rect 117038 230772 117044 230784
rect 109000 230744 117044 230772
rect 109000 230732 109006 230744
rect 117038 230732 117044 230744
rect 117096 230732 117102 230784
rect 117222 230732 117228 230784
rect 117280 230772 117286 230784
rect 132402 230772 132408 230784
rect 117280 230744 132408 230772
rect 117280 230732 117286 230744
rect 132402 230732 132408 230744
rect 132460 230732 132466 230784
rect 181254 230664 181260 230716
rect 181312 230704 181318 230716
rect 183094 230704 183100 230716
rect 181312 230676 183100 230704
rect 181312 230664 181318 230676
rect 183094 230664 183100 230676
rect 183152 230664 183158 230716
rect 474642 230664 474648 230716
rect 474700 230704 474706 230716
rect 478046 230704 478052 230716
rect 474700 230676 478052 230704
rect 474700 230664 474706 230676
rect 478046 230664 478052 230676
rect 478104 230664 478110 230716
rect 481266 230664 481272 230716
rect 481324 230704 481330 230716
rect 507486 230704 507492 230716
rect 481324 230676 507492 230704
rect 481324 230664 481330 230676
rect 507486 230664 507492 230676
rect 507544 230664 507550 230716
rect 89622 230596 89628 230648
rect 89680 230636 89686 230648
rect 171226 230636 171232 230648
rect 89680 230608 171232 230636
rect 89680 230596 89686 230608
rect 171226 230596 171232 230608
rect 171284 230596 171290 230648
rect 184474 230568 184480 230580
rect 176626 230540 184480 230568
rect 79962 230460 79968 230512
rect 80020 230500 80026 230512
rect 116854 230500 116860 230512
rect 80020 230472 116860 230500
rect 80020 230460 80026 230472
rect 116854 230460 116860 230472
rect 116912 230460 116918 230512
rect 117038 230460 117044 230512
rect 117096 230500 117102 230512
rect 176626 230500 176654 230540
rect 184474 230528 184480 230540
rect 184532 230528 184538 230580
rect 189166 230568 189172 230580
rect 187252 230540 189172 230568
rect 117096 230472 176654 230500
rect 117096 230460 117102 230472
rect 42150 230392 42156 230444
rect 42208 230432 42214 230444
rect 43162 230432 43168 230444
rect 42208 230404 43168 230432
rect 42208 230392 42214 230404
rect 43162 230392 43168 230404
rect 43220 230392 43226 230444
rect 176838 230392 176844 230444
rect 176896 230432 176902 230444
rect 181254 230432 181260 230444
rect 176896 230404 181260 230432
rect 176896 230392 176902 230404
rect 181254 230392 181260 230404
rect 181312 230392 181318 230444
rect 181438 230392 181444 230444
rect 181496 230432 181502 230444
rect 187252 230432 187280 230540
rect 189166 230528 189172 230540
rect 189224 230528 189230 230580
rect 191742 230528 191748 230580
rect 191800 230568 191806 230580
rect 193582 230568 193588 230580
rect 191800 230540 193588 230568
rect 191800 230528 191806 230540
rect 193582 230528 193588 230540
rect 193640 230528 193646 230580
rect 204714 230528 204720 230580
rect 204772 230568 204778 230580
rect 438026 230568 438032 230580
rect 204772 230540 205036 230568
rect 204772 230528 204778 230540
rect 181496 230404 187280 230432
rect 181496 230392 181502 230404
rect 187418 230392 187424 230444
rect 187476 230432 187482 230444
rect 190270 230432 190276 230444
rect 187476 230404 190276 230432
rect 187476 230392 187482 230404
rect 190270 230392 190276 230404
rect 190328 230392 190334 230444
rect 190454 230392 190460 230444
rect 190512 230432 190518 230444
rect 205008 230432 205036 230540
rect 437584 230540 438032 230568
rect 205450 230432 205456 230444
rect 190512 230404 204944 230432
rect 205008 230404 205456 230432
rect 190512 230392 190518 230404
rect 107562 230256 107568 230308
rect 107620 230296 107626 230308
rect 182818 230296 182824 230308
rect 107620 230268 182824 230296
rect 107620 230256 107626 230268
rect 182818 230256 182824 230268
rect 182876 230256 182882 230308
rect 183462 230256 183468 230308
rect 183520 230296 183526 230308
rect 203242 230296 203248 230308
rect 183520 230268 203248 230296
rect 183520 230256 183526 230268
rect 203242 230256 203248 230268
rect 203300 230256 203306 230308
rect 82906 230120 82912 230172
rect 82964 230160 82970 230172
rect 153746 230160 153752 230172
rect 82964 230132 153752 230160
rect 82964 230120 82970 230132
rect 153746 230120 153752 230132
rect 153804 230120 153810 230172
rect 153930 230120 153936 230172
rect 153988 230160 153994 230172
rect 156322 230160 156328 230172
rect 153988 230132 156328 230160
rect 153988 230120 153994 230132
rect 156322 230120 156328 230132
rect 156380 230120 156386 230172
rect 166810 230160 166816 230172
rect 157306 230132 166816 230160
rect 88242 229984 88248 230036
rect 88300 230024 88306 230036
rect 157306 230024 157334 230132
rect 166810 230120 166816 230132
rect 166868 230120 166874 230172
rect 166994 230120 167000 230172
rect 167052 230160 167058 230172
rect 204714 230160 204720 230172
rect 167052 230132 204720 230160
rect 167052 230120 167058 230132
rect 204714 230120 204720 230132
rect 204772 230120 204778 230172
rect 204916 230160 204944 230404
rect 205450 230392 205456 230404
rect 205508 230392 205514 230444
rect 206002 230392 206008 230444
rect 206060 230432 206066 230444
rect 244642 230432 244648 230444
rect 206060 230404 244648 230432
rect 206060 230392 206066 230404
rect 244642 230392 244648 230404
rect 244700 230392 244706 230444
rect 256326 230392 256332 230444
rect 256384 230432 256390 230444
rect 279970 230432 279976 230444
rect 256384 230404 279976 230432
rect 256384 230392 256390 230404
rect 279970 230392 279976 230404
rect 280028 230392 280034 230444
rect 290458 230392 290464 230444
rect 290516 230432 290522 230444
rect 295426 230432 295432 230444
rect 290516 230404 295432 230432
rect 290516 230392 290522 230404
rect 295426 230392 295432 230404
rect 295484 230392 295490 230444
rect 388162 230392 388168 230444
rect 388220 230432 388226 230444
rect 390738 230432 390744 230444
rect 388220 230404 390744 230432
rect 388220 230392 388226 230404
rect 390738 230392 390744 230404
rect 390796 230392 390802 230444
rect 403250 230432 403256 230444
rect 398576 230404 403256 230432
rect 284938 230324 284944 230376
rect 284996 230364 285002 230376
rect 286594 230364 286600 230376
rect 284996 230336 286600 230364
rect 284996 230324 285002 230336
rect 286594 230324 286600 230336
rect 286652 230324 286658 230376
rect 296714 230324 296720 230376
rect 296772 230364 296778 230376
rect 299290 230364 299296 230376
rect 296772 230336 299296 230364
rect 296772 230324 296778 230336
rect 299290 230324 299296 230336
rect 299348 230324 299354 230376
rect 300486 230324 300492 230376
rect 300544 230364 300550 230376
rect 301498 230364 301504 230376
rect 300544 230336 301504 230364
rect 300544 230324 300550 230336
rect 301498 230324 301504 230336
rect 301556 230324 301562 230376
rect 319438 230324 319444 230376
rect 319496 230364 319502 230376
rect 320266 230364 320272 230376
rect 319496 230336 320272 230364
rect 319496 230324 319502 230336
rect 320266 230324 320272 230336
rect 320324 230324 320330 230376
rect 331858 230324 331864 230376
rect 331916 230364 331922 230376
rect 333054 230364 333060 230376
rect 331916 230336 333060 230364
rect 331916 230324 331922 230336
rect 333054 230324 333060 230336
rect 333112 230324 333118 230376
rect 333514 230324 333520 230376
rect 333572 230364 333578 230376
rect 334526 230364 334532 230376
rect 333572 230336 334532 230364
rect 333572 230324 333578 230336
rect 334526 230324 334532 230336
rect 334584 230324 334590 230376
rect 339586 230324 339592 230376
rect 339644 230364 339650 230376
rect 340966 230364 340972 230376
rect 339644 230336 340972 230364
rect 339644 230324 339650 230336
rect 340966 230324 340972 230336
rect 341024 230324 341030 230376
rect 353386 230324 353392 230376
rect 353444 230364 353450 230376
rect 354582 230364 354588 230376
rect 353444 230336 354588 230364
rect 353444 230324 353450 230336
rect 354582 230324 354588 230336
rect 354640 230324 354646 230376
rect 355042 230324 355048 230376
rect 355100 230364 355106 230376
rect 356698 230364 356704 230376
rect 355100 230336 356704 230364
rect 355100 230324 355106 230336
rect 356698 230324 356704 230336
rect 356756 230324 356762 230376
rect 359458 230324 359464 230376
rect 359516 230364 359522 230376
rect 361482 230364 361488 230376
rect 359516 230336 361488 230364
rect 359516 230324 359522 230336
rect 361482 230324 361488 230336
rect 361540 230324 361546 230376
rect 364426 230324 364432 230376
rect 364484 230364 364490 230376
rect 365622 230364 365628 230376
rect 364484 230336 365628 230364
rect 364484 230324 364490 230336
rect 365622 230324 365628 230336
rect 365680 230324 365686 230376
rect 371602 230324 371608 230376
rect 371660 230364 371666 230376
rect 373626 230364 373632 230376
rect 371660 230336 373632 230364
rect 371660 230324 371666 230336
rect 373626 230324 373632 230336
rect 373684 230324 373690 230376
rect 376570 230324 376576 230376
rect 376628 230364 376634 230376
rect 377858 230364 377864 230376
rect 376628 230336 377864 230364
rect 376628 230324 376634 230336
rect 377858 230324 377864 230336
rect 377916 230324 377922 230376
rect 378226 230324 378232 230376
rect 378284 230364 378290 230376
rect 379146 230364 379152 230376
rect 378284 230336 379152 230364
rect 378284 230324 378290 230336
rect 379146 230324 379152 230336
rect 379204 230324 379210 230376
rect 391474 230324 391480 230376
rect 391532 230364 391538 230376
rect 392578 230364 392584 230376
rect 391532 230336 392584 230364
rect 391532 230324 391538 230336
rect 392578 230324 392584 230336
rect 392636 230324 392642 230376
rect 395890 230324 395896 230376
rect 395948 230364 395954 230376
rect 396718 230364 396724 230376
rect 395948 230336 396724 230364
rect 395948 230324 395954 230336
rect 396718 230324 396724 230336
rect 396776 230324 396782 230376
rect 205082 230256 205088 230308
rect 205140 230296 205146 230308
rect 240226 230296 240232 230308
rect 205140 230268 240232 230296
rect 205140 230256 205146 230268
rect 240226 230256 240232 230268
rect 240284 230256 240290 230308
rect 247770 230256 247776 230308
rect 247828 230296 247834 230308
rect 275554 230296 275560 230308
rect 247828 230268 275560 230296
rect 247828 230256 247834 230268
rect 275554 230256 275560 230268
rect 275612 230256 275618 230308
rect 380986 230256 380992 230308
rect 381044 230296 381050 230308
rect 389082 230296 389088 230308
rect 381044 230268 389088 230296
rect 381044 230256 381050 230268
rect 389082 230256 389088 230268
rect 389140 230256 389146 230308
rect 338022 230188 338028 230240
rect 338080 230228 338086 230240
rect 341426 230228 341432 230240
rect 338080 230200 341432 230228
rect 338080 230188 338086 230200
rect 341426 230188 341432 230200
rect 341484 230188 341490 230240
rect 341794 230188 341800 230240
rect 341852 230228 341858 230240
rect 343726 230228 343732 230240
rect 341852 230200 343732 230228
rect 341852 230188 341858 230200
rect 343726 230188 343732 230200
rect 343784 230188 343790 230240
rect 345658 230188 345664 230240
rect 345716 230228 345722 230240
rect 349706 230228 349712 230240
rect 345716 230200 349712 230228
rect 345716 230188 345722 230200
rect 349706 230188 349712 230200
rect 349764 230188 349770 230240
rect 357250 230188 357256 230240
rect 357308 230228 357314 230240
rect 359734 230228 359740 230240
rect 357308 230200 359740 230228
rect 357308 230188 357314 230200
rect 359734 230188 359740 230200
rect 359792 230188 359798 230240
rect 369394 230188 369400 230240
rect 369452 230228 369458 230240
rect 371878 230228 371884 230240
rect 369452 230200 371884 230228
rect 369452 230188 369458 230200
rect 371878 230188 371884 230200
rect 371936 230188 371942 230240
rect 394050 230228 394056 230240
rect 392964 230200 394056 230228
rect 235810 230160 235816 230172
rect 204916 230132 235816 230160
rect 235810 230120 235816 230132
rect 235868 230120 235874 230172
rect 235994 230120 236000 230172
rect 236052 230160 236058 230172
rect 238570 230160 238576 230172
rect 236052 230132 238576 230160
rect 236052 230120 236058 230132
rect 238570 230120 238576 230132
rect 238628 230120 238634 230172
rect 240962 230120 240968 230172
rect 241020 230160 241026 230172
rect 271138 230160 271144 230172
rect 241020 230132 271144 230160
rect 241020 230120 241026 230132
rect 271138 230120 271144 230132
rect 271196 230120 271202 230172
rect 279878 230120 279884 230172
rect 279936 230160 279942 230172
rect 297634 230160 297640 230172
rect 279936 230132 297640 230160
rect 279936 230120 279942 230132
rect 297634 230120 297640 230132
rect 297692 230120 297698 230172
rect 335722 230120 335728 230172
rect 335780 230160 335786 230172
rect 337286 230160 337292 230172
rect 335780 230132 337292 230160
rect 335780 230120 335786 230132
rect 337286 230120 337292 230132
rect 337344 230120 337350 230172
rect 361114 230120 361120 230172
rect 361172 230160 361178 230172
rect 363966 230160 363972 230172
rect 361172 230132 363972 230160
rect 361172 230120 361178 230132
rect 363966 230120 363972 230132
rect 364024 230120 364030 230172
rect 374914 230120 374920 230172
rect 374972 230160 374978 230172
rect 381170 230160 381176 230172
rect 374972 230132 381176 230160
rect 374972 230120 374978 230132
rect 381170 230120 381176 230132
rect 381228 230120 381234 230172
rect 298738 230052 298744 230104
rect 298796 230092 298802 230104
rect 299842 230092 299848 230104
rect 298796 230064 299848 230092
rect 298796 230052 298802 230064
rect 299842 230052 299848 230064
rect 299900 230052 299906 230104
rect 338482 230052 338488 230104
rect 338540 230092 338546 230104
rect 342714 230092 342720 230104
rect 338540 230064 342720 230092
rect 338540 230052 338546 230064
rect 342714 230052 342720 230064
rect 342772 230052 342778 230104
rect 383194 230052 383200 230104
rect 383252 230092 383258 230104
rect 390002 230092 390008 230104
rect 383252 230064 390008 230092
rect 383252 230052 383258 230064
rect 390002 230052 390008 230064
rect 390060 230052 390066 230104
rect 390370 230052 390376 230104
rect 390428 230092 390434 230104
rect 392964 230092 392992 230200
rect 394050 230188 394056 230200
rect 394108 230188 394114 230240
rect 394234 230188 394240 230240
rect 394292 230228 394298 230240
rect 397178 230228 397184 230240
rect 394292 230200 397184 230228
rect 394292 230188 394298 230200
rect 397178 230188 397184 230200
rect 397236 230188 397242 230240
rect 390428 230064 392992 230092
rect 390428 230052 390434 230064
rect 88300 229996 157334 230024
rect 88300 229984 88306 229996
rect 159726 229984 159732 230036
rect 159784 230024 159790 230036
rect 168834 230024 168840 230036
rect 159784 229996 168840 230024
rect 159784 229984 159790 229996
rect 168834 229984 168840 229996
rect 168892 229984 168898 230036
rect 169018 229984 169024 230036
rect 169076 230024 169082 230036
rect 170122 230024 170128 230036
rect 169076 229996 170128 230024
rect 169076 229984 169082 229996
rect 170122 229984 170128 229996
rect 170180 229984 170186 230036
rect 171134 229984 171140 230036
rect 171192 230024 171198 230036
rect 174538 230024 174544 230036
rect 171192 229996 174544 230024
rect 171192 229984 171198 229996
rect 174538 229984 174544 229996
rect 174596 229984 174602 230036
rect 174998 229984 175004 230036
rect 175056 230024 175062 230036
rect 191742 230024 191748 230036
rect 175056 229996 191748 230024
rect 175056 229984 175062 229996
rect 191742 229984 191748 229996
rect 191800 229984 191806 230036
rect 192110 229984 192116 230036
rect 192168 230024 192174 230036
rect 193306 230024 193312 230036
rect 192168 229996 193312 230024
rect 192168 229984 192174 229996
rect 193306 229984 193312 229996
rect 193364 229984 193370 230036
rect 195238 229984 195244 230036
rect 195296 230024 195302 230036
rect 231394 230024 231400 230036
rect 195296 229996 231400 230024
rect 195296 229984 195302 229996
rect 231394 229984 231400 229996
rect 231452 229984 231458 230036
rect 243538 229984 243544 230036
rect 243596 230024 243602 230036
rect 266722 230024 266728 230036
rect 243596 229996 266728 230024
rect 243596 229984 243602 229996
rect 266722 229984 266728 229996
rect 266780 229984 266786 230036
rect 275646 229984 275652 230036
rect 275704 230024 275710 230036
rect 293218 230024 293224 230036
rect 275704 229996 293224 230024
rect 275704 229984 275710 229996
rect 293218 229984 293224 229996
rect 293276 229984 293282 230036
rect 305638 229984 305644 230036
rect 305696 230024 305702 230036
rect 313090 230024 313096 230036
rect 305696 229996 313096 230024
rect 305696 229984 305702 229996
rect 313090 229984 313096 229996
rect 313148 229984 313154 230036
rect 344002 229984 344008 230036
rect 344060 230024 344066 230036
rect 348234 230024 348240 230036
rect 344060 229996 348240 230024
rect 344060 229984 344066 229996
rect 348234 229984 348240 229996
rect 348292 229984 348298 230036
rect 349522 229984 349528 230036
rect 349580 230024 349586 230036
rect 356330 230024 356336 230036
rect 349580 229996 356336 230024
rect 349580 229984 349586 229996
rect 356330 229984 356336 229996
rect 356388 229984 356394 230036
rect 363322 229984 363328 230036
rect 363380 230024 363386 230036
rect 368382 230024 368388 230036
rect 363380 229996 368388 230024
rect 363380 229984 363386 229996
rect 368382 229984 368388 229996
rect 368440 229984 368446 230036
rect 372706 229984 372712 230036
rect 372764 230024 372770 230036
rect 382274 230024 382280 230036
rect 372764 229996 382280 230024
rect 372764 229984 372770 229996
rect 382274 229984 382280 229996
rect 382332 229984 382338 230036
rect 397914 230024 397920 230036
rect 393056 229996 397920 230024
rect 339034 229916 339040 229968
rect 339092 229956 339098 229968
rect 340138 229956 340144 229968
rect 339092 229928 340144 229956
rect 339092 229916 339098 229928
rect 340138 229916 340144 229928
rect 340196 229916 340202 229968
rect 390738 229916 390744 229968
rect 390796 229956 390802 229968
rect 393056 229956 393084 229996
rect 397914 229984 397920 229996
rect 397972 229984 397978 230036
rect 390796 229928 393084 229956
rect 390796 229916 390802 229928
rect 69658 229848 69664 229900
rect 69716 229888 69722 229900
rect 153930 229888 153936 229900
rect 69716 229860 153936 229888
rect 69716 229848 69722 229860
rect 153930 229848 153936 229860
rect 153988 229848 153994 229900
rect 154114 229848 154120 229900
rect 154172 229888 154178 229900
rect 154172 229860 159956 229888
rect 154172 229848 154178 229860
rect 66898 229712 66904 229764
rect 66956 229752 66962 229764
rect 144638 229752 144644 229764
rect 66956 229724 144644 229752
rect 66956 229712 66962 229724
rect 144638 229712 144644 229724
rect 144696 229712 144702 229764
rect 144822 229712 144828 229764
rect 144880 229752 144886 229764
rect 150250 229752 150256 229764
rect 144880 229724 150256 229752
rect 144880 229712 144886 229724
rect 150250 229712 150256 229724
rect 150308 229712 150314 229764
rect 150434 229712 150440 229764
rect 150492 229752 150498 229764
rect 159726 229752 159732 229764
rect 150492 229724 159732 229752
rect 150492 229712 150498 229724
rect 159726 229712 159732 229724
rect 159784 229712 159790 229764
rect 159928 229752 159956 229860
rect 160738 229848 160744 229900
rect 160796 229888 160802 229900
rect 214098 229888 214104 229900
rect 160796 229860 214104 229888
rect 160796 229848 160802 229860
rect 214098 229848 214104 229860
rect 214156 229848 214162 229900
rect 214466 229848 214472 229900
rect 214524 229888 214530 229900
rect 216490 229888 216496 229900
rect 214524 229860 216496 229888
rect 214524 229848 214530 229860
rect 216490 229848 216496 229860
rect 216548 229848 216554 229900
rect 220446 229848 220452 229900
rect 220504 229888 220510 229900
rect 257890 229888 257896 229900
rect 220504 229860 257896 229888
rect 220504 229848 220510 229860
rect 257890 229848 257896 229860
rect 257948 229848 257954 229900
rect 266998 229848 267004 229900
rect 267056 229888 267062 229900
rect 288802 229888 288808 229900
rect 267056 229860 288808 229888
rect 267056 229848 267062 229860
rect 288802 229848 288808 229860
rect 288860 229848 288866 229900
rect 297358 229848 297364 229900
rect 297416 229888 297422 229900
rect 308674 229888 308680 229900
rect 297416 229860 308680 229888
rect 297416 229848 297422 229860
rect 308674 229848 308680 229860
rect 308732 229848 308738 229900
rect 308858 229848 308864 229900
rect 308916 229888 308922 229900
rect 317506 229888 317512 229900
rect 308916 229860 317512 229888
rect 308916 229848 308922 229860
rect 317506 229848 317512 229860
rect 317564 229848 317570 229900
rect 341242 229848 341248 229900
rect 341300 229888 341306 229900
rect 344094 229888 344100 229900
rect 341300 229860 344100 229888
rect 341300 229848 341306 229860
rect 344094 229848 344100 229860
rect 344152 229848 344158 229900
rect 358906 229848 358912 229900
rect 358964 229888 358970 229900
rect 362402 229888 362408 229900
rect 358964 229860 362408 229888
rect 358964 229848 358970 229860
rect 362402 229848 362408 229860
rect 362460 229848 362466 229900
rect 365806 229848 365812 229900
rect 365864 229888 365870 229900
rect 378042 229888 378048 229900
rect 365864 229860 378048 229888
rect 365864 229848 365870 229860
rect 378042 229848 378048 229860
rect 378100 229848 378106 229900
rect 389266 229848 389272 229900
rect 389324 229888 389330 229900
rect 390462 229888 390468 229900
rect 389324 229860 390468 229888
rect 389324 229848 389330 229860
rect 390462 229848 390468 229860
rect 390520 229848 390526 229900
rect 395154 229848 395160 229900
rect 395212 229888 395218 229900
rect 398576 229888 398604 230404
rect 403250 230392 403256 230404
rect 403308 230392 403314 230444
rect 408770 230392 408776 230444
rect 408828 230432 408834 230444
rect 416038 230432 416044 230444
rect 408828 230404 416044 230432
rect 408828 230392 408834 230404
rect 416038 230392 416044 230404
rect 416096 230392 416102 230444
rect 421282 230392 421288 230444
rect 421340 230432 421346 230444
rect 422202 230432 422208 230444
rect 421340 230404 422208 230432
rect 421340 230392 421346 230404
rect 422202 230392 422208 230404
rect 422260 230392 422266 230444
rect 422386 230392 422392 230444
rect 422444 230432 422450 230444
rect 437584 230432 437612 230540
rect 438026 230528 438032 230540
rect 438084 230528 438090 230580
rect 472618 230528 472624 230580
rect 472676 230568 472682 230580
rect 472676 230540 480254 230568
rect 472676 230528 472682 230540
rect 480226 230500 480254 230540
rect 544378 230500 544384 230512
rect 480226 230472 544384 230500
rect 544378 230460 544384 230472
rect 544436 230460 544442 230512
rect 442258 230432 442264 230444
rect 422444 230404 437612 230432
rect 437676 230404 442264 230432
rect 422444 230392 422450 230404
rect 403618 230324 403624 230376
rect 403676 230364 403682 230376
rect 404998 230364 405004 230376
rect 403676 230336 405004 230364
rect 403676 230324 403682 230336
rect 404998 230324 405004 230336
rect 405056 230324 405062 230376
rect 406378 230324 406384 230376
rect 406436 230364 406442 230376
rect 408402 230364 408408 230376
rect 406436 230336 408408 230364
rect 406436 230324 406442 230336
rect 408402 230324 408408 230336
rect 408460 230324 408466 230376
rect 414106 230256 414112 230308
rect 414164 230296 414170 230308
rect 427722 230296 427728 230308
rect 414164 230268 427728 230296
rect 414164 230256 414170 230268
rect 427722 230256 427728 230268
rect 427780 230256 427786 230308
rect 429562 230256 429568 230308
rect 429620 230296 429626 230308
rect 432138 230296 432144 230308
rect 429620 230268 432144 230296
rect 429620 230256 429626 230268
rect 432138 230256 432144 230268
rect 432196 230256 432202 230308
rect 432322 230256 432328 230308
rect 432380 230296 432386 230308
rect 437676 230296 437704 230404
rect 442258 230392 442264 230404
rect 442316 230392 442322 230444
rect 443914 230392 443920 230444
rect 443972 230432 443978 230444
rect 445938 230432 445944 230444
rect 443972 230404 445944 230432
rect 443972 230392 443978 230404
rect 445938 230392 445944 230404
rect 445996 230392 446002 230444
rect 447226 230392 447232 230444
rect 447284 230432 447290 230444
rect 448054 230432 448060 230444
rect 447284 230404 448060 230432
rect 447284 230392 447290 230404
rect 448054 230392 448060 230404
rect 448112 230392 448118 230444
rect 453298 230392 453304 230444
rect 453356 230432 453362 230444
rect 454494 230432 454500 230444
rect 453356 230404 454500 230432
rect 453356 230392 453362 230404
rect 454494 230392 454500 230404
rect 454552 230392 454558 230444
rect 456610 230392 456616 230444
rect 456668 230432 456674 230444
rect 465810 230432 465816 230444
rect 456668 230404 465816 230432
rect 456668 230392 456674 230404
rect 465810 230392 465816 230404
rect 465868 230392 465874 230444
rect 466546 230392 466552 230444
rect 466604 230432 466610 230444
rect 467742 230432 467748 230444
rect 466604 230404 467748 230432
rect 466604 230392 466610 230404
rect 467742 230392 467748 230404
rect 467800 230392 467806 230444
rect 476482 230392 476488 230444
rect 476540 230432 476546 230444
rect 477402 230432 477408 230444
rect 476540 230404 477408 230432
rect 476540 230392 476546 230404
rect 477402 230392 477408 230404
rect 477460 230392 477466 230444
rect 478046 230392 478052 230444
rect 478104 230432 478110 230444
rect 480070 230432 480076 230444
rect 478104 230404 480076 230432
rect 478104 230392 478110 230404
rect 480070 230392 480076 230404
rect 480128 230392 480134 230444
rect 480898 230324 480904 230376
rect 480956 230364 480962 230376
rect 483290 230364 483296 230376
rect 480956 230336 483296 230364
rect 480956 230324 480962 230336
rect 483290 230324 483296 230336
rect 483348 230324 483354 230376
rect 432380 230268 437704 230296
rect 432380 230256 432386 230268
rect 437842 230256 437848 230308
rect 437900 230296 437906 230308
rect 480530 230296 480536 230308
rect 437900 230268 480536 230296
rect 437900 230256 437906 230268
rect 480530 230256 480536 230268
rect 480588 230256 480594 230308
rect 483750 230256 483756 230308
rect 483808 230296 483814 230308
rect 488074 230296 488080 230308
rect 483808 230268 488080 230296
rect 483808 230256 483814 230268
rect 488074 230256 488080 230268
rect 488132 230256 488138 230308
rect 542446 230296 542452 230308
rect 488276 230268 542452 230296
rect 398742 230120 398748 230172
rect 398800 230160 398806 230172
rect 413186 230160 413192 230172
rect 398800 230132 413192 230160
rect 398800 230120 398806 230132
rect 413186 230120 413192 230132
rect 413244 230120 413250 230172
rect 420730 230120 420736 230172
rect 420788 230160 420794 230172
rect 451458 230160 451464 230172
rect 420788 230132 451464 230160
rect 420788 230120 420794 230132
rect 451458 230120 451464 230132
rect 451516 230120 451522 230172
rect 454954 230120 454960 230172
rect 455012 230160 455018 230172
rect 459554 230160 459560 230172
rect 455012 230132 459560 230160
rect 455012 230120 455018 230132
rect 459554 230120 459560 230132
rect 459612 230120 459618 230172
rect 463234 230120 463240 230172
rect 463292 230160 463298 230172
rect 463292 230132 482416 230160
rect 463292 230120 463298 230132
rect 399202 229984 399208 230036
rect 399260 230024 399266 230036
rect 406654 230024 406660 230036
rect 399260 229996 406660 230024
rect 399260 229984 399266 229996
rect 406654 229984 406660 229996
rect 406712 229984 406718 230036
rect 409782 229984 409788 230036
rect 409840 230024 409846 230036
rect 427538 230024 427544 230036
rect 409840 229996 427544 230024
rect 409840 229984 409846 229996
rect 427538 229984 427544 229996
rect 427596 229984 427602 230036
rect 431862 229984 431868 230036
rect 431920 230024 431926 230036
rect 481818 230024 481824 230036
rect 431920 229996 481824 230024
rect 431920 229984 431926 229996
rect 481818 229984 481824 229996
rect 481876 229984 481882 230036
rect 482388 230024 482416 230132
rect 482554 230120 482560 230172
rect 482612 230160 482618 230172
rect 488276 230160 488304 230268
rect 542446 230256 542452 230268
rect 542504 230256 542510 230308
rect 482612 230132 488304 230160
rect 482612 230120 482618 230132
rect 488442 230120 488448 230172
rect 488500 230160 488506 230172
rect 542078 230160 542084 230172
rect 488500 230132 542084 230160
rect 488500 230120 488506 230132
rect 542078 230120 542084 230132
rect 542136 230120 542142 230172
rect 483290 230024 483296 230036
rect 482388 229996 483296 230024
rect 483290 229984 483296 229996
rect 483348 229984 483354 230036
rect 484210 229984 484216 230036
rect 484268 230024 484274 230036
rect 549898 230024 549904 230036
rect 484268 229996 549904 230024
rect 484268 229984 484274 229996
rect 549898 229984 549904 229996
rect 549956 229984 549962 230036
rect 395212 229860 398604 229888
rect 395212 229848 395218 229860
rect 400858 229848 400864 229900
rect 400916 229888 400922 229900
rect 400916 229860 412634 229888
rect 400916 229848 400922 229860
rect 336274 229780 336280 229832
rect 336332 229820 336338 229832
rect 339770 229820 339776 229832
rect 336332 229792 339776 229820
rect 336332 229780 336338 229792
rect 339770 229780 339776 229792
rect 339828 229780 339834 229832
rect 392210 229780 392216 229832
rect 392268 229820 392274 229832
rect 394694 229820 394700 229832
rect 392268 229792 394700 229820
rect 392268 229780 392274 229792
rect 394694 229780 394700 229792
rect 394752 229780 394758 229832
rect 213362 229752 213368 229764
rect 159928 229724 213368 229752
rect 213362 229712 213368 229724
rect 213420 229712 213426 229764
rect 213546 229712 213552 229764
rect 213604 229752 213610 229764
rect 253474 229752 253480 229764
rect 213604 229724 253480 229752
rect 213604 229712 213610 229724
rect 253474 229712 253480 229724
rect 253532 229712 253538 229764
rect 259086 229712 259092 229764
rect 259144 229752 259150 229764
rect 284386 229752 284392 229764
rect 259144 229724 284392 229752
rect 259144 229712 259150 229724
rect 284386 229712 284392 229724
rect 284444 229712 284450 229764
rect 293862 229712 293868 229764
rect 293920 229752 293926 229764
rect 304258 229752 304264 229764
rect 293920 229724 304264 229752
rect 293920 229712 293926 229724
rect 304258 229712 304264 229724
rect 304316 229712 304322 229764
rect 340506 229712 340512 229764
rect 340564 229752 340570 229764
rect 343910 229752 343916 229764
rect 340564 229724 343916 229752
rect 340564 229712 340570 229724
rect 343910 229712 343916 229724
rect 343968 229712 343974 229764
rect 361666 229712 361672 229764
rect 361724 229752 361730 229764
rect 369578 229752 369584 229764
rect 361724 229724 369584 229752
rect 361724 229712 361730 229724
rect 369578 229712 369584 229724
rect 369636 229712 369642 229764
rect 377122 229712 377128 229764
rect 377180 229752 377186 229764
rect 377180 229724 391980 229752
rect 377180 229712 377186 229724
rect 321830 229644 321836 229696
rect 321888 229684 321894 229696
rect 323578 229684 323584 229696
rect 321888 229656 323584 229684
rect 321888 229644 321894 229656
rect 323578 229644 323584 229656
rect 323636 229644 323642 229696
rect 391952 229684 391980 229724
rect 396442 229712 396448 229764
rect 396500 229752 396506 229764
rect 401686 229752 401692 229764
rect 396500 229724 401692 229752
rect 396500 229712 396506 229724
rect 401686 229712 401692 229724
rect 401744 229712 401750 229764
rect 405826 229712 405832 229764
rect 405884 229752 405890 229764
rect 409782 229752 409788 229764
rect 405884 229724 409788 229752
rect 405884 229712 405890 229724
rect 409782 229712 409788 229724
rect 409840 229712 409846 229764
rect 412606 229752 412634 229860
rect 417234 229848 417240 229900
rect 417292 229888 417298 229900
rect 424226 229888 424232 229900
rect 417292 229860 424232 229888
rect 417292 229848 417298 229860
rect 424226 229848 424232 229860
rect 424284 229848 424290 229900
rect 427354 229848 427360 229900
rect 427412 229888 427418 229900
rect 432598 229888 432604 229900
rect 427412 229860 432604 229888
rect 427412 229848 427418 229860
rect 432598 229848 432604 229860
rect 432656 229848 432662 229900
rect 432874 229848 432880 229900
rect 432932 229888 432938 229900
rect 437842 229888 437848 229900
rect 432932 229860 437848 229888
rect 432932 229848 432938 229860
rect 437842 229848 437848 229860
rect 437900 229848 437906 229900
rect 438026 229848 438032 229900
rect 438084 229888 438090 229900
rect 441890 229888 441896 229900
rect 438084 229860 441896 229888
rect 438084 229848 438090 229860
rect 441890 229848 441896 229860
rect 441948 229848 441954 229900
rect 442258 229848 442264 229900
rect 442316 229888 442322 229900
rect 484854 229888 484860 229900
rect 442316 229860 484860 229888
rect 442316 229848 442322 229860
rect 484854 229848 484860 229860
rect 484912 229848 484918 229900
rect 485866 229848 485872 229900
rect 485924 229888 485930 229900
rect 558178 229888 558184 229900
rect 485924 229860 558184 229888
rect 485924 229848 485930 229860
rect 558178 229848 558184 229860
rect 558236 229848 558242 229900
rect 420914 229752 420920 229764
rect 412606 229724 420920 229752
rect 420914 229712 420920 229724
rect 420972 229712 420978 229764
rect 425514 229752 425520 229764
rect 421116 229724 425520 229752
rect 395154 229684 395160 229696
rect 391952 229656 395160 229684
rect 395154 229644 395160 229656
rect 395212 229644 395218 229696
rect 117222 229576 117228 229628
rect 117280 229616 117286 229628
rect 181438 229616 181444 229628
rect 117280 229588 181444 229616
rect 117280 229576 117286 229588
rect 181438 229576 181444 229588
rect 181496 229576 181502 229628
rect 182082 229576 182088 229628
rect 182140 229616 182146 229628
rect 182140 229588 191420 229616
rect 182140 229576 182146 229588
rect 126882 229440 126888 229492
rect 126940 229480 126946 229492
rect 190914 229480 190920 229492
rect 126940 229452 190920 229480
rect 126940 229440 126946 229452
rect 190914 229440 190920 229452
rect 190972 229440 190978 229492
rect 191392 229480 191420 229588
rect 191558 229576 191564 229628
rect 191616 229616 191622 229628
rect 192754 229616 192760 229628
rect 191616 229588 192760 229616
rect 191616 229576 191622 229588
rect 192754 229576 192760 229588
rect 192812 229576 192818 229628
rect 194226 229576 194232 229628
rect 194284 229616 194290 229628
rect 194284 229588 195468 229616
rect 194284 229576 194290 229588
rect 195238 229480 195244 229492
rect 191392 229452 195244 229480
rect 195238 229440 195244 229452
rect 195296 229440 195302 229492
rect 195440 229480 195468 229588
rect 195882 229576 195888 229628
rect 195940 229616 195946 229628
rect 202782 229616 202788 229628
rect 195940 229588 202788 229616
rect 195940 229576 195946 229588
rect 202782 229576 202788 229588
rect 202840 229576 202846 229628
rect 205082 229616 205088 229628
rect 203352 229588 205088 229616
rect 203352 229480 203380 229588
rect 205082 229576 205088 229588
rect 205140 229576 205146 229628
rect 205450 229576 205456 229628
rect 205508 229616 205514 229628
rect 209314 229616 209320 229628
rect 205508 229588 209320 229616
rect 205508 229576 205514 229588
rect 209314 229576 209320 229588
rect 209372 229576 209378 229628
rect 211706 229576 211712 229628
rect 211764 229616 211770 229628
rect 249058 229616 249064 229628
rect 211764 229588 249064 229616
rect 211764 229576 211770 229588
rect 249058 229576 249064 229588
rect 249116 229576 249122 229628
rect 342346 229576 342352 229628
rect 342404 229616 342410 229628
rect 343542 229616 343548 229628
rect 342404 229588 343548 229616
rect 342404 229576 342410 229588
rect 343542 229576 343548 229588
rect 343600 229576 343606 229628
rect 349062 229576 349068 229628
rect 349120 229616 349126 229628
rect 353018 229616 353024 229628
rect 349120 229588 353024 229616
rect 349120 229576 349126 229588
rect 353018 229576 353024 229588
rect 353076 229576 353082 229628
rect 356146 229576 356152 229628
rect 356204 229616 356210 229628
rect 363138 229616 363144 229628
rect 356204 229588 363144 229616
rect 356204 229576 356210 229588
rect 363138 229576 363144 229588
rect 363196 229576 363202 229628
rect 387702 229576 387708 229628
rect 387760 229616 387766 229628
rect 391750 229616 391756 229628
rect 387760 229588 391756 229616
rect 387760 229576 387766 229588
rect 391750 229576 391756 229588
rect 391808 229576 391814 229628
rect 404722 229576 404728 229628
rect 404780 229616 404786 229628
rect 408770 229616 408776 229628
rect 404780 229588 408776 229616
rect 404780 229576 404786 229588
rect 408770 229576 408776 229588
rect 408828 229576 408834 229628
rect 416866 229576 416872 229628
rect 416924 229616 416930 229628
rect 421116 229616 421144 229724
rect 425514 229712 425520 229724
rect 425572 229712 425578 229764
rect 429010 229712 429016 229764
rect 429068 229752 429074 229764
rect 430022 229752 430028 229764
rect 429068 229724 430028 229752
rect 429068 229712 429074 229724
rect 430022 229712 430028 229724
rect 430080 229712 430086 229764
rect 430206 229712 430212 229764
rect 430264 229752 430270 229764
rect 433610 229752 433616 229764
rect 430264 229724 433616 229752
rect 430264 229712 430270 229724
rect 433610 229712 433616 229724
rect 433668 229712 433674 229764
rect 433794 229712 433800 229764
rect 433852 229752 433858 229764
rect 436186 229752 436192 229764
rect 433852 229724 436192 229752
rect 433852 229712 433858 229724
rect 436186 229712 436192 229724
rect 436244 229712 436250 229764
rect 438026 229712 438032 229764
rect 438084 229752 438090 229764
rect 487338 229752 487344 229764
rect 438084 229724 487344 229752
rect 438084 229712 438090 229724
rect 487338 229712 487344 229724
rect 487396 229712 487402 229764
rect 487522 229712 487528 229764
rect 487580 229752 487586 229764
rect 565078 229752 565084 229764
rect 487580 229724 565084 229752
rect 487580 229712 487586 229724
rect 565078 229712 565084 229724
rect 565136 229712 565142 229764
rect 416924 229588 421144 229616
rect 416924 229576 416930 229588
rect 421834 229576 421840 229628
rect 421892 229616 421898 229628
rect 438578 229616 438584 229628
rect 421892 229588 438584 229616
rect 421892 229576 421898 229588
rect 438578 229576 438584 229588
rect 438636 229576 438642 229628
rect 438946 229576 438952 229628
rect 439004 229616 439010 229628
rect 439004 229588 441016 229616
rect 439004 229576 439010 229588
rect 287698 229508 287704 229560
rect 287756 229548 287762 229560
rect 291010 229548 291016 229560
rect 287756 229520 291016 229548
rect 287756 229508 287762 229520
rect 291010 229508 291016 229520
rect 291068 229508 291074 229560
rect 343726 229508 343732 229560
rect 343784 229548 343790 229560
rect 345382 229548 345388 229560
rect 343784 229520 345388 229548
rect 343784 229508 343790 229520
rect 345382 229508 345388 229520
rect 345440 229508 345446 229560
rect 394050 229508 394056 229560
rect 394108 229548 394114 229560
rect 399478 229548 399484 229560
rect 394108 229520 399484 229548
rect 394108 229508 394114 229520
rect 399478 229508 399484 229520
rect 399536 229508 399542 229560
rect 195440 229452 203380 229480
rect 203518 229440 203524 229492
rect 203576 229480 203582 229492
rect 222562 229480 222568 229492
rect 203576 229452 222568 229480
rect 203576 229440 203582 229452
rect 222562 229440 222568 229452
rect 222620 229440 222626 229492
rect 227346 229440 227352 229492
rect 227404 229480 227410 229492
rect 262306 229480 262312 229492
rect 227404 229452 262312 229480
rect 227404 229440 227410 229452
rect 262306 229440 262312 229452
rect 262364 229440 262370 229492
rect 317506 229440 317512 229492
rect 317564 229480 317570 229492
rect 319714 229480 319720 229492
rect 317564 229452 319720 229480
rect 317564 229440 317570 229452
rect 319714 229440 319720 229452
rect 319772 229440 319778 229492
rect 384850 229440 384856 229492
rect 384908 229480 384914 229492
rect 388438 229480 388444 229492
rect 384908 229452 388444 229480
rect 384908 229440 384914 229452
rect 388438 229440 388444 229452
rect 388496 229440 388502 229492
rect 392210 229480 392216 229492
rect 391860 229452 392216 229480
rect 343358 229372 343364 229424
rect 343416 229412 343422 229424
rect 346670 229412 346676 229424
rect 343416 229384 346676 229412
rect 343416 229372 343422 229384
rect 346670 229372 346676 229384
rect 346728 229372 346734 229424
rect 378778 229372 378784 229424
rect 378836 229412 378842 229424
rect 383930 229412 383936 229424
rect 378836 229384 383936 229412
rect 378836 229372 378842 229384
rect 383930 229372 383936 229384
rect 383988 229372 383994 229424
rect 133782 229304 133788 229356
rect 133840 229344 133846 229356
rect 200482 229344 200488 229356
rect 133840 229316 200488 229344
rect 133840 229304 133846 229316
rect 200482 229304 200488 229316
rect 200540 229304 200546 229356
rect 202598 229344 202604 229356
rect 200684 229316 202604 229344
rect 140682 229168 140688 229220
rect 140740 229208 140746 229220
rect 200684 229208 200712 229316
rect 202598 229304 202604 229316
rect 202656 229304 202662 229356
rect 202782 229304 202788 229356
rect 202840 229344 202846 229356
rect 205266 229344 205272 229356
rect 202840 229316 205272 229344
rect 202840 229304 202846 229316
rect 205266 229304 205272 229316
rect 205324 229304 205330 229356
rect 205542 229304 205548 229356
rect 205600 229344 205606 229356
rect 214282 229344 214288 229356
rect 205600 229316 214288 229344
rect 205600 229304 205606 229316
rect 214282 229304 214288 229316
rect 214340 229304 214346 229356
rect 214650 229304 214656 229356
rect 214708 229344 214714 229356
rect 218146 229344 218152 229356
rect 214708 229316 218152 229344
rect 214708 229304 214714 229316
rect 218146 229304 218152 229316
rect 218204 229304 218210 229356
rect 220906 229344 220912 229356
rect 219406 229316 220912 229344
rect 140740 229180 200712 229208
rect 140740 229168 140746 229180
rect 200850 229168 200856 229220
rect 200908 229208 200914 229220
rect 206002 229208 206008 229220
rect 200908 229180 206008 229208
rect 200908 229168 200914 229180
rect 206002 229168 206008 229180
rect 206060 229168 206066 229220
rect 211154 229168 211160 229220
rect 211212 229208 211218 229220
rect 219406 229208 219434 229316
rect 220906 229304 220912 229316
rect 220964 229304 220970 229356
rect 222194 229304 222200 229356
rect 222252 229344 222258 229356
rect 227530 229344 227536 229356
rect 222252 229316 227536 229344
rect 222252 229304 222258 229316
rect 227530 229304 227536 229316
rect 227588 229304 227594 229356
rect 229186 229304 229192 229356
rect 229244 229344 229250 229356
rect 250162 229344 250168 229356
rect 229244 229316 250168 229344
rect 229244 229304 229250 229316
rect 250162 229304 250168 229316
rect 250220 229304 250226 229356
rect 320082 229304 320088 229356
rect 320140 229344 320146 229356
rect 321370 229344 321376 229356
rect 320140 229316 321376 229344
rect 320140 229304 320146 229316
rect 321370 229304 321376 229316
rect 321428 229304 321434 229356
rect 385954 229304 385960 229356
rect 386012 229344 386018 229356
rect 391860 229344 391888 229452
rect 392210 229440 392216 229452
rect 392268 229440 392274 229492
rect 403066 229440 403072 229492
rect 403124 229480 403130 229492
rect 417234 229480 417240 229492
rect 403124 229452 417240 229480
rect 403124 229440 403130 229452
rect 417234 229440 417240 229452
rect 417292 229440 417298 229492
rect 419074 229440 419080 229492
rect 419132 229480 419138 229492
rect 429838 229480 429844 229492
rect 419132 229452 429844 229480
rect 419132 229440 419138 229452
rect 429838 229440 429844 229452
rect 429896 229440 429902 229492
rect 430022 229440 430028 229492
rect 430080 229480 430086 229492
rect 432414 229480 432420 229492
rect 430080 229452 432420 229480
rect 430080 229440 430086 229452
rect 432414 229440 432420 229452
rect 432472 229440 432478 229492
rect 440786 229480 440792 229492
rect 432616 229452 440792 229480
rect 386012 229316 391888 229344
rect 386012 229304 386018 229316
rect 392026 229304 392032 229356
rect 392084 229344 392090 229356
rect 394050 229344 394056 229356
rect 392084 229316 394056 229344
rect 392084 229304 392090 229316
rect 394050 229304 394056 229316
rect 394108 229304 394114 229356
rect 413554 229304 413560 229356
rect 413612 229344 413618 229356
rect 418798 229344 418804 229356
rect 413612 229316 418804 229344
rect 413612 229304 413618 229316
rect 418798 229304 418804 229316
rect 418856 229304 418862 229356
rect 426802 229304 426808 229356
rect 426860 229344 426866 229356
rect 432616 229344 432644 229452
rect 440786 229440 440792 229452
rect 440844 229440 440850 229492
rect 440988 229480 441016 229588
rect 441154 229576 441160 229628
rect 441212 229616 441218 229628
rect 490374 229616 490380 229628
rect 441212 229588 490380 229616
rect 441212 229576 441218 229588
rect 490374 229576 490380 229588
rect 490432 229576 490438 229628
rect 490558 229576 490564 229628
rect 490616 229616 490622 229628
rect 510614 229616 510620 229628
rect 490616 229588 510620 229616
rect 490616 229576 490622 229588
rect 510614 229576 510620 229588
rect 510672 229576 510678 229628
rect 494698 229480 494704 229492
rect 440988 229452 494704 229480
rect 494698 229440 494704 229452
rect 494756 229440 494762 229492
rect 433794 229344 433800 229356
rect 426860 229316 432644 229344
rect 433260 229316 433800 229344
rect 426860 229304 426866 229316
rect 250438 229236 250444 229288
rect 250496 229276 250502 229288
rect 255682 229276 255688 229288
rect 250496 229248 255688 229276
rect 250496 229236 250502 229248
rect 255682 229236 255688 229248
rect 255740 229236 255746 229288
rect 334066 229236 334072 229288
rect 334124 229276 334130 229288
rect 335538 229276 335544 229288
rect 334124 229248 335544 229276
rect 334124 229236 334130 229248
rect 335538 229236 335544 229248
rect 335596 229236 335602 229288
rect 350626 229236 350632 229288
rect 350684 229276 350690 229288
rect 355318 229276 355324 229288
rect 350684 229248 355324 229276
rect 350684 229236 350690 229248
rect 355318 229236 355324 229248
rect 355376 229236 355382 229288
rect 367738 229236 367744 229288
rect 367796 229276 367802 229288
rect 422938 229276 422944 229288
rect 367796 229248 374868 229276
rect 367796 229236 367802 229248
rect 211212 229180 219434 229208
rect 211212 229168 211218 229180
rect 220814 229168 220820 229220
rect 220872 229208 220878 229220
rect 225322 229208 225328 229220
rect 220872 229180 225328 229208
rect 220872 229168 220878 229180
rect 225322 229168 225328 229180
rect 225380 229168 225386 229220
rect 233878 229168 233884 229220
rect 233936 229208 233942 229220
rect 243538 229208 243544 229220
rect 233936 229180 243544 229208
rect 233936 229168 233942 229180
rect 243538 229168 243544 229180
rect 243596 229168 243602 229220
rect 229738 229140 229744 229152
rect 227732 229112 229744 229140
rect 109770 229032 109776 229084
rect 109828 229072 109834 229084
rect 176838 229072 176844 229084
rect 109828 229044 176844 229072
rect 109828 229032 109834 229044
rect 176838 229032 176844 229044
rect 176896 229032 176902 229084
rect 222194 229072 222200 229084
rect 181640 229044 222200 229072
rect 181640 229004 181668 229044
rect 222194 229032 222200 229044
rect 222252 229032 222258 229084
rect 227732 229072 227760 229112
rect 229738 229100 229744 229112
rect 229796 229100 229802 229152
rect 321370 229100 321376 229152
rect 321428 229140 321434 229152
rect 325786 229140 325792 229152
rect 321428 229112 325792 229140
rect 321428 229100 321434 229112
rect 325786 229100 325792 229112
rect 325844 229100 325850 229152
rect 373810 229100 373816 229152
rect 373868 229140 373874 229152
rect 374638 229140 374644 229152
rect 373868 229112 374644 229140
rect 373868 229100 373874 229112
rect 374638 229100 374644 229112
rect 374696 229100 374702 229152
rect 223592 229044 227760 229072
rect 181456 228976 181668 229004
rect 99834 228896 99840 228948
rect 99892 228936 99898 228948
rect 99892 228908 171824 228936
rect 99892 228896 99898 228908
rect 96522 228760 96528 228812
rect 96580 228800 96586 228812
rect 171134 228800 171140 228812
rect 96580 228772 171140 228800
rect 96580 228760 96586 228772
rect 171134 228760 171140 228772
rect 171192 228760 171198 228812
rect 171796 228800 171824 228908
rect 176470 228896 176476 228948
rect 176528 228936 176534 228948
rect 181456 228936 181484 228976
rect 223592 228936 223620 229044
rect 233694 229032 233700 229084
rect 233752 229072 233758 229084
rect 261754 229072 261760 229084
rect 233752 229044 261760 229072
rect 233752 229032 233758 229044
rect 261754 229032 261760 229044
rect 261812 229032 261818 229084
rect 374840 229072 374868 229248
rect 422266 229248 422944 229276
rect 389818 229168 389824 229220
rect 389876 229208 389882 229220
rect 392854 229208 392860 229220
rect 389876 229180 392860 229208
rect 389876 229168 389882 229180
rect 392854 229168 392860 229180
rect 392912 229168 392918 229220
rect 410242 229168 410248 229220
rect 410300 229208 410306 229220
rect 412726 229208 412732 229220
rect 410300 229180 412732 229208
rect 410300 229168 410306 229180
rect 412726 229168 412732 229180
rect 412784 229168 412790 229220
rect 418522 229168 418528 229220
rect 418580 229208 418586 229220
rect 422266 229208 422294 229248
rect 422938 229236 422944 229248
rect 422996 229236 423002 229288
rect 418580 229180 422294 229208
rect 418580 229168 418586 229180
rect 424594 229168 424600 229220
rect 424652 229208 424658 229220
rect 430206 229208 430212 229220
rect 424652 229180 430212 229208
rect 424652 229168 424658 229180
rect 430206 229168 430212 229180
rect 430264 229168 430270 229220
rect 430666 229168 430672 229220
rect 430724 229208 430730 229220
rect 431586 229208 431592 229220
rect 430724 229180 431592 229208
rect 430724 229168 430730 229180
rect 431586 229168 431592 229180
rect 431644 229168 431650 229220
rect 432414 229168 432420 229220
rect 432472 229208 432478 229220
rect 433260 229208 433288 229316
rect 433794 229304 433800 229316
rect 433852 229304 433858 229356
rect 434530 229304 434536 229356
rect 434588 229344 434594 229356
rect 438026 229344 438032 229356
rect 434588 229316 438032 229344
rect 434588 229304 434594 229316
rect 438026 229304 438032 229316
rect 438084 229304 438090 229356
rect 438578 229304 438584 229356
rect 438636 229344 438642 229356
rect 439590 229344 439596 229356
rect 438636 229316 439596 229344
rect 438636 229304 438642 229316
rect 439590 229304 439596 229316
rect 439648 229304 439654 229356
rect 440602 229304 440608 229356
rect 440660 229344 440666 229356
rect 441430 229344 441436 229356
rect 440660 229316 441436 229344
rect 440660 229304 440666 229316
rect 441430 229304 441436 229316
rect 441488 229304 441494 229356
rect 444466 229304 444472 229356
rect 444524 229344 444530 229356
rect 445662 229344 445668 229356
rect 444524 229316 445668 229344
rect 444524 229304 444530 229316
rect 445662 229304 445668 229316
rect 445720 229304 445726 229356
rect 488902 229344 488908 229356
rect 447106 229316 488908 229344
rect 432472 229180 433288 229208
rect 432472 229168 432478 229180
rect 433426 229168 433432 229220
rect 433484 229208 433490 229220
rect 434346 229208 434352 229220
rect 433484 229180 434352 229208
rect 433484 229168 433490 229180
rect 434346 229168 434352 229180
rect 434404 229168 434410 229220
rect 435082 229168 435088 229220
rect 435140 229208 435146 229220
rect 436002 229208 436008 229220
rect 435140 229180 436008 229208
rect 435140 229168 435146 229180
rect 436002 229168 436008 229180
rect 436060 229168 436066 229220
rect 436738 229168 436744 229220
rect 436796 229208 436802 229220
rect 447106 229208 447134 229316
rect 488902 229304 488908 229316
rect 488960 229304 488966 229356
rect 490374 229304 490380 229356
rect 490432 229344 490438 229356
rect 497458 229344 497464 229356
rect 490432 229316 497464 229344
rect 490432 229304 490438 229316
rect 497458 229304 497464 229316
rect 497516 229304 497522 229356
rect 436796 229180 447134 229208
rect 436796 229168 436802 229180
rect 465994 229168 466000 229220
rect 466052 229208 466058 229220
rect 474642 229208 474648 229220
rect 466052 229180 474648 229208
rect 466052 229168 466058 229180
rect 474642 229168 474648 229180
rect 474700 229168 474706 229220
rect 474826 229168 474832 229220
rect 474884 229208 474890 229220
rect 477218 229208 477224 229220
rect 474884 229180 477224 229208
rect 474884 229168 474890 229180
rect 477218 229168 477224 229180
rect 477276 229168 477282 229220
rect 479242 229168 479248 229220
rect 479300 229208 479306 229220
rect 522574 229208 522580 229220
rect 479300 229180 522580 229208
rect 479300 229168 479306 229180
rect 522574 229168 522580 229180
rect 522632 229168 522638 229220
rect 382458 229072 382464 229084
rect 374840 229044 382464 229072
rect 382458 229032 382464 229044
rect 382516 229032 382522 229084
rect 384298 229032 384304 229084
rect 384356 229072 384362 229084
rect 410426 229072 410432 229084
rect 384356 229044 410432 229072
rect 384356 229032 384362 229044
rect 410426 229032 410432 229044
rect 410484 229032 410490 229084
rect 442258 229072 442264 229084
rect 422496 229044 442264 229072
rect 419626 228964 419632 229016
rect 419684 229004 419690 229016
rect 422496 229004 422524 229044
rect 442258 229032 442264 229044
rect 442316 229032 442322 229084
rect 451274 229032 451280 229084
rect 451332 229072 451338 229084
rect 453942 229072 453948 229084
rect 451332 229044 453948 229072
rect 451332 229032 451338 229044
rect 453942 229032 453948 229044
rect 454000 229032 454006 229084
rect 458818 229032 458824 229084
rect 458876 229072 458882 229084
rect 524046 229072 524052 229084
rect 458876 229044 524052 229072
rect 458876 229032 458882 229044
rect 524046 229032 524052 229044
rect 524104 229032 524110 229084
rect 419684 228976 422524 229004
rect 419684 228964 419690 228976
rect 176528 228908 181484 228936
rect 181732 228908 223620 228936
rect 176528 228896 176534 228908
rect 181732 228868 181760 228908
rect 229002 228896 229008 228948
rect 229060 228936 229066 228948
rect 262858 228936 262864 228948
rect 229060 228908 262864 228936
rect 229060 228896 229066 228908
rect 262858 228896 262864 228908
rect 262916 228896 262922 228948
rect 275370 228896 275376 228948
rect 275428 228936 275434 228948
rect 293494 228936 293500 228948
rect 275428 228908 293500 228936
rect 275428 228896 275434 228908
rect 293494 228896 293500 228908
rect 293552 228896 293558 228948
rect 390922 228896 390928 228948
rect 390980 228936 390986 228948
rect 419442 228936 419448 228948
rect 390980 228908 419448 228936
rect 390980 228896 390986 228908
rect 419442 228896 419448 228908
rect 419500 228896 419506 228948
rect 424042 228896 424048 228948
rect 424100 228936 424106 228948
rect 457070 228936 457076 228948
rect 424100 228908 457076 228936
rect 424100 228896 424106 228908
rect 457070 228896 457076 228908
rect 457128 228896 457134 228948
rect 458266 228896 458272 228948
rect 458324 228936 458330 228948
rect 523126 228936 523132 228948
rect 458324 228908 523132 228936
rect 458324 228896 458330 228908
rect 523126 228896 523132 228908
rect 523184 228896 523190 228948
rect 181548 228840 181760 228868
rect 176608 228800 176614 228812
rect 171796 228772 176614 228800
rect 176608 228760 176614 228772
rect 176666 228760 176672 228812
rect 179230 228760 179236 228812
rect 179288 228800 179294 228812
rect 181548 228800 181576 228840
rect 179288 228772 181576 228800
rect 179288 228760 179294 228772
rect 182358 228760 182364 228812
rect 182416 228800 182422 228812
rect 220814 228800 220820 228812
rect 182416 228772 220820 228800
rect 182416 228760 182422 228772
rect 220814 228760 220820 228772
rect 220872 228760 220878 228812
rect 222102 228760 222108 228812
rect 222160 228800 222166 228812
rect 258442 228800 258448 228812
rect 222160 228772 258448 228800
rect 222160 228760 222166 228772
rect 258442 228760 258448 228772
rect 258500 228760 258506 228812
rect 265434 228760 265440 228812
rect 265492 228800 265498 228812
rect 287146 228800 287152 228812
rect 265492 228772 287152 228800
rect 265492 228760 265498 228772
rect 287146 228760 287152 228772
rect 287204 228760 287210 228812
rect 291930 228760 291936 228812
rect 291988 228800 291994 228812
rect 304810 228800 304816 228812
rect 291988 228772 304816 228800
rect 291988 228760 291994 228772
rect 304810 228760 304816 228772
rect 304868 228760 304874 228812
rect 360562 228760 360568 228812
rect 360620 228800 360626 228812
rect 375650 228800 375656 228812
rect 360620 228772 375656 228800
rect 360620 228760 360626 228772
rect 375650 228760 375656 228772
rect 375708 228760 375714 228812
rect 382274 228760 382280 228812
rect 382332 228800 382338 228812
rect 390738 228800 390744 228812
rect 382332 228772 390744 228800
rect 382332 228760 382338 228772
rect 390738 228760 390744 228772
rect 390796 228760 390802 228812
rect 401962 228760 401968 228812
rect 402020 228800 402026 228812
rect 434714 228800 434720 228812
rect 402020 228772 434720 228800
rect 402020 228760 402026 228772
rect 434714 228760 434720 228772
rect 434772 228760 434778 228812
rect 442258 228760 442264 228812
rect 442316 228800 442322 228812
rect 451274 228800 451280 228812
rect 442316 228772 451280 228800
rect 442316 228760 442322 228772
rect 451274 228760 451280 228772
rect 451332 228760 451338 228812
rect 451642 228760 451648 228812
rect 451700 228800 451706 228812
rect 456242 228800 456248 228812
rect 451700 228772 456248 228800
rect 451700 228760 451706 228772
rect 456242 228760 456248 228772
rect 456300 228760 456306 228812
rect 464890 228760 464896 228812
rect 464948 228800 464954 228812
rect 532694 228800 532700 228812
rect 464948 228772 532700 228800
rect 464948 228760 464954 228772
rect 532694 228760 532700 228772
rect 532752 228760 532758 228812
rect 93210 228624 93216 228676
rect 93268 228664 93274 228676
rect 150434 228664 150440 228676
rect 93268 228636 150440 228664
rect 93268 228624 93274 228636
rect 150434 228624 150440 228636
rect 150492 228624 150498 228676
rect 150618 228624 150624 228676
rect 150676 228664 150682 228676
rect 178954 228664 178960 228676
rect 150676 228636 178960 228664
rect 150676 228624 150682 228636
rect 178954 228624 178960 228636
rect 179012 228624 179018 228676
rect 182174 228624 182180 228676
rect 182232 228664 182238 228676
rect 233050 228664 233056 228676
rect 182232 228636 233056 228664
rect 182232 228624 182238 228636
rect 233050 228624 233056 228636
rect 233108 228624 233114 228676
rect 245470 228624 245476 228676
rect 245528 228664 245534 228676
rect 273898 228664 273904 228676
rect 245528 228636 273904 228664
rect 245528 228624 245534 228636
rect 273898 228624 273904 228636
rect 273956 228624 273962 228676
rect 276290 228624 276296 228676
rect 276348 228664 276354 228676
rect 294874 228664 294880 228676
rect 276348 228636 294880 228664
rect 276348 228624 276354 228636
rect 294874 228624 294880 228636
rect 294932 228624 294938 228676
rect 295242 228624 295248 228676
rect 295300 228664 295306 228676
rect 307018 228664 307024 228676
rect 295300 228636 307024 228664
rect 295300 228624 295306 228636
rect 307018 228624 307024 228636
rect 307076 228624 307082 228676
rect 360010 228624 360016 228676
rect 360068 228664 360074 228676
rect 374178 228664 374184 228676
rect 360068 228636 374184 228664
rect 360068 228624 360074 228636
rect 374178 228624 374184 228636
rect 374236 228624 374242 228676
rect 377674 228624 377680 228676
rect 377732 228664 377738 228676
rect 400490 228664 400496 228676
rect 377732 228636 400496 228664
rect 377732 228624 377738 228636
rect 400490 228624 400496 228636
rect 400548 228624 400554 228676
rect 404170 228624 404176 228676
rect 404228 228664 404234 228676
rect 440418 228664 440424 228676
rect 404228 228636 440424 228664
rect 404228 228624 404234 228636
rect 440418 228624 440424 228636
rect 440476 228624 440482 228676
rect 441890 228624 441896 228676
rect 441948 228664 441954 228676
rect 468386 228664 468392 228676
rect 441948 228636 468392 228664
rect 441948 228624 441954 228636
rect 468386 228624 468392 228636
rect 468444 228624 468450 228676
rect 471882 228624 471888 228676
rect 471940 228664 471946 228676
rect 471940 228636 540560 228664
rect 471940 228624 471946 228636
rect 75822 228488 75828 228540
rect 75880 228528 75886 228540
rect 162394 228528 162400 228540
rect 75880 228500 162400 228528
rect 75880 228488 75886 228500
rect 162394 228488 162400 228500
rect 162452 228488 162458 228540
rect 166258 228488 166264 228540
rect 166316 228528 166322 228540
rect 211154 228528 211160 228540
rect 166316 228500 211160 228528
rect 166316 228488 166322 228500
rect 211154 228488 211160 228500
rect 211212 228488 211218 228540
rect 212258 228488 212264 228540
rect 212316 228528 212322 228540
rect 251818 228528 251824 228540
rect 212316 228500 251824 228528
rect 212316 228488 212322 228500
rect 251818 228488 251824 228500
rect 251876 228488 251882 228540
rect 253750 228488 253756 228540
rect 253808 228528 253814 228540
rect 278866 228528 278872 228540
rect 253808 228500 278872 228528
rect 253808 228488 253814 228500
rect 278866 228488 278872 228500
rect 278924 228488 278930 228540
rect 286962 228488 286968 228540
rect 287020 228528 287026 228540
rect 300946 228528 300952 228540
rect 287020 228500 300952 228528
rect 287020 228488 287026 228500
rect 300946 228488 300952 228500
rect 301004 228488 301010 228540
rect 347314 228488 347320 228540
rect 347372 228528 347378 228540
rect 356146 228528 356152 228540
rect 347372 228500 356152 228528
rect 347372 228488 347378 228500
rect 356146 228488 356152 228500
rect 356204 228488 356210 228540
rect 369946 228488 369952 228540
rect 370004 228528 370010 228540
rect 386598 228528 386604 228540
rect 370004 228500 386604 228528
rect 370004 228488 370010 228500
rect 386598 228488 386604 228500
rect 386656 228488 386662 228540
rect 393222 228488 393228 228540
rect 393280 228528 393286 228540
rect 423950 228528 423956 228540
rect 393280 228500 423956 228528
rect 393280 228488 393286 228500
rect 423950 228488 423956 228500
rect 424008 228488 424014 228540
rect 432598 228488 432604 228540
rect 432656 228528 432662 228540
rect 472802 228528 472808 228540
rect 432656 228500 472808 228528
rect 432656 228488 432662 228500
rect 472802 228488 472808 228500
rect 472860 228488 472866 228540
rect 473722 228488 473728 228540
rect 473780 228528 473786 228540
rect 540330 228528 540336 228540
rect 473780 228500 540336 228528
rect 473780 228488 473786 228500
rect 540330 228488 540336 228500
rect 540388 228488 540394 228540
rect 540532 228528 540560 228636
rect 542446 228624 542452 228676
rect 542504 228664 542510 228676
rect 559466 228664 559472 228676
rect 542504 228636 559472 228664
rect 542504 228624 542510 228636
rect 559466 228624 559472 228636
rect 559524 228624 559530 228676
rect 542814 228528 542820 228540
rect 540532 228500 542820 228528
rect 542814 228488 542820 228500
rect 542872 228488 542878 228540
rect 68922 228352 68928 228404
rect 68980 228392 68986 228404
rect 157978 228392 157984 228404
rect 68980 228364 157984 228392
rect 68980 228352 68986 228364
rect 157978 228352 157984 228364
rect 158036 228352 158042 228404
rect 159726 228352 159732 228404
rect 159784 228392 159790 228404
rect 214466 228392 214472 228404
rect 159784 228364 214472 228392
rect 159784 228352 159790 228364
rect 214466 228352 214472 228364
rect 214524 228352 214530 228404
rect 214926 228352 214932 228404
rect 214984 228392 214990 228404
rect 255130 228392 255136 228404
rect 214984 228364 255136 228392
rect 214984 228352 214990 228364
rect 255130 228352 255136 228364
rect 255188 228352 255194 228404
rect 256510 228352 256516 228404
rect 256568 228392 256574 228404
rect 281626 228392 281632 228404
rect 256568 228364 281632 228392
rect 256568 228352 256574 228364
rect 281626 228352 281632 228364
rect 281684 228352 281690 228404
rect 281994 228352 282000 228404
rect 282052 228392 282058 228404
rect 298186 228392 298192 228404
rect 282052 228364 298192 228392
rect 282052 228352 282058 228364
rect 298186 228352 298192 228364
rect 298244 228352 298250 228404
rect 304350 228352 304356 228404
rect 304408 228392 304414 228404
rect 314746 228392 314752 228404
rect 304408 228364 314752 228392
rect 304408 228352 304414 228364
rect 314746 228352 314752 228364
rect 314804 228352 314810 228404
rect 351178 228352 351184 228404
rect 351236 228392 351242 228404
rect 360746 228392 360752 228404
rect 351236 228364 360752 228392
rect 351236 228352 351242 228364
rect 360746 228352 360752 228364
rect 360804 228352 360810 228404
rect 363966 228352 363972 228404
rect 364024 228392 364030 228404
rect 373074 228392 373080 228404
rect 364024 228364 373080 228392
rect 364024 228352 364030 228364
rect 373074 228352 373080 228364
rect 373132 228352 373138 228404
rect 373258 228352 373264 228404
rect 373316 228392 373322 228404
rect 393314 228392 393320 228404
rect 373316 228364 393320 228392
rect 373316 228352 373322 228364
rect 393314 228352 393320 228364
rect 393372 228352 393378 228404
rect 397546 228352 397552 228404
rect 397604 228392 397610 228404
rect 430574 228392 430580 228404
rect 397604 228364 430580 228392
rect 397604 228352 397610 228364
rect 430574 228352 430580 228364
rect 430632 228352 430638 228404
rect 433610 228352 433616 228404
rect 433668 228392 433674 228404
rect 433668 228364 463740 228392
rect 433668 228352 433674 228364
rect 118786 228216 118792 228268
rect 118844 228256 118850 228268
rect 150618 228256 150624 228268
rect 118844 228228 150624 228256
rect 118844 228216 118850 228228
rect 150618 228216 150624 228228
rect 150676 228216 150682 228268
rect 150802 228216 150808 228268
rect 150860 228256 150866 228268
rect 195882 228256 195888 228268
rect 150860 228228 195888 228256
rect 150860 228216 150866 228228
rect 195882 228216 195888 228228
rect 195940 228216 195946 228268
rect 249334 228256 249340 228268
rect 219406 228228 249340 228256
rect 149514 228080 149520 228132
rect 149572 228120 149578 228132
rect 209682 228120 209688 228132
rect 149572 228092 209688 228120
rect 149572 228080 149578 228092
rect 209682 228080 209688 228092
rect 209740 228080 209746 228132
rect 65978 227944 65984 227996
rect 66036 227984 66042 227996
rect 155770 227984 155776 227996
rect 66036 227956 155776 227984
rect 66036 227944 66042 227956
rect 155770 227944 155776 227956
rect 155828 227944 155834 227996
rect 155954 227944 155960 227996
rect 156012 227984 156018 227996
rect 205542 227984 205548 227996
rect 156012 227956 205548 227984
rect 156012 227944 156018 227956
rect 205542 227944 205548 227956
rect 205600 227944 205606 227996
rect 208946 227944 208952 227996
rect 209004 227984 209010 227996
rect 219406 227984 219434 228228
rect 249334 228216 249340 228228
rect 249392 228216 249398 228268
rect 276106 228256 276112 228268
rect 258046 228228 276112 228256
rect 226610 228080 226616 228132
rect 226668 228120 226674 228132
rect 233694 228120 233700 228132
rect 226668 228092 233700 228120
rect 226668 228080 226674 228092
rect 233694 228080 233700 228092
rect 233752 228080 233758 228132
rect 248874 228080 248880 228132
rect 248932 228120 248938 228132
rect 258046 228120 258074 228228
rect 276106 228216 276112 228228
rect 276164 228216 276170 228268
rect 428458 228216 428464 228268
rect 428516 228256 428522 228268
rect 455690 228256 455696 228268
rect 428516 228228 455696 228256
rect 428516 228216 428522 228228
rect 455690 228216 455696 228228
rect 455748 228216 455754 228268
rect 463326 228256 463332 228268
rect 456076 228228 463332 228256
rect 248932 228092 258074 228120
rect 248932 228080 248938 228092
rect 440786 228080 440792 228132
rect 440844 228120 440850 228132
rect 456076 228120 456104 228228
rect 463326 228216 463332 228228
rect 463384 228216 463390 228268
rect 463712 228256 463740 228364
rect 463878 228352 463884 228404
rect 463936 228392 463942 228404
rect 474918 228392 474924 228404
rect 463936 228364 474924 228392
rect 463936 228352 463942 228364
rect 474918 228352 474924 228364
rect 474976 228352 474982 228404
rect 477586 228352 477592 228404
rect 477644 228392 477650 228404
rect 552290 228392 552296 228404
rect 477644 228364 552296 228392
rect 477644 228352 477650 228364
rect 552290 228352 552296 228364
rect 552348 228352 552354 228404
rect 471974 228256 471980 228268
rect 463712 228228 471980 228256
rect 471974 228216 471980 228228
rect 472032 228216 472038 228268
rect 474642 228216 474648 228268
rect 474700 228256 474706 228268
rect 534718 228256 534724 228268
rect 474700 228228 534724 228256
rect 474700 228216 474706 228228
rect 534718 228216 534724 228228
rect 534776 228216 534782 228268
rect 540330 228216 540336 228268
rect 540388 228256 540394 228268
rect 546494 228256 546500 228268
rect 540388 228228 546500 228256
rect 540388 228216 540394 228228
rect 546494 228216 546500 228228
rect 546552 228216 546558 228268
rect 440844 228092 456104 228120
rect 440844 228080 440850 228092
rect 456242 228080 456248 228132
rect 456300 228120 456306 228132
rect 513190 228120 513196 228132
rect 456300 228092 513196 228120
rect 456300 228080 456306 228092
rect 513190 228080 513196 228092
rect 513248 228080 513254 228132
rect 209004 227956 219434 227984
rect 209004 227944 209010 227956
rect 356330 227944 356336 227996
rect 356388 227984 356394 227996
rect 359090 227984 359096 227996
rect 356388 227956 359096 227984
rect 356388 227944 356394 227956
rect 359090 227944 359096 227956
rect 359148 227944 359154 227996
rect 454494 227944 454500 227996
rect 454552 227984 454558 227996
rect 514754 227984 514760 227996
rect 454552 227956 514760 227984
rect 454552 227944 454558 227956
rect 514754 227944 514760 227956
rect 514812 227944 514818 227996
rect 127066 227808 127072 227860
rect 127124 227848 127130 227860
rect 181714 227848 181720 227860
rect 127124 227820 181720 227848
rect 127124 227808 127130 227820
rect 181714 227808 181720 227820
rect 181772 227808 181778 227860
rect 204530 227808 204536 227860
rect 204588 227848 204594 227860
rect 211522 227848 211528 227860
rect 204588 227820 211528 227848
rect 204588 227808 204594 227820
rect 211522 227808 211528 227820
rect 211580 227808 211586 227860
rect 455690 227808 455696 227860
rect 455748 227848 455754 227860
rect 455748 227820 459416 227848
rect 455748 227808 455754 227820
rect 262122 227740 262128 227792
rect 262180 227780 262186 227792
rect 268930 227780 268936 227792
rect 262180 227752 268936 227780
rect 262180 227740 262186 227752
rect 268930 227740 268936 227752
rect 268988 227740 268994 227792
rect 308490 227740 308496 227792
rect 308548 227780 308554 227792
rect 315850 227780 315856 227792
rect 308548 227752 315856 227780
rect 308548 227740 308554 227752
rect 315850 227740 315856 227752
rect 315908 227740 315914 227792
rect 316954 227780 316960 227792
rect 316006 227752 316960 227780
rect 42518 227672 42524 227724
rect 42576 227712 42582 227724
rect 47210 227712 47216 227724
rect 42576 227684 47216 227712
rect 42576 227672 42582 227684
rect 47210 227672 47216 227684
rect 47268 227672 47274 227724
rect 118602 227672 118608 227724
rect 118660 227712 118666 227724
rect 118660 227684 127480 227712
rect 118660 227672 118666 227684
rect 127452 227644 127480 227684
rect 127802 227672 127808 227724
rect 127860 227712 127866 227724
rect 137094 227712 137100 227724
rect 127860 227684 137100 227712
rect 127860 227672 127866 227684
rect 137094 227672 137100 227684
rect 137152 227672 137158 227724
rect 137278 227672 137284 227724
rect 137336 227712 137342 227724
rect 197722 227712 197728 227724
rect 137336 227684 197728 227712
rect 137336 227672 137342 227684
rect 197722 227672 197728 227684
rect 197780 227672 197786 227724
rect 199378 227672 199384 227724
rect 199436 227712 199442 227724
rect 242986 227712 242992 227724
rect 199436 227684 242992 227712
rect 199436 227672 199442 227684
rect 242986 227672 242992 227684
rect 243044 227672 243050 227724
rect 272518 227672 272524 227724
rect 272576 227712 272582 227724
rect 285490 227712 285496 227724
rect 272576 227684 285496 227712
rect 272576 227672 272582 227684
rect 285490 227672 285496 227684
rect 285548 227672 285554 227724
rect 127452 227616 127664 227644
rect 127250 227576 127256 227588
rect 103486 227548 127256 227576
rect 97350 227400 97356 227452
rect 97408 227440 97414 227452
rect 103486 227440 103514 227548
rect 127250 227536 127256 227548
rect 127308 227536 127314 227588
rect 127636 227576 127664 227616
rect 315850 227604 315856 227656
rect 315908 227644 315914 227656
rect 316006 227644 316034 227752
rect 316954 227740 316960 227752
rect 317012 227740 317018 227792
rect 317322 227740 317328 227792
rect 317380 227780 317386 227792
rect 321830 227780 321836 227792
rect 317380 227752 321836 227780
rect 317380 227740 317386 227752
rect 321830 227740 321836 227752
rect 321888 227740 321894 227792
rect 408402 227672 408408 227724
rect 408460 227712 408466 227724
rect 443546 227712 443552 227724
rect 408460 227684 443552 227712
rect 408460 227672 408466 227684
rect 443546 227672 443552 227684
rect 443604 227672 443610 227724
rect 459388 227712 459416 227820
rect 459554 227808 459560 227860
rect 459612 227848 459618 227860
rect 518066 227848 518072 227860
rect 459612 227820 518072 227848
rect 459612 227808 459618 227820
rect 518066 227808 518072 227820
rect 518124 227808 518130 227860
rect 459738 227712 459744 227724
rect 459388 227684 459744 227712
rect 459738 227672 459744 227684
rect 459796 227672 459802 227724
rect 461026 227672 461032 227724
rect 461084 227712 461090 227724
rect 527818 227712 527824 227724
rect 461084 227684 527824 227712
rect 461084 227672 461090 227684
rect 527818 227672 527824 227684
rect 527876 227672 527882 227724
rect 315908 227616 316034 227644
rect 315908 227604 315914 227616
rect 191098 227576 191104 227588
rect 127636 227548 191104 227576
rect 191098 227536 191104 227548
rect 191156 227536 191162 227588
rect 192662 227536 192668 227588
rect 192720 227576 192726 227588
rect 235994 227576 236000 227588
rect 192720 227548 236000 227576
rect 192720 227536 192726 227548
rect 235994 227536 236000 227548
rect 236052 227536 236058 227588
rect 249702 227536 249708 227588
rect 249760 227576 249766 227588
rect 277210 227576 277216 227588
rect 249760 227548 277216 227576
rect 249760 227536 249766 227548
rect 277210 227536 277216 227548
rect 277268 227536 277274 227588
rect 383930 227536 383936 227588
rect 383988 227576 383994 227588
rect 398834 227576 398840 227588
rect 383988 227548 398840 227576
rect 383988 227536 383994 227548
rect 398834 227536 398840 227548
rect 398892 227536 398898 227588
rect 415210 227536 415216 227588
rect 415268 227576 415274 227588
rect 452562 227576 452568 227588
rect 415268 227548 452568 227576
rect 415268 227536 415274 227548
rect 452562 227536 452568 227548
rect 452620 227536 452626 227588
rect 468202 227536 468208 227588
rect 468260 227576 468266 227588
rect 538214 227576 538220 227588
rect 468260 227548 538220 227576
rect 468260 227536 468266 227548
rect 538214 227536 538220 227548
rect 538272 227536 538278 227588
rect 97408 227412 103514 227440
rect 97408 227400 97414 227412
rect 115658 227400 115664 227452
rect 115716 227440 115722 227452
rect 188890 227440 188896 227452
rect 115716 227412 188896 227440
rect 115716 227400 115722 227412
rect 188890 227400 188896 227412
rect 188948 227400 188954 227452
rect 189074 227400 189080 227452
rect 189132 227440 189138 227452
rect 236362 227440 236368 227452
rect 189132 227412 236368 227440
rect 189132 227400 189138 227412
rect 236362 227400 236368 227412
rect 236420 227400 236426 227452
rect 242250 227400 242256 227452
rect 242308 227440 242314 227452
rect 271690 227440 271696 227452
rect 242308 227412 271696 227440
rect 242308 227400 242314 227412
rect 271690 227400 271696 227412
rect 271748 227400 271754 227452
rect 372154 227400 372160 227452
rect 372212 227440 372218 227452
rect 389726 227440 389732 227452
rect 372212 227412 389732 227440
rect 372212 227400 372218 227412
rect 389726 227400 389732 227412
rect 389784 227400 389790 227452
rect 395338 227400 395344 227452
rect 395396 227440 395402 227452
rect 426434 227440 426440 227452
rect 395396 227412 426440 227440
rect 395396 227400 395402 227412
rect 426434 227400 426440 227412
rect 426492 227400 426498 227452
rect 432138 227400 432144 227452
rect 432196 227440 432202 227452
rect 476206 227440 476212 227452
rect 432196 227412 476212 227440
rect 432196 227400 432202 227412
rect 476206 227400 476212 227412
rect 476264 227400 476270 227452
rect 477218 227400 477224 227452
rect 477276 227440 477282 227452
rect 547966 227440 547972 227452
rect 477276 227412 547972 227440
rect 477276 227400 477282 227412
rect 547966 227400 547972 227412
rect 548024 227400 548030 227452
rect 82538 227264 82544 227316
rect 82596 227304 82602 227316
rect 157426 227304 157432 227316
rect 82596 227276 157432 227304
rect 82596 227264 82602 227276
rect 157426 227264 157432 227276
rect 157484 227264 157490 227316
rect 175826 227304 175832 227316
rect 164206 227276 175832 227304
rect 157702 227196 157708 227248
rect 157760 227236 157766 227248
rect 164206 227236 164234 227276
rect 175826 227264 175832 227276
rect 175884 227264 175890 227316
rect 179046 227264 179052 227316
rect 179104 227304 179110 227316
rect 192110 227304 192116 227316
rect 179104 227276 192116 227304
rect 179104 227264 179110 227276
rect 192110 227264 192116 227276
rect 192168 227264 192174 227316
rect 234154 227304 234160 227316
rect 195256 227276 234160 227304
rect 157760 227208 164234 227236
rect 157760 227196 157766 227208
rect 72510 227128 72516 227180
rect 72568 227168 72574 227180
rect 156598 227168 156604 227180
rect 72568 227140 156604 227168
rect 72568 227128 72574 227140
rect 156598 227128 156604 227140
rect 156656 227128 156662 227180
rect 165154 227128 165160 227180
rect 165212 227168 165218 227180
rect 187234 227168 187240 227180
rect 165212 227140 187240 227168
rect 165212 227128 165218 227140
rect 187234 227128 187240 227140
rect 187292 227128 187298 227180
rect 195256 227168 195284 227276
rect 234154 227264 234160 227276
rect 234212 227264 234218 227316
rect 235994 227264 236000 227316
rect 236052 227304 236058 227316
rect 266170 227304 266176 227316
rect 236052 227276 266176 227304
rect 236052 227264 236058 227276
rect 266170 227264 266176 227276
rect 266228 227264 266234 227316
rect 267550 227264 267556 227316
rect 267608 227304 267614 227316
rect 287422 227304 287428 227316
rect 267608 227276 287428 227304
rect 267608 227264 267614 227276
rect 287422 227264 287428 227276
rect 287480 227264 287486 227316
rect 367186 227264 367192 227316
rect 367244 227304 367250 227316
rect 385586 227304 385592 227316
rect 367244 227276 385592 227304
rect 367244 227264 367250 227276
rect 385586 227264 385592 227276
rect 385644 227264 385650 227316
rect 415762 227264 415768 227316
rect 415820 227304 415826 227316
rect 458450 227304 458456 227316
rect 415820 227276 458456 227304
rect 415820 227264 415826 227276
rect 458450 227264 458456 227276
rect 458508 227264 458514 227316
rect 465258 227304 465264 227316
rect 460906 227276 465264 227304
rect 187528 227140 195284 227168
rect 63586 226992 63592 227044
rect 63644 227032 63650 227044
rect 142108 227032 142114 227044
rect 63644 227004 142114 227032
rect 63644 226992 63650 227004
rect 142108 226992 142114 227004
rect 142166 226992 142172 227044
rect 142246 226992 142252 227044
rect 142304 227032 142310 227044
rect 157518 227032 157524 227044
rect 142304 227004 157524 227032
rect 142304 226992 142310 227004
rect 157518 226992 157524 227004
rect 157576 226992 157582 227044
rect 157794 226992 157800 227044
rect 157852 227032 157858 227044
rect 157852 227004 179276 227032
rect 157852 226992 157858 227004
rect 122190 226856 122196 226908
rect 122248 226896 122254 226908
rect 179046 226896 179052 226908
rect 122248 226868 179052 226896
rect 122248 226856 122254 226868
rect 179046 226856 179052 226868
rect 179104 226856 179110 226908
rect 179248 226896 179276 227004
rect 182818 226992 182824 227044
rect 182876 227032 182882 227044
rect 185946 227032 185952 227044
rect 182876 227004 185952 227032
rect 182876 226992 182882 227004
rect 185946 226992 185952 227004
rect 186004 226992 186010 227044
rect 186130 226992 186136 227044
rect 186188 227032 186194 227044
rect 187528 227032 187556 227140
rect 197446 227128 197452 227180
rect 197504 227168 197510 227180
rect 204898 227168 204904 227180
rect 197504 227140 204904 227168
rect 197504 227128 197510 227140
rect 204898 227128 204904 227140
rect 204956 227128 204962 227180
rect 205082 227128 205088 227180
rect 205140 227168 205146 227180
rect 212626 227168 212632 227180
rect 205140 227140 212632 227168
rect 205140 227128 205146 227140
rect 212626 227128 212632 227140
rect 212684 227128 212690 227180
rect 235718 227128 235724 227180
rect 235776 227168 235782 227180
rect 267182 227168 267188 227180
rect 235776 227140 267188 227168
rect 235776 227128 235782 227140
rect 267182 227128 267188 227140
rect 267240 227128 267246 227180
rect 267366 227128 267372 227180
rect 267424 227168 267430 227180
rect 290182 227168 290188 227180
rect 267424 227140 290188 227168
rect 267424 227128 267430 227140
rect 290182 227128 290188 227140
rect 290240 227128 290246 227180
rect 293678 227128 293684 227180
rect 293736 227168 293742 227180
rect 305362 227168 305368 227180
rect 293736 227140 305368 227168
rect 293736 227128 293742 227140
rect 305362 227128 305368 227140
rect 305420 227128 305426 227180
rect 361482 227128 361488 227180
rect 361540 227168 361546 227180
rect 371510 227168 371516 227180
rect 361540 227140 371516 227168
rect 361540 227128 361546 227140
rect 371510 227128 371516 227140
rect 371568 227128 371574 227180
rect 382090 227128 382096 227180
rect 382148 227168 382154 227180
rect 407298 227168 407304 227180
rect 382148 227140 407304 227168
rect 382148 227128 382154 227140
rect 407298 227128 407304 227140
rect 407356 227128 407362 227180
rect 420178 227128 420184 227180
rect 420236 227168 420242 227180
rect 460906 227168 460934 227276
rect 465258 227264 465264 227276
rect 465316 227264 465322 227316
rect 475378 227264 475384 227316
rect 475436 227304 475442 227316
rect 548702 227304 548708 227316
rect 475436 227276 548708 227304
rect 475436 227264 475442 227276
rect 548702 227264 548708 227276
rect 548760 227264 548766 227316
rect 420236 227140 460934 227168
rect 420236 227128 420242 227140
rect 464982 227128 464988 227180
rect 465040 227168 465046 227180
rect 478322 227168 478328 227180
rect 465040 227140 478328 227168
rect 465040 227128 465046 227140
rect 478322 227128 478328 227140
rect 478380 227128 478386 227180
rect 479794 227128 479800 227180
rect 479852 227168 479858 227180
rect 554774 227168 554780 227180
rect 479852 227140 554780 227168
rect 479852 227128 479858 227140
rect 554774 227128 554780 227140
rect 554832 227128 554838 227180
rect 186188 227004 187556 227032
rect 186188 226992 186194 227004
rect 187970 226992 187976 227044
rect 188028 227032 188034 227044
rect 231946 227032 231952 227044
rect 188028 227004 231952 227032
rect 188028 226992 188034 227004
rect 231946 226992 231952 227004
rect 232004 226992 232010 227044
rect 237282 226992 237288 227044
rect 237340 227032 237346 227044
rect 237340 227004 258074 227032
rect 237340 226992 237346 227004
rect 179248 226868 204760 226896
rect 128814 226720 128820 226772
rect 128872 226760 128878 226772
rect 137278 226760 137284 226772
rect 128872 226732 137284 226760
rect 128872 226720 128878 226732
rect 137278 226720 137284 226732
rect 137336 226720 137342 226772
rect 137462 226720 137468 226772
rect 137520 226760 137526 226772
rect 142108 226760 142114 226772
rect 137520 226732 142114 226760
rect 137520 226720 137526 226732
rect 142108 226720 142114 226732
rect 142166 226720 142172 226772
rect 142246 226720 142252 226772
rect 142304 226760 142310 226772
rect 204732 226760 204760 226868
rect 204898 226856 204904 226908
rect 204956 226896 204962 226908
rect 240778 226896 240784 226908
rect 204956 226868 240784 226896
rect 204956 226856 204962 226868
rect 240778 226856 240784 226868
rect 240836 226856 240842 226908
rect 258046 226896 258074 227004
rect 263410 226992 263416 227044
rect 263468 227032 263474 227044
rect 272518 227032 272524 227044
rect 263468 227004 272524 227032
rect 263468 226992 263474 227004
rect 272518 226992 272524 227004
rect 272576 226992 272582 227044
rect 283650 226992 283656 227044
rect 283708 227032 283714 227044
rect 298462 227032 298468 227044
rect 283708 227004 298468 227032
rect 283708 226992 283714 227004
rect 298462 226992 298468 227004
rect 298520 226992 298526 227044
rect 299382 226992 299388 227044
rect 299440 227032 299446 227044
rect 310330 227032 310336 227044
rect 299440 227004 310336 227032
rect 299440 226992 299446 227004
rect 310330 226992 310336 227004
rect 310388 226992 310394 227044
rect 311066 226992 311072 227044
rect 311124 227032 311130 227044
rect 319162 227032 319168 227044
rect 311124 227004 319168 227032
rect 311124 226992 311130 227004
rect 319162 226992 319168 227004
rect 319220 226992 319226 227044
rect 353938 226992 353944 227044
rect 353996 227032 354002 227044
rect 365806 227032 365812 227044
rect 353996 227004 365812 227032
rect 353996 226992 354002 227004
rect 365806 226992 365812 227004
rect 365864 226992 365870 227044
rect 366818 226992 366824 227044
rect 366876 227032 366882 227044
rect 383930 227032 383936 227044
rect 366876 227004 383936 227032
rect 366876 226992 366882 227004
rect 383930 226992 383936 227004
rect 383988 226992 383994 227044
rect 388714 226992 388720 227044
rect 388772 227032 388778 227044
rect 417050 227032 417056 227044
rect 388772 227004 417056 227032
rect 388772 226992 388778 227004
rect 417050 226992 417056 227004
rect 417108 226992 417114 227044
rect 426250 226992 426256 227044
rect 426308 227032 426314 227044
rect 473538 227032 473544 227044
rect 426308 227004 473544 227032
rect 426308 226992 426314 227004
rect 473538 226992 473544 227004
rect 473596 226992 473602 227044
rect 480530 226992 480536 227044
rect 480588 227032 480594 227044
rect 484670 227032 484676 227044
rect 480588 227004 484676 227032
rect 480588 226992 480594 227004
rect 484670 226992 484676 227004
rect 484728 226992 484734 227044
rect 485314 226992 485320 227044
rect 485372 227032 485378 227044
rect 563882 227032 563888 227044
rect 485372 227004 563888 227032
rect 485372 226992 485378 227004
rect 563882 226992 563888 227004
rect 563940 226992 563946 227044
rect 267826 226896 267832 226908
rect 258046 226868 267832 226896
rect 267826 226856 267832 226868
rect 267884 226856 267890 226908
rect 399754 226856 399760 226908
rect 399812 226896 399818 226908
rect 433610 226896 433616 226908
rect 399812 226868 433616 226896
rect 399812 226856 399818 226868
rect 433610 226856 433616 226868
rect 433668 226856 433674 226908
rect 436186 226856 436192 226908
rect 436244 226896 436250 226908
rect 464982 226896 464988 226908
rect 436244 226868 464988 226896
rect 436244 226856 436250 226868
rect 464982 226856 464988 226868
rect 465040 226856 465046 226908
rect 465718 226856 465724 226908
rect 465776 226896 465782 226908
rect 519170 226896 519176 226908
rect 465776 226868 519176 226896
rect 465776 226856 465782 226868
rect 519170 226856 519176 226868
rect 519228 226856 519234 226908
rect 248506 226828 248512 226840
rect 248386 226800 248512 226828
rect 205082 226760 205088 226772
rect 142304 226732 200114 226760
rect 204732 226732 205088 226760
rect 142304 226720 142310 226732
rect 132218 226584 132224 226636
rect 132276 226624 132282 226636
rect 199654 226624 199660 226636
rect 132276 226596 199660 226624
rect 132276 226584 132282 226596
rect 199654 226584 199660 226596
rect 199712 226584 199718 226636
rect 200086 226624 200114 226732
rect 205082 226720 205088 226732
rect 205140 226720 205146 226772
rect 205634 226720 205640 226772
rect 205692 226760 205698 226772
rect 248386 226760 248414 226800
rect 248506 226788 248512 226800
rect 248564 226788 248570 226840
rect 205692 226732 248414 226760
rect 205692 226720 205698 226732
rect 427722 226720 427728 226772
rect 427780 226760 427786 226772
rect 427780 226720 427814 226760
rect 452746 226720 452752 226772
rect 452804 226760 452810 226772
rect 513374 226760 513380 226772
rect 452804 226732 513380 226760
rect 452804 226720 452810 226732
rect 513374 226720 513380 226732
rect 513432 226720 513438 226772
rect 206554 226624 206560 226636
rect 200086 226596 206560 226624
rect 206554 226584 206560 226596
rect 206612 226584 206618 226636
rect 241882 226624 241888 226636
rect 209746 226596 241888 226624
rect 141878 226448 141884 226500
rect 141936 226488 141942 226500
rect 142154 226488 142160 226500
rect 141936 226460 142160 226488
rect 141936 226448 141942 226460
rect 142154 226448 142160 226460
rect 142212 226448 142218 226500
rect 142338 226448 142344 226500
rect 142396 226488 142402 226500
rect 204346 226488 204352 226500
rect 142396 226460 204352 226488
rect 142396 226448 142402 226460
rect 204346 226448 204352 226460
rect 204404 226448 204410 226500
rect 138750 226380 138756 226432
rect 138808 226420 138814 226432
rect 141694 226420 141700 226432
rect 138808 226392 141700 226420
rect 138808 226380 138814 226392
rect 141694 226380 141700 226392
rect 141752 226380 141758 226432
rect 209746 226420 209774 226596
rect 241882 226584 241888 226596
rect 241940 226584 241946 226636
rect 427786 226624 427814 226720
rect 452746 226624 452752 226636
rect 427786 226596 452752 226624
rect 452746 226584 452752 226596
rect 452804 226584 452810 226636
rect 456058 226584 456064 226636
rect 456116 226624 456122 226636
rect 465718 226624 465724 226636
rect 456116 226596 465724 226624
rect 456116 226584 456122 226596
rect 465718 226584 465724 226596
rect 465776 226584 465782 226636
rect 465902 226584 465908 226636
rect 465960 226624 465966 226636
rect 520550 226624 520556 226636
rect 465960 226596 520556 226624
rect 465960 226584 465966 226596
rect 520550 226584 520556 226596
rect 520608 226584 520614 226636
rect 450538 226448 450544 226500
rect 450596 226488 450602 226500
rect 489868 226488 489874 226500
rect 450596 226460 489874 226488
rect 450596 226448 450602 226460
rect 489868 226448 489874 226460
rect 489926 226448 489932 226500
rect 490926 226448 490932 226500
rect 490984 226488 490990 226500
rect 495526 226488 495532 226500
rect 490984 226460 495532 226488
rect 490984 226448 490990 226460
rect 495526 226448 495532 226460
rect 495584 226448 495590 226500
rect 204640 226392 209774 226420
rect 201954 226312 201960 226364
rect 202012 226352 202018 226364
rect 204640 226352 204668 226392
rect 243354 226380 243360 226432
rect 243412 226420 243418 226432
rect 246850 226420 246856 226432
rect 243412 226392 246856 226420
rect 243412 226380 243418 226392
rect 246850 226380 246856 226392
rect 246908 226380 246914 226432
rect 202012 226324 204668 226352
rect 202012 226312 202018 226324
rect 289538 226312 289544 226364
rect 289596 226352 289602 226364
rect 293862 226352 293868 226364
rect 289596 226324 293868 226352
rect 289596 226312 289602 226324
rect 293862 226312 293868 226324
rect 293920 226312 293926 226364
rect 97902 226244 97908 226296
rect 97960 226284 97966 226296
rect 166994 226284 167000 226296
rect 97960 226256 167000 226284
rect 97960 226244 97966 226256
rect 166994 226244 167000 226256
rect 167052 226244 167058 226296
rect 167178 226244 167184 226296
rect 167236 226284 167242 226296
rect 173434 226284 173440 226296
rect 167236 226256 173440 226284
rect 167236 226244 167242 226256
rect 173434 226244 173440 226256
rect 173492 226244 173498 226296
rect 173618 226244 173624 226296
rect 173676 226284 173682 226296
rect 175642 226284 175648 226296
rect 173676 226256 175648 226284
rect 173676 226244 173682 226256
rect 175642 226244 175648 226256
rect 175700 226244 175706 226296
rect 175826 226244 175832 226296
rect 175884 226284 175890 226296
rect 175884 226256 176654 226284
rect 175884 226244 175890 226256
rect 42426 226176 42432 226228
rect 42484 226216 42490 226228
rect 45554 226216 45560 226228
rect 42484 226188 45560 226216
rect 42484 226176 42490 226188
rect 45554 226176 45560 226188
rect 45612 226176 45618 226228
rect 84930 226108 84936 226160
rect 84988 226148 84994 226160
rect 84988 226120 162256 226148
rect 84988 226108 84994 226120
rect 92382 225972 92388 226024
rect 92440 226012 92446 226024
rect 162228 226012 162256 226120
rect 162394 226108 162400 226160
rect 162452 226148 162458 226160
rect 162452 226120 171824 226148
rect 162452 226108 162458 226120
rect 165982 226012 165988 226024
rect 92440 225984 162164 226012
rect 162228 225984 165988 226012
rect 92440 225972 92446 225984
rect 88058 225836 88064 225888
rect 88116 225876 88122 225888
rect 162136 225876 162164 225984
rect 165982 225972 165988 225984
rect 166040 225972 166046 226024
rect 166442 225972 166448 226024
rect 166500 226012 166506 226024
rect 167362 226012 167368 226024
rect 166500 225984 167368 226012
rect 166500 225972 166506 225984
rect 167362 225972 167368 225984
rect 167420 225972 167426 226024
rect 168466 226012 168472 226024
rect 167656 225984 168472 226012
rect 167178 225876 167184 225888
rect 88116 225848 162072 225876
rect 162136 225848 167184 225876
rect 88116 225836 88122 225848
rect 78398 225700 78404 225752
rect 78456 225740 78462 225752
rect 161842 225740 161848 225752
rect 78456 225712 161848 225740
rect 78456 225700 78462 225712
rect 161842 225700 161848 225712
rect 161900 225700 161906 225752
rect 162044 225740 162072 225848
rect 167178 225836 167184 225848
rect 167236 225836 167242 225888
rect 167656 225740 167684 225984
rect 168466 225972 168472 225984
rect 168524 225972 168530 226024
rect 171796 226012 171824 226120
rect 173250 226108 173256 226160
rect 173308 226148 173314 226160
rect 176470 226148 176476 226160
rect 173308 226120 176476 226148
rect 173308 226108 173314 226120
rect 176470 226108 176476 226120
rect 176528 226108 176534 226160
rect 176626 226148 176654 226256
rect 176746 226244 176752 226296
rect 176804 226284 176810 226296
rect 190270 226284 190276 226296
rect 176804 226256 190276 226284
rect 176804 226244 176810 226256
rect 190270 226244 190276 226256
rect 190328 226244 190334 226296
rect 190408 226244 190414 226296
rect 190466 226284 190472 226296
rect 195054 226284 195060 226296
rect 190466 226256 195060 226284
rect 190466 226244 190472 226256
rect 195054 226244 195060 226256
rect 195112 226244 195118 226296
rect 195238 226244 195244 226296
rect 195296 226284 195302 226296
rect 201770 226284 201776 226296
rect 195296 226256 201776 226284
rect 195296 226244 195302 226256
rect 201770 226244 201776 226256
rect 201828 226244 201834 226296
rect 205450 226244 205456 226296
rect 205508 226284 205514 226296
rect 247402 226284 247408 226296
rect 205508 226256 247408 226284
rect 205508 226244 205514 226256
rect 247402 226244 247408 226256
rect 247460 226244 247466 226296
rect 413002 226244 413008 226296
rect 413060 226284 413066 226296
rect 449066 226284 449072 226296
rect 413060 226256 449072 226284
rect 413060 226244 413066 226256
rect 449066 226244 449072 226256
rect 449124 226244 449130 226296
rect 469306 226244 469312 226296
rect 469364 226284 469370 226296
rect 540330 226284 540336 226296
rect 469364 226256 540336 226284
rect 469364 226244 469370 226256
rect 540330 226244 540336 226256
rect 540388 226244 540394 226296
rect 176626 226120 181208 226148
rect 181180 226012 181208 226120
rect 181346 226108 181352 226160
rect 181404 226148 181410 226160
rect 224218 226148 224224 226160
rect 181404 226120 224224 226148
rect 181404 226108 181410 226120
rect 224218 226108 224224 226120
rect 224276 226108 224282 226160
rect 225690 226108 225696 226160
rect 225748 226148 225754 226160
rect 260650 226148 260656 226160
rect 225748 226120 260656 226148
rect 225748 226108 225754 226120
rect 260650 226108 260656 226120
rect 260708 226108 260714 226160
rect 273714 226108 273720 226160
rect 273772 226148 273778 226160
rect 292114 226148 292120 226160
rect 273772 226120 292120 226148
rect 273772 226108 273778 226120
rect 292114 226108 292120 226120
rect 292172 226108 292178 226160
rect 379882 226108 379888 226160
rect 379940 226148 379946 226160
rect 402974 226148 402980 226160
rect 379940 226120 402980 226148
rect 379940 226108 379946 226120
rect 402974 226108 402980 226120
rect 403032 226108 403038 226160
rect 408586 226108 408592 226160
rect 408644 226148 408650 226160
rect 447042 226148 447048 226160
rect 408644 226120 447048 226148
rect 408644 226108 408650 226120
rect 447042 226108 447048 226120
rect 447100 226108 447106 226160
rect 478690 226108 478696 226160
rect 478748 226148 478754 226160
rect 553670 226148 553676 226160
rect 478748 226120 553676 226148
rect 478748 226108 478754 226120
rect 553670 226108 553676 226120
rect 553728 226108 553734 226160
rect 226426 226012 226432 226024
rect 171796 225984 181116 226012
rect 181180 225984 226432 226012
rect 168282 225836 168288 225888
rect 168340 225876 168346 225888
rect 180794 225876 180800 225888
rect 168340 225848 180800 225876
rect 168340 225836 168346 225848
rect 180794 225836 180800 225848
rect 180852 225836 180858 225888
rect 181088 225876 181116 225984
rect 226426 225972 226432 225984
rect 226484 225972 226490 226024
rect 255222 225972 255228 226024
rect 255280 226012 255286 226024
rect 280522 226012 280528 226024
rect 255280 225984 280528 226012
rect 255280 225972 255286 225984
rect 280522 225972 280528 225984
rect 280580 225972 280586 226024
rect 381170 225972 381176 226024
rect 381228 226012 381234 226024
rect 394878 226012 394884 226024
rect 381228 225984 394884 226012
rect 381228 225972 381234 225984
rect 394878 225972 394884 225984
rect 394936 225972 394942 226024
rect 400674 225972 400680 226024
rect 400732 226012 400738 226024
rect 400732 225984 412634 226012
rect 400732 225972 400738 225984
rect 219802 225876 219808 225888
rect 181088 225848 219808 225876
rect 219802 225836 219808 225848
rect 219860 225836 219866 225888
rect 224218 225836 224224 225888
rect 224276 225876 224282 225888
rect 230842 225876 230848 225888
rect 224276 225848 230848 225876
rect 224276 225836 224282 225848
rect 230842 225836 230848 225848
rect 230900 225836 230906 225888
rect 252738 225836 252744 225888
rect 252796 225876 252802 225888
rect 279418 225876 279424 225888
rect 252796 225848 279424 225876
rect 252796 225836 252802 225848
rect 279418 225836 279424 225848
rect 279476 225836 279482 225888
rect 382642 225836 382648 225888
rect 382700 225876 382706 225888
rect 408770 225876 408776 225888
rect 382700 225848 408776 225876
rect 382700 225836 382706 225848
rect 408770 225836 408776 225848
rect 408828 225836 408834 225888
rect 412606 225876 412634 225984
rect 425146 225972 425152 226024
rect 425204 226012 425210 226024
rect 469306 226012 469312 226024
rect 425204 225984 469312 226012
rect 425204 225972 425210 225984
rect 469306 225972 469312 225984
rect 469364 225972 469370 226024
rect 475102 225972 475108 226024
rect 475160 226012 475166 226024
rect 483566 226012 483572 226024
rect 475160 225984 483572 226012
rect 475160 225972 475166 225984
rect 483566 225972 483572 225984
rect 483624 225972 483630 226024
rect 484026 225972 484032 226024
rect 484084 226012 484090 226024
rect 489546 226012 489552 226024
rect 484084 225984 489552 226012
rect 484084 225972 484090 225984
rect 489546 225972 489552 225984
rect 489604 225972 489610 226024
rect 489730 225972 489736 226024
rect 489788 226012 489794 226024
rect 556154 226012 556160 226024
rect 489788 225984 556160 226012
rect 489788 225972 489794 225984
rect 556154 225972 556160 225984
rect 556212 225972 556218 226024
rect 425790 225876 425796 225888
rect 412606 225848 425796 225876
rect 425790 225836 425796 225848
rect 425848 225836 425854 225888
rect 427906 225836 427912 225888
rect 427964 225876 427970 225888
rect 474182 225876 474188 225888
rect 427964 225848 474188 225876
rect 427964 225836 427970 225848
rect 474182 225836 474188 225848
rect 474240 225836 474246 225888
rect 482002 225836 482008 225888
rect 482060 225876 482066 225888
rect 558914 225876 558920 225888
rect 482060 225848 558920 225876
rect 482060 225836 482066 225848
rect 558914 225836 558920 225848
rect 558972 225836 558978 225888
rect 162044 225712 167684 225740
rect 167822 225700 167828 225752
rect 167880 225740 167886 225752
rect 214374 225740 214380 225752
rect 167880 225712 214380 225740
rect 167880 225700 167886 225712
rect 214374 225700 214380 225712
rect 214432 225700 214438 225752
rect 214558 225700 214564 225752
rect 214616 225740 214622 225752
rect 226978 225740 226984 225752
rect 214616 225712 226984 225740
rect 214616 225700 214622 225712
rect 226978 225700 226984 225712
rect 227036 225700 227042 225752
rect 227162 225700 227168 225752
rect 227220 225740 227226 225752
rect 259546 225740 259552 225752
rect 227220 225712 259552 225740
rect 227220 225700 227226 225712
rect 259546 225700 259552 225712
rect 259604 225700 259610 225752
rect 260558 225700 260564 225752
rect 260616 225740 260622 225752
rect 283282 225740 283288 225752
rect 260616 225712 283288 225740
rect 260616 225700 260622 225712
rect 283282 225700 283288 225712
rect 283340 225700 283346 225752
rect 290274 225700 290280 225752
rect 290332 225740 290338 225752
rect 303154 225740 303160 225752
rect 290332 225712 303160 225740
rect 290332 225700 290338 225712
rect 303154 225700 303160 225712
rect 303212 225700 303218 225752
rect 303338 225700 303344 225752
rect 303396 225740 303402 225752
rect 310882 225740 310888 225752
rect 303396 225712 310888 225740
rect 303396 225700 303402 225712
rect 310882 225700 310888 225712
rect 310940 225700 310946 225752
rect 312722 225700 312728 225752
rect 312780 225740 312786 225752
rect 317506 225740 317512 225752
rect 312780 225712 317512 225740
rect 312780 225700 312786 225712
rect 317506 225700 317512 225712
rect 317564 225700 317570 225752
rect 352282 225700 352288 225752
rect 352340 225740 352346 225752
rect 357618 225740 357624 225752
rect 352340 225712 357624 225740
rect 352340 225700 352346 225712
rect 357618 225700 357624 225712
rect 357676 225700 357682 225752
rect 362770 225700 362776 225752
rect 362828 225740 362834 225752
rect 378962 225740 378968 225752
rect 362828 225712 378968 225740
rect 362828 225700 362834 225712
rect 378962 225700 378968 225712
rect 379020 225700 379026 225752
rect 386874 225700 386880 225752
rect 386932 225740 386938 225752
rect 414014 225740 414020 225752
rect 386932 225712 414020 225740
rect 386932 225700 386938 225712
rect 414014 225700 414020 225712
rect 414072 225700 414078 225752
rect 438210 225700 438216 225752
rect 438268 225740 438274 225752
rect 489868 225740 489874 225752
rect 438268 225712 489874 225740
rect 438268 225700 438274 225712
rect 489868 225700 489874 225712
rect 489926 225700 489932 225752
rect 490006 225700 490012 225752
rect 490064 225740 490070 225752
rect 561214 225740 561220 225752
rect 490064 225712 561220 225740
rect 490064 225700 490070 225712
rect 561214 225700 561220 225712
rect 561272 225700 561278 225752
rect 62114 225564 62120 225616
rect 62172 225604 62178 225616
rect 149698 225604 149704 225616
rect 62172 225576 149704 225604
rect 62172 225564 62178 225576
rect 149698 225564 149704 225576
rect 149756 225564 149762 225616
rect 151170 225564 151176 225616
rect 151228 225604 151234 225616
rect 213178 225604 213184 225616
rect 151228 225576 213184 225604
rect 151228 225564 151234 225576
rect 213178 225564 213184 225576
rect 213236 225564 213242 225616
rect 214190 225564 214196 225616
rect 214248 225604 214254 225616
rect 224218 225604 224224 225616
rect 214248 225576 224224 225604
rect 214248 225564 214254 225576
rect 224218 225564 224224 225576
rect 224276 225564 224282 225616
rect 246758 225564 246764 225616
rect 246816 225604 246822 225616
rect 274174 225604 274180 225616
rect 246816 225576 274180 225604
rect 246816 225564 246822 225576
rect 274174 225564 274180 225576
rect 274232 225564 274238 225616
rect 279602 225564 279608 225616
rect 279660 225604 279666 225616
rect 297082 225604 297088 225616
rect 279660 225576 297088 225604
rect 279660 225564 279666 225576
rect 297082 225564 297088 225576
rect 297140 225564 297146 225616
rect 298002 225564 298008 225616
rect 298060 225604 298066 225616
rect 308122 225604 308128 225616
rect 298060 225576 308128 225604
rect 298060 225564 298066 225576
rect 308122 225564 308128 225576
rect 308180 225564 308186 225616
rect 357066 225564 357072 225616
rect 357124 225604 357130 225616
rect 365254 225604 365260 225616
rect 357124 225576 365260 225604
rect 357124 225564 357130 225576
rect 365254 225564 365260 225576
rect 365312 225564 365318 225616
rect 365438 225564 365444 225616
rect 365496 225604 365502 225616
rect 382642 225604 382648 225616
rect 365496 225576 382648 225604
rect 365496 225564 365502 225576
rect 382642 225564 382648 225576
rect 382700 225564 382706 225616
rect 393682 225564 393688 225616
rect 393740 225604 393746 225616
rect 423030 225604 423036 225616
rect 393740 225576 423036 225604
rect 393740 225564 393746 225576
rect 423030 225564 423036 225576
rect 423088 225564 423094 225616
rect 433978 225564 433984 225616
rect 434036 225604 434042 225616
rect 475102 225604 475108 225616
rect 434036 225576 475108 225604
rect 434036 225564 434042 225576
rect 475102 225564 475108 225576
rect 475160 225564 475166 225616
rect 480346 225564 480352 225616
rect 480404 225604 480410 225616
rect 486786 225604 486792 225616
rect 480404 225576 486792 225604
rect 480404 225564 480410 225576
rect 486786 225564 486792 225576
rect 486844 225564 486850 225616
rect 486970 225564 486976 225616
rect 487028 225604 487034 225616
rect 566090 225604 566096 225616
rect 487028 225576 566096 225604
rect 487028 225564 487034 225576
rect 566090 225564 566096 225576
rect 566148 225564 566154 225616
rect 81342 225428 81348 225480
rect 81400 225468 81406 225480
rect 158438 225468 158444 225480
rect 81400 225440 158444 225468
rect 81400 225428 81406 225440
rect 158438 225428 158444 225440
rect 158496 225428 158502 225480
rect 158622 225428 158628 225480
rect 158680 225468 158686 225480
rect 212350 225468 212356 225480
rect 158680 225440 212356 225468
rect 158680 225428 158686 225440
rect 212350 225428 212356 225440
rect 212408 225428 212414 225480
rect 212534 225428 212540 225480
rect 212592 225468 212598 225480
rect 215386 225468 215392 225480
rect 212592 225440 215392 225468
rect 212592 225428 212598 225440
rect 215386 225428 215392 225440
rect 215444 225428 215450 225480
rect 215570 225428 215576 225480
rect 215628 225468 215634 225480
rect 215628 225440 217824 225468
rect 215628 225428 215634 225440
rect 104802 225292 104808 225344
rect 104860 225332 104866 225344
rect 178126 225332 178132 225344
rect 104860 225304 178132 225332
rect 104860 225292 104866 225304
rect 178126 225292 178132 225304
rect 178184 225292 178190 225344
rect 178494 225292 178500 225344
rect 178552 225332 178558 225344
rect 214190 225332 214196 225344
rect 178552 225304 214196 225332
rect 178552 225292 178558 225304
rect 214190 225292 214196 225304
rect 214248 225292 214254 225344
rect 214742 225292 214748 225344
rect 214800 225332 214806 225344
rect 217594 225332 217600 225344
rect 214800 225304 217600 225332
rect 214800 225292 214806 225304
rect 217594 225292 217600 225304
rect 217652 225292 217658 225344
rect 217796 225332 217824 225440
rect 219158 225428 219164 225480
rect 219216 225468 219222 225480
rect 255958 225468 255964 225480
rect 219216 225440 255964 225468
rect 219216 225428 219222 225440
rect 255958 225428 255964 225440
rect 256016 225428 256022 225480
rect 410794 225428 410800 225480
rect 410852 225468 410858 225480
rect 437474 225468 437480 225480
rect 410852 225440 437480 225468
rect 410852 225428 410858 225440
rect 437474 225428 437480 225440
rect 437532 225428 437538 225480
rect 448882 225428 448888 225480
rect 448940 225468 448946 225480
rect 509510 225468 509516 225480
rect 448940 225440 509516 225468
rect 448940 225428 448946 225440
rect 509510 225428 509516 225440
rect 509568 225428 509574 225480
rect 252922 225332 252928 225344
rect 217796 225304 252928 225332
rect 252922 225292 252928 225304
rect 252980 225292 252986 225344
rect 417418 225292 417424 225344
rect 417476 225332 417482 225344
rect 436738 225332 436744 225344
rect 417476 225304 436744 225332
rect 417476 225292 417482 225304
rect 436738 225292 436744 225304
rect 436796 225292 436802 225344
rect 442626 225292 442632 225344
rect 442684 225332 442690 225344
rect 489868 225332 489874 225344
rect 442684 225304 489874 225332
rect 442684 225292 442690 225304
rect 489868 225292 489874 225304
rect 489926 225292 489932 225344
rect 490006 225292 490012 225344
rect 490064 225332 490070 225344
rect 492582 225332 492588 225344
rect 490064 225304 492588 225332
rect 490064 225292 490070 225304
rect 492582 225292 492588 225304
rect 492640 225292 492646 225344
rect 492766 225292 492772 225344
rect 492824 225332 492830 225344
rect 499022 225332 499028 225344
rect 492824 225304 499028 225332
rect 492824 225292 492830 225304
rect 499022 225292 499028 225304
rect 499080 225292 499086 225344
rect 134978 225156 134984 225208
rect 135036 225196 135042 225208
rect 195238 225196 195244 225208
rect 135036 225168 195244 225196
rect 135036 225156 135042 225168
rect 195238 225156 195244 225168
rect 195296 225156 195302 225208
rect 195422 225156 195428 225208
rect 195480 225196 195486 225208
rect 214558 225196 214564 225208
rect 195480 225168 214564 225196
rect 195480 225156 195486 225168
rect 214558 225156 214564 225168
rect 214616 225156 214622 225208
rect 215754 225156 215760 225208
rect 215812 225196 215818 225208
rect 254026 225196 254032 225208
rect 215812 225168 254032 225196
rect 215812 225156 215818 225168
rect 254026 225156 254032 225168
rect 254084 225156 254090 225208
rect 407482 225156 407488 225208
rect 407540 225196 407546 225208
rect 421098 225196 421104 225208
rect 407540 225168 421104 225196
rect 407540 225156 407546 225168
rect 421098 225156 421104 225168
rect 421156 225156 421162 225208
rect 440050 225156 440056 225208
rect 440108 225196 440114 225208
rect 495710 225196 495716 225208
rect 440108 225168 495716 225196
rect 440108 225156 440114 225168
rect 495710 225156 495716 225168
rect 495768 225156 495774 225208
rect 120074 225020 120080 225072
rect 120132 225060 120138 225072
rect 151630 225060 151636 225072
rect 120132 225032 151636 225060
rect 120132 225020 120138 225032
rect 151630 225020 151636 225032
rect 151688 225020 151694 225072
rect 151768 225020 151774 225072
rect 151826 225060 151832 225072
rect 161290 225060 161296 225072
rect 151826 225032 161296 225060
rect 151826 225020 151832 225032
rect 161290 225020 161296 225032
rect 161348 225020 161354 225072
rect 161474 225020 161480 225072
rect 161532 225060 161538 225072
rect 212534 225060 212540 225072
rect 161532 225032 212540 225060
rect 161532 225020 161538 225032
rect 212534 225020 212540 225032
rect 212592 225020 212598 225072
rect 214374 225020 214380 225072
rect 214432 225060 214438 225072
rect 221458 225060 221464 225072
rect 214432 225032 221464 225060
rect 214432 225020 214438 225032
rect 221458 225020 221464 225032
rect 221516 225020 221522 225072
rect 222286 225020 222292 225072
rect 222344 225060 222350 225072
rect 227162 225060 227168 225072
rect 222344 225032 227168 225060
rect 222344 225020 222350 225032
rect 227162 225020 227168 225032
rect 227220 225020 227226 225072
rect 231670 225020 231676 225072
rect 231728 225060 231734 225072
rect 238018 225060 238024 225072
rect 231728 225032 238024 225060
rect 231728 225020 231734 225032
rect 238018 225020 238024 225032
rect 238076 225020 238082 225072
rect 445938 225020 445944 225072
rect 445996 225060 446002 225072
rect 501506 225060 501512 225072
rect 445996 225032 501512 225060
rect 445996 225020 446002 225032
rect 501506 225020 501512 225032
rect 501564 225020 501570 225072
rect 378042 224952 378048 225004
rect 378100 224992 378106 225004
rect 379790 224992 379796 225004
rect 378100 224964 379796 224992
rect 378100 224952 378106 224964
rect 379790 224952 379796 224964
rect 379848 224952 379854 225004
rect 42610 224884 42616 224936
rect 42668 224924 42674 224936
rect 45738 224924 45744 224936
rect 42668 224896 45744 224924
rect 42668 224884 42674 224896
rect 45738 224884 45744 224896
rect 45796 224884 45802 224936
rect 121362 224884 121368 224936
rect 121420 224924 121426 224936
rect 121420 224896 184704 224924
rect 121420 224884 121426 224896
rect 77018 224748 77024 224800
rect 77076 224788 77082 224800
rect 151446 224788 151452 224800
rect 77076 224760 151452 224788
rect 77076 224748 77082 224760
rect 151446 224748 151452 224760
rect 151504 224748 151510 224800
rect 151722 224748 151728 224800
rect 151780 224788 151786 224800
rect 159358 224788 159364 224800
rect 151780 224760 159364 224788
rect 151780 224748 151786 224760
rect 159358 224748 159364 224760
rect 159416 224748 159422 224800
rect 159726 224748 159732 224800
rect 159784 224788 159790 224800
rect 180610 224788 180616 224800
rect 159784 224760 180616 224788
rect 159784 224748 159790 224760
rect 180610 224748 180616 224760
rect 180668 224748 180674 224800
rect 180794 224748 180800 224800
rect 180852 224788 180858 224800
rect 181898 224788 181904 224800
rect 180852 224760 181904 224788
rect 180852 224748 180858 224760
rect 181898 224748 181904 224760
rect 181956 224748 181962 224800
rect 184676 224788 184704 224896
rect 184842 224884 184848 224936
rect 184900 224924 184906 224936
rect 194410 224924 194416 224936
rect 184900 224896 194416 224924
rect 184900 224884 184906 224896
rect 194410 224884 194416 224896
rect 194468 224884 194474 224936
rect 194870 224884 194876 224936
rect 194928 224924 194934 224936
rect 198274 224924 198280 224936
rect 194928 224896 198280 224924
rect 194928 224884 194934 224896
rect 198274 224884 198280 224896
rect 198332 224884 198338 224936
rect 198458 224884 198464 224936
rect 198516 224924 198522 224936
rect 243722 224924 243728 224936
rect 198516 224896 243728 224924
rect 198516 224884 198522 224896
rect 243722 224884 243728 224896
rect 243780 224884 243786 224936
rect 244550 224884 244556 224936
rect 244608 224924 244614 224936
rect 272794 224924 272800 224936
rect 244608 224896 272800 224924
rect 244608 224884 244614 224896
rect 272794 224884 272800 224896
rect 272852 224884 272858 224936
rect 370498 224884 370504 224936
rect 370556 224924 370562 224936
rect 376110 224924 376116 224936
rect 370556 224896 376116 224924
rect 370556 224884 370562 224896
rect 376110 224884 376116 224896
rect 376168 224884 376174 224936
rect 409782 224884 409788 224936
rect 409840 224924 409846 224936
rect 441062 224924 441068 224936
rect 409840 224896 441068 224924
rect 409840 224884 409846 224896
rect 441062 224884 441068 224896
rect 441120 224884 441126 224936
rect 442810 224884 442816 224936
rect 442868 224924 442874 224936
rect 442868 224896 463188 224924
rect 442868 224884 442874 224896
rect 187050 224788 187056 224800
rect 184676 224760 187056 224788
rect 187050 224748 187056 224760
rect 187108 224748 187114 224800
rect 187234 224748 187240 224800
rect 187292 224788 187298 224800
rect 234706 224788 234712 224800
rect 187292 224760 234712 224788
rect 187292 224748 187298 224760
rect 234706 224748 234712 224760
rect 234764 224748 234770 224800
rect 240594 224748 240600 224800
rect 240652 224788 240658 224800
rect 270034 224788 270040 224800
rect 240652 224760 270040 224788
rect 240652 224748 240658 224760
rect 270034 224748 270040 224760
rect 270092 224748 270098 224800
rect 347866 224748 347872 224800
rect 347924 224788 347930 224800
rect 353478 224788 353484 224800
rect 347924 224760 353484 224788
rect 347924 224748 347930 224760
rect 353478 224748 353484 224760
rect 353536 224748 353542 224800
rect 394694 224748 394700 224800
rect 394752 224788 394758 224800
rect 411254 224788 411260 224800
rect 394752 224760 411260 224788
rect 394752 224748 394758 224760
rect 411254 224748 411260 224760
rect 411312 224748 411318 224800
rect 412450 224748 412456 224800
rect 412508 224788 412514 224800
rect 451274 224788 451280 224800
rect 412508 224760 451280 224788
rect 412508 224748 412514 224760
rect 451274 224748 451280 224760
rect 451332 224748 451338 224800
rect 451458 224748 451464 224800
rect 451516 224788 451522 224800
rect 462958 224788 462964 224800
rect 451516 224760 462964 224788
rect 451516 224748 451522 224760
rect 462958 224748 462964 224760
rect 463016 224748 463022 224800
rect 463160 224788 463188 224896
rect 464338 224884 464344 224936
rect 464396 224924 464402 224936
rect 471790 224924 471796 224936
rect 464396 224896 471796 224924
rect 464396 224884 464402 224896
rect 471790 224884 471796 224896
rect 471848 224884 471854 224936
rect 472250 224884 472256 224936
rect 472308 224924 472314 224936
rect 534166 224924 534172 224936
rect 472308 224896 534172 224924
rect 472308 224884 472314 224896
rect 534166 224884 534172 224896
rect 534224 224884 534230 224936
rect 465074 224788 465080 224800
rect 463160 224760 465080 224788
rect 465074 224748 465080 224760
rect 465132 224748 465138 224800
rect 467098 224748 467104 224800
rect 467156 224788 467162 224800
rect 536374 224788 536380 224800
rect 467156 224760 536380 224788
rect 467156 224748 467162 224760
rect 536374 224748 536380 224760
rect 536432 224748 536438 224800
rect 99098 224612 99104 224664
rect 99156 224652 99162 224664
rect 177850 224652 177856 224664
rect 99156 224624 177856 224652
rect 99156 224612 99162 224624
rect 177850 224612 177856 224624
rect 177908 224612 177914 224664
rect 178034 224612 178040 224664
rect 178092 224652 178098 224664
rect 194870 224652 194876 224664
rect 178092 224624 194876 224652
rect 178092 224612 178098 224624
rect 194870 224612 194876 224624
rect 194928 224612 194934 224664
rect 197262 224612 197268 224664
rect 197320 224652 197326 224664
rect 204530 224652 204536 224664
rect 197320 224624 204536 224652
rect 197320 224612 197326 224624
rect 204530 224612 204536 224624
rect 204588 224612 204594 224664
rect 204714 224612 204720 224664
rect 204772 224652 204778 224664
rect 210694 224652 210700 224664
rect 204772 224624 210700 224652
rect 204772 224612 204778 224624
rect 210694 224612 210700 224624
rect 210752 224612 210758 224664
rect 210878 224612 210884 224664
rect 210936 224652 210942 224664
rect 229186 224652 229192 224664
rect 210936 224624 229192 224652
rect 210936 224612 210942 224624
rect 229186 224612 229192 224624
rect 229244 224612 229250 224664
rect 231854 224612 231860 224664
rect 231912 224652 231918 224664
rect 236914 224652 236920 224664
rect 231912 224624 236920 224652
rect 231912 224612 231918 224624
rect 236914 224612 236920 224624
rect 236972 224612 236978 224664
rect 238570 224612 238576 224664
rect 238628 224652 238634 224664
rect 269482 224652 269488 224664
rect 238628 224624 269488 224652
rect 238628 224612 238634 224624
rect 269482 224612 269488 224624
rect 269540 224612 269546 224664
rect 281258 224612 281264 224664
rect 281316 224652 281322 224664
rect 296714 224652 296720 224664
rect 281316 224624 296720 224652
rect 281316 224612 281322 224624
rect 296714 224612 296720 224624
rect 296772 224612 296778 224664
rect 375834 224612 375840 224664
rect 375892 224652 375898 224664
rect 397546 224652 397552 224664
rect 375892 224624 397552 224652
rect 375892 224612 375898 224624
rect 397546 224612 397552 224624
rect 397604 224612 397610 224664
rect 397914 224612 397920 224664
rect 397972 224652 397978 224664
rect 414566 224652 414572 224664
rect 397972 224624 414572 224652
rect 397972 224612 397978 224624
rect 414566 224612 414572 224624
rect 414624 224612 414630 224664
rect 414750 224612 414756 224664
rect 414808 224652 414814 224664
rect 454310 224652 454316 224664
rect 414808 224624 454316 224652
rect 414808 224612 414814 224624
rect 454310 224612 454316 224624
rect 454368 224612 454374 224664
rect 460474 224612 460480 224664
rect 460532 224652 460538 224664
rect 524230 224652 524236 224664
rect 460532 224624 524236 224652
rect 460532 224612 460538 224624
rect 524230 224612 524236 224624
rect 524288 224612 524294 224664
rect 524368 224612 524374 224664
rect 524426 224652 524432 224664
rect 533338 224652 533344 224664
rect 524426 224624 533344 224652
rect 524426 224612 524432 224624
rect 533338 224612 533344 224624
rect 533396 224612 533402 224664
rect 74994 224476 75000 224528
rect 75052 224516 75058 224528
rect 151722 224516 151728 224528
rect 75052 224488 151728 224516
rect 75052 224476 75058 224488
rect 151722 224476 151728 224488
rect 151780 224476 151786 224528
rect 152090 224476 152096 224528
rect 152148 224516 152154 224528
rect 155034 224516 155040 224528
rect 152148 224488 155040 224516
rect 152148 224476 152154 224488
rect 155034 224476 155040 224488
rect 155092 224476 155098 224528
rect 155402 224476 155408 224528
rect 155460 224516 155466 224528
rect 157288 224516 157294 224528
rect 155460 224488 157294 224516
rect 155460 224476 155466 224488
rect 157288 224476 157294 224488
rect 157346 224476 157352 224528
rect 157426 224476 157432 224528
rect 157484 224516 157490 224528
rect 159726 224516 159732 224528
rect 157484 224488 159732 224516
rect 157484 224476 157490 224488
rect 159726 224476 159732 224488
rect 159784 224476 159790 224528
rect 159910 224476 159916 224528
rect 159968 224516 159974 224528
rect 162946 224516 162952 224528
rect 159968 224488 162952 224516
rect 159968 224476 159974 224488
rect 162946 224476 162952 224488
rect 163004 224476 163010 224528
rect 163130 224476 163136 224528
rect 163188 224516 163194 224528
rect 218698 224516 218704 224528
rect 163188 224488 218704 224516
rect 163188 224476 163194 224488
rect 218698 224476 218704 224488
rect 218756 224476 218762 224528
rect 232314 224476 232320 224528
rect 232372 224516 232378 224528
rect 265066 224516 265072 224528
rect 232372 224488 265072 224516
rect 232372 224476 232378 224488
rect 265066 224476 265072 224488
rect 265124 224476 265130 224528
rect 270218 224476 270224 224528
rect 270276 224516 270282 224528
rect 288250 224516 288256 224528
rect 270276 224488 288256 224516
rect 270276 224476 270282 224488
rect 288250 224476 288256 224488
rect 288308 224476 288314 224528
rect 304994 224476 305000 224528
rect 305052 224516 305058 224528
rect 312538 224516 312544 224528
rect 305052 224488 312544 224516
rect 305052 224476 305058 224488
rect 312538 224476 312544 224488
rect 312596 224476 312602 224528
rect 368382 224476 368388 224528
rect 368440 224516 368446 224528
rect 376754 224516 376760 224528
rect 368440 224488 376760 224516
rect 368440 224476 368446 224488
rect 376754 224476 376760 224488
rect 376812 224476 376818 224528
rect 384114 224476 384120 224528
rect 384172 224516 384178 224528
rect 407942 224516 407948 224528
rect 384172 224488 407948 224516
rect 384172 224476 384178 224488
rect 407942 224476 407948 224488
rect 408000 224476 408006 224528
rect 423398 224476 423404 224528
rect 423456 224516 423462 224528
rect 445294 224516 445300 224528
rect 423456 224488 445300 224516
rect 423456 224476 423462 224488
rect 445294 224476 445300 224488
rect 445352 224476 445358 224528
rect 446122 224476 446128 224528
rect 446180 224516 446186 224528
rect 461578 224516 461584 224528
rect 446180 224488 461584 224516
rect 446180 224476 446186 224488
rect 461578 224476 461584 224488
rect 461636 224476 461642 224528
rect 465442 224476 465448 224528
rect 465500 224516 465506 224528
rect 472250 224516 472256 224528
rect 465500 224488 472256 224516
rect 465500 224476 465506 224488
rect 472250 224476 472256 224488
rect 472308 224476 472314 224528
rect 475378 224516 475384 224528
rect 472452 224488 475384 224516
rect 61838 224340 61844 224392
rect 61896 224380 61902 224392
rect 146018 224380 146024 224392
rect 61896 224352 146024 224380
rect 61896 224340 61902 224352
rect 146018 224340 146024 224352
rect 146076 224340 146082 224392
rect 146202 224340 146208 224392
rect 146260 224380 146266 224392
rect 206830 224380 206836 224392
rect 146260 224352 206836 224380
rect 146260 224340 146266 224352
rect 206830 224340 206836 224352
rect 206888 224340 206894 224392
rect 207014 224340 207020 224392
rect 207072 224380 207078 224392
rect 207934 224380 207940 224392
rect 207072 224352 207940 224380
rect 207072 224340 207078 224352
rect 207934 224340 207940 224352
rect 207992 224340 207998 224392
rect 210418 224340 210424 224392
rect 210476 224380 210482 224392
rect 212074 224380 212080 224392
rect 210476 224352 212080 224380
rect 210476 224340 210482 224352
rect 212074 224340 212080 224352
rect 212132 224340 212138 224392
rect 214558 224340 214564 224392
rect 214616 224380 214622 224392
rect 250714 224380 250720 224392
rect 214616 224352 250720 224380
rect 214616 224340 214622 224352
rect 250714 224340 250720 224352
rect 250772 224340 250778 224392
rect 271598 224340 271604 224392
rect 271656 224380 271662 224392
rect 291562 224380 291568 224392
rect 271656 224352 291568 224380
rect 271656 224340 271662 224352
rect 291562 224340 291568 224352
rect 291620 224340 291626 224392
rect 296622 224340 296628 224392
rect 296680 224380 296686 224392
rect 307570 224380 307576 224392
rect 296680 224352 307576 224380
rect 296680 224340 296686 224352
rect 307570 224340 307576 224352
rect 307628 224340 307634 224392
rect 359734 224340 359740 224392
rect 359792 224380 359798 224392
rect 368474 224380 368480 224392
rect 359792 224352 368480 224380
rect 359792 224340 359798 224352
rect 368474 224340 368480 224352
rect 368532 224340 368538 224392
rect 376386 224340 376392 224392
rect 376444 224380 376450 224392
rect 399018 224380 399024 224392
rect 376444 224352 399024 224380
rect 376444 224340 376450 224352
rect 399018 224340 399024 224352
rect 399076 224340 399082 224392
rect 423674 224340 423680 224392
rect 423732 224380 423738 224392
rect 467926 224380 467932 224392
rect 423732 224352 467932 224380
rect 423732 224340 423738 224352
rect 467926 224340 467932 224352
rect 467984 224340 467990 224392
rect 470410 224340 470416 224392
rect 470468 224380 470474 224392
rect 472452 224380 472480 224488
rect 475378 224476 475384 224488
rect 475436 224476 475442 224528
rect 475562 224476 475568 224528
rect 475620 224516 475626 224528
rect 543918 224516 543924 224528
rect 475620 224488 543924 224516
rect 475620 224476 475626 224488
rect 543918 224476 543924 224488
rect 543976 224476 543982 224528
rect 470468 224352 472480 224380
rect 470468 224340 470474 224352
rect 472618 224340 472624 224392
rect 472676 224380 472682 224392
rect 533154 224380 533160 224392
rect 472676 224352 533160 224380
rect 472676 224340 472682 224352
rect 533154 224340 533160 224352
rect 533212 224340 533218 224392
rect 533338 224340 533344 224392
rect 533396 224380 533402 224392
rect 541342 224380 541348 224392
rect 533396 224352 541348 224380
rect 533396 224340 533402 224352
rect 541342 224340 541348 224352
rect 541400 224340 541406 224392
rect 542078 224340 542084 224392
rect 542136 224380 542142 224392
rect 557350 224380 557356 224392
rect 542136 224352 557356 224380
rect 542136 224340 542142 224352
rect 557350 224340 557356 224352
rect 557408 224340 557414 224392
rect 68462 224204 68468 224256
rect 68520 224244 68526 224256
rect 155218 224244 155224 224256
rect 68520 224216 155224 224244
rect 68520 224204 68526 224216
rect 155218 224204 155224 224216
rect 155276 224204 155282 224256
rect 155586 224204 155592 224256
rect 155644 224244 155650 224256
rect 204714 224244 204720 224256
rect 155644 224216 204720 224244
rect 155644 224204 155650 224216
rect 204714 224204 204720 224216
rect 204772 224204 204778 224256
rect 204898 224204 204904 224256
rect 204956 224244 204962 224256
rect 204956 224216 232084 224244
rect 204956 224204 204962 224216
rect 124674 224068 124680 224120
rect 124732 224108 124738 224120
rect 190362 224108 190368 224120
rect 124732 224080 190368 224108
rect 124732 224068 124738 224080
rect 190362 224068 190368 224080
rect 190420 224068 190426 224120
rect 191742 224068 191748 224120
rect 191800 224108 191806 224120
rect 231854 224108 231860 224120
rect 191800 224080 231860 224108
rect 191800 224068 191806 224080
rect 231854 224068 231860 224080
rect 231912 224068 231918 224120
rect 232056 224108 232084 224216
rect 234614 224204 234620 224256
rect 234672 224244 234678 224256
rect 268378 224244 268384 224256
rect 234672 224216 268384 224244
rect 234672 224204 234678 224216
rect 268378 224204 268384 224216
rect 268436 224204 268442 224256
rect 270402 224204 270408 224256
rect 270460 224244 270466 224256
rect 289906 224244 289912 224256
rect 270460 224216 289912 224244
rect 270460 224204 270466 224216
rect 289906 224204 289912 224216
rect 289964 224204 289970 224256
rect 291194 224204 291200 224256
rect 291252 224244 291258 224256
rect 305914 224244 305920 224256
rect 291252 224216 305920 224244
rect 291252 224204 291258 224216
rect 305914 224204 305920 224216
rect 305972 224204 305978 224256
rect 307478 224204 307484 224256
rect 307536 224244 307542 224256
rect 315022 224244 315028 224256
rect 307536 224216 315028 224244
rect 307536 224204 307542 224216
rect 315022 224204 315028 224216
rect 315080 224204 315086 224256
rect 358354 224204 358360 224256
rect 358412 224244 358418 224256
rect 372706 224244 372712 224256
rect 358412 224216 372712 224244
rect 358412 224204 358418 224216
rect 372706 224204 372712 224216
rect 372764 224204 372770 224256
rect 380434 224204 380440 224256
rect 380492 224244 380498 224256
rect 405734 224244 405740 224256
rect 380492 224216 405740 224244
rect 380492 224204 380498 224216
rect 405734 224204 405740 224216
rect 405792 224204 405798 224256
rect 406654 224204 406660 224256
rect 406712 224244 406718 224256
rect 431126 224244 431132 224256
rect 406712 224216 431132 224244
rect 406712 224204 406718 224216
rect 431126 224204 431132 224216
rect 431184 224204 431190 224256
rect 435634 224204 435640 224256
rect 435692 224244 435698 224256
rect 485222 224244 485228 224256
rect 435692 224216 485228 224244
rect 435692 224204 435698 224216
rect 485222 224204 485228 224216
rect 485280 224204 485286 224256
rect 499482 224244 499488 224256
rect 485608 224216 499488 224244
rect 485608 224176 485636 224216
rect 499482 224204 499488 224216
rect 499540 224204 499546 224256
rect 505186 224204 505192 224256
rect 505244 224244 505250 224256
rect 547414 224244 547420 224256
rect 505244 224216 547420 224244
rect 505244 224204 505250 224216
rect 547414 224204 547420 224216
rect 547472 224204 547478 224256
rect 562318 224204 562324 224256
rect 562376 224244 562382 224256
rect 571334 224244 571340 224256
rect 562376 224216 571340 224244
rect 562376 224204 562382 224216
rect 571334 224204 571340 224216
rect 571392 224204 571398 224256
rect 485378 224148 485636 224176
rect 234982 224108 234988 224120
rect 232056 224080 234988 224108
rect 234982 224068 234988 224080
rect 235040 224068 235046 224120
rect 399478 224068 399484 224120
rect 399536 224108 399542 224120
rect 418154 224108 418160 224120
rect 399536 224080 418160 224108
rect 399536 224068 399542 224080
rect 418154 224068 418160 224080
rect 418212 224068 418218 224120
rect 429838 224068 429844 224120
rect 429896 224108 429902 224120
rect 461026 224108 461032 224120
rect 429896 224080 461032 224108
rect 429896 224068 429902 224080
rect 461026 224068 461032 224080
rect 461084 224068 461090 224120
rect 461578 224068 461584 224120
rect 461636 224108 461642 224120
rect 466454 224108 466460 224120
rect 461636 224080 466460 224108
rect 461636 224068 461642 224080
rect 466454 224068 466460 224080
rect 466512 224068 466518 224120
rect 468754 224068 468760 224120
rect 468812 224108 468818 224120
rect 472618 224108 472624 224120
rect 468812 224080 472624 224108
rect 468812 224068 468818 224080
rect 472618 224068 472624 224080
rect 472676 224068 472682 224120
rect 475378 224068 475384 224120
rect 475436 224108 475442 224120
rect 480898 224108 480904 224120
rect 475436 224080 480904 224108
rect 475436 224068 475442 224080
rect 480898 224068 480904 224080
rect 480956 224068 480962 224120
rect 481082 224068 481088 224120
rect 481140 224108 481146 224120
rect 485378 224108 485406 224148
rect 499666 224136 499672 224188
rect 499724 224176 499730 224188
rect 504910 224176 504916 224188
rect 499724 224148 504916 224176
rect 499724 224136 499730 224148
rect 504910 224136 504916 224148
rect 504968 224136 504974 224188
rect 481140 224080 485406 224108
rect 481140 224068 481146 224080
rect 485774 224068 485780 224120
rect 485832 224108 485838 224120
rect 499482 224108 499488 224120
rect 485832 224080 499488 224108
rect 485832 224068 485838 224080
rect 499482 224068 499488 224080
rect 499540 224068 499546 224120
rect 509878 224068 509884 224120
rect 509936 224108 509942 224120
rect 551278 224108 551284 224120
rect 509936 224080 551284 224108
rect 509936 224068 509942 224080
rect 551278 224068 551284 224080
rect 551336 224068 551342 224120
rect 131022 223932 131028 223984
rect 131080 223972 131086 223984
rect 131080 223944 193720 223972
rect 131080 223932 131086 223944
rect 134702 223796 134708 223848
rect 134760 223836 134766 223848
rect 193490 223836 193496 223848
rect 134760 223808 193496 223836
rect 134760 223796 134766 223808
rect 193490 223796 193496 223808
rect 193548 223796 193554 223848
rect 193692 223836 193720 223944
rect 194410 223932 194416 223984
rect 194468 223972 194474 223984
rect 204898 223972 204904 223984
rect 194468 223944 204904 223972
rect 194468 223932 194474 223944
rect 204898 223932 204904 223944
rect 204956 223932 204962 223984
rect 241146 223972 241152 223984
rect 205100 223944 241152 223972
rect 196894 223836 196900 223848
rect 193692 223808 196900 223836
rect 196894 223796 196900 223808
rect 196952 223796 196958 223848
rect 200850 223796 200856 223848
rect 200908 223836 200914 223848
rect 200908 223808 204024 223836
rect 200908 223796 200914 223808
rect 141234 223660 141240 223712
rect 141292 223700 141298 223712
rect 203794 223700 203800 223712
rect 141292 223672 203800 223700
rect 141292 223660 141298 223672
rect 203794 223660 203800 223672
rect 203852 223660 203858 223712
rect 203996 223700 204024 223808
rect 204530 223796 204536 223848
rect 204588 223836 204594 223848
rect 205100 223836 205128 223944
rect 241146 223932 241152 223944
rect 241204 223932 241210 223984
rect 272978 223932 272984 223984
rect 273036 223972 273042 223984
rect 275646 223972 275652 223984
rect 273036 223944 275652 223972
rect 273036 223932 273042 223944
rect 275646 223932 275652 223944
rect 275704 223932 275710 223984
rect 403250 223932 403256 223984
rect 403308 223972 403314 223984
rect 424686 223972 424692 223984
rect 403308 223944 424692 223972
rect 403308 223932 403314 223944
rect 424686 223932 424692 223944
rect 424744 223932 424750 223984
rect 425514 223932 425520 223984
rect 425572 223972 425578 223984
rect 457714 223972 457720 223984
rect 425572 223944 457720 223972
rect 425572 223932 425578 223944
rect 457714 223932 457720 223944
rect 457772 223932 457778 223984
rect 462130 223932 462136 223984
rect 462188 223972 462194 223984
rect 528830 223972 528836 223984
rect 462188 223944 528836 223972
rect 462188 223932 462194 223944
rect 528830 223932 528836 223944
rect 528888 223932 528894 223984
rect 533154 223932 533160 223984
rect 533212 223972 533218 223984
rect 538858 223972 538864 223984
rect 533212 223944 538864 223972
rect 533212 223932 533218 223944
rect 538858 223932 538864 223944
rect 538916 223932 538922 223984
rect 243170 223836 243176 223848
rect 204588 223808 205128 223836
rect 205284 223808 243176 223836
rect 204588 223796 204594 223808
rect 205284 223700 205312 223808
rect 243170 223796 243176 223808
rect 243228 223796 243234 223848
rect 412726 223796 412732 223848
rect 412784 223836 412790 223848
rect 447686 223836 447692 223848
rect 412784 223808 447692 223836
rect 412784 223796 412790 223808
rect 447686 223796 447692 223808
rect 447744 223796 447750 223848
rect 454770 223796 454776 223848
rect 454828 223836 454834 223848
rect 454828 223808 499804 223836
rect 454828 223796 454834 223808
rect 203996 223672 205312 223700
rect 208394 223660 208400 223712
rect 208452 223700 208458 223712
rect 214558 223700 214564 223712
rect 208452 223672 214564 223700
rect 208452 223660 208458 223672
rect 214558 223660 214564 223672
rect 214616 223660 214622 223712
rect 416314 223660 416320 223712
rect 416372 223700 416378 223712
rect 429194 223700 429200 223712
rect 416372 223672 429200 223700
rect 416372 223660 416378 223672
rect 429194 223660 429200 223672
rect 429252 223660 429258 223712
rect 472434 223660 472440 223712
rect 472492 223700 472498 223712
rect 475562 223700 475568 223712
rect 472492 223672 475568 223700
rect 472492 223660 472498 223672
rect 475562 223660 475568 223672
rect 475620 223660 475626 223712
rect 477034 223660 477040 223712
rect 477092 223700 477098 223712
rect 477092 223672 480760 223700
rect 477092 223660 477098 223672
rect 242894 223592 242900 223644
rect 242952 223632 242958 223644
rect 245194 223632 245200 223644
rect 242952 223604 245200 223632
rect 242952 223592 242958 223604
rect 245194 223592 245200 223604
rect 245252 223592 245258 223644
rect 94958 223524 94964 223576
rect 95016 223564 95022 223576
rect 95016 223536 171134 223564
rect 95016 223524 95022 223536
rect 91554 223388 91560 223440
rect 91612 223428 91618 223440
rect 161934 223428 161940 223440
rect 91612 223400 161940 223428
rect 91612 223388 91618 223400
rect 161934 223388 161940 223400
rect 161992 223388 161998 223440
rect 167638 223428 167644 223440
rect 162136 223400 167644 223428
rect 86678 223252 86684 223304
rect 86736 223292 86742 223304
rect 162136 223292 162164 223400
rect 167638 223388 167644 223400
rect 167696 223388 167702 223440
rect 171106 223428 171134 223536
rect 173802 223524 173808 223576
rect 173860 223564 173866 223576
rect 173860 223536 177252 223564
rect 173860 223524 173866 223536
rect 172606 223428 172612 223440
rect 171106 223400 172612 223428
rect 172606 223388 172612 223400
rect 172664 223388 172670 223440
rect 173526 223388 173532 223440
rect 173584 223428 173590 223440
rect 177022 223428 177028 223440
rect 173584 223400 177028 223428
rect 173584 223388 173590 223400
rect 177022 223388 177028 223400
rect 177080 223388 177086 223440
rect 177224 223428 177252 223536
rect 180702 223524 180708 223576
rect 180760 223564 180766 223576
rect 230290 223564 230296 223576
rect 180760 223536 230296 223564
rect 180760 223524 180766 223536
rect 230290 223524 230296 223536
rect 230348 223524 230354 223576
rect 250530 223524 250536 223576
rect 250588 223564 250594 223576
rect 276474 223564 276480 223576
rect 250588 223536 276480 223564
rect 250588 223524 250594 223536
rect 276474 223524 276480 223536
rect 276532 223524 276538 223576
rect 277118 223524 277124 223576
rect 277176 223564 277182 223576
rect 294322 223564 294328 223576
rect 277176 223536 294328 223564
rect 277176 223524 277182 223536
rect 294322 223524 294328 223536
rect 294380 223524 294386 223576
rect 313090 223524 313096 223576
rect 313148 223564 313154 223576
rect 318610 223564 318616 223576
rect 313148 223536 318616 223564
rect 313148 223524 313154 223536
rect 318610 223524 318616 223536
rect 318668 223524 318674 223576
rect 350166 223524 350172 223576
rect 350224 223564 350230 223576
rect 355686 223564 355692 223576
rect 350224 223536 355692 223564
rect 350224 223524 350230 223536
rect 355686 223524 355692 223536
rect 355744 223524 355750 223576
rect 369578 223524 369584 223576
rect 369636 223564 369642 223576
rect 373994 223564 374000 223576
rect 369636 223536 374000 223564
rect 369636 223524 369642 223536
rect 373994 223524 374000 223536
rect 374052 223524 374058 223576
rect 387242 223564 387248 223576
rect 378796 223536 387248 223564
rect 223114 223428 223120 223440
rect 177224 223400 223120 223428
rect 223114 223388 223120 223400
rect 223172 223388 223178 223440
rect 226058 223388 226064 223440
rect 226116 223428 226122 223440
rect 227346 223428 227352 223440
rect 226116 223400 227352 223428
rect 226116 223388 226122 223400
rect 227346 223388 227352 223400
rect 227404 223388 227410 223440
rect 227622 223388 227628 223440
rect 227680 223428 227686 223440
rect 258626 223428 258632 223440
rect 227680 223400 258632 223428
rect 227680 223388 227686 223400
rect 258626 223388 258632 223400
rect 258684 223388 258690 223440
rect 258810 223388 258816 223440
rect 258868 223428 258874 223440
rect 282454 223428 282460 223440
rect 258868 223400 282460 223428
rect 258868 223388 258874 223400
rect 282454 223388 282460 223400
rect 282512 223388 282518 223440
rect 310606 223388 310612 223440
rect 310664 223428 310670 223440
rect 314194 223428 314200 223440
rect 310664 223400 314200 223428
rect 310664 223388 310670 223400
rect 314194 223388 314200 223400
rect 314252 223388 314258 223440
rect 345106 223388 345112 223440
rect 345164 223428 345170 223440
rect 352466 223428 352472 223440
rect 345164 223400 352472 223428
rect 345164 223388 345170 223400
rect 352466 223388 352472 223400
rect 352524 223388 352530 223440
rect 368842 223388 368848 223440
rect 368900 223428 368906 223440
rect 378796 223428 378824 223536
rect 387242 223524 387248 223536
rect 387300 223524 387306 223576
rect 392854 223524 392860 223576
rect 392912 223564 392918 223576
rect 416222 223564 416228 223576
rect 392912 223536 416228 223564
rect 392912 223524 392918 223536
rect 416222 223524 416228 223536
rect 416280 223524 416286 223576
rect 424226 223524 424232 223576
rect 424284 223564 424290 223576
rect 436186 223564 436192 223576
rect 424284 223536 436192 223564
rect 424284 223524 424290 223536
rect 436186 223524 436192 223536
rect 436244 223524 436250 223576
rect 443730 223524 443736 223576
rect 443788 223564 443794 223576
rect 444190 223564 444196 223576
rect 443788 223536 444196 223564
rect 443788 223524 443794 223536
rect 444190 223524 444196 223536
rect 444248 223524 444254 223576
rect 480732 223564 480760 223672
rect 480898 223660 480904 223712
rect 480956 223700 480962 223712
rect 499298 223700 499304 223712
rect 480956 223672 499304 223700
rect 480956 223660 480962 223672
rect 499298 223660 499304 223672
rect 499356 223660 499362 223712
rect 499776 223700 499804 223808
rect 499942 223796 499948 223848
rect 500000 223836 500006 223848
rect 509878 223836 509884 223848
rect 500000 223808 509884 223836
rect 500000 223796 500006 223808
rect 509878 223796 509884 223808
rect 509936 223796 509942 223848
rect 510062 223796 510068 223848
rect 510120 223836 510126 223848
rect 514570 223836 514576 223848
rect 510120 223808 514576 223836
rect 510120 223796 510126 223808
rect 514570 223796 514576 223808
rect 514628 223796 514634 223848
rect 516778 223796 516784 223848
rect 516836 223836 516842 223848
rect 524230 223836 524236 223848
rect 516836 223808 524236 223836
rect 516836 223796 516842 223808
rect 524230 223796 524236 223808
rect 524288 223796 524294 223848
rect 524368 223796 524374 223848
rect 524426 223836 524432 223848
rect 617702 223836 617708 223848
rect 524426 223808 617708 223836
rect 524426 223796 524432 223808
rect 617702 223796 617708 223808
rect 617760 223796 617766 223848
rect 504726 223700 504732 223712
rect 499776 223672 504732 223700
rect 504726 223660 504732 223672
rect 504784 223660 504790 223712
rect 511966 223672 521654 223700
rect 499528 223632 499534 223644
rect 499487 223604 499534 223632
rect 499528 223592 499534 223604
rect 499586 223632 499592 223644
rect 511966 223632 511994 223672
rect 499586 223592 499620 223632
rect 485222 223564 485228 223576
rect 480732 223536 485228 223564
rect 485222 223524 485228 223536
rect 485280 223524 485286 223576
rect 485866 223524 485872 223576
rect 485924 223564 485930 223576
rect 499298 223564 499304 223576
rect 485924 223536 499304 223564
rect 485924 223524 485930 223536
rect 499298 223524 499304 223536
rect 499356 223524 499362 223576
rect 499592 223564 499620 223592
rect 505204 223604 511994 223632
rect 521626 223632 521654 223672
rect 629846 223632 629852 223644
rect 521626 223604 629852 223632
rect 505204 223564 505232 223604
rect 629846 223592 629852 223604
rect 629904 223592 629910 223644
rect 499592 223536 505232 223564
rect 505370 223456 505376 223508
rect 505428 223496 505434 223508
rect 516778 223496 516784 223508
rect 505428 223468 516784 223496
rect 505428 223456 505434 223468
rect 516778 223456 516784 223468
rect 516836 223456 516842 223508
rect 368900 223400 378824 223428
rect 368900 223388 368906 223400
rect 379330 223388 379336 223440
rect 379388 223428 379394 223440
rect 393498 223428 393504 223440
rect 379388 223400 393504 223428
rect 379388 223388 379394 223400
rect 393498 223388 393504 223400
rect 393556 223388 393562 223440
rect 401686 223388 401692 223440
rect 401744 223428 401750 223440
rect 426618 223428 426624 223440
rect 401744 223400 426624 223428
rect 401744 223388 401750 223400
rect 426618 223388 426624 223400
rect 426676 223388 426682 223440
rect 436554 223388 436560 223440
rect 436612 223428 436618 223440
rect 449894 223428 449900 223440
rect 436612 223400 449900 223428
rect 436612 223388 436618 223400
rect 449894 223388 449900 223400
rect 449952 223388 449958 223440
rect 452194 223388 452200 223440
rect 452252 223428 452258 223440
rect 505186 223428 505192 223440
rect 452252 223400 505192 223428
rect 452252 223388 452258 223400
rect 505186 223388 505192 223400
rect 505244 223388 505250 223440
rect 522574 223388 522580 223440
rect 522632 223428 522638 223440
rect 554958 223428 554964 223440
rect 522632 223400 554964 223428
rect 522632 223388 522638 223400
rect 554958 223388 554964 223400
rect 555016 223388 555022 223440
rect 170674 223292 170680 223304
rect 86736 223264 162164 223292
rect 162228 223264 170680 223292
rect 86736 223252 86742 223264
rect 74258 223116 74264 223168
rect 74316 223156 74322 223168
rect 82906 223156 82912 223168
rect 74316 223128 82912 223156
rect 74316 223116 74322 223128
rect 82906 223116 82912 223128
rect 82964 223116 82970 223168
rect 83274 223116 83280 223168
rect 83332 223156 83338 223168
rect 157288 223156 157294 223168
rect 83332 223128 157294 223156
rect 83332 223116 83338 223128
rect 157288 223116 157294 223128
rect 157346 223116 157352 223168
rect 157426 223116 157432 223168
rect 157484 223156 157490 223168
rect 161106 223156 161112 223168
rect 157484 223128 161112 223156
rect 157484 223116 157490 223128
rect 161106 223116 161112 223128
rect 161164 223116 161170 223168
rect 161934 223116 161940 223168
rect 161992 223156 161998 223168
rect 162228 223156 162256 223264
rect 170674 223252 170680 223264
rect 170732 223252 170738 223304
rect 170858 223252 170864 223304
rect 170916 223292 170922 223304
rect 223666 223292 223672 223304
rect 170916 223264 223672 223292
rect 170916 223252 170922 223264
rect 223666 223252 223672 223264
rect 223724 223252 223730 223304
rect 227438 223252 227444 223304
rect 227496 223292 227502 223304
rect 261110 223292 261116 223304
rect 227496 223264 261116 223292
rect 227496 223252 227502 223264
rect 261110 223252 261116 223264
rect 261168 223252 261174 223304
rect 261294 223252 261300 223304
rect 261352 223292 261358 223304
rect 286042 223292 286048 223304
rect 261352 223264 286048 223292
rect 261352 223252 261358 223264
rect 286042 223252 286048 223264
rect 286100 223252 286106 223304
rect 293954 223252 293960 223304
rect 294012 223292 294018 223304
rect 302050 223292 302056 223304
rect 294012 223264 302056 223292
rect 294012 223252 294018 223264
rect 302050 223252 302056 223264
rect 302108 223252 302114 223304
rect 362402 223252 362408 223304
rect 362460 223292 362466 223304
rect 362460 223264 364334 223292
rect 362460 223252 362466 223264
rect 161992 223128 162256 223156
rect 161992 223116 161998 223128
rect 165246 223116 165252 223168
rect 165304 223156 165310 223168
rect 173066 223156 173072 223168
rect 165304 223128 173072 223156
rect 165304 223116 165310 223128
rect 173066 223116 173072 223128
rect 173124 223116 173130 223168
rect 185578 223156 185584 223168
rect 173636 223128 185584 223156
rect 79778 222980 79784 223032
rect 79836 223020 79842 223032
rect 163498 223020 163504 223032
rect 79836 222992 163504 223020
rect 79836 222980 79842 222992
rect 163498 222980 163504 222992
rect 163556 222980 163562 223032
rect 164142 222980 164148 223032
rect 164200 223020 164206 223032
rect 173636 223020 173664 223128
rect 185578 223116 185584 223128
rect 185636 223116 185642 223168
rect 185762 223116 185768 223168
rect 185820 223156 185826 223168
rect 185820 223128 219434 223156
rect 185820 223116 185826 223128
rect 164200 222992 173664 223020
rect 164200 222980 164206 222992
rect 174078 222980 174084 223032
rect 174136 223020 174142 223032
rect 214558 223020 214564 223032
rect 174136 222992 214564 223020
rect 174136 222980 174142 222992
rect 214558 222980 214564 222992
rect 214616 222980 214622 223032
rect 214742 222980 214748 223032
rect 214800 223020 214806 223032
rect 218974 223020 218980 223032
rect 214800 222992 218980 223020
rect 214800 222980 214806 222992
rect 218974 222980 218980 222992
rect 219032 222980 219038 223032
rect 219406 223020 219434 223128
rect 224218 223116 224224 223168
rect 224276 223156 224282 223168
rect 227622 223156 227628 223168
rect 224276 223128 227628 223156
rect 224276 223116 224282 223128
rect 227622 223116 227628 223128
rect 227680 223116 227686 223168
rect 228634 223156 228640 223168
rect 227824 223128 228640 223156
rect 227824 223020 227852 223128
rect 228634 223116 228640 223128
rect 228692 223116 228698 223168
rect 252278 223116 252284 223168
rect 252336 223156 252342 223168
rect 278314 223156 278320 223168
rect 252336 223128 278320 223156
rect 252336 223116 252342 223128
rect 278314 223116 278320 223128
rect 278372 223116 278378 223168
rect 288342 223116 288348 223168
rect 288400 223156 288406 223168
rect 302602 223156 302608 223168
rect 288400 223128 302608 223156
rect 288400 223116 288406 223128
rect 302602 223116 302608 223128
rect 302660 223116 302666 223168
rect 353018 223116 353024 223168
rect 353076 223156 353082 223168
rect 357434 223156 357440 223168
rect 353076 223128 357440 223156
rect 353076 223116 353082 223128
rect 357434 223116 357440 223128
rect 357492 223116 357498 223168
rect 363138 223116 363144 223168
rect 363196 223156 363202 223168
rect 364306 223156 364334 223264
rect 377858 223252 377864 223304
rect 377916 223292 377922 223304
rect 396350 223292 396356 223304
rect 377916 223264 396356 223292
rect 377916 223252 377922 223264
rect 396350 223252 396356 223264
rect 396408 223252 396414 223304
rect 397178 223252 397184 223304
rect 397236 223292 397242 223304
rect 422846 223292 422852 223304
rect 397236 223264 422852 223292
rect 397236 223252 397242 223264
rect 422846 223252 422852 223264
rect 422904 223252 422910 223304
rect 427538 223252 427544 223304
rect 427596 223292 427602 223304
rect 446030 223292 446036 223304
rect 427596 223264 446036 223292
rect 427596 223252 427602 223264
rect 446030 223252 446036 223264
rect 446088 223252 446094 223304
rect 447870 223252 447876 223304
rect 447928 223292 447934 223304
rect 455690 223292 455696 223304
rect 447928 223264 455696 223292
rect 447928 223252 447934 223264
rect 455690 223252 455696 223264
rect 455748 223252 455754 223304
rect 455874 223252 455880 223304
rect 455932 223292 455938 223304
rect 518986 223292 518992 223304
rect 455932 223264 518992 223292
rect 455932 223252 455938 223264
rect 518986 223252 518992 223264
rect 519044 223252 519050 223304
rect 519538 223252 519544 223304
rect 519596 223292 519602 223304
rect 531314 223292 531320 223304
rect 519596 223264 531320 223292
rect 519596 223252 519602 223264
rect 531314 223252 531320 223264
rect 531372 223252 531378 223304
rect 369854 223156 369860 223168
rect 363196 223128 363552 223156
rect 364306 223128 369860 223156
rect 363196 223116 363202 223128
rect 219406 222992 227852 223020
rect 228174 222980 228180 223032
rect 228232 223020 228238 223032
rect 263962 223020 263968 223032
rect 228232 222992 263968 223020
rect 228232 222980 228238 222992
rect 263962 222980 263968 222992
rect 264020 222980 264026 223032
rect 278682 222980 278688 223032
rect 278740 223020 278746 223032
rect 295978 223020 295984 223032
rect 278740 222992 295984 223020
rect 278740 222980 278746 222992
rect 295978 222980 295984 222992
rect 296036 222980 296042 223032
rect 302234 222980 302240 223032
rect 302292 223020 302298 223032
rect 311434 223020 311440 223032
rect 302292 222992 311440 223020
rect 302292 222980 302298 222992
rect 311434 222980 311440 222992
rect 311492 222980 311498 223032
rect 354398 222980 354404 223032
rect 354456 223020 354462 223032
rect 363230 223020 363236 223032
rect 354456 222992 363236 223020
rect 354456 222980 354462 222992
rect 363230 222980 363236 222992
rect 363288 222980 363294 223032
rect 363524 223020 363552 223128
rect 369854 223116 369860 223128
rect 369912 223116 369918 223168
rect 374362 223116 374368 223168
rect 374420 223156 374426 223168
rect 379330 223156 379336 223168
rect 374420 223128 379336 223156
rect 374420 223116 374426 223128
rect 379330 223116 379336 223128
rect 379388 223116 379394 223168
rect 385770 223116 385776 223168
rect 385828 223156 385834 223168
rect 409966 223156 409972 223168
rect 385828 223128 409972 223156
rect 385828 223116 385834 223128
rect 409966 223116 409972 223128
rect 410024 223116 410030 223168
rect 411898 223116 411904 223168
rect 411956 223156 411962 223168
rect 444006 223156 444012 223168
rect 411956 223128 444012 223156
rect 411956 223116 411962 223128
rect 444006 223116 444012 223128
rect 444064 223116 444070 223168
rect 444190 223116 444196 223168
rect 444248 223156 444254 223168
rect 485728 223156 485734 223168
rect 444248 223128 485734 223156
rect 444248 223116 444254 223128
rect 485728 223116 485734 223128
rect 485786 223116 485792 223168
rect 485866 223116 485872 223168
rect 485924 223156 485930 223168
rect 560386 223156 560392 223168
rect 485924 223128 560392 223156
rect 485924 223116 485930 223128
rect 560386 223116 560392 223128
rect 560444 223116 560450 223168
rect 369026 223020 369032 223032
rect 363524 222992 369032 223020
rect 369026 222980 369032 222992
rect 369084 222980 369090 223032
rect 373626 222980 373632 223032
rect 373684 223020 373690 223032
rect 392210 223020 392216 223032
rect 373684 222992 392216 223020
rect 373684 222980 373690 222992
rect 392210 222980 392216 222992
rect 392268 222980 392274 223032
rect 394050 222980 394056 223032
rect 394108 223020 394114 223032
rect 419718 223020 419724 223032
rect 394108 222992 419724 223020
rect 394108 222980 394114 222992
rect 419718 222980 419724 222992
rect 419776 222980 419782 223032
rect 426066 222980 426072 223032
rect 426124 223020 426130 223032
rect 463878 223020 463884 223032
rect 426124 222992 463884 223020
rect 426124 222980 426130 222992
rect 463878 222980 463884 222992
rect 463936 222980 463942 223032
rect 464154 222980 464160 223032
rect 464212 223020 464218 223032
rect 464212 222992 491248 223020
rect 464212 222980 464218 222992
rect 60366 222844 60372 222896
rect 60424 222884 60430 222896
rect 142108 222884 142114 222896
rect 60424 222856 142114 222884
rect 60424 222844 60430 222856
rect 142108 222844 142114 222856
rect 142166 222844 142172 222896
rect 142430 222844 142436 222896
rect 142488 222884 142494 222896
rect 152458 222884 152464 222896
rect 142488 222856 152464 222884
rect 142488 222844 142494 222856
rect 152458 222844 152464 222856
rect 152516 222844 152522 222896
rect 152642 222844 152648 222896
rect 152700 222884 152706 222896
rect 157150 222884 157156 222896
rect 152700 222856 157156 222884
rect 152700 222844 152706 222856
rect 157150 222844 157156 222856
rect 157208 222844 157214 222896
rect 157334 222844 157340 222896
rect 157392 222884 157398 222896
rect 158162 222884 158168 222896
rect 157392 222856 158168 222884
rect 157392 222844 157398 222856
rect 158162 222844 158168 222856
rect 158220 222844 158226 222896
rect 158346 222844 158352 222896
rect 158404 222884 158410 222896
rect 165522 222884 165528 222896
rect 158404 222856 165528 222884
rect 158404 222844 158410 222856
rect 165522 222844 165528 222856
rect 165580 222844 165586 222896
rect 165706 222844 165712 222896
rect 165764 222884 165770 222896
rect 215202 222884 215208 222896
rect 165764 222856 215208 222884
rect 165764 222844 165770 222856
rect 215202 222844 215208 222856
rect 215260 222844 215266 222896
rect 218054 222844 218060 222896
rect 218112 222884 218118 222896
rect 257338 222884 257344 222896
rect 218112 222856 257344 222884
rect 218112 222844 218118 222856
rect 257338 222844 257344 222856
rect 257396 222844 257402 222896
rect 257982 222844 257988 222896
rect 258040 222884 258046 222896
rect 283834 222884 283840 222896
rect 258040 222856 283840 222884
rect 258040 222844 258046 222856
rect 283834 222844 283840 222856
rect 283892 222844 283898 222896
rect 284018 222844 284024 222896
rect 284076 222884 284082 222896
rect 300486 222884 300492 222896
rect 284076 222856 300492 222884
rect 284076 222844 284082 222856
rect 300486 222844 300492 222856
rect 300544 222844 300550 222896
rect 303522 222844 303528 222896
rect 303580 222884 303586 222896
rect 311986 222884 311992 222896
rect 303580 222856 311992 222884
rect 303580 222844 303586 222856
rect 311986 222844 311992 222856
rect 312044 222844 312050 222896
rect 314378 222844 314384 222896
rect 314436 222884 314442 222896
rect 320082 222884 320088 222896
rect 314436 222856 320088 222884
rect 314436 222844 314442 222856
rect 320082 222844 320088 222856
rect 320140 222844 320146 222896
rect 342898 222844 342904 222896
rect 342956 222884 342962 222896
rect 349246 222884 349252 222896
rect 342956 222856 349252 222884
rect 342956 222844 342962 222856
rect 349246 222844 349252 222856
rect 349304 222844 349310 222896
rect 355962 222844 355968 222896
rect 356020 222884 356026 222896
rect 367370 222884 367376 222896
rect 356020 222856 367376 222884
rect 356020 222844 356026 222856
rect 367370 222844 367376 222856
rect 367428 222844 367434 222896
rect 371050 222844 371056 222896
rect 371108 222884 371114 222896
rect 390922 222884 390928 222896
rect 371108 222856 390928 222884
rect 371108 222844 371114 222856
rect 390922 222844 390928 222856
rect 390980 222844 390986 222896
rect 405274 222844 405280 222896
rect 405332 222884 405338 222896
rect 439406 222884 439412 222896
rect 405332 222856 439412 222884
rect 405332 222844 405338 222856
rect 439406 222844 439412 222856
rect 439464 222844 439470 222896
rect 439866 222844 439872 222896
rect 439924 222884 439930 222896
rect 485866 222884 485872 222896
rect 439924 222856 485872 222884
rect 439924 222844 439930 222856
rect 485866 222844 485872 222856
rect 485924 222844 485930 222896
rect 488902 222776 488908 222828
rect 488960 222816 488966 222828
rect 490926 222816 490932 222828
rect 488960 222788 490932 222816
rect 488960 222776 488966 222788
rect 490926 222776 490932 222788
rect 490984 222776 490990 222828
rect 114462 222708 114468 222760
rect 114520 222748 114526 222760
rect 185026 222748 185032 222760
rect 114520 222720 185032 222748
rect 114520 222708 114526 222720
rect 185026 222708 185032 222720
rect 185084 222708 185090 222760
rect 185762 222748 185768 222760
rect 185412 222720 185768 222748
rect 102134 222572 102140 222624
rect 102192 222612 102198 222624
rect 152274 222612 152280 222624
rect 102192 222584 152280 222612
rect 102192 222572 102198 222584
rect 152274 222572 152280 222584
rect 152332 222572 152338 222624
rect 152458 222572 152464 222624
rect 152516 222612 152522 222624
rect 173526 222612 173532 222624
rect 152516 222584 173532 222612
rect 152516 222572 152522 222584
rect 173526 222572 173532 222584
rect 173584 222572 173590 222624
rect 175182 222572 175188 222624
rect 175240 222612 175246 222624
rect 185412 222612 185440 222720
rect 185762 222708 185768 222720
rect 185820 222708 185826 222760
rect 191558 222708 191564 222760
rect 191616 222748 191622 222760
rect 239674 222748 239680 222760
rect 191616 222720 239680 222748
rect 191616 222708 191622 222720
rect 239674 222708 239680 222720
rect 239732 222708 239738 222760
rect 391750 222708 391756 222760
rect 391808 222748 391814 222760
rect 412910 222748 412916 222760
rect 391808 222720 412916 222748
rect 391808 222708 391814 222720
rect 412910 222708 412916 222720
rect 412968 222708 412974 222760
rect 413186 222708 413192 222760
rect 413244 222748 413250 222760
rect 429470 222748 429476 222760
rect 413244 222720 429476 222748
rect 413244 222708 413250 222720
rect 429470 222708 429476 222720
rect 429528 222708 429534 222760
rect 442074 222708 442080 222760
rect 442132 222748 442138 222760
rect 486418 222748 486424 222760
rect 442132 222720 486424 222748
rect 442132 222708 442138 222720
rect 486418 222708 486424 222720
rect 486476 222708 486482 222760
rect 491220 222748 491248 222992
rect 491386 222980 491392 223032
rect 491444 223020 491450 223032
rect 563606 223020 563612 223032
rect 491444 222992 563612 223020
rect 491444 222980 491450 222992
rect 563606 222980 563612 222992
rect 563664 222980 563670 223032
rect 491570 222844 491576 222896
rect 491628 222884 491634 222896
rect 565722 222884 565728 222896
rect 491628 222856 565728 222884
rect 491628 222844 491634 222856
rect 565722 222844 565728 222856
rect 565780 222844 565786 222896
rect 519538 222748 519544 222760
rect 491220 222720 519544 222748
rect 519538 222708 519544 222720
rect 519596 222708 519602 222760
rect 668394 222748 668400 222760
rect 563026 222720 615494 222748
rect 175240 222584 185440 222612
rect 175240 222572 175246 222584
rect 185578 222572 185584 222624
rect 185636 222612 185642 222624
rect 213362 222612 213368 222624
rect 185636 222584 213368 222612
rect 185636 222572 185642 222584
rect 213362 222572 213368 222584
rect 213420 222572 213426 222624
rect 213730 222572 213736 222624
rect 213788 222612 213794 222624
rect 252094 222612 252100 222624
rect 213788 222584 252100 222612
rect 213788 222572 213794 222584
rect 252094 222572 252100 222584
rect 252152 222572 252158 222624
rect 299750 222572 299756 222624
rect 299808 222612 299814 222624
rect 306466 222612 306472 222624
rect 299808 222584 306472 222612
rect 299808 222572 299814 222584
rect 306466 222572 306472 222584
rect 306524 222572 306530 222624
rect 390002 222572 390008 222624
rect 390060 222612 390066 222624
rect 406286 222612 406292 222624
rect 390060 222584 406292 222612
rect 390060 222572 390066 222584
rect 406286 222572 406292 222584
rect 406344 222572 406350 222624
rect 406930 222572 406936 222624
rect 406988 222612 406994 222624
rect 423766 222612 423772 222624
rect 406988 222584 423772 222612
rect 406988 222572 406994 222584
rect 423766 222572 423772 222584
rect 423824 222572 423830 222624
rect 448330 222572 448336 222624
rect 448388 222612 448394 222624
rect 499482 222612 499488 222624
rect 448388 222584 499488 222612
rect 448388 222572 448394 222584
rect 499482 222572 499488 222584
rect 499540 222572 499546 222624
rect 499666 222572 499672 222624
rect 499724 222612 499730 222624
rect 500862 222612 500868 222624
rect 499724 222584 500868 222612
rect 499724 222572 499730 222584
rect 500862 222572 500868 222584
rect 500920 222572 500926 222624
rect 501046 222572 501052 222624
rect 501104 222612 501110 222624
rect 503438 222612 503444 222624
rect 501104 222584 503444 222612
rect 501104 222572 501110 222584
rect 503438 222572 503444 222584
rect 503496 222572 503502 222624
rect 505186 222572 505192 222624
rect 505244 222612 505250 222624
rect 514018 222612 514024 222624
rect 505244 222584 514024 222612
rect 505244 222572 505250 222584
rect 514018 222572 514024 222584
rect 514076 222572 514082 222624
rect 554774 222572 554780 222624
rect 554832 222612 554838 222624
rect 555418 222612 555424 222624
rect 554832 222584 555424 222612
rect 554832 222572 554838 222584
rect 555418 222572 555424 222584
rect 555476 222572 555482 222624
rect 557350 222572 557356 222624
rect 557408 222612 557414 222624
rect 563026 222612 563054 222720
rect 557408 222584 563054 222612
rect 557408 222572 557414 222584
rect 565722 222572 565728 222624
rect 565780 222612 565786 222624
rect 611354 222612 611360 222624
rect 565780 222584 611360 222612
rect 565780 222572 565786 222584
rect 611354 222572 611360 222584
rect 611412 222572 611418 222624
rect 615466 222612 615494 222720
rect 663766 222720 668400 222748
rect 626534 222612 626540 222624
rect 615466 222584 626540 222612
rect 626534 222572 626540 222584
rect 626592 222572 626598 222624
rect 661678 222572 661684 222624
rect 661736 222612 661742 222624
rect 663766 222612 663794 222720
rect 668394 222708 668400 222720
rect 668452 222708 668458 222760
rect 675110 222680 675116 222692
rect 673472 222652 675116 222680
rect 673472 222612 673500 222652
rect 675110 222640 675116 222652
rect 675168 222640 675174 222692
rect 661736 222584 663794 222612
rect 667124 222584 673500 222612
rect 661736 222572 661742 222584
rect 101490 222436 101496 222488
rect 101548 222476 101554 222488
rect 101548 222448 122834 222476
rect 101548 222436 101554 222448
rect 122806 222340 122834 222448
rect 125318 222436 125324 222488
rect 125376 222476 125382 222488
rect 125376 222448 194824 222476
rect 125376 222436 125382 222448
rect 142108 222340 142114 222352
rect 122806 222312 142114 222340
rect 142108 222300 142114 222312
rect 142166 222300 142172 222352
rect 142614 222300 142620 222352
rect 142672 222340 142678 222352
rect 194594 222340 194600 222352
rect 142672 222312 194600 222340
rect 142672 222300 142678 222312
rect 194594 222300 194600 222312
rect 194652 222300 194658 222352
rect 194796 222340 194824 222448
rect 194962 222436 194968 222488
rect 195020 222476 195026 222488
rect 195020 222448 203656 222476
rect 195020 222436 195026 222448
rect 195606 222340 195612 222352
rect 194796 222312 195612 222340
rect 195606 222300 195612 222312
rect 195664 222300 195670 222352
rect 203628 222340 203656 222448
rect 207198 222436 207204 222488
rect 207256 222476 207262 222488
rect 215938 222476 215944 222488
rect 207256 222448 215944 222476
rect 207256 222436 207262 222448
rect 215938 222436 215944 222448
rect 215996 222436 216002 222488
rect 220630 222436 220636 222488
rect 220688 222476 220694 222488
rect 256786 222476 256792 222488
rect 220688 222448 256792 222476
rect 220688 222436 220694 222448
rect 256786 222436 256792 222448
rect 256844 222436 256850 222488
rect 389082 222436 389088 222488
rect 389140 222476 389146 222488
rect 403158 222476 403164 222488
rect 389140 222448 403164 222476
rect 389140 222436 389146 222448
rect 403158 222436 403164 222448
rect 403216 222436 403222 222488
rect 411714 222436 411720 222488
rect 411772 222476 411778 222488
rect 428090 222476 428096 222488
rect 411772 222448 428096 222476
rect 411772 222436 411778 222448
rect 428090 222436 428096 222448
rect 428148 222436 428154 222488
rect 450078 222436 450084 222488
rect 450136 222476 450142 222488
rect 505002 222476 505008 222488
rect 450136 222448 505008 222476
rect 450136 222436 450142 222448
rect 505002 222436 505008 222448
rect 505060 222436 505066 222488
rect 505186 222436 505192 222488
rect 505244 222476 505250 222488
rect 510706 222476 510712 222488
rect 505244 222448 510712 222476
rect 505244 222436 505250 222448
rect 510706 222436 510712 222448
rect 510764 222436 510770 222488
rect 555418 222436 555424 222488
rect 555476 222476 555482 222488
rect 608594 222476 608600 222488
rect 555476 222448 608600 222476
rect 555476 222436 555482 222448
rect 608594 222436 608600 222448
rect 608652 222436 608658 222488
rect 663058 222436 663064 222488
rect 663116 222476 663122 222488
rect 667124 222476 667152 222584
rect 675478 222544 675484 222556
rect 673564 222516 675484 222544
rect 663116 222448 667152 222476
rect 663116 222436 663122 222448
rect 668394 222436 668400 222488
rect 668452 222476 668458 222488
rect 673564 222476 673592 222516
rect 675478 222504 675484 222516
rect 675536 222504 675542 222556
rect 668452 222448 673592 222476
rect 668452 222436 668458 222448
rect 438394 222368 438400 222420
rect 438452 222408 438458 222420
rect 442902 222408 442908 222420
rect 438452 222380 442908 222408
rect 438452 222368 438458 222380
rect 442902 222368 442908 222380
rect 442960 222368 442966 222420
rect 523126 222368 523132 222420
rect 523184 222408 523190 222420
rect 523678 222408 523684 222420
rect 523184 222380 523684 222408
rect 523184 222368 523190 222380
rect 523678 222368 523684 222380
rect 523736 222408 523742 222420
rect 675294 222408 675300 222420
rect 523736 222380 534074 222408
rect 523736 222368 523742 222380
rect 207382 222340 207388 222352
rect 203628 222312 207388 222340
rect 207382 222300 207388 222312
rect 207440 222300 207446 222352
rect 214558 222300 214564 222352
rect 214616 222340 214622 222352
rect 221734 222340 221740 222352
rect 214616 222312 221740 222340
rect 214616 222300 214622 222312
rect 221734 222300 221740 222312
rect 221792 222300 221798 222352
rect 420914 222300 420920 222352
rect 420972 222340 420978 222352
rect 432782 222340 432788 222352
rect 420972 222312 432788 222340
rect 420972 222300 420978 222312
rect 432782 222300 432788 222312
rect 432840 222300 432846 222352
rect 444834 222300 444840 222352
rect 444892 222340 444898 222352
rect 503162 222340 503168 222352
rect 444892 222312 503168 222340
rect 444892 222300 444898 222312
rect 503162 222300 503168 222312
rect 503220 222300 503226 222352
rect 503438 222300 503444 222352
rect 503496 222340 503502 222352
rect 508498 222340 508504 222352
rect 503496 222312 508504 222340
rect 503496 222300 503502 222312
rect 508498 222300 508504 222312
rect 508556 222300 508562 222352
rect 201586 222272 201592 222284
rect 201052 222244 201592 222272
rect 181162 222204 181168 222216
rect 180766 222176 181168 222204
rect 119706 222096 119712 222148
rect 119764 222136 119770 222148
rect 180766 222136 180794 222176
rect 181162 222164 181168 222176
rect 181220 222164 181226 222216
rect 119764 222108 180794 222136
rect 119764 222096 119770 222108
rect 181438 222096 181444 222148
rect 181496 222136 181502 222148
rect 183462 222136 183468 222148
rect 181496 222108 183468 222136
rect 181496 222096 181502 222108
rect 183462 222096 183468 222108
rect 183520 222096 183526 222148
rect 184290 222096 184296 222148
rect 184348 222136 184354 222148
rect 184348 222108 185992 222136
rect 184348 222096 184354 222108
rect 116394 221960 116400 222012
rect 116452 222000 116458 222012
rect 181990 222000 181996 222012
rect 116452 221972 181996 222000
rect 116452 221960 116458 221972
rect 181990 221960 181996 221972
rect 182048 221960 182054 222012
rect 182174 221960 182180 222012
rect 182232 222000 182238 222012
rect 185762 222000 185768 222012
rect 182232 221972 185768 222000
rect 182232 221960 182238 221972
rect 185762 221960 185768 221972
rect 185820 221960 185826 222012
rect 185964 222000 185992 222108
rect 188982 222096 188988 222148
rect 189040 222136 189046 222148
rect 189040 222108 192708 222136
rect 189040 222096 189046 222108
rect 192478 222000 192484 222012
rect 185964 221972 192484 222000
rect 192478 221960 192484 221972
rect 192536 221960 192542 222012
rect 80790 221824 80796 221876
rect 80848 221864 80854 221876
rect 111058 221864 111064 221876
rect 80848 221836 111064 221864
rect 80848 221824 80854 221836
rect 111058 221824 111064 221836
rect 111116 221824 111122 221876
rect 111426 221824 111432 221876
rect 111484 221864 111490 221876
rect 183830 221864 183836 221876
rect 111484 221836 183836 221864
rect 111484 221824 111490 221836
rect 183830 221824 183836 221836
rect 183888 221824 183894 221876
rect 185578 221824 185584 221876
rect 185636 221864 185642 221876
rect 191926 221864 191932 221876
rect 185636 221836 191932 221864
rect 185636 221824 185642 221836
rect 191926 221824 191932 221836
rect 191984 221824 191990 221876
rect 192680 221864 192708 222108
rect 195146 222096 195152 222148
rect 195204 222136 195210 222148
rect 201052 222136 201080 222244
rect 201586 222232 201592 222244
rect 201644 222232 201650 222284
rect 519722 222272 519728 222284
rect 519372 222244 519728 222272
rect 195204 222108 201080 222136
rect 195204 222096 195210 222108
rect 201218 222096 201224 222148
rect 201276 222136 201282 222148
rect 245930 222136 245936 222148
rect 201276 222108 245936 222136
rect 201276 222096 201282 222108
rect 245930 222096 245936 222108
rect 245988 222096 245994 222148
rect 248138 222096 248144 222148
rect 248196 222136 248202 222148
rect 251266 222136 251272 222148
rect 248196 222108 251272 222136
rect 248196 222096 248202 222108
rect 251266 222096 251272 222108
rect 251324 222096 251330 222148
rect 261662 222096 261668 222148
rect 261720 222136 261726 222148
rect 265250 222136 265256 222148
rect 261720 222108 265256 222136
rect 261720 222096 261726 222108
rect 265250 222096 265256 222108
rect 265308 222096 265314 222148
rect 266262 222096 266268 222148
rect 266320 222136 266326 222148
rect 266998 222136 267004 222148
rect 266320 222108 267004 222136
rect 266320 222096 266326 222108
rect 266998 222096 267004 222108
rect 267056 222096 267062 222148
rect 267182 222096 267188 222148
rect 267240 222136 267246 222148
rect 284570 222136 284576 222148
rect 267240 222108 284576 222136
rect 267240 222096 267246 222108
rect 284570 222096 284576 222108
rect 284628 222096 284634 222148
rect 347130 222096 347136 222148
rect 347188 222136 347194 222148
rect 354214 222136 354220 222148
rect 347188 222108 354220 222136
rect 347188 222096 347194 222108
rect 354214 222096 354220 222108
rect 354272 222096 354278 222148
rect 381906 222096 381912 222148
rect 381964 222136 381970 222148
rect 388438 222136 388444 222148
rect 381964 222108 388444 222136
rect 381964 222096 381970 222108
rect 388438 222096 388444 222108
rect 388496 222096 388502 222148
rect 402698 222096 402704 222148
rect 402756 222136 402762 222148
rect 438854 222136 438860 222148
rect 402756 222108 438860 222136
rect 402756 222096 402762 222108
rect 438854 222096 438860 222108
rect 438912 222096 438918 222148
rect 446858 222096 446864 222148
rect 446916 222136 446922 222148
rect 499574 222136 499580 222148
rect 446916 222108 499580 222136
rect 446916 222096 446922 222108
rect 499574 222096 499580 222108
rect 499632 222096 499638 222148
rect 499758 222096 499764 222148
rect 499816 222136 499822 222148
rect 519372 222136 519400 222244
rect 519722 222232 519728 222244
rect 519780 222232 519786 222284
rect 534046 222204 534074 222380
rect 673656 222380 675300 222408
rect 547414 222300 547420 222352
rect 547472 222340 547478 222352
rect 623958 222340 623964 222352
rect 547472 222312 623964 222340
rect 547472 222300 547478 222312
rect 623958 222300 623964 222312
rect 624016 222300 624022 222352
rect 664622 222300 664628 222352
rect 664680 222340 664686 222352
rect 673656 222340 673684 222380
rect 675294 222368 675300 222380
rect 675352 222368 675358 222420
rect 664680 222312 673684 222340
rect 664680 222300 664686 222312
rect 675478 222272 675484 222284
rect 673748 222244 675484 222272
rect 601694 222204 601700 222216
rect 534046 222176 601700 222204
rect 601694 222164 601700 222176
rect 601752 222164 601758 222216
rect 664438 222164 664444 222216
rect 664496 222204 664502 222216
rect 664496 222176 673500 222204
rect 664496 222164 664502 222176
rect 499816 222108 519400 222136
rect 499816 222096 499822 222108
rect 519538 222096 519544 222148
rect 519596 222136 519602 222148
rect 530762 222136 530768 222148
rect 519596 222108 530768 222136
rect 519596 222096 519602 222108
rect 530762 222096 530768 222108
rect 530820 222096 530826 222148
rect 673472 222136 673500 222176
rect 673748 222136 673776 222244
rect 675478 222232 675484 222244
rect 675536 222232 675542 222284
rect 673472 222108 673776 222136
rect 192846 222028 192852 222080
rect 192904 222068 192910 222080
rect 194226 222068 194232 222080
rect 192904 222040 194232 222068
rect 192904 222028 192910 222040
rect 194226 222028 194232 222040
rect 194284 222028 194290 222080
rect 246390 222028 246396 222080
rect 246448 222068 246454 222080
rect 247770 222068 247776 222080
rect 246448 222040 247776 222068
rect 246448 222028 246454 222040
rect 247770 222028 247776 222040
rect 247828 222028 247834 222080
rect 194410 221960 194416 222012
rect 194468 222000 194474 222012
rect 238938 222000 238944 222012
rect 194468 221972 238944 222000
rect 194468 221960 194474 221972
rect 238938 221960 238944 221972
rect 238996 221960 239002 222012
rect 247954 221960 247960 222012
rect 248012 222000 248018 222012
rect 274726 222000 274732 222012
rect 248012 221972 274732 222000
rect 248012 221960 248018 221972
rect 274726 221960 274732 221972
rect 274784 221960 274790 222012
rect 288986 222000 288992 222012
rect 277366 221972 288992 222000
rect 237466 221864 237472 221876
rect 192680 221836 237472 221864
rect 237466 221824 237472 221836
rect 237524 221824 237530 221876
rect 243906 221824 243912 221876
rect 243964 221864 243970 221876
rect 272058 221864 272064 221876
rect 243964 221836 272064 221864
rect 243964 221824 243970 221836
rect 272058 221824 272064 221836
rect 272116 221824 272122 221876
rect 97718 221688 97724 221740
rect 97776 221728 97782 221740
rect 171042 221728 171048 221740
rect 97776 221700 171048 221728
rect 97776 221688 97782 221700
rect 171042 221688 171048 221700
rect 171100 221688 171106 221740
rect 171226 221688 171232 221740
rect 171284 221728 171290 221740
rect 181254 221728 181260 221740
rect 171284 221700 181260 221728
rect 171284 221688 171290 221700
rect 181254 221688 181260 221700
rect 181312 221688 181318 221740
rect 181438 221688 181444 221740
rect 181496 221728 181502 221740
rect 225506 221728 225512 221740
rect 181496 221700 225512 221728
rect 181496 221688 181502 221700
rect 225506 221688 225512 221700
rect 225564 221688 225570 221740
rect 231854 221688 231860 221740
rect 231912 221728 231918 221740
rect 233418 221728 233424 221740
rect 231912 221700 233424 221728
rect 231912 221688 231918 221700
rect 233418 221688 233424 221700
rect 233476 221688 233482 221740
rect 233694 221688 233700 221740
rect 233752 221728 233758 221740
rect 261662 221728 261668 221740
rect 233752 221700 261668 221728
rect 233752 221688 233758 221700
rect 261662 221688 261668 221700
rect 261720 221688 261726 221740
rect 261938 221688 261944 221740
rect 261996 221728 262002 221740
rect 267182 221728 267188 221740
rect 261996 221700 267188 221728
rect 261996 221688 262002 221700
rect 267182 221688 267188 221700
rect 267240 221688 267246 221740
rect 59814 221552 59820 221604
rect 59872 221592 59878 221604
rect 144362 221592 144368 221604
rect 59872 221564 144368 221592
rect 59872 221552 59878 221564
rect 144362 221552 144368 221564
rect 144420 221552 144426 221604
rect 144546 221552 144552 221604
rect 144604 221592 144610 221604
rect 200068 221592 200074 221604
rect 144604 221564 200074 221592
rect 144604 221552 144610 221564
rect 200068 221552 200074 221564
rect 200126 221552 200132 221604
rect 200298 221552 200304 221604
rect 200356 221592 200362 221604
rect 202322 221592 202328 221604
rect 200356 221564 202328 221592
rect 200356 221552 200362 221564
rect 202322 221552 202328 221564
rect 202380 221552 202386 221604
rect 204714 221552 204720 221604
rect 204772 221592 204778 221604
rect 227898 221592 227904 221604
rect 204772 221564 227904 221592
rect 204772 221552 204778 221564
rect 227898 221552 227904 221564
rect 227956 221552 227962 221604
rect 230382 221552 230388 221604
rect 230440 221592 230446 221604
rect 263134 221592 263140 221604
rect 230440 221564 263140 221592
rect 230440 221552 230446 221564
rect 263134 221552 263140 221564
rect 263192 221552 263198 221604
rect 268746 221552 268752 221604
rect 268804 221592 268810 221604
rect 277366 221592 277394 221972
rect 288986 221960 288992 221972
rect 289044 221960 289050 222012
rect 388622 221960 388628 222012
rect 388680 222000 388686 222012
rect 412174 222000 412180 222012
rect 388680 221972 412180 222000
rect 388680 221960 388686 221972
rect 412174 221960 412180 221972
rect 412232 221960 412238 222012
rect 417786 221960 417792 222012
rect 417844 222000 417850 222012
rect 461854 222000 461860 222012
rect 417844 221972 461860 222000
rect 417844 221960 417850 221972
rect 461854 221960 461860 221972
rect 461912 221960 461918 222012
rect 473170 221960 473176 222012
rect 473228 222000 473234 222012
rect 545758 222000 545764 222012
rect 473228 221972 545764 222000
rect 473228 221960 473234 221972
rect 545758 221960 545764 221972
rect 545816 221960 545822 222012
rect 549898 221960 549904 222012
rect 549956 222000 549962 222012
rect 560570 222000 560576 222012
rect 549956 221972 560576 222000
rect 549956 221960 549962 221972
rect 560570 221960 560576 221972
rect 560628 221960 560634 222012
rect 285306 221824 285312 221876
rect 285364 221864 285370 221876
rect 300118 221864 300124 221876
rect 285364 221836 300124 221864
rect 285364 221824 285370 221836
rect 300118 221824 300124 221836
rect 300176 221824 300182 221876
rect 362586 221824 362592 221876
rect 362644 221864 362650 221876
rect 377398 221864 377404 221876
rect 362644 221836 377404 221864
rect 362644 221824 362650 221836
rect 377398 221824 377404 221836
rect 377456 221824 377462 221876
rect 379146 221824 379152 221876
rect 379204 221864 379210 221876
rect 402238 221864 402244 221876
rect 379204 221836 402244 221864
rect 379204 221824 379210 221836
rect 402238 221824 402244 221836
rect 402296 221824 402302 221876
rect 409598 221824 409604 221876
rect 409656 221864 409662 221876
rect 448606 221864 448612 221876
rect 409656 221836 448612 221864
rect 409656 221824 409662 221836
rect 448606 221824 448612 221836
rect 448664 221824 448670 221876
rect 477402 221824 477408 221876
rect 477460 221864 477466 221876
rect 550634 221864 550640 221876
rect 477460 221836 550640 221864
rect 477460 221824 477466 221836
rect 550634 221824 550640 221836
rect 550692 221824 550698 221876
rect 558178 221824 558184 221876
rect 558236 221864 558242 221876
rect 564710 221864 564716 221876
rect 558236 221836 564716 221864
rect 558236 221824 558242 221836
rect 564710 221824 564716 221836
rect 564768 221824 564774 221876
rect 280062 221688 280068 221740
rect 280120 221728 280126 221740
rect 296162 221728 296168 221740
rect 280120 221700 296168 221728
rect 280120 221688 280126 221700
rect 296162 221688 296168 221700
rect 296220 221688 296226 221740
rect 300118 221688 300124 221740
rect 300176 221728 300182 221740
rect 309502 221728 309508 221740
rect 300176 221700 309508 221728
rect 300176 221688 300182 221700
rect 309502 221688 309508 221700
rect 309560 221688 309566 221740
rect 310054 221688 310060 221740
rect 310112 221728 310118 221740
rect 316126 221728 316132 221740
rect 310112 221700 316132 221728
rect 310112 221688 310118 221700
rect 316126 221688 316132 221700
rect 316184 221688 316190 221740
rect 343542 221688 343548 221740
rect 343600 221728 343606 221740
rect 347866 221728 347872 221740
rect 343600 221700 347872 221728
rect 343600 221688 343606 221700
rect 347866 221688 347872 221700
rect 347924 221688 347930 221740
rect 351730 221688 351736 221740
rect 351788 221728 351794 221740
rect 362494 221728 362500 221740
rect 351788 221700 362500 221728
rect 351788 221688 351794 221700
rect 362494 221688 362500 221700
rect 362552 221688 362558 221740
rect 371878 221688 371884 221740
rect 371936 221728 371942 221740
rect 389174 221728 389180 221740
rect 371936 221700 389180 221728
rect 371936 221688 371942 221700
rect 389174 221688 389180 221700
rect 389232 221688 389238 221740
rect 390462 221688 390468 221740
rect 390520 221728 390526 221740
rect 418798 221728 418804 221740
rect 390520 221700 418804 221728
rect 390520 221688 390526 221700
rect 418798 221688 418804 221700
rect 418856 221688 418862 221740
rect 422202 221688 422208 221740
rect 422260 221728 422266 221740
rect 464338 221728 464344 221740
rect 422260 221700 464344 221728
rect 422260 221688 422266 221700
rect 464338 221688 464344 221700
rect 464396 221688 464402 221740
rect 475930 221688 475936 221740
rect 475988 221728 475994 221740
rect 549990 221728 549996 221740
rect 475988 221700 549996 221728
rect 475988 221688 475994 221700
rect 549990 221688 549996 221700
rect 550048 221688 550054 221740
rect 565078 221688 565084 221740
rect 565136 221728 565142 221740
rect 567378 221728 567384 221740
rect 565136 221700 567384 221728
rect 565136 221688 565142 221700
rect 567378 221688 567384 221700
rect 567436 221728 567442 221740
rect 567436 221700 576854 221728
rect 567436 221688 567442 221700
rect 268804 221564 277394 221592
rect 268804 221552 268810 221564
rect 288618 221552 288624 221604
rect 288676 221592 288682 221604
rect 303706 221592 303712 221604
rect 288676 221564 303712 221592
rect 288676 221552 288682 221564
rect 303706 221552 303712 221564
rect 303764 221552 303770 221604
rect 315114 221552 315120 221604
rect 315172 221592 315178 221604
rect 319438 221592 319444 221604
rect 315172 221564 319444 221592
rect 315172 221552 315178 221564
rect 319438 221552 319444 221564
rect 319496 221552 319502 221604
rect 344830 221552 344836 221604
rect 344888 221592 344894 221604
rect 350902 221592 350908 221604
rect 344888 221564 350908 221592
rect 344888 221552 344894 221564
rect 350902 221552 350908 221564
rect 350960 221552 350966 221604
rect 354582 221552 354588 221604
rect 354640 221592 354646 221604
rect 364334 221592 364340 221604
rect 354640 221564 364340 221592
rect 354640 221552 354646 221564
rect 364334 221552 364340 221564
rect 364392 221552 364398 221604
rect 365622 221552 365628 221604
rect 365680 221592 365686 221604
rect 380894 221592 380900 221604
rect 365680 221564 380900 221592
rect 365680 221552 365686 221564
rect 380894 221552 380900 221564
rect 380952 221552 380958 221604
rect 387518 221552 387524 221604
rect 387576 221592 387582 221604
rect 415578 221592 415584 221604
rect 387576 221564 415584 221592
rect 387576 221552 387582 221564
rect 415578 221552 415584 221564
rect 415636 221552 415642 221604
rect 445662 221552 445668 221604
rect 445720 221592 445726 221604
rect 475378 221592 475384 221604
rect 445720 221564 475384 221592
rect 445720 221552 445726 221564
rect 475378 221552 475384 221564
rect 475436 221552 475442 221604
rect 477862 221552 477868 221604
rect 477920 221592 477926 221604
rect 477920 221564 553394 221592
rect 477920 221552 477926 221564
rect 70026 221416 70032 221468
rect 70084 221456 70090 221468
rect 151630 221456 151636 221468
rect 70084 221428 151636 221456
rect 70084 221416 70090 221428
rect 151630 221416 151636 221428
rect 151688 221416 151694 221468
rect 151814 221416 151820 221468
rect 151872 221456 151878 221468
rect 159818 221456 159824 221468
rect 151872 221428 159824 221456
rect 151872 221416 151878 221428
rect 159818 221416 159824 221428
rect 159876 221416 159882 221468
rect 160002 221416 160008 221468
rect 160060 221456 160066 221468
rect 160738 221456 160744 221468
rect 160060 221428 160744 221456
rect 160060 221416 160066 221428
rect 160738 221416 160744 221428
rect 160796 221416 160802 221468
rect 160922 221416 160928 221468
rect 160980 221456 160986 221468
rect 166810 221456 166816 221468
rect 160980 221428 166816 221456
rect 160980 221416 160986 221428
rect 166810 221416 166816 221428
rect 166868 221416 166874 221468
rect 166948 221416 166954 221468
rect 167006 221456 167012 221468
rect 213270 221456 213276 221468
rect 167006 221428 213276 221456
rect 167006 221416 167012 221428
rect 213270 221416 213276 221428
rect 213328 221416 213334 221468
rect 232130 221456 232136 221468
rect 214576 221428 232136 221456
rect 122558 221280 122564 221332
rect 122616 221320 122622 221332
rect 185578 221320 185584 221332
rect 122616 221292 185584 221320
rect 122616 221280 122622 221292
rect 185578 221280 185584 221292
rect 185636 221280 185642 221332
rect 185762 221280 185768 221332
rect 185820 221320 185826 221332
rect 204714 221320 204720 221332
rect 185820 221292 204720 221320
rect 185820 221280 185826 221292
rect 204714 221280 204720 221292
rect 204772 221280 204778 221332
rect 214576 221320 214604 221428
rect 232130 221416 232136 221428
rect 232188 221416 232194 221468
rect 240042 221416 240048 221468
rect 240100 221456 240106 221468
rect 270586 221456 270592 221468
rect 240100 221428 270592 221456
rect 240100 221416 240106 221428
rect 270586 221416 270592 221428
rect 270644 221416 270650 221468
rect 271230 221416 271236 221468
rect 271288 221456 271294 221468
rect 292666 221456 292672 221468
rect 271288 221428 292672 221456
rect 271288 221416 271294 221428
rect 292666 221416 292672 221428
rect 292724 221416 292730 221468
rect 298554 221416 298560 221468
rect 298612 221456 298618 221468
rect 309226 221456 309232 221468
rect 298612 221428 309232 221456
rect 298612 221416 298618 221428
rect 309226 221416 309232 221428
rect 309284 221416 309290 221468
rect 316034 221416 316040 221468
rect 316092 221456 316098 221468
rect 321646 221456 321652 221468
rect 316092 221428 321652 221456
rect 316092 221416 316098 221428
rect 321646 221416 321652 221428
rect 321704 221416 321710 221468
rect 358170 221416 358176 221468
rect 358228 221456 358234 221468
rect 370774 221456 370780 221468
rect 358228 221428 370780 221456
rect 358228 221416 358234 221428
rect 370774 221416 370780 221428
rect 370832 221416 370838 221468
rect 374638 221416 374644 221468
rect 374696 221456 374702 221468
rect 395614 221456 395620 221468
rect 374696 221428 395620 221456
rect 374696 221416 374702 221428
rect 395614 221416 395620 221428
rect 395672 221416 395678 221468
rect 398558 221416 398564 221468
rect 398616 221456 398622 221468
rect 432046 221456 432052 221468
rect 398616 221428 432052 221456
rect 398616 221416 398622 221428
rect 432046 221416 432052 221428
rect 432104 221416 432110 221468
rect 436002 221416 436008 221468
rect 436060 221456 436066 221468
rect 485728 221456 485734 221468
rect 436060 221428 485734 221456
rect 436060 221416 436066 221428
rect 485728 221416 485734 221428
rect 485786 221416 485792 221468
rect 485866 221416 485872 221468
rect 485924 221456 485930 221468
rect 495250 221456 495256 221468
rect 485924 221428 495256 221456
rect 485924 221416 485930 221428
rect 495250 221416 495256 221428
rect 495308 221416 495314 221468
rect 495388 221416 495394 221468
rect 495446 221456 495452 221468
rect 519538 221456 519544 221468
rect 495446 221428 519544 221456
rect 495446 221416 495452 221428
rect 519538 221416 519544 221428
rect 519596 221416 519602 221468
rect 519722 221416 519728 221468
rect 519780 221456 519786 221468
rect 519780 221428 543734 221456
rect 519780 221416 519786 221428
rect 204916 221292 214604 221320
rect 129458 221144 129464 221196
rect 129516 221184 129522 221196
rect 192294 221184 192300 221196
rect 129516 221156 192300 221184
rect 129516 221144 129522 221156
rect 192294 221144 192300 221156
rect 192352 221144 192358 221196
rect 192478 221144 192484 221196
rect 192536 221184 192542 221196
rect 204916 221184 204944 221292
rect 214742 221280 214748 221332
rect 214800 221320 214806 221332
rect 245746 221320 245752 221332
rect 214800 221292 245752 221320
rect 214800 221280 214806 221292
rect 245746 221280 245752 221292
rect 245804 221280 245810 221332
rect 257154 221280 257160 221332
rect 257212 221320 257218 221332
rect 280706 221320 280712 221332
rect 257212 221292 280712 221320
rect 257212 221280 257218 221292
rect 280706 221280 280712 221292
rect 280764 221280 280770 221332
rect 392578 221280 392584 221332
rect 392636 221320 392642 221332
rect 422294 221320 422300 221332
rect 392636 221292 422300 221320
rect 392636 221280 392642 221292
rect 422294 221280 422300 221292
rect 422352 221280 422358 221332
rect 423214 221280 423220 221332
rect 423272 221320 423278 221332
rect 459554 221320 459560 221332
rect 423272 221292 459560 221320
rect 423272 221280 423278 221292
rect 459554 221280 459560 221292
rect 459612 221280 459618 221332
rect 470226 221280 470232 221332
rect 470284 221320 470290 221332
rect 540514 221320 540520 221332
rect 470284 221292 540520 221320
rect 470284 221280 470290 221292
rect 540514 221280 540520 221292
rect 540572 221280 540578 221332
rect 192536 221156 204944 221184
rect 192536 221144 192542 221156
rect 207474 221144 207480 221196
rect 207532 221184 207538 221196
rect 247586 221184 247592 221196
rect 207532 221156 247592 221184
rect 207532 221144 207538 221156
rect 247586 221144 247592 221156
rect 247644 221144 247650 221196
rect 396718 221144 396724 221196
rect 396776 221184 396782 221196
rect 428734 221184 428740 221196
rect 396776 221156 428740 221184
rect 396776 221144 396782 221156
rect 428734 221144 428740 221156
rect 428792 221144 428798 221196
rect 439590 221144 439596 221196
rect 439648 221184 439654 221196
rect 466822 221184 466828 221196
rect 439648 221156 466828 221184
rect 439648 221144 439654 221156
rect 466822 221144 466828 221156
rect 466880 221144 466886 221196
rect 467742 221144 467748 221196
rect 467800 221184 467806 221196
rect 535546 221184 535552 221196
rect 467800 221156 535552 221184
rect 467800 221144 467806 221156
rect 535546 221144 535552 221156
rect 535604 221144 535610 221196
rect 543706 221184 543734 221428
rect 553366 221332 553394 221564
rect 564710 221552 564716 221604
rect 564768 221592 564774 221604
rect 576826 221592 576854 221700
rect 596726 221688 596732 221740
rect 596784 221728 596790 221740
rect 603442 221728 603448 221740
rect 596784 221700 603448 221728
rect 596784 221688 596790 221700
rect 603442 221688 603448 221700
rect 603500 221688 603506 221740
rect 564768 221564 572714 221592
rect 576826 221564 605834 221592
rect 564768 221552 564774 221564
rect 568574 221416 568580 221468
rect 568632 221456 568638 221468
rect 569494 221456 569500 221468
rect 568632 221428 569500 221456
rect 568632 221416 568638 221428
rect 569494 221416 569500 221428
rect 569552 221416 569558 221468
rect 572686 221456 572714 221564
rect 605806 221456 605834 221564
rect 620278 221456 620284 221468
rect 572686 221428 598796 221456
rect 605806 221428 620284 221456
rect 553302 221280 553308 221332
rect 553360 221320 553394 221332
rect 553360 221292 558224 221320
rect 553360 221280 553366 221292
rect 557994 221184 558000 221196
rect 543706 221156 558000 221184
rect 557994 221144 558000 221156
rect 558052 221144 558058 221196
rect 558196 221184 558224 221292
rect 558362 221280 558368 221332
rect 558420 221320 558426 221332
rect 597094 221320 597100 221332
rect 558420 221292 597100 221320
rect 558420 221280 558426 221292
rect 597094 221280 597100 221292
rect 597152 221280 597158 221332
rect 598768 221320 598796 221428
rect 620278 221416 620284 221428
rect 620336 221416 620342 221468
rect 628190 221320 628196 221332
rect 598768 221292 628196 221320
rect 628190 221280 628196 221292
rect 628248 221280 628254 221332
rect 608962 221184 608968 221196
rect 558196 221156 608968 221184
rect 608962 221144 608968 221156
rect 609020 221144 609026 221196
rect 620278 221144 620284 221196
rect 620336 221184 620342 221196
rect 628006 221184 628012 221196
rect 620336 221156 628012 221184
rect 620336 221144 620342 221156
rect 628006 221144 628012 221156
rect 628064 221144 628070 221196
rect 664254 221076 664260 221128
rect 664312 221116 664318 221128
rect 675478 221116 675484 221128
rect 664312 221088 675484 221116
rect 664312 221076 664318 221088
rect 675478 221076 675484 221088
rect 675536 221076 675542 221128
rect 139118 221008 139124 221060
rect 139176 221048 139182 221060
rect 171042 221048 171048 221060
rect 139176 221020 171048 221048
rect 139176 221008 139182 221020
rect 171042 221008 171048 221020
rect 171100 221008 171106 221060
rect 171226 221008 171232 221060
rect 171284 221048 171290 221060
rect 210142 221048 210148 221060
rect 171284 221020 210148 221048
rect 171284 221008 171290 221020
rect 210142 221008 210148 221020
rect 210200 221008 210206 221060
rect 213270 221008 213276 221060
rect 213328 221048 213334 221060
rect 216858 221048 216864 221060
rect 213328 221020 216864 221048
rect 213328 221008 213334 221020
rect 216858 221008 216864 221020
rect 216916 221008 216922 221060
rect 217410 221008 217416 221060
rect 217468 221048 217474 221060
rect 254302 221048 254308 221060
rect 217468 221020 254308 221048
rect 217468 221008 217474 221020
rect 254302 221008 254308 221020
rect 254360 221008 254366 221060
rect 416038 221008 416044 221060
rect 416096 221048 416102 221060
rect 441982 221048 441988 221060
rect 416096 221020 441988 221048
rect 416096 221008 416102 221020
rect 441982 221008 441988 221020
rect 442040 221008 442046 221060
rect 459922 221008 459928 221060
rect 459980 221048 459986 221060
rect 526162 221048 526168 221060
rect 459980 221020 526168 221048
rect 459980 221008 459986 221020
rect 526162 221008 526168 221020
rect 526220 221048 526226 221060
rect 526220 221020 596956 221048
rect 526220 221008 526226 221020
rect 126146 220872 126152 220924
rect 126204 220912 126210 220924
rect 127066 220912 127072 220924
rect 126204 220884 127072 220912
rect 126204 220872 126210 220884
rect 127066 220872 127072 220884
rect 127124 220872 127130 220924
rect 137922 220872 137928 220924
rect 137980 220912 137986 220924
rect 195146 220912 195152 220924
rect 137980 220884 195152 220912
rect 137980 220872 137986 220884
rect 195146 220872 195152 220884
rect 195204 220872 195210 220924
rect 195330 220872 195336 220924
rect 195388 220912 195394 220924
rect 199470 220912 199476 220924
rect 195388 220884 199476 220912
rect 195388 220872 195394 220884
rect 199470 220872 199476 220884
rect 199528 220872 199534 220924
rect 204162 220872 204168 220924
rect 204220 220912 204226 220924
rect 214742 220912 214748 220924
rect 204220 220884 214748 220912
rect 204220 220872 204226 220884
rect 214742 220872 214748 220884
rect 214800 220872 214806 220924
rect 277578 220912 277584 220924
rect 274652 220884 277584 220912
rect 63954 220804 63960 220856
rect 64012 220844 64018 220856
rect 66898 220844 66904 220856
rect 64012 220816 66904 220844
rect 64012 220804 64018 220816
rect 66898 220804 66904 220816
rect 66956 220804 66962 220856
rect 199838 220804 199844 220856
rect 199896 220844 199902 220856
rect 201034 220844 201040 220856
rect 199896 220816 201040 220844
rect 199896 220804 199902 220816
rect 201034 220804 201040 220816
rect 201092 220804 201098 220856
rect 57606 220736 57612 220788
rect 57664 220776 57670 220788
rect 62114 220776 62120 220788
rect 57664 220748 62120 220776
rect 57664 220736 57670 220748
rect 62114 220736 62120 220748
rect 62172 220736 62178 220788
rect 67358 220736 67364 220788
rect 67416 220776 67422 220788
rect 69658 220776 69664 220788
rect 67416 220748 69664 220776
rect 67416 220736 67422 220748
rect 69658 220736 69664 220748
rect 69716 220736 69722 220788
rect 79134 220736 79140 220788
rect 79192 220776 79198 220788
rect 79962 220776 79968 220788
rect 79192 220748 79968 220776
rect 79192 220736 79198 220748
rect 79962 220736 79968 220748
rect 80020 220736 80026 220788
rect 80146 220736 80152 220788
rect 80204 220776 80210 220788
rect 102134 220776 102140 220788
rect 80204 220748 102140 220776
rect 80204 220736 80210 220748
rect 102134 220736 102140 220748
rect 102192 220736 102198 220788
rect 108114 220736 108120 220788
rect 108172 220776 108178 220788
rect 108172 220748 122834 220776
rect 108172 220736 108178 220748
rect 63402 220600 63408 220652
rect 63460 220640 63466 220652
rect 120074 220640 120080 220652
rect 63460 220612 120080 220640
rect 63460 220600 63466 220612
rect 120074 220600 120080 220612
rect 120132 220600 120138 220652
rect 122806 220640 122834 220748
rect 123846 220736 123852 220788
rect 123904 220776 123910 220788
rect 127802 220776 127808 220788
rect 123904 220748 127808 220776
rect 123904 220736 123910 220748
rect 127802 220736 127808 220748
rect 127860 220736 127866 220788
rect 127986 220736 127992 220788
rect 128044 220776 128050 220788
rect 136542 220776 136548 220788
rect 128044 220748 136548 220776
rect 128044 220736 128050 220748
rect 136542 220736 136548 220748
rect 136600 220736 136606 220788
rect 136910 220736 136916 220788
rect 136968 220776 136974 220788
rect 152458 220776 152464 220788
rect 136968 220748 152464 220776
rect 136968 220736 136974 220748
rect 152458 220736 152464 220748
rect 152516 220736 152522 220788
rect 153654 220736 153660 220788
rect 153712 220776 153718 220788
rect 154114 220776 154120 220788
rect 153712 220748 154120 220776
rect 153712 220736 153718 220748
rect 154114 220736 154120 220748
rect 154172 220736 154178 220788
rect 154482 220736 154488 220788
rect 154540 220776 154546 220788
rect 194962 220776 194968 220788
rect 154540 220748 194968 220776
rect 154540 220736 154546 220748
rect 194962 220736 194968 220748
rect 195020 220736 195026 220788
rect 195146 220736 195152 220788
rect 195204 220776 195210 220788
rect 199654 220776 199660 220788
rect 195204 220748 199660 220776
rect 195204 220736 195210 220748
rect 199654 220736 199660 220748
rect 199712 220736 199718 220788
rect 203426 220736 203432 220788
rect 203484 220776 203490 220788
rect 203484 220748 205036 220776
rect 203484 220736 203490 220748
rect 126146 220640 126152 220652
rect 122806 220612 126152 220640
rect 126146 220600 126152 220612
rect 126204 220600 126210 220652
rect 126330 220600 126336 220652
rect 126388 220640 126394 220652
rect 192478 220640 192484 220652
rect 126388 220612 192484 220640
rect 126388 220600 126394 220612
rect 192478 220600 192484 220612
rect 192536 220600 192542 220652
rect 193030 220600 193036 220652
rect 193088 220640 193094 220652
rect 205008 220640 205036 220748
rect 205266 220736 205272 220788
rect 205324 220776 205330 220788
rect 239582 220776 239588 220788
rect 205324 220748 239588 220776
rect 205324 220736 205330 220748
rect 239582 220736 239588 220748
rect 239640 220736 239646 220788
rect 239766 220736 239772 220788
rect 239824 220776 239830 220788
rect 240962 220776 240968 220788
rect 239824 220748 240968 220776
rect 239824 220736 239830 220748
rect 240962 220736 240968 220748
rect 241020 220736 241026 220788
rect 241238 220736 241244 220788
rect 241296 220776 241302 220788
rect 244550 220776 244556 220788
rect 241296 220748 244556 220776
rect 241296 220736 241302 220748
rect 244550 220736 244556 220748
rect 244608 220736 244614 220788
rect 251082 220736 251088 220788
rect 251140 220776 251146 220788
rect 252738 220776 252744 220788
rect 251140 220748 252744 220776
rect 251140 220736 251146 220748
rect 252738 220736 252744 220748
rect 252796 220736 252802 220788
rect 253014 220736 253020 220788
rect 253072 220776 253078 220788
rect 256326 220776 256332 220788
rect 253072 220748 256332 220776
rect 253072 220736 253078 220748
rect 256326 220736 256332 220748
rect 256384 220736 256390 220788
rect 267090 220736 267096 220788
rect 267148 220776 267154 220788
rect 267550 220776 267556 220788
rect 267148 220748 267556 220776
rect 267148 220736 267154 220748
rect 267550 220736 267556 220748
rect 267608 220736 267614 220788
rect 244734 220668 244740 220720
rect 244792 220708 244798 220720
rect 247954 220708 247960 220720
rect 244792 220680 247960 220708
rect 244792 220668 244798 220680
rect 247954 220668 247960 220680
rect 248012 220668 248018 220720
rect 214558 220640 214564 220652
rect 193088 220612 204944 220640
rect 205008 220612 214564 220640
rect 193088 220600 193094 220612
rect 55950 220464 55956 220516
rect 56008 220504 56014 220516
rect 56870 220504 56876 220516
rect 56008 220476 56876 220504
rect 56008 220464 56014 220476
rect 56870 220464 56876 220476
rect 56928 220464 56934 220516
rect 76650 220464 76656 220516
rect 76708 220504 76714 220516
rect 80146 220504 80152 220516
rect 76708 220476 80152 220504
rect 76708 220464 76714 220476
rect 80146 220464 80152 220476
rect 80204 220464 80210 220516
rect 87414 220464 87420 220516
rect 87472 220504 87478 220516
rect 88242 220504 88248 220516
rect 87472 220476 88248 220504
rect 87472 220464 87478 220476
rect 88242 220464 88248 220476
rect 88300 220464 88306 220516
rect 89070 220464 89076 220516
rect 89128 220504 89134 220516
rect 89622 220504 89628 220516
rect 89128 220476 89628 220504
rect 89128 220464 89134 220476
rect 89622 220464 89628 220476
rect 89680 220464 89686 220516
rect 95694 220464 95700 220516
rect 95752 220504 95758 220516
rect 97902 220504 97908 220516
rect 95752 220476 97908 220504
rect 95752 220464 95758 220476
rect 97902 220464 97908 220476
rect 97960 220464 97966 220516
rect 120534 220464 120540 220516
rect 120592 220504 120598 220516
rect 127618 220504 127624 220516
rect 120592 220476 127624 220504
rect 120592 220464 120598 220476
rect 127618 220464 127624 220476
rect 127676 220464 127682 220516
rect 127802 220464 127808 220516
rect 127860 220504 127866 220516
rect 161750 220504 161756 220516
rect 127860 220476 161756 220504
rect 127860 220464 127866 220476
rect 161750 220464 161756 220476
rect 161808 220464 161814 220516
rect 161934 220464 161940 220516
rect 161992 220504 161998 220516
rect 162394 220504 162400 220516
rect 161992 220476 162400 220504
rect 161992 220464 161998 220476
rect 162394 220464 162400 220476
rect 162452 220464 162458 220516
rect 162578 220464 162584 220516
rect 162636 220504 162642 220516
rect 165062 220504 165068 220516
rect 162636 220476 165068 220504
rect 162636 220464 162642 220476
rect 165062 220464 165068 220476
rect 165120 220464 165126 220516
rect 165614 220464 165620 220516
rect 165672 220504 165678 220516
rect 166442 220504 166448 220516
rect 165672 220476 166448 220504
rect 165672 220464 165678 220476
rect 166442 220464 166448 220476
rect 166500 220464 166506 220516
rect 166626 220464 166632 220516
rect 166684 220504 166690 220516
rect 203610 220504 203616 220516
rect 166684 220476 203616 220504
rect 166684 220464 166690 220476
rect 203610 220464 203616 220476
rect 203668 220464 203674 220516
rect 204916 220504 204944 220612
rect 214558 220600 214564 220612
rect 214616 220600 214622 220652
rect 216306 220600 216312 220652
rect 216364 220640 216370 220652
rect 219710 220640 219716 220652
rect 216364 220612 219716 220640
rect 216364 220600 216370 220612
rect 219710 220600 219716 220612
rect 219768 220600 219774 220652
rect 219894 220600 219900 220652
rect 219952 220640 219958 220652
rect 220446 220640 220452 220652
rect 219952 220612 220452 220640
rect 219952 220600 219958 220612
rect 220446 220600 220452 220612
rect 220504 220600 220510 220652
rect 221550 220600 221556 220652
rect 221608 220640 221614 220652
rect 222286 220640 222292 220652
rect 221608 220612 222292 220640
rect 221608 220600 221614 220612
rect 222286 220600 222292 220612
rect 222344 220600 222350 220652
rect 222470 220600 222476 220652
rect 222528 220640 222534 220652
rect 223850 220640 223856 220652
rect 222528 220612 223856 220640
rect 222528 220600 222534 220612
rect 223850 220600 223856 220612
rect 223908 220600 223914 220652
rect 224034 220600 224040 220652
rect 224092 220640 224098 220652
rect 224092 220612 224356 220640
rect 224092 220600 224098 220612
rect 224328 220504 224356 220612
rect 224494 220600 224500 220652
rect 224552 220640 224558 220652
rect 232682 220640 232688 220652
rect 224552 220612 232688 220640
rect 224552 220600 224558 220612
rect 232682 220600 232688 220612
rect 232740 220600 232746 220652
rect 232866 220600 232872 220652
rect 232924 220640 232930 220652
rect 233878 220640 233884 220652
rect 232924 220612 233884 220640
rect 232924 220600 232930 220612
rect 233878 220600 233884 220612
rect 233936 220600 233942 220652
rect 236454 220600 236460 220652
rect 236512 220640 236518 220652
rect 243722 220640 243728 220652
rect 236512 220612 243728 220640
rect 236512 220600 236518 220612
rect 243722 220600 243728 220612
rect 243780 220600 243786 220652
rect 249518 220600 249524 220652
rect 249576 220640 249582 220652
rect 274652 220640 274680 220884
rect 277578 220872 277584 220884
rect 277636 220872 277642 220924
rect 418982 220872 418988 220924
rect 419040 220912 419046 220924
rect 455414 220912 455420 220924
rect 419040 220884 455420 220912
rect 419040 220872 419046 220884
rect 455414 220872 455420 220884
rect 455472 220872 455478 220924
rect 596928 220912 596956 221020
rect 597094 221008 597100 221060
rect 597152 221048 597158 221060
rect 608778 221048 608784 221060
rect 597152 221020 608784 221048
rect 597152 221008 597158 221020
rect 608778 221008 608784 221020
rect 608836 221008 608842 221060
rect 673270 220940 673276 220992
rect 673328 220980 673334 220992
rect 675110 220980 675116 220992
rect 673328 220952 675116 220980
rect 673328 220940 673334 220952
rect 675110 220940 675116 220952
rect 675168 220940 675174 220992
rect 602246 220912 602252 220924
rect 596928 220884 602252 220912
rect 602246 220872 602252 220884
rect 602304 220872 602310 220924
rect 296070 220804 296076 220856
rect 296128 220844 296134 220856
rect 297358 220844 297364 220856
rect 296128 220816 297364 220844
rect 296128 220804 296134 220816
rect 297358 220804 297364 220816
rect 297416 220804 297422 220856
rect 313458 220844 313464 220856
rect 309152 220816 313464 220844
rect 275646 220736 275652 220788
rect 275704 220776 275710 220788
rect 290458 220776 290464 220788
rect 275704 220748 290464 220776
rect 275704 220736 275710 220748
rect 290458 220736 290464 220748
rect 290516 220736 290522 220788
rect 302694 220736 302700 220788
rect 302752 220776 302758 220788
rect 305638 220776 305644 220788
rect 302752 220748 305644 220776
rect 302752 220736 302758 220748
rect 305638 220736 305644 220748
rect 305696 220736 305702 220788
rect 249576 220612 274680 220640
rect 249576 220600 249582 220612
rect 277854 220600 277860 220652
rect 277912 220640 277918 220652
rect 279602 220640 279608 220652
rect 277912 220612 279608 220640
rect 277912 220600 277918 220612
rect 279602 220600 279608 220612
rect 279660 220600 279666 220652
rect 304626 220600 304632 220652
rect 304684 220640 304690 220652
rect 309152 220640 309180 220816
rect 313458 220804 313464 220816
rect 313516 220804 313522 220856
rect 461210 220804 461216 220856
rect 461268 220844 461274 220856
rect 528370 220844 528376 220856
rect 461268 220816 528376 220844
rect 461268 220804 461274 220816
rect 528370 220804 528376 220816
rect 528428 220844 528434 220856
rect 596726 220844 596732 220856
rect 528428 220816 596732 220844
rect 528428 220804 528434 220816
rect 596726 220804 596732 220816
rect 596784 220804 596790 220856
rect 667842 220804 667848 220856
rect 667900 220844 667906 220856
rect 675294 220844 675300 220856
rect 667900 220816 675300 220844
rect 667900 220804 667906 220816
rect 675294 220804 675300 220816
rect 675352 220804 675358 220856
rect 316770 220736 316776 220788
rect 316828 220776 316834 220788
rect 320542 220776 320548 220788
rect 316828 220748 320548 220776
rect 316828 220736 316834 220748
rect 320542 220736 320548 220748
rect 320600 220736 320606 220788
rect 320910 220736 320916 220788
rect 320968 220776 320974 220788
rect 321370 220776 321376 220788
rect 320968 220748 321376 220776
rect 320968 220736 320974 220748
rect 321370 220736 321376 220748
rect 321428 220736 321434 220788
rect 323394 220736 323400 220788
rect 323452 220776 323458 220788
rect 324958 220776 324964 220788
rect 323452 220748 324964 220776
rect 323452 220736 323458 220748
rect 324958 220736 324964 220748
rect 325016 220736 325022 220788
rect 326706 220736 326712 220788
rect 326764 220776 326770 220788
rect 327350 220776 327356 220788
rect 326764 220748 327356 220776
rect 326764 220736 326770 220748
rect 327350 220736 327356 220748
rect 327408 220736 327414 220788
rect 328178 220736 328184 220788
rect 328236 220776 328242 220788
rect 328914 220776 328920 220788
rect 328236 220748 328920 220776
rect 328236 220736 328242 220748
rect 328914 220736 328920 220748
rect 328972 220736 328978 220788
rect 329098 220736 329104 220788
rect 329156 220776 329162 220788
rect 330478 220776 330484 220788
rect 329156 220748 330484 220776
rect 329156 220736 329162 220748
rect 330478 220736 330484 220748
rect 330536 220736 330542 220788
rect 330846 220736 330852 220788
rect 330904 220776 330910 220788
rect 332134 220776 332140 220788
rect 330904 220748 332140 220776
rect 330904 220736 330910 220748
rect 332134 220736 332140 220748
rect 332192 220736 332198 220788
rect 333882 220736 333888 220788
rect 333940 220776 333946 220788
rect 334342 220776 334348 220788
rect 333940 220748 334348 220776
rect 333940 220736 333946 220748
rect 334342 220736 334348 220748
rect 334400 220736 334406 220788
rect 346210 220736 346216 220788
rect 346268 220776 346274 220788
rect 351914 220776 351920 220788
rect 346268 220748 351920 220776
rect 346268 220736 346274 220748
rect 351914 220736 351920 220748
rect 351972 220736 351978 220788
rect 355318 220736 355324 220788
rect 355376 220776 355382 220788
rect 358354 220776 358360 220788
rect 355376 220748 358360 220776
rect 355376 220736 355382 220748
rect 358354 220736 358360 220748
rect 358412 220736 358418 220788
rect 365254 220736 365260 220788
rect 365312 220776 365318 220788
rect 366634 220776 366640 220788
rect 365312 220748 366640 220776
rect 365312 220736 365318 220748
rect 366634 220736 366640 220748
rect 366692 220736 366698 220788
rect 395154 220736 395160 220788
rect 395212 220776 395218 220788
rect 398098 220776 398104 220788
rect 395212 220748 398104 220776
rect 395212 220736 395218 220748
rect 398098 220736 398104 220748
rect 398156 220736 398162 220788
rect 423030 220736 423036 220788
rect 423088 220776 423094 220788
rect 425422 220776 425428 220788
rect 423088 220748 425428 220776
rect 423088 220736 423094 220748
rect 425422 220736 425428 220748
rect 425480 220736 425486 220788
rect 429194 220736 429200 220788
rect 429252 220776 429258 220788
rect 456058 220776 456064 220788
rect 429252 220748 456064 220776
rect 429252 220736 429258 220748
rect 456058 220736 456064 220748
rect 456116 220736 456122 220788
rect 591298 220668 591304 220720
rect 591356 220708 591362 220720
rect 591356 220680 596174 220708
rect 591356 220668 591362 220680
rect 304684 220612 309180 220640
rect 304684 220600 304690 220612
rect 321186 220600 321192 220652
rect 321244 220640 321250 220652
rect 324682 220640 324688 220652
rect 321244 220612 324688 220640
rect 321244 220600 321250 220612
rect 324682 220600 324688 220612
rect 324740 220600 324746 220652
rect 327534 220600 327540 220652
rect 327592 220640 327598 220652
rect 330202 220640 330208 220652
rect 327592 220612 330208 220640
rect 327592 220600 327598 220612
rect 330202 220600 330208 220612
rect 330260 220600 330266 220652
rect 355686 220600 355692 220652
rect 355744 220640 355750 220652
rect 356698 220640 356704 220652
rect 355744 220612 356704 220640
rect 355744 220600 355750 220612
rect 356698 220600 356704 220612
rect 356756 220600 356762 220652
rect 357618 220600 357624 220652
rect 357676 220640 357682 220652
rect 360194 220640 360200 220652
rect 357676 220612 360200 220640
rect 357676 220600 357682 220612
rect 360194 220600 360200 220612
rect 360252 220600 360258 220652
rect 393038 220600 393044 220652
rect 393096 220640 393102 220652
rect 421282 220640 421288 220652
rect 393096 220612 421288 220640
rect 393096 220600 393102 220612
rect 421282 220600 421288 220612
rect 421340 220600 421346 220652
rect 425790 220600 425796 220652
rect 425848 220640 425854 220652
rect 435542 220640 435548 220652
rect 425848 220612 435548 220640
rect 425848 220600 425854 220612
rect 435542 220600 435548 220612
rect 435600 220600 435606 220652
rect 444006 220600 444012 220652
rect 444064 220640 444070 220652
rect 449434 220640 449440 220652
rect 444064 220612 449440 220640
rect 444064 220600 444070 220612
rect 449434 220600 449440 220612
rect 449492 220600 449498 220652
rect 449710 220600 449716 220652
rect 449768 220640 449774 220652
rect 449768 220612 451274 220640
rect 449768 220600 449774 220612
rect 250346 220504 250352 220516
rect 204916 220476 224264 220504
rect 224328 220476 250352 220504
rect 60642 220396 60648 220448
rect 60700 220436 60706 220448
rect 61378 220436 61384 220448
rect 60700 220408 61384 220436
rect 60700 220396 60706 220408
rect 61378 220396 61384 220408
rect 61436 220396 61442 220448
rect 89438 220328 89444 220380
rect 89496 220368 89502 220380
rect 165982 220368 165988 220380
rect 89496 220340 165988 220368
rect 89496 220328 89502 220340
rect 165982 220328 165988 220340
rect 166040 220328 166046 220380
rect 170030 220368 170036 220380
rect 166828 220340 170036 220368
rect 62574 220192 62580 220244
rect 62632 220232 62638 220244
rect 63586 220232 63592 220244
rect 62632 220204 63592 220232
rect 62632 220192 62638 220204
rect 63586 220192 63592 220204
rect 63644 220192 63650 220244
rect 77202 220192 77208 220244
rect 77260 220232 77266 220244
rect 156874 220232 156880 220244
rect 77260 220204 156880 220232
rect 77260 220192 77266 220204
rect 156874 220192 156880 220204
rect 156932 220192 156938 220244
rect 161290 220232 161296 220244
rect 157168 220204 161296 220232
rect 157168 220164 157196 220204
rect 161290 220192 161296 220204
rect 161348 220192 161354 220244
rect 161750 220192 161756 220244
rect 161808 220232 161814 220244
rect 166828 220232 166856 220340
rect 170030 220328 170036 220340
rect 170088 220328 170094 220380
rect 170214 220328 170220 220380
rect 170272 220368 170278 220380
rect 219526 220368 219532 220380
rect 170272 220340 219532 220368
rect 170272 220328 170278 220340
rect 219526 220328 219532 220340
rect 219584 220328 219590 220380
rect 219710 220328 219716 220380
rect 219768 220368 219774 220380
rect 224034 220368 224040 220380
rect 219768 220340 224040 220368
rect 219768 220328 219774 220340
rect 224034 220328 224040 220340
rect 224092 220328 224098 220380
rect 224236 220368 224264 220476
rect 250346 220464 250352 220476
rect 250404 220464 250410 220516
rect 252830 220464 252836 220516
rect 252888 220504 252894 220516
rect 253566 220504 253572 220516
rect 252888 220476 253572 220504
rect 252888 220464 252894 220476
rect 253566 220464 253572 220476
rect 253624 220464 253630 220516
rect 256326 220464 256332 220516
rect 256384 220504 256390 220516
rect 281810 220504 281816 220516
rect 256384 220476 281816 220504
rect 256384 220464 256390 220476
rect 281810 220464 281816 220476
rect 281868 220464 281874 220516
rect 297726 220464 297732 220516
rect 297784 220504 297790 220516
rect 299382 220504 299388 220516
rect 297784 220476 299388 220504
rect 297784 220464 297790 220476
rect 299382 220464 299388 220476
rect 299440 220464 299446 220516
rect 306834 220464 306840 220516
rect 306892 220504 306898 220516
rect 310606 220504 310612 220516
rect 306892 220476 310612 220504
rect 306892 220464 306898 220476
rect 310606 220464 310612 220476
rect 310664 220464 310670 220516
rect 320082 220464 320088 220516
rect 320140 220504 320146 220516
rect 323210 220504 323216 220516
rect 320140 220476 323216 220504
rect 320140 220464 320146 220476
rect 323210 220464 323216 220476
rect 323268 220464 323274 220516
rect 376110 220464 376116 220516
rect 376168 220504 376174 220516
rect 388162 220504 388168 220516
rect 376168 220476 388168 220504
rect 376168 220464 376174 220476
rect 388162 220464 388168 220476
rect 388220 220464 388226 220516
rect 397362 220464 397368 220516
rect 397420 220504 397426 220516
rect 427906 220504 427912 220516
rect 397420 220476 427912 220504
rect 397420 220464 397426 220476
rect 427906 220464 427912 220476
rect 427964 220464 427970 220516
rect 434714 220464 434720 220516
rect 434772 220504 434778 220516
rect 437014 220504 437020 220516
rect 434772 220476 437020 220504
rect 434772 220464 434778 220476
rect 437014 220464 437020 220476
rect 437072 220464 437078 220516
rect 445294 220464 445300 220516
rect 445352 220504 445358 220516
rect 445662 220504 445668 220516
rect 445352 220476 445668 220504
rect 445352 220464 445358 220476
rect 445662 220464 445668 220476
rect 445720 220464 445726 220516
rect 451246 220504 451274 220612
rect 452562 220600 452568 220652
rect 452620 220640 452626 220652
rect 456978 220640 456984 220652
rect 452620 220612 456984 220640
rect 452620 220600 452626 220612
rect 456978 220600 456984 220612
rect 457036 220600 457042 220652
rect 457162 220600 457168 220652
rect 457220 220640 457226 220652
rect 470134 220640 470140 220652
rect 457220 220612 470140 220640
rect 457220 220600 457226 220612
rect 470134 220600 470140 220612
rect 470192 220600 470198 220652
rect 480346 220640 480352 220652
rect 470566 220612 480352 220640
rect 470566 220504 470594 220612
rect 480346 220600 480352 220612
rect 480404 220600 480410 220652
rect 502334 220640 502340 220652
rect 480916 220612 502340 220640
rect 451246 220476 470594 220504
rect 471790 220464 471796 220516
rect 471848 220504 471854 220516
rect 475194 220504 475200 220516
rect 471848 220476 475200 220504
rect 471848 220464 471854 220476
rect 475194 220464 475200 220476
rect 475252 220464 475258 220516
rect 475378 220464 475384 220516
rect 475436 220504 475442 220516
rect 480916 220504 480944 220612
rect 502334 220600 502340 220612
rect 502392 220600 502398 220652
rect 504358 220600 504364 220652
rect 504416 220640 504422 220652
rect 506014 220640 506020 220652
rect 504416 220612 506020 220640
rect 504416 220600 504422 220612
rect 506014 220600 506020 220612
rect 506072 220600 506078 220652
rect 506198 220600 506204 220652
rect 506256 220640 506262 220652
rect 528554 220640 528560 220652
rect 506256 220612 528560 220640
rect 506256 220600 506262 220612
rect 528554 220600 528560 220612
rect 528612 220600 528618 220652
rect 548334 220600 548340 220652
rect 548392 220640 548398 220652
rect 562502 220640 562508 220652
rect 548392 220612 562508 220640
rect 548392 220600 548398 220612
rect 562502 220600 562508 220612
rect 562560 220600 562566 220652
rect 562962 220600 562968 220652
rect 563020 220640 563026 220652
rect 596146 220640 596174 220680
rect 596266 220640 596272 220652
rect 563020 220612 591160 220640
rect 596146 220612 596272 220640
rect 563020 220600 563026 220612
rect 591132 220572 591160 220612
rect 596266 220600 596272 220612
rect 596324 220600 596330 220652
rect 591132 220544 591344 220572
rect 475436 220476 480944 220504
rect 475436 220464 475442 220476
rect 481082 220464 481088 220516
rect 481140 220504 481146 220516
rect 481140 220476 528554 220504
rect 481140 220464 481146 220476
rect 229462 220368 229468 220380
rect 224236 220340 229468 220368
rect 229462 220328 229468 220340
rect 229520 220328 229526 220380
rect 231486 220328 231492 220380
rect 231544 220368 231550 220380
rect 235994 220368 236000 220380
rect 231544 220340 236000 220368
rect 231544 220328 231550 220340
rect 235994 220328 236000 220340
rect 236052 220328 236058 220380
rect 239582 220328 239588 220380
rect 239640 220368 239646 220380
rect 239640 220340 242296 220368
rect 239640 220328 239646 220340
rect 161808 220204 166856 220232
rect 161808 220192 161814 220204
rect 166948 220192 166954 220244
rect 167006 220232 167012 220244
rect 171042 220232 171048 220244
rect 167006 220204 171048 220232
rect 167006 220192 167012 220204
rect 171042 220192 171048 220204
rect 171100 220192 171106 220244
rect 171870 220192 171876 220244
rect 171928 220232 171934 220244
rect 173434 220232 173440 220244
rect 171928 220204 173440 220232
rect 171928 220192 171934 220204
rect 173434 220192 173440 220204
rect 173492 220192 173498 220244
rect 173618 220192 173624 220244
rect 173676 220232 173682 220244
rect 181070 220232 181076 220244
rect 173676 220204 181076 220232
rect 173676 220192 173682 220204
rect 181070 220192 181076 220204
rect 181128 220192 181134 220244
rect 186866 220192 186872 220244
rect 186924 220232 186930 220244
rect 187418 220232 187424 220244
rect 186924 220204 187424 220232
rect 186924 220192 186930 220204
rect 187418 220192 187424 220204
rect 187476 220192 187482 220244
rect 187602 220192 187608 220244
rect 187660 220232 187666 220244
rect 187660 220204 204944 220232
rect 187660 220192 187666 220204
rect 157076 220136 157196 220164
rect 58434 220056 58440 220108
rect 58492 220096 58498 220108
rect 60366 220096 60372 220108
rect 58492 220068 60372 220096
rect 58492 220056 58498 220068
rect 60366 220056 60372 220068
rect 60424 220056 60430 220108
rect 64782 220056 64788 220108
rect 64840 220096 64846 220108
rect 77018 220096 77024 220108
rect 64840 220068 77024 220096
rect 64840 220056 64846 220068
rect 77018 220056 77024 220068
rect 77076 220056 77082 220108
rect 103974 220056 103980 220108
rect 104032 220096 104038 220108
rect 147628 220096 147634 220108
rect 104032 220068 147634 220096
rect 104032 220056 104038 220068
rect 147628 220056 147634 220068
rect 147686 220056 147692 220108
rect 147766 220056 147772 220108
rect 147824 220096 147830 220108
rect 148962 220096 148968 220108
rect 147824 220068 148968 220096
rect 147824 220056 147830 220068
rect 148962 220056 148968 220068
rect 149020 220056 149026 220108
rect 149146 220056 149152 220108
rect 149204 220096 149210 220108
rect 150158 220096 150164 220108
rect 149204 220068 150164 220096
rect 149204 220056 149210 220068
rect 150158 220056 150164 220068
rect 150216 220056 150222 220108
rect 151078 220056 151084 220108
rect 151136 220096 151142 220108
rect 151814 220096 151820 220108
rect 151136 220068 151820 220096
rect 151136 220056 151142 220068
rect 151814 220056 151820 220068
rect 151872 220056 151878 220108
rect 152458 220056 152464 220108
rect 152516 220096 152522 220108
rect 157076 220096 157104 220136
rect 152516 220068 157104 220096
rect 152516 220056 152522 220068
rect 157334 220056 157340 220108
rect 157392 220096 157398 220108
rect 204622 220096 204628 220108
rect 157392 220068 204628 220096
rect 157392 220056 157398 220068
rect 204622 220056 204628 220068
rect 204680 220056 204686 220108
rect 204916 220096 204944 220204
rect 205082 220192 205088 220244
rect 205140 220232 205146 220244
rect 242066 220232 242072 220244
rect 205140 220204 242072 220232
rect 205140 220192 205146 220204
rect 242066 220192 242072 220204
rect 242124 220192 242130 220244
rect 242268 220232 242296 220340
rect 242618 220328 242624 220380
rect 242676 220368 242682 220380
rect 273530 220368 273536 220380
rect 242676 220340 273536 220368
rect 242676 220328 242682 220340
rect 273530 220328 273536 220340
rect 273588 220328 273594 220380
rect 274358 220328 274364 220380
rect 274416 220368 274422 220380
rect 276290 220368 276296 220380
rect 274416 220340 276296 220368
rect 274416 220328 274422 220340
rect 276290 220328 276296 220340
rect 276348 220328 276354 220380
rect 282546 220328 282552 220380
rect 282604 220368 282610 220380
rect 298738 220368 298744 220380
rect 282604 220340 298744 220368
rect 282604 220328 282610 220340
rect 298738 220328 298744 220340
rect 298796 220328 298802 220380
rect 300762 220328 300768 220380
rect 300820 220368 300826 220380
rect 304994 220368 305000 220380
rect 300820 220340 305000 220368
rect 300820 220328 300826 220340
rect 304994 220328 305000 220340
rect 305052 220328 305058 220380
rect 318426 220328 318432 220380
rect 318484 220368 318490 220380
rect 322198 220368 322204 220380
rect 318484 220340 322204 220368
rect 318484 220328 318490 220340
rect 322198 220328 322204 220340
rect 322256 220328 322262 220380
rect 325602 220328 325608 220380
rect 325660 220368 325666 220380
rect 328730 220368 328736 220380
rect 325660 220340 328736 220368
rect 325660 220328 325666 220340
rect 328730 220328 328736 220340
rect 328788 220328 328794 220380
rect 366450 220328 366456 220380
rect 366508 220368 366514 220380
rect 381538 220368 381544 220380
rect 366508 220340 381544 220368
rect 366508 220328 366514 220340
rect 381538 220328 381544 220340
rect 381596 220328 381602 220380
rect 388438 220328 388444 220380
rect 388496 220368 388502 220380
rect 404722 220368 404728 220380
rect 388496 220340 404728 220368
rect 388496 220328 388502 220340
rect 404722 220328 404728 220340
rect 404780 220328 404786 220380
rect 404998 220328 405004 220380
rect 405056 220368 405062 220380
rect 437842 220368 437848 220380
rect 405056 220340 437848 220368
rect 405056 220328 405062 220340
rect 437842 220328 437848 220340
rect 437900 220328 437906 220380
rect 441430 220328 441436 220380
rect 441488 220368 441494 220380
rect 495250 220368 495256 220380
rect 441488 220340 495256 220368
rect 441488 220328 441494 220340
rect 495250 220328 495256 220340
rect 495308 220328 495314 220380
rect 495388 220328 495394 220380
rect 495446 220368 495452 220380
rect 504358 220368 504364 220380
rect 495446 220340 504364 220368
rect 495446 220328 495452 220340
rect 504358 220328 504364 220340
rect 504416 220328 504422 220380
rect 504542 220328 504548 220380
rect 504600 220368 504606 220380
rect 511534 220368 511540 220380
rect 504600 220340 511540 220368
rect 504600 220328 504606 220340
rect 511534 220328 511540 220340
rect 511592 220328 511598 220380
rect 513374 220328 513380 220380
rect 513432 220368 513438 220380
rect 515582 220368 515588 220380
rect 513432 220340 515588 220368
rect 513432 220328 513438 220340
rect 515582 220328 515588 220340
rect 515640 220328 515646 220380
rect 528526 220368 528554 220476
rect 534718 220464 534724 220516
rect 534776 220504 534782 220516
rect 542538 220504 542544 220516
rect 534776 220476 542544 220504
rect 534776 220464 534782 220476
rect 542538 220464 542544 220476
rect 542596 220464 542602 220516
rect 544562 220464 544568 220516
rect 544620 220504 544626 220516
rect 548150 220504 548156 220516
rect 544620 220476 548156 220504
rect 544620 220464 544626 220476
rect 548150 220464 548156 220476
rect 548208 220464 548214 220516
rect 548518 220464 548524 220516
rect 548576 220504 548582 220516
rect 572530 220504 572536 220516
rect 548576 220476 572536 220504
rect 548576 220464 548582 220476
rect 572530 220464 572536 220476
rect 572588 220464 572594 220516
rect 572668 220464 572674 220516
rect 572726 220504 572732 220516
rect 590930 220504 590936 220516
rect 572726 220476 590936 220504
rect 572726 220464 572732 220476
rect 590930 220464 590936 220476
rect 590988 220464 590994 220516
rect 591316 220504 591344 220544
rect 602890 220504 602896 220516
rect 591316 220476 602896 220504
rect 602890 220464 602896 220476
rect 602948 220464 602954 220516
rect 532510 220368 532516 220380
rect 528526 220340 532516 220368
rect 532510 220328 532516 220340
rect 532568 220368 532574 220380
rect 607214 220368 607220 220380
rect 532568 220340 607220 220368
rect 532568 220328 532574 220340
rect 607214 220328 607220 220340
rect 607272 220328 607278 220380
rect 307662 220260 307668 220312
rect 307720 220300 307726 220312
rect 315850 220300 315856 220312
rect 307720 220272 315856 220300
rect 307720 220260 307726 220272
rect 315850 220260 315856 220272
rect 315908 220260 315914 220312
rect 242894 220232 242900 220244
rect 242268 220204 242900 220232
rect 242894 220192 242900 220204
rect 242952 220192 242958 220244
rect 243538 220192 243544 220244
rect 243596 220232 243602 220244
rect 252830 220232 252836 220244
rect 243596 220204 252836 220232
rect 243596 220192 243602 220204
rect 252830 220192 252836 220204
rect 252888 220192 252894 220244
rect 259822 220232 259828 220244
rect 253124 220204 259828 220232
rect 219342 220096 219348 220108
rect 204916 220068 219348 220096
rect 219342 220056 219348 220068
rect 219400 220056 219406 220108
rect 219526 220056 219532 220108
rect 219584 220096 219590 220108
rect 222470 220096 222476 220108
rect 219584 220068 222476 220096
rect 219584 220056 219590 220068
rect 222470 220056 222476 220068
rect 222528 220056 222534 220108
rect 223206 220056 223212 220108
rect 223264 220096 223270 220108
rect 224494 220096 224500 220108
rect 223264 220068 224500 220096
rect 223264 220056 223270 220068
rect 224494 220056 224500 220068
rect 224552 220056 224558 220108
rect 224678 220056 224684 220108
rect 224736 220096 224742 220108
rect 226610 220096 226616 220108
rect 224736 220068 226616 220096
rect 224736 220056 224742 220068
rect 226610 220056 226616 220068
rect 226668 220056 226674 220108
rect 231854 220096 231860 220108
rect 229066 220068 231860 220096
rect 101858 219920 101864 219972
rect 101916 219960 101922 219972
rect 104802 219960 104808 219972
rect 101916 219932 104808 219960
rect 101916 219920 101922 219932
rect 104802 219920 104808 219932
rect 104860 219920 104866 219972
rect 113910 219920 113916 219972
rect 113968 219960 113974 219972
rect 113968 219932 122834 219960
rect 113968 219920 113974 219932
rect 83918 219784 83924 219836
rect 83976 219824 83982 219836
rect 88886 219824 88892 219836
rect 83976 219796 88892 219824
rect 83976 219784 83982 219796
rect 88886 219784 88892 219796
rect 88944 219784 88950 219836
rect 103146 219784 103152 219836
rect 103204 219824 103210 219836
rect 118786 219824 118792 219836
rect 103204 219796 118792 219824
rect 103204 219784 103210 219796
rect 118786 219784 118792 219796
rect 118844 219784 118850 219836
rect 122806 219824 122834 219932
rect 127618 219920 127624 219972
rect 127676 219960 127682 219972
rect 166810 219960 166816 219972
rect 127676 219932 166816 219960
rect 127676 219920 127682 219932
rect 166810 219920 166816 219932
rect 166868 219920 166874 219972
rect 166948 219920 166954 219972
rect 167006 219960 167012 219972
rect 187602 219960 187608 219972
rect 167006 219932 187608 219960
rect 167006 219920 167012 219932
rect 187602 219920 187608 219932
rect 187660 219920 187666 219972
rect 187786 219920 187792 219972
rect 187844 219960 187850 219972
rect 229066 219960 229094 220068
rect 231854 220056 231860 220068
rect 231912 220056 231918 220108
rect 232682 220056 232688 220108
rect 232740 220096 232746 220108
rect 253124 220096 253152 220204
rect 259822 220192 259828 220204
rect 259880 220192 259886 220244
rect 262950 220192 262956 220244
rect 263008 220232 263014 220244
rect 284938 220232 284944 220244
rect 263008 220204 284944 220232
rect 263008 220192 263014 220204
rect 284938 220192 284944 220204
rect 284996 220192 285002 220244
rect 286134 220192 286140 220244
rect 286192 220232 286198 220244
rect 293954 220232 293960 220244
rect 286192 220204 293960 220232
rect 286192 220192 286198 220204
rect 293954 220192 293960 220204
rect 294012 220192 294018 220244
rect 299198 220192 299204 220244
rect 299256 220232 299262 220244
rect 303338 220232 303344 220244
rect 299256 220204 303344 220232
rect 299256 220192 299262 220204
rect 303338 220192 303344 220204
rect 303396 220192 303402 220244
rect 356882 220192 356888 220244
rect 356940 220232 356946 220244
rect 365162 220232 365168 220244
rect 356940 220204 365168 220232
rect 356940 220192 356946 220204
rect 365162 220192 365168 220204
rect 365220 220192 365226 220244
rect 368106 220192 368112 220244
rect 368164 220232 368170 220244
rect 385034 220232 385040 220244
rect 368164 220204 385040 220232
rect 368164 220192 368170 220204
rect 385034 220192 385040 220204
rect 385092 220192 385098 220244
rect 401410 220192 401416 220244
rect 401468 220232 401474 220244
rect 434806 220232 434812 220244
rect 401468 220204 434812 220232
rect 401468 220192 401474 220204
rect 434806 220192 434812 220204
rect 434864 220192 434870 220244
rect 437474 220192 437480 220244
rect 437532 220232 437538 220244
rect 450262 220232 450268 220244
rect 437532 220204 450268 220232
rect 437532 220192 437538 220204
rect 450262 220192 450268 220204
rect 450320 220192 450326 220244
rect 450906 220192 450912 220244
rect 450964 220232 450970 220244
rect 511994 220232 512000 220244
rect 450964 220204 512000 220232
rect 450964 220192 450970 220204
rect 511994 220192 512000 220204
rect 512052 220192 512058 220244
rect 540330 220192 540336 220244
rect 540388 220232 540394 220244
rect 622670 220232 622676 220244
rect 540388 220204 622676 220232
rect 540388 220192 540394 220204
rect 622670 220192 622676 220204
rect 622728 220192 622734 220244
rect 232740 220068 253152 220096
rect 232740 220056 232746 220068
rect 253566 220056 253572 220108
rect 253624 220096 253630 220108
rect 264238 220096 264244 220108
rect 253624 220068 264244 220096
rect 253624 220056 253630 220068
rect 264238 220056 264244 220068
rect 264296 220056 264302 220108
rect 269574 220056 269580 220108
rect 269632 220096 269638 220108
rect 287606 220096 287612 220108
rect 269632 220068 287612 220096
rect 269632 220056 269638 220068
rect 287606 220056 287612 220068
rect 287664 220056 287670 220108
rect 287790 220056 287796 220108
rect 287848 220096 287854 220108
rect 288618 220096 288624 220108
rect 287848 220068 288624 220096
rect 287848 220056 287854 220068
rect 288618 220056 288624 220068
rect 288676 220056 288682 220108
rect 292298 220056 292304 220108
rect 292356 220096 292362 220108
rect 299750 220096 299756 220108
rect 292356 220068 299756 220096
rect 292356 220056 292362 220068
rect 299750 220056 299756 220068
rect 299808 220056 299814 220108
rect 319254 220056 319260 220108
rect 319312 220096 319318 220108
rect 323854 220096 323860 220108
rect 319312 220068 323860 220096
rect 319312 220056 319318 220068
rect 323854 220056 323860 220068
rect 323912 220056 323918 220108
rect 353202 220056 353208 220108
rect 353260 220096 353266 220108
rect 361666 220096 361672 220108
rect 353260 220068 361672 220096
rect 353260 220056 353266 220068
rect 361666 220056 361672 220068
rect 361724 220056 361730 220108
rect 364150 220056 364156 220108
rect 364208 220096 364214 220108
rect 378226 220096 378232 220108
rect 364208 220068 378232 220096
rect 364208 220056 364214 220068
rect 378226 220056 378232 220068
rect 378284 220056 378290 220108
rect 379514 220056 379520 220108
rect 379572 220096 379578 220108
rect 401594 220096 401600 220108
rect 379572 220068 401600 220096
rect 379572 220056 379578 220068
rect 401594 220056 401600 220068
rect 401652 220056 401658 220108
rect 408126 220056 408132 220108
rect 408184 220096 408190 220108
rect 444558 220096 444564 220108
rect 408184 220068 444564 220096
rect 408184 220056 408190 220068
rect 444558 220056 444564 220068
rect 444616 220056 444622 220108
rect 453942 220056 453948 220108
rect 454000 220096 454006 220108
rect 463694 220096 463700 220108
rect 454000 220068 463700 220096
rect 454000 220056 454006 220068
rect 463694 220056 463700 220068
rect 463752 220056 463758 220108
rect 465074 220056 465080 220108
rect 465132 220096 465138 220108
rect 475562 220096 475568 220108
rect 465132 220068 475568 220096
rect 465132 220056 465138 220068
rect 475562 220056 475568 220068
rect 475620 220056 475626 220108
rect 475746 220056 475752 220108
rect 475804 220096 475810 220108
rect 480530 220096 480536 220108
rect 475804 220068 480536 220096
rect 475804 220056 475810 220068
rect 480530 220056 480536 220068
rect 480588 220056 480594 220108
rect 480714 220056 480720 220108
rect 480772 220096 480778 220108
rect 481266 220096 481272 220108
rect 480772 220068 481272 220096
rect 480772 220056 480778 220068
rect 481266 220056 481272 220068
rect 481324 220056 481330 220108
rect 481450 220056 481456 220108
rect 481508 220096 481514 220108
rect 542354 220096 542360 220108
rect 481508 220068 542360 220096
rect 481508 220056 481514 220068
rect 542354 220056 542360 220068
rect 542412 220056 542418 220108
rect 542538 219988 542544 220040
rect 542596 220028 542602 220040
rect 548518 220028 548524 220040
rect 542596 220000 548524 220028
rect 542596 219988 542602 220000
rect 548518 219988 548524 220000
rect 548576 219988 548582 220040
rect 548886 219988 548892 220040
rect 548944 220028 548950 220040
rect 601510 220028 601516 220040
rect 548944 220000 601516 220028
rect 548944 219988 548950 220000
rect 601510 219988 601516 220000
rect 601568 219988 601574 220040
rect 187844 219932 229094 219960
rect 187844 219920 187850 219932
rect 229830 219920 229836 219972
rect 229888 219960 229894 219972
rect 243538 219960 243544 219972
rect 229888 219932 243544 219960
rect 229888 219920 229894 219932
rect 243538 219920 243544 219932
rect 243596 219920 243602 219972
rect 243722 219920 243728 219972
rect 243780 219960 243786 219972
rect 262122 219960 262128 219972
rect 243780 219932 262128 219960
rect 243780 219920 243786 219932
rect 262122 219920 262128 219932
rect 262180 219920 262186 219972
rect 428090 219920 428096 219972
rect 428148 219960 428154 219972
rect 451918 219960 451924 219972
rect 428148 219932 451924 219960
rect 428148 219920 428154 219932
rect 451918 219920 451924 219932
rect 451976 219920 451982 219972
rect 455690 219920 455696 219972
rect 455748 219960 455754 219972
rect 507762 219960 507768 219972
rect 455748 219932 507768 219960
rect 455748 219920 455754 219932
rect 507762 219920 507768 219932
rect 507820 219920 507826 219972
rect 530394 219852 530400 219904
rect 530452 219892 530458 219904
rect 562318 219892 562324 219904
rect 530452 219864 562324 219892
rect 530452 219852 530458 219864
rect 562318 219852 562324 219864
rect 562376 219852 562382 219904
rect 562502 219852 562508 219904
rect 562560 219892 562566 219904
rect 562870 219892 562876 219904
rect 562560 219864 562876 219892
rect 562560 219852 562566 219864
rect 562870 219852 562876 219864
rect 562928 219852 562934 219904
rect 563054 219852 563060 219904
rect 563112 219892 563118 219904
rect 567930 219892 567936 219904
rect 563112 219864 567936 219892
rect 563112 219852 563118 219864
rect 567930 219852 567936 219864
rect 567988 219852 567994 219904
rect 574922 219892 574928 219904
rect 568132 219864 574928 219892
rect 136910 219824 136916 219836
rect 122806 219796 136916 219824
rect 136910 219784 136916 219796
rect 136968 219784 136974 219836
rect 137094 219784 137100 219836
rect 137152 219824 137158 219836
rect 142062 219824 142068 219836
rect 137152 219796 142068 219824
rect 137152 219784 137158 219796
rect 142062 219784 142068 219796
rect 142120 219784 142126 219836
rect 142246 219784 142252 219836
rect 142304 219824 142310 219836
rect 195330 219824 195336 219836
rect 142304 219796 195336 219824
rect 142304 219784 142310 219796
rect 195330 219784 195336 219796
rect 195388 219784 195394 219836
rect 195882 219784 195888 219836
rect 195940 219824 195946 219836
rect 197446 219824 197452 219836
rect 195940 219796 197452 219824
rect 195940 219784 195946 219796
rect 197446 219784 197452 219796
rect 197504 219784 197510 219836
rect 201586 219784 201592 219836
rect 201644 219824 201650 219836
rect 205082 219824 205088 219836
rect 201644 219796 205088 219824
rect 201644 219784 201650 219796
rect 205082 219784 205088 219796
rect 205140 219784 205146 219836
rect 206646 219784 206652 219836
rect 206704 219824 206710 219836
rect 209682 219824 209688 219836
rect 206704 219796 209688 219824
rect 206704 219784 206710 219796
rect 209682 219784 209688 219796
rect 209740 219784 209746 219836
rect 209866 219784 209872 219836
rect 209924 219824 209930 219836
rect 211430 219824 211436 219836
rect 209924 219796 211436 219824
rect 209924 219784 209930 219796
rect 211430 219784 211436 219796
rect 211488 219784 211494 219836
rect 211614 219784 211620 219836
rect 211672 219824 211678 219836
rect 214374 219824 214380 219836
rect 211672 219796 214380 219824
rect 211672 219784 211678 219796
rect 214374 219784 214380 219796
rect 214432 219784 214438 219836
rect 214558 219784 214564 219836
rect 214616 219824 214622 219836
rect 243354 219824 243360 219836
rect 214616 219796 243360 219824
rect 214616 219784 214622 219796
rect 243354 219784 243360 219796
rect 243412 219784 243418 219836
rect 442994 219824 443000 219836
rect 431926 219796 443000 219824
rect 322566 219716 322572 219768
rect 322624 219756 322630 219768
rect 325970 219756 325976 219768
rect 322624 219728 325976 219756
rect 322624 219716 322630 219728
rect 325970 219716 325976 219728
rect 326028 219716 326034 219768
rect 70854 219648 70860 219700
rect 70912 219688 70918 219700
rect 143074 219688 143080 219700
rect 70912 219660 143080 219688
rect 70912 219648 70918 219660
rect 143074 219648 143080 219660
rect 143132 219648 143138 219700
rect 143258 219648 143264 219700
rect 143316 219688 143322 219700
rect 154482 219688 154488 219700
rect 143316 219660 154488 219688
rect 143316 219648 143322 219660
rect 154482 219648 154488 219660
rect 154540 219648 154546 219700
rect 154666 219648 154672 219700
rect 154724 219688 154730 219700
rect 156782 219688 156788 219700
rect 154724 219660 156788 219688
rect 154724 219648 154730 219660
rect 156782 219648 156788 219660
rect 156840 219648 156846 219700
rect 156966 219648 156972 219700
rect 157024 219688 157030 219700
rect 202322 219688 202328 219700
rect 157024 219660 202328 219688
rect 157024 219648 157030 219660
rect 202322 219648 202328 219660
rect 202380 219648 202386 219700
rect 202506 219648 202512 219700
rect 202564 219688 202570 219700
rect 205266 219688 205272 219700
rect 202564 219660 205272 219688
rect 202564 219648 202570 219660
rect 205266 219648 205272 219660
rect 205324 219648 205330 219700
rect 205910 219648 205916 219700
rect 205968 219688 205974 219700
rect 207198 219688 207204 219700
rect 205968 219660 207204 219688
rect 205968 219648 205974 219660
rect 207198 219648 207204 219660
rect 207256 219648 207262 219700
rect 209682 219648 209688 219700
rect 209740 219688 209746 219700
rect 248138 219688 248144 219700
rect 209740 219660 248144 219688
rect 209740 219648 209746 219660
rect 248138 219648 248144 219660
rect 248196 219648 248202 219700
rect 254670 219648 254676 219700
rect 254728 219688 254734 219700
rect 256510 219688 256516 219700
rect 254728 219660 256516 219688
rect 254728 219648 254734 219660
rect 256510 219648 256516 219660
rect 256568 219648 256574 219700
rect 421098 219648 421104 219700
rect 421156 219688 421162 219700
rect 431926 219688 431954 219796
rect 442994 219784 443000 219796
rect 443052 219784 443058 219836
rect 460198 219824 460204 219836
rect 446416 219796 460204 219824
rect 421156 219660 431954 219688
rect 421156 219648 421162 219660
rect 436738 219648 436744 219700
rect 436796 219688 436802 219700
rect 446416 219688 446444 219796
rect 460198 219784 460204 219796
rect 460256 219784 460262 219836
rect 463878 219784 463884 219836
rect 463936 219824 463942 219836
rect 470962 219824 470968 219836
rect 463936 219796 470968 219824
rect 463936 219784 463942 219796
rect 470962 219784 470968 219796
rect 471020 219784 471026 219836
rect 471422 219784 471428 219836
rect 471480 219824 471486 219836
rect 474458 219824 474464 219836
rect 471480 219796 474464 219824
rect 471480 219784 471486 219796
rect 474458 219784 474464 219796
rect 474516 219784 474522 219836
rect 505094 219824 505100 219836
rect 475396 219796 505100 219824
rect 465994 219688 466000 219700
rect 436796 219660 446444 219688
rect 446508 219660 466000 219688
rect 436796 219648 436802 219660
rect 264606 219580 264612 219632
rect 264664 219620 264670 219632
rect 270218 219620 270224 219632
rect 264664 219592 270224 219620
rect 264664 219580 264670 219592
rect 270218 219580 270224 219592
rect 270276 219580 270282 219632
rect 311618 219580 311624 219632
rect 311676 219620 311682 219632
rect 317782 219620 317788 219632
rect 311676 219592 317788 219620
rect 311676 219580 311682 219592
rect 317782 219580 317788 219592
rect 317840 219580 317846 219632
rect 324222 219580 324228 219632
rect 324280 219620 324286 219632
rect 327718 219620 327724 219632
rect 324280 219592 327724 219620
rect 324280 219580 324286 219592
rect 327718 219580 327724 219592
rect 327776 219580 327782 219632
rect 88886 219512 88892 219564
rect 88944 219552 88950 219564
rect 160922 219552 160928 219564
rect 88944 219524 160928 219552
rect 88944 219512 88950 219524
rect 160922 219512 160928 219524
rect 160980 219512 160986 219564
rect 161290 219512 161296 219564
rect 161348 219552 161354 219564
rect 162578 219552 162584 219564
rect 161348 219524 162584 219552
rect 161348 219512 161354 219524
rect 162578 219512 162584 219524
rect 162636 219512 162642 219564
rect 163590 219512 163596 219564
rect 163648 219552 163654 219564
rect 166902 219552 166908 219564
rect 163648 219524 166908 219552
rect 163648 219512 163654 219524
rect 166902 219512 166908 219524
rect 166960 219512 166966 219564
rect 169386 219512 169392 219564
rect 169444 219552 169450 219564
rect 173802 219552 173808 219564
rect 169444 219524 173808 219552
rect 169444 219512 169450 219524
rect 173802 219512 173808 219524
rect 173860 219512 173866 219564
rect 174170 219512 174176 219564
rect 174228 219552 174234 219564
rect 176562 219552 176568 219564
rect 174228 219524 176568 219552
rect 174228 219512 174234 219524
rect 176562 219512 176568 219524
rect 176620 219512 176626 219564
rect 177666 219512 177672 219564
rect 177724 219552 177730 219564
rect 180518 219552 180524 219564
rect 177724 219524 180524 219552
rect 177724 219512 177730 219524
rect 180518 219512 180524 219524
rect 180576 219512 180582 219564
rect 181162 219512 181168 219564
rect 181220 219552 181226 219564
rect 183278 219552 183284 219564
rect 181220 219524 183284 219552
rect 181220 219512 181226 219524
rect 183278 219512 183284 219524
rect 183336 219512 183342 219564
rect 183462 219512 183468 219564
rect 183520 219552 183526 219564
rect 187786 219552 187792 219564
rect 183520 219524 187792 219552
rect 183520 219512 183526 219524
rect 187786 219512 187792 219524
rect 187844 219512 187850 219564
rect 187970 219512 187976 219564
rect 188028 219552 188034 219564
rect 193030 219552 193036 219564
rect 188028 219524 193036 219552
rect 188028 219512 188034 219524
rect 193030 219512 193036 219524
rect 193088 219512 193094 219564
rect 193186 219524 223896 219552
rect 118050 219376 118056 219428
rect 118108 219416 118114 219428
rect 188154 219416 188160 219428
rect 118108 219388 188160 219416
rect 118108 219376 118114 219388
rect 188154 219376 188160 219388
rect 188212 219376 188218 219428
rect 190086 219376 190092 219428
rect 190144 219416 190150 219428
rect 193186 219416 193214 219524
rect 190144 219388 193214 219416
rect 190144 219376 190150 219388
rect 196710 219376 196716 219428
rect 196768 219416 196774 219428
rect 201586 219416 201592 219428
rect 196768 219388 201592 219416
rect 196768 219376 196774 219388
rect 201586 219376 201592 219388
rect 201644 219376 201650 219428
rect 204622 219376 204628 219428
rect 204680 219416 204686 219428
rect 210418 219416 210424 219428
rect 204680 219388 210424 219416
rect 204680 219376 204686 219388
rect 210418 219376 210424 219388
rect 210476 219376 210482 219428
rect 223868 219348 223896 219524
rect 423766 219512 423772 219564
rect 423824 219552 423830 219564
rect 445294 219552 445300 219564
rect 423824 219524 445300 219552
rect 423824 219512 423830 219524
rect 445294 219512 445300 219524
rect 445352 219512 445358 219564
rect 445662 219512 445668 219564
rect 445720 219552 445726 219564
rect 446508 219552 446536 219660
rect 465994 219648 466000 219660
rect 466052 219648 466058 219700
rect 466454 219648 466460 219700
rect 466512 219688 466518 219700
rect 475396 219688 475424 219796
rect 505094 219784 505100 219796
rect 505152 219784 505158 219836
rect 506566 219784 506572 219836
rect 506624 219824 506630 219836
rect 509970 219824 509976 219836
rect 506624 219796 509976 219824
rect 506624 219784 506630 219796
rect 509970 219784 509976 219796
rect 510028 219784 510034 219836
rect 521654 219716 521660 219768
rect 521712 219756 521718 219768
rect 522574 219756 522580 219768
rect 521712 219728 522580 219756
rect 521712 219716 521718 219728
rect 522574 219716 522580 219728
rect 522632 219756 522638 219768
rect 568132 219756 568160 219864
rect 574922 219852 574928 219864
rect 574980 219852 574986 219904
rect 575290 219852 575296 219904
rect 575348 219892 575354 219904
rect 610342 219892 610348 219904
rect 575348 219864 610348 219892
rect 575348 219852 575354 219864
rect 610342 219852 610348 219864
rect 610400 219852 610406 219904
rect 522632 219728 568160 219756
rect 522632 219716 522638 219728
rect 568298 219716 568304 219768
rect 568356 219756 568362 219768
rect 575658 219756 575664 219768
rect 568356 219728 575664 219756
rect 568356 219716 568362 219728
rect 575658 219716 575664 219728
rect 575716 219716 575722 219768
rect 575842 219716 575848 219768
rect 575900 219756 575906 219768
rect 597554 219756 597560 219768
rect 575900 219728 597560 219756
rect 575900 219716 575906 219728
rect 597554 219716 597560 219728
rect 597612 219716 597618 219768
rect 666002 219716 666008 219768
rect 666060 219756 666066 219768
rect 675294 219756 675300 219768
rect 666060 219728 675300 219756
rect 666060 219716 666066 219728
rect 675294 219716 675300 219728
rect 675352 219716 675358 219768
rect 466512 219660 475424 219688
rect 466512 219648 466518 219660
rect 475562 219648 475568 219700
rect 475620 219688 475626 219700
rect 475620 219660 495434 219688
rect 475620 219648 475626 219660
rect 445720 219524 446536 219552
rect 445720 219512 445726 219524
rect 449066 219512 449072 219564
rect 449124 219552 449130 219564
rect 453574 219552 453580 219564
rect 449124 219524 453580 219552
rect 449124 219512 449130 219524
rect 453574 219512 453580 219524
rect 453632 219512 453638 219564
rect 459738 219512 459744 219564
rect 459796 219552 459802 219564
rect 459796 219524 476436 219552
rect 459796 219512 459802 219524
rect 231670 219484 231676 219496
rect 226444 219456 228036 219484
rect 226444 219348 226472 219456
rect 223868 219320 226472 219348
rect 228008 219348 228036 219456
rect 229020 219456 231676 219484
rect 229020 219348 229048 219456
rect 231670 219444 231676 219456
rect 231728 219444 231734 219496
rect 238110 219444 238116 219496
rect 238168 219484 238174 219496
rect 240042 219484 240048 219496
rect 238168 219456 240048 219484
rect 238168 219444 238174 219456
rect 240042 219444 240048 219456
rect 240100 219444 240106 219496
rect 248046 219444 248052 219496
rect 248104 219484 248110 219496
rect 249702 219484 249708 219496
rect 248104 219456 249708 219484
rect 248104 219444 248110 219456
rect 249702 219444 249708 219456
rect 249760 219444 249766 219496
rect 294414 219444 294420 219496
rect 294472 219484 294478 219496
rect 298002 219484 298008 219496
rect 294472 219456 298008 219484
rect 294472 219444 294478 219456
rect 298002 219444 298008 219456
rect 298060 219444 298066 219496
rect 306006 219444 306012 219496
rect 306064 219484 306070 219496
rect 307478 219484 307484 219496
rect 306064 219456 307484 219484
rect 306064 219444 306070 219456
rect 307478 219444 307484 219456
rect 307536 219444 307542 219496
rect 325050 219444 325056 219496
rect 325108 219484 325114 219496
rect 326522 219484 326528 219496
rect 325108 219456 326528 219484
rect 325108 219444 325114 219456
rect 326522 219444 326528 219456
rect 326580 219444 326586 219496
rect 340690 219444 340696 219496
rect 340748 219484 340754 219496
rect 345934 219484 345940 219496
rect 340748 219456 345940 219484
rect 340748 219444 340754 219456
rect 345934 219444 345940 219456
rect 345992 219444 345998 219496
rect 348878 219444 348884 219496
rect 348936 219484 348942 219496
rect 355042 219484 355048 219496
rect 348936 219456 355048 219484
rect 348936 219444 348942 219456
rect 355042 219444 355048 219456
rect 355100 219444 355106 219496
rect 430390 219376 430396 219428
rect 430448 219416 430454 219428
rect 475930 219416 475936 219428
rect 430448 219388 475936 219416
rect 430448 219376 430454 219388
rect 475930 219376 475936 219388
rect 475988 219376 475994 219428
rect 476408 219416 476436 219524
rect 476574 219512 476580 219564
rect 476632 219552 476638 219564
rect 481450 219552 481456 219564
rect 476632 219524 481456 219552
rect 476632 219512 476638 219524
rect 481450 219512 481456 219524
rect 481508 219512 481514 219564
rect 485866 219512 485872 219564
rect 485924 219552 485930 219564
rect 495250 219552 495256 219564
rect 485924 219524 495256 219552
rect 485924 219512 485930 219524
rect 495250 219512 495256 219524
rect 495308 219512 495314 219564
rect 495406 219552 495434 219660
rect 495526 219648 495532 219700
rect 495584 219688 495590 219700
rect 504542 219688 504548 219700
rect 495584 219660 504548 219688
rect 495584 219648 495590 219660
rect 504542 219648 504548 219660
rect 504600 219648 504606 219700
rect 504726 219648 504732 219700
rect 504784 219688 504790 219700
rect 504784 219660 505094 219688
rect 504784 219648 504790 219660
rect 505066 219620 505094 219660
rect 506198 219620 506204 219632
rect 505066 219592 506204 219620
rect 506198 219580 506204 219592
rect 506256 219580 506262 219632
rect 527818 219580 527824 219632
rect 527876 219620 527882 219632
rect 563054 219620 563060 219632
rect 527876 219592 563060 219620
rect 527876 219580 527882 219592
rect 563054 219580 563060 219592
rect 563112 219580 563118 219632
rect 563348 219592 576854 219620
rect 499942 219552 499948 219564
rect 495406 219524 499948 219552
rect 499942 219512 499948 219524
rect 500000 219512 500006 219564
rect 563348 219552 563376 219592
rect 563256 219524 563376 219552
rect 535362 219484 535368 219496
rect 481652 219456 485774 219484
rect 476758 219416 476764 219428
rect 476408 219388 476764 219416
rect 476758 219376 476764 219388
rect 476816 219376 476822 219428
rect 479886 219376 479892 219428
rect 479944 219416 479950 219428
rect 481652 219416 481680 219456
rect 479944 219388 481680 219416
rect 485746 219416 485774 219456
rect 501248 219456 535368 219484
rect 490098 219416 490104 219428
rect 485746 219388 490104 219416
rect 479944 219376 479950 219388
rect 490098 219376 490104 219388
rect 490156 219376 490162 219428
rect 228008 219320 229048 219348
rect 496814 219308 496820 219360
rect 496872 219348 496878 219360
rect 501248 219348 501276 219456
rect 535362 219444 535368 219456
rect 535420 219444 535426 219496
rect 537478 219444 537484 219496
rect 537536 219484 537542 219496
rect 548334 219484 548340 219496
rect 537536 219456 548340 219484
rect 537536 219444 537542 219456
rect 548334 219444 548340 219456
rect 548392 219444 548398 219496
rect 549990 219444 549996 219496
rect 550048 219484 550054 219496
rect 563256 219484 563284 219524
rect 572162 219484 572168 219496
rect 550048 219456 563284 219484
rect 563532 219456 572168 219484
rect 550048 219444 550054 219456
rect 496872 219320 501276 219348
rect 496872 219308 496878 219320
rect 112898 219240 112904 219292
rect 112956 219280 112962 219292
rect 185394 219280 185400 219292
rect 112956 219252 185400 219280
rect 112956 219240 112962 219252
rect 185394 219240 185400 219252
rect 185452 219240 185458 219292
rect 431586 219240 431592 219292
rect 431644 219280 431650 219292
rect 475746 219280 475752 219292
rect 431644 219252 475752 219280
rect 431644 219240 431650 219252
rect 475746 219240 475752 219252
rect 475804 219240 475810 219292
rect 483566 219240 483572 219292
rect 483624 219280 483630 219292
rect 485774 219280 485780 219292
rect 483624 219252 485780 219280
rect 483624 219240 483630 219252
rect 485774 219240 485780 219252
rect 485832 219240 485838 219292
rect 515582 219240 515588 219292
rect 515640 219280 515646 219292
rect 563054 219280 563060 219292
rect 515640 219252 563060 219280
rect 515640 219240 515646 219252
rect 563054 219240 563060 219252
rect 563112 219240 563118 219292
rect 563238 219240 563244 219292
rect 563296 219280 563302 219292
rect 563532 219280 563560 219456
rect 572162 219444 572168 219456
rect 572220 219444 572226 219496
rect 575290 219484 575296 219496
rect 572548 219456 575296 219484
rect 572548 219416 572576 219456
rect 575290 219444 575296 219456
rect 575348 219444 575354 219496
rect 576826 219484 576854 219592
rect 665082 219580 665088 219632
rect 665140 219620 665146 219632
rect 675478 219620 675484 219632
rect 665140 219592 675484 219620
rect 665140 219580 665146 219592
rect 675478 219580 675484 219592
rect 675536 219580 675542 219632
rect 624142 219484 624148 219496
rect 576826 219456 624148 219484
rect 624142 219444 624148 219456
rect 624200 219444 624206 219496
rect 572318 219388 572576 219416
rect 564066 219308 564072 219360
rect 564124 219348 564130 219360
rect 572318 219348 572346 219388
rect 564124 219320 572346 219348
rect 564124 219308 564130 219320
rect 563296 219252 563560 219280
rect 563296 219240 563302 219252
rect 572990 219240 572996 219292
rect 573048 219280 573054 219292
rect 609238 219280 609244 219292
rect 573048 219252 609244 219280
rect 573048 219240 573054 219252
rect 609238 219240 609244 219252
rect 609296 219240 609302 219292
rect 486418 219172 486424 219224
rect 486476 219212 486482 219224
rect 498286 219212 498292 219224
rect 486476 219184 498292 219212
rect 486476 219172 486482 219184
rect 498286 219172 498292 219184
rect 498344 219172 498350 219224
rect 112254 219104 112260 219156
rect 112312 219144 112318 219156
rect 186590 219144 186596 219156
rect 112312 219116 186596 219144
rect 112312 219104 112318 219116
rect 186590 219104 186596 219116
rect 186648 219104 186654 219156
rect 431770 219104 431776 219156
rect 431828 219144 431834 219156
rect 476068 219144 476074 219156
rect 431828 219116 476074 219144
rect 431828 219104 431834 219116
rect 476068 219104 476074 219116
rect 476126 219104 476132 219156
rect 484670 219104 484676 219156
rect 484728 219144 484734 219156
rect 485038 219144 485044 219156
rect 484728 219116 485044 219144
rect 484728 219104 484734 219116
rect 485038 219104 485044 219116
rect 485096 219104 485102 219156
rect 501046 219104 501052 219156
rect 501104 219144 501110 219156
rect 596082 219144 596088 219156
rect 501104 219116 596088 219144
rect 501104 219104 501110 219116
rect 596082 219104 596088 219116
rect 596140 219104 596146 219156
rect 596266 219104 596272 219156
rect 596324 219144 596330 219156
rect 627822 219144 627828 219156
rect 596324 219116 627828 219144
rect 596324 219104 596330 219116
rect 627822 219104 627828 219116
rect 627880 219104 627886 219156
rect 628006 219104 628012 219156
rect 628064 219144 628070 219156
rect 628834 219144 628840 219156
rect 628064 219116 628840 219144
rect 628064 219104 628070 219116
rect 628834 219104 628840 219116
rect 628892 219104 628898 219156
rect 486142 219036 486148 219088
rect 486200 219076 486206 219088
rect 494054 219076 494060 219088
rect 486200 219048 494060 219076
rect 486200 219036 486206 219048
rect 494054 219036 494060 219048
rect 494112 219036 494118 219088
rect 104802 218968 104808 219020
rect 104860 219008 104866 219020
rect 176194 219008 176200 219020
rect 104860 218980 176200 219008
rect 104860 218968 104866 218980
rect 176194 218968 176200 218980
rect 176252 218968 176258 219020
rect 176562 218968 176568 219020
rect 176620 219008 176626 219020
rect 181162 219008 181168 219020
rect 176620 218980 181168 219008
rect 176620 218968 176626 218980
rect 181162 218968 181168 218980
rect 181220 218968 181226 219020
rect 434346 218968 434352 219020
rect 434404 219008 434410 219020
rect 485958 219008 485964 219020
rect 434404 218980 485964 219008
rect 434404 218968 434410 218980
rect 485958 218968 485964 218980
rect 486016 218968 486022 219020
rect 503162 218968 503168 219020
rect 503220 219008 503226 219020
rect 503622 219008 503628 219020
rect 503220 218980 503628 219008
rect 503220 218968 503226 218980
rect 503622 218968 503628 218980
rect 503680 219008 503686 219020
rect 587894 219008 587900 219020
rect 503680 218980 587900 219008
rect 503680 218968 503686 218980
rect 587894 218968 587900 218980
rect 587952 218968 587958 219020
rect 591298 218968 591304 219020
rect 591356 219008 591362 219020
rect 617242 219008 617248 219020
rect 591356 218980 617248 219008
rect 591356 218968 591362 218980
rect 617242 218968 617248 218980
rect 617300 218968 617306 219020
rect 106182 218832 106188 218884
rect 106240 218872 106246 218884
rect 180978 218872 180984 218884
rect 106240 218844 180984 218872
rect 106240 218832 106246 218844
rect 180978 218832 180984 218844
rect 181036 218832 181042 218884
rect 448054 218832 448060 218884
rect 448112 218872 448118 218884
rect 506566 218872 506572 218884
rect 448112 218844 506572 218872
rect 448112 218832 448118 218844
rect 506566 218832 506572 218844
rect 506624 218832 506630 218884
rect 539594 218832 539600 218884
rect 539652 218872 539658 218884
rect 546126 218872 546132 218884
rect 539652 218844 546132 218872
rect 539652 218832 539658 218844
rect 546126 218832 546132 218844
rect 546184 218832 546190 218884
rect 546310 218832 546316 218884
rect 546368 218872 546374 218884
rect 548518 218872 548524 218884
rect 546368 218844 548524 218872
rect 546368 218832 546374 218844
rect 548518 218832 548524 218844
rect 548576 218832 548582 218884
rect 552290 218832 552296 218884
rect 552348 218872 552354 218884
rect 625522 218872 625528 218884
rect 552348 218844 625528 218872
rect 552348 218832 552354 218844
rect 625522 218832 625528 218844
rect 625580 218832 625586 218884
rect 105630 218696 105636 218748
rect 105688 218736 105694 218748
rect 175826 218736 175832 218748
rect 105688 218708 175832 218736
rect 105688 218696 105694 218708
rect 175826 218696 175832 218708
rect 175884 218696 175890 218748
rect 176194 218696 176200 218748
rect 176252 218736 176258 218748
rect 179690 218736 179696 218748
rect 176252 218708 179696 218736
rect 176252 218696 176258 218708
rect 179690 218696 179696 218708
rect 179748 218696 179754 218748
rect 445478 218696 445484 218748
rect 445536 218736 445542 218748
rect 445536 218708 476114 218736
rect 445536 218696 445542 218708
rect 132954 218560 132960 218612
rect 133012 218600 133018 218612
rect 199010 218600 199016 218612
rect 133012 218572 199016 218600
rect 133012 218560 133018 218572
rect 199010 218560 199016 218572
rect 199068 218560 199074 218612
rect 136266 218424 136272 218476
rect 136324 218464 136330 218476
rect 200390 218464 200396 218476
rect 136324 218436 200396 218464
rect 136324 218424 136330 218436
rect 200390 218424 200396 218436
rect 200448 218424 200454 218476
rect 476086 218464 476114 218708
rect 476390 218696 476396 218748
rect 476448 218736 476454 218748
rect 481726 218736 481732 218748
rect 476448 218708 481732 218736
rect 476448 218696 476454 218708
rect 481726 218696 481732 218708
rect 481784 218696 481790 218748
rect 504358 218736 504364 218748
rect 485746 218708 504364 218736
rect 485746 218464 485774 218708
rect 504358 218696 504364 218708
rect 504416 218696 504422 218748
rect 528554 218696 528560 218748
rect 528612 218736 528618 218748
rect 597370 218736 597376 218748
rect 528612 218708 597376 218736
rect 528612 218696 528618 218708
rect 597370 218696 597376 218708
rect 597428 218696 597434 218748
rect 597554 218696 597560 218748
rect 597612 218736 597618 218748
rect 621658 218736 621664 218748
rect 597612 218708 621664 218736
rect 597612 218696 597618 218708
rect 621658 218696 621664 218708
rect 621716 218696 621722 218748
rect 508498 218560 508504 218612
rect 508556 218600 508562 218612
rect 598474 218600 598480 218612
rect 508556 218572 598480 218600
rect 508556 218560 508562 218572
rect 598474 218560 598480 218572
rect 598532 218560 598538 218612
rect 476086 218436 485774 218464
rect 498286 218424 498292 218476
rect 498344 218464 498350 218476
rect 587526 218464 587532 218476
rect 498344 218436 587532 218464
rect 498344 218424 498350 218436
rect 587526 218424 587532 218436
rect 587584 218424 587590 218476
rect 591298 218464 591304 218476
rect 587728 218436 591304 218464
rect 146202 218288 146208 218340
rect 146260 218328 146266 218340
rect 207750 218328 207756 218340
rect 146260 218300 207756 218328
rect 146260 218288 146266 218300
rect 207750 218288 207756 218300
rect 207808 218288 207814 218340
rect 494054 218288 494060 218340
rect 494112 218328 494118 218340
rect 495250 218328 495256 218340
rect 494112 218300 495256 218328
rect 494112 218288 494118 218300
rect 495250 218288 495256 218300
rect 495308 218328 495314 218340
rect 571794 218328 571800 218340
rect 495308 218300 571800 218328
rect 495308 218288 495314 218300
rect 571794 218288 571800 218300
rect 571852 218288 571858 218340
rect 572438 218288 572444 218340
rect 572496 218328 572502 218340
rect 580350 218328 580356 218340
rect 572496 218300 580356 218328
rect 572496 218288 572502 218300
rect 580350 218288 580356 218300
rect 580408 218288 580414 218340
rect 581638 218288 581644 218340
rect 581696 218328 581702 218340
rect 587728 218328 587756 218436
rect 591298 218424 591304 218436
rect 591356 218424 591362 218476
rect 597370 218424 597376 218476
rect 597428 218464 597434 218476
rect 597922 218464 597928 218476
rect 597428 218436 597928 218464
rect 597428 218424 597434 218436
rect 597922 218424 597928 218436
rect 597980 218424 597986 218476
rect 581696 218300 587756 218328
rect 581696 218288 581702 218300
rect 587894 218288 587900 218340
rect 587952 218328 587958 218340
rect 597554 218328 597560 218340
rect 587952 218300 597560 218328
rect 587952 218288 587958 218300
rect 597554 218288 597560 218300
rect 597612 218288 597618 218340
rect 147582 218152 147588 218204
rect 147640 218192 147646 218204
rect 207014 218192 207020 218204
rect 147640 218164 207020 218192
rect 147640 218152 147646 218164
rect 207014 218152 207020 218164
rect 207072 218152 207078 218204
rect 510706 218152 510712 218204
rect 510764 218192 510770 218204
rect 599026 218192 599032 218204
rect 510764 218164 599032 218192
rect 510764 218152 510770 218164
rect 599026 218152 599032 218164
rect 599084 218152 599090 218204
rect 175826 218016 175832 218068
rect 175884 218056 175890 218068
rect 182542 218056 182548 218068
rect 175884 218028 182548 218056
rect 175884 218016 175890 218028
rect 182542 218016 182548 218028
rect 182600 218016 182606 218068
rect 491662 218016 491668 218068
rect 491720 218056 491726 218068
rect 563008 218056 563014 218068
rect 491720 218028 563014 218056
rect 491720 218016 491726 218028
rect 563008 218016 563014 218028
rect 563066 218016 563072 218068
rect 563146 218016 563152 218068
rect 563204 218056 563210 218068
rect 573358 218056 573364 218068
rect 563204 218028 573364 218056
rect 563204 218016 563210 218028
rect 573358 218016 573364 218028
rect 573416 218016 573422 218068
rect 574462 218016 574468 218068
rect 574520 218056 574526 218068
rect 581638 218056 581644 218068
rect 574520 218028 581644 218056
rect 574520 218016 574526 218028
rect 581638 218016 581644 218028
rect 581696 218016 581702 218068
rect 587526 218016 587532 218068
rect 587584 218056 587590 218068
rect 595346 218056 595352 218068
rect 587584 218028 595352 218056
rect 587584 218016 587590 218028
rect 595346 218016 595352 218028
rect 595404 218016 595410 218068
rect 596174 218016 596180 218068
rect 596232 218056 596238 218068
rect 596818 218056 596824 218068
rect 596232 218028 596824 218056
rect 596232 218016 596238 218028
rect 596818 218016 596824 218028
rect 596876 218016 596882 218068
rect 488534 217880 488540 217932
rect 488592 217920 488598 217932
rect 594794 217920 594800 217932
rect 488592 217892 594800 217920
rect 488592 217880 488598 217892
rect 594794 217880 594800 217892
rect 594852 217880 594858 217932
rect 188430 217812 188436 217864
rect 188488 217852 188494 217864
rect 188982 217852 188988 217864
rect 188488 217824 188988 217852
rect 188488 217812 188494 217824
rect 188982 217812 188988 217824
rect 189040 217812 189046 217864
rect 190914 217812 190920 217864
rect 190972 217852 190978 217864
rect 191742 217852 191748 217864
rect 190972 217824 191748 217852
rect 190972 217812 190978 217824
rect 191742 217812 191748 217824
rect 191800 217812 191806 217864
rect 340966 217812 340972 217864
rect 341024 217852 341030 217864
rect 341794 217852 341800 217864
rect 341024 217824 341800 217852
rect 341024 217812 341030 217824
rect 341794 217812 341800 217824
rect 341852 217812 341858 217864
rect 343910 217812 343916 217864
rect 343968 217852 343974 217864
rect 344278 217852 344284 217864
rect 343968 217824 344284 217852
rect 343968 217812 343974 217824
rect 344278 217812 344284 217824
rect 344336 217812 344342 217864
rect 373994 217812 374000 217864
rect 374052 217852 374058 217864
rect 374914 217852 374920 217864
rect 374052 217824 374920 217852
rect 374052 217812 374058 217824
rect 374914 217812 374920 217824
rect 374972 217812 374978 217864
rect 382458 217812 382464 217864
rect 382516 217852 382522 217864
rect 383194 217852 383200 217864
rect 382516 217824 383200 217852
rect 382516 217812 382522 217824
rect 383194 217812 383200 217824
rect 383252 217812 383258 217864
rect 390738 217812 390744 217864
rect 390796 217852 390802 217864
rect 391474 217852 391480 217864
rect 390796 217824 391480 217852
rect 390796 217812 390802 217824
rect 391474 217812 391480 217824
rect 391532 217812 391538 217864
rect 393314 217812 393320 217864
rect 393372 217852 393378 217864
rect 393958 217852 393964 217864
rect 393372 217824 393964 217852
rect 393372 217812 393378 217824
rect 393958 217812 393964 217824
rect 394016 217812 394022 217864
rect 398834 217812 398840 217864
rect 398892 217852 398898 217864
rect 399754 217852 399760 217864
rect 398892 217824 399760 217852
rect 398892 217812 398898 217824
rect 399754 217812 399760 217824
rect 399812 217812 399818 217864
rect 402974 217812 402980 217864
rect 403032 217852 403038 217864
rect 403894 217852 403900 217864
rect 403032 217824 403900 217852
rect 403032 217812 403038 217824
rect 403894 217812 403900 217824
rect 403952 217812 403958 217864
rect 419534 217812 419540 217864
rect 419592 217852 419598 217864
rect 420454 217852 420460 217864
rect 419592 217824 420460 217852
rect 419592 217812 419598 217824
rect 420454 217812 420460 217824
rect 420512 217812 420518 217864
rect 426434 217812 426440 217864
rect 426492 217852 426498 217864
rect 427078 217852 427084 217864
rect 426492 217824 427084 217852
rect 426492 217812 426498 217824
rect 427078 217812 427084 217824
rect 427136 217812 427142 217864
rect 541710 217744 541716 217796
rect 541768 217784 541774 217796
rect 542722 217784 542728 217796
rect 541768 217756 542728 217784
rect 541768 217744 541774 217756
rect 542722 217744 542728 217756
rect 542780 217744 542786 217796
rect 543090 217744 543096 217796
rect 543148 217784 543154 217796
rect 544378 217784 544384 217796
rect 543148 217756 544384 217784
rect 543148 217744 543154 217756
rect 544378 217744 544384 217756
rect 544436 217744 544442 217796
rect 546310 217784 546316 217796
rect 545086 217756 546316 217784
rect 475930 217608 475936 217660
rect 475988 217648 475994 217660
rect 477908 217648 477914 217660
rect 475988 217620 477914 217648
rect 475988 217608 475994 217620
rect 477908 217608 477914 217620
rect 477966 217608 477972 217660
rect 514754 217608 514760 217660
rect 514812 217648 514818 217660
rect 515996 217648 516002 217660
rect 514812 217620 516002 217648
rect 514812 217608 514818 217620
rect 515996 217608 516002 217620
rect 516054 217608 516060 217660
rect 519170 217608 519176 217660
rect 519228 217648 519234 217660
rect 520136 217648 520142 217660
rect 519228 217620 520142 217648
rect 519228 217608 519234 217620
rect 520136 217608 520142 217620
rect 520194 217608 520200 217660
rect 537662 217608 537668 217660
rect 537720 217648 537726 217660
rect 545086 217648 545114 217756
rect 546310 217744 546316 217756
rect 546368 217744 546374 217796
rect 548518 217744 548524 217796
rect 548576 217784 548582 217796
rect 553486 217784 553492 217796
rect 548576 217756 553492 217784
rect 548576 217744 548582 217756
rect 553486 217744 553492 217756
rect 553544 217744 553550 217796
rect 556798 217744 556804 217796
rect 556856 217784 556862 217796
rect 607858 217784 607864 217796
rect 556856 217756 607864 217784
rect 556856 217744 556862 217756
rect 607858 217744 607864 217756
rect 607916 217744 607922 217796
rect 537720 217620 545114 217648
rect 537720 217608 537726 217620
rect 545574 217608 545580 217660
rect 545632 217648 545638 217660
rect 570414 217648 570420 217660
rect 545632 217620 570420 217648
rect 545632 217608 545638 217620
rect 570414 217608 570420 217620
rect 570472 217608 570478 217660
rect 573358 217608 573364 217660
rect 573416 217648 573422 217660
rect 609882 217648 609888 217660
rect 573416 217620 609888 217648
rect 573416 217608 573422 217620
rect 609882 217608 609888 217620
rect 609940 217608 609946 217660
rect 475746 217472 475752 217524
rect 475804 217512 475810 217524
rect 481220 217512 481226 217524
rect 475804 217484 481226 217512
rect 475804 217472 475810 217484
rect 481220 217472 481226 217484
rect 481278 217472 481284 217524
rect 538674 217472 538680 217524
rect 538732 217512 538738 217524
rect 541710 217512 541716 217524
rect 538732 217484 541716 217512
rect 538732 217472 538738 217484
rect 541710 217472 541716 217484
rect 541768 217472 541774 217524
rect 542170 217472 542176 217524
rect 542228 217512 542234 217524
rect 543090 217512 543096 217524
rect 542228 217484 543096 217512
rect 542228 217472 542234 217484
rect 543090 217472 543096 217484
rect 543148 217472 543154 217524
rect 543320 217472 543326 217524
rect 543378 217512 543384 217524
rect 605282 217512 605288 217524
rect 543378 217484 545896 217512
rect 543378 217472 543384 217484
rect 545574 217376 545580 217388
rect 532666 217348 545580 217376
rect 42058 217268 42064 217320
rect 42116 217308 42122 217320
rect 62758 217308 62764 217320
rect 42116 217280 62764 217308
rect 42116 217268 42122 217280
rect 62758 217268 62764 217280
rect 62816 217268 62822 217320
rect 33042 217200 33048 217252
rect 33100 217240 33106 217252
rect 41506 217240 41512 217252
rect 33100 217212 41512 217240
rect 33100 217200 33106 217212
rect 41506 217200 41512 217212
rect 41564 217200 41570 217252
rect 110414 217200 110420 217252
rect 110472 217240 110478 217252
rect 185210 217240 185216 217252
rect 110472 217212 185216 217240
rect 110472 217200 110478 217212
rect 185210 217200 185216 217212
rect 185268 217200 185274 217252
rect 532666 217240 532694 217348
rect 545574 217336 545580 217348
rect 545632 217336 545638 217388
rect 545868 217376 545896 217484
rect 546466 217484 605288 217512
rect 546466 217376 546494 217484
rect 605282 217472 605288 217484
rect 605340 217472 605346 217524
rect 607398 217444 607404 217456
rect 605806 217416 607404 217444
rect 545868 217348 546494 217376
rect 548518 217336 548524 217388
rect 548576 217376 548582 217388
rect 605806 217376 605834 217416
rect 607398 217404 607404 217416
rect 607456 217404 607462 217456
rect 610342 217404 610348 217456
rect 610400 217444 610406 217456
rect 620554 217444 620560 217456
rect 610400 217416 620560 217444
rect 610400 217404 610406 217416
rect 620554 217404 620560 217416
rect 620612 217404 620618 217456
rect 548576 217348 605834 217376
rect 548576 217336 548582 217348
rect 607214 217268 607220 217320
rect 607272 217308 607278 217320
rect 621106 217308 621112 217320
rect 607272 217280 621112 217308
rect 607272 217268 607278 217280
rect 621106 217268 621112 217280
rect 621164 217268 621170 217320
rect 525766 217212 532694 217240
rect 100662 217064 100668 217116
rect 100720 217104 100726 217116
rect 178034 217104 178040 217116
rect 100720 217076 178040 217104
rect 100720 217064 100726 217076
rect 178034 217064 178040 217076
rect 178092 217064 178098 217116
rect 510338 217064 510344 217116
rect 510396 217104 510402 217116
rect 525766 217104 525794 217212
rect 538214 217200 538220 217252
rect 538272 217240 538278 217252
rect 602062 217240 602068 217252
rect 538272 217212 602068 217240
rect 538272 217200 538278 217212
rect 602062 217200 602068 217212
rect 602120 217200 602126 217252
rect 510396 217076 525794 217104
rect 510396 217064 510402 217076
rect 526438 217064 526444 217116
rect 526496 217104 526502 217116
rect 531222 217104 531228 217116
rect 526496 217076 531228 217104
rect 526496 217064 526502 217076
rect 531222 217064 531228 217076
rect 531280 217064 531286 217116
rect 536190 217064 536196 217116
rect 536248 217104 536254 217116
rect 567838 217104 567844 217116
rect 536248 217076 567844 217104
rect 536248 217064 536254 217076
rect 567838 217064 567844 217076
rect 567896 217064 567902 217116
rect 570414 217064 570420 217116
rect 570472 217104 570478 217116
rect 616138 217104 616144 217116
rect 570472 217076 616144 217104
rect 570472 217064 570478 217076
rect 616138 217064 616144 217076
rect 616196 217064 616202 217116
rect 93854 216928 93860 216980
rect 93912 216968 93918 216980
rect 174354 216968 174360 216980
rect 93912 216940 174360 216968
rect 93912 216928 93918 216940
rect 174354 216928 174360 216940
rect 174412 216928 174418 216980
rect 453390 216928 453396 216980
rect 453448 216968 453454 216980
rect 516502 216968 516508 216980
rect 453448 216940 516508 216968
rect 453448 216928 453454 216940
rect 516502 216928 516508 216940
rect 516560 216928 516566 216980
rect 531222 216928 531228 216980
rect 531280 216968 531286 216980
rect 573542 216968 573548 216980
rect 531280 216940 573548 216968
rect 531280 216928 531286 216940
rect 573542 216928 573548 216940
rect 573600 216928 573606 216980
rect 573726 216928 573732 216980
rect 573784 216968 573790 216980
rect 575290 216968 575296 216980
rect 573784 216940 575296 216968
rect 573784 216928 573790 216940
rect 575290 216928 575296 216940
rect 575348 216928 575354 216980
rect 90726 216792 90732 216844
rect 90784 216832 90790 216844
rect 171134 216832 171140 216844
rect 90784 216804 171140 216832
rect 90784 216792 90790 216804
rect 171134 216792 171140 216804
rect 171192 216792 171198 216844
rect 457530 216792 457536 216844
rect 457588 216832 457594 216844
rect 521654 216832 521660 216844
rect 457588 216804 521660 216832
rect 457588 216792 457594 216804
rect 521654 216792 521660 216804
rect 521712 216792 521718 216844
rect 525426 216792 525432 216844
rect 525484 216832 525490 216844
rect 531866 216832 531872 216844
rect 525484 216804 531872 216832
rect 525484 216792 525490 216804
rect 531866 216792 531872 216804
rect 531924 216792 531930 216844
rect 538030 216792 538036 216844
rect 538088 216832 538094 216844
rect 539778 216832 539784 216844
rect 538088 216804 539784 216832
rect 538088 216792 538094 216804
rect 539778 216792 539784 216804
rect 539836 216792 539842 216844
rect 540974 216792 540980 216844
rect 541032 216832 541038 216844
rect 603074 216832 603080 216844
rect 541032 216804 603080 216832
rect 541032 216792 541038 216804
rect 603074 216792 603080 216804
rect 603132 216792 603138 216844
rect 614022 216792 614028 216844
rect 614080 216832 614086 216844
rect 614482 216832 614488 216844
rect 614080 216804 614488 216832
rect 614080 216792 614086 216804
rect 614482 216792 614488 216804
rect 614540 216792 614546 216844
rect 671982 216792 671988 216844
rect 672040 216832 672046 216844
rect 675294 216832 675300 216844
rect 672040 216804 675300 216832
rect 672040 216792 672046 216804
rect 675294 216792 675300 216804
rect 675352 216792 675358 216844
rect 85574 216656 85580 216708
rect 85632 216696 85638 216708
rect 168650 216696 168656 216708
rect 85632 216668 168656 216696
rect 85632 216656 85638 216668
rect 168650 216656 168656 216668
rect 168708 216656 168714 216708
rect 516134 216656 516140 216708
rect 516192 216696 516198 216708
rect 518618 216696 518624 216708
rect 516192 216668 518624 216696
rect 516192 216656 516198 216668
rect 518618 216656 518624 216668
rect 518676 216656 518682 216708
rect 520274 216656 520280 216708
rect 520332 216696 520338 216708
rect 520332 216668 559788 216696
rect 520332 216656 520338 216668
rect 525426 216560 525432 216572
rect 516014 216532 525432 216560
rect 516014 216492 516042 216532
rect 525426 216520 525432 216532
rect 525484 216520 525490 216572
rect 531406 216560 531412 216572
rect 531056 216532 531412 216560
rect 511966 216464 516042 216492
rect 485498 216384 485504 216436
rect 485556 216424 485562 216436
rect 485556 216396 485774 216424
rect 485556 216384 485562 216396
rect 485746 215472 485774 216396
rect 500586 216384 500592 216436
rect 500644 216424 500650 216436
rect 500644 216396 505094 216424
rect 500644 216384 500650 216396
rect 505066 216288 505094 216396
rect 511966 216288 511994 216464
rect 516134 216384 516140 216436
rect 516192 216384 516198 216436
rect 516318 216384 516324 216436
rect 516376 216424 516382 216436
rect 516376 216396 518296 216424
rect 516376 216384 516382 216396
rect 505066 216260 511994 216288
rect 516152 215472 516180 216384
rect 485746 215444 516180 215472
rect 48958 215296 48964 215348
rect 49016 215336 49022 215348
rect 49016 215308 516134 215336
rect 49016 215296 49022 215308
rect 35802 214820 35808 214872
rect 35860 214860 35866 214872
rect 41506 214860 41512 214872
rect 35860 214832 41512 214860
rect 35860 214820 35866 214832
rect 41506 214820 41512 214832
rect 41564 214820 41570 214872
rect 43162 214752 43168 214804
rect 43220 214792 43226 214804
rect 49326 214792 49332 214804
rect 43220 214764 49332 214792
rect 43220 214752 43226 214764
rect 49326 214752 49332 214764
rect 49384 214752 49390 214804
rect 516106 214656 516134 215308
rect 518268 215294 518296 216396
rect 518618 216384 518624 216436
rect 518676 216384 518682 216436
rect 518802 216384 518808 216436
rect 518860 216384 518866 216436
rect 520642 216384 520648 216436
rect 520700 216384 520706 216436
rect 521194 216384 521200 216436
rect 521252 216384 521258 216436
rect 526070 216424 526076 216436
rect 521626 216396 526076 216424
rect 518636 215608 518664 216384
rect 518820 215744 518848 216384
rect 520660 215880 520688 216384
rect 521212 216016 521240 216384
rect 521626 216016 521654 216396
rect 526070 216384 526076 216396
rect 526128 216384 526134 216436
rect 526438 216384 526444 216436
rect 526496 216384 526502 216436
rect 521212 215988 521654 216016
rect 526456 215880 526484 216384
rect 531056 215948 531084 216532
rect 531406 216520 531412 216532
rect 531464 216520 531470 216572
rect 532694 216520 532700 216572
rect 532752 216560 532758 216572
rect 533706 216560 533712 216572
rect 532752 216532 533712 216560
rect 532752 216520 532758 216532
rect 533706 216520 533712 216532
rect 533764 216560 533770 216572
rect 539594 216560 539600 216572
rect 533764 216532 539600 216560
rect 533764 216520 533770 216532
rect 539594 216520 539600 216532
rect 539652 216520 539658 216572
rect 539778 216520 539784 216572
rect 539836 216560 539842 216572
rect 542170 216560 542176 216572
rect 539836 216532 542176 216560
rect 539836 216520 539842 216532
rect 542170 216520 542176 216532
rect 542228 216520 542234 216572
rect 545316 216532 545988 216560
rect 542722 216452 542728 216504
rect 542780 216452 542786 216504
rect 531222 216384 531228 216436
rect 531280 216424 531286 216436
rect 531280 216384 531314 216424
rect 531866 216384 531872 216436
rect 531924 216424 531930 216436
rect 537386 216424 537392 216436
rect 531924 216396 537392 216424
rect 531924 216384 531930 216396
rect 537386 216384 537392 216396
rect 537444 216384 537450 216436
rect 537662 216384 537668 216436
rect 537720 216384 537726 216436
rect 538030 216384 538036 216436
rect 538088 216384 538094 216436
rect 538674 216384 538680 216436
rect 538732 216384 538738 216436
rect 541158 216424 541164 216436
rect 539566 216396 541164 216424
rect 531286 216288 531314 216384
rect 531286 216260 534074 216288
rect 534046 216084 534074 216260
rect 537680 216152 537708 216384
rect 536806 216124 537708 216152
rect 536806 216084 536834 216124
rect 534046 216056 536834 216084
rect 531056 215920 534074 215948
rect 520660 215852 526484 215880
rect 534046 215880 534074 215920
rect 538048 215880 538076 216384
rect 534046 215852 538076 215880
rect 538692 215744 538720 216384
rect 518820 215716 538720 215744
rect 518636 215580 524414 215608
rect 524386 215540 524414 215580
rect 524386 215512 525794 215540
rect 525766 215472 525794 215512
rect 535426 215512 538214 215540
rect 525766 215444 527174 215472
rect 527146 215404 527174 215444
rect 527146 215376 532694 215404
rect 532666 215336 532694 215376
rect 535426 215336 535454 215512
rect 532666 215308 535454 215336
rect 538186 215336 538214 215512
rect 539566 215336 539594 216396
rect 541158 216384 541164 216396
rect 541216 216384 541222 216436
rect 541986 216384 541992 216436
rect 542044 216384 542050 216436
rect 542004 215540 542032 216384
rect 538186 215308 539594 215336
rect 539704 215512 542032 215540
rect 518176 215266 518296 215294
rect 518176 215200 518204 215266
rect 539704 215200 539732 215512
rect 518176 215172 527174 215200
rect 527146 214928 527174 215172
rect 535426 215172 539732 215200
rect 535426 214928 535454 215172
rect 527146 214900 535454 214928
rect 516106 214628 539594 214656
rect 539566 214520 539594 214628
rect 542740 214520 542768 216452
rect 542998 216384 543004 216436
rect 543056 216384 543062 216436
rect 543458 216384 543464 216436
rect 543516 216384 543522 216436
rect 543642 216384 543648 216436
rect 543700 216384 543706 216436
rect 545114 216384 545120 216436
rect 545172 216384 545178 216436
rect 543016 214588 543044 216384
rect 543476 215948 543504 216384
rect 543660 216084 543688 216384
rect 545132 216084 545160 216384
rect 545316 216152 545344 216532
rect 545482 216384 545488 216436
rect 545540 216384 545546 216436
rect 545666 216384 545672 216436
rect 545724 216424 545730 216436
rect 545724 216396 545896 216424
rect 545724 216384 545730 216396
rect 545500 216288 545528 216384
rect 545500 216260 545804 216288
rect 543660 216056 545160 216084
rect 545224 216124 545344 216152
rect 543476 215920 543734 215948
rect 543706 215880 543734 215920
rect 545224 215880 545252 216124
rect 543706 215852 545252 215880
rect 545776 215812 545804 216260
rect 545868 216084 545896 216396
rect 545960 216288 545988 216532
rect 547966 216520 547972 216572
rect 548024 216560 548030 216572
rect 548024 216532 553808 216560
rect 548024 216520 548030 216532
rect 546770 216384 546776 216436
rect 546828 216424 546834 216436
rect 546828 216396 552014 216424
rect 546828 216384 546834 216396
rect 551986 216356 552014 216396
rect 552658 216384 552664 216436
rect 552716 216424 552722 216436
rect 552716 216396 553256 216424
rect 552716 216384 552722 216396
rect 551986 216328 552244 216356
rect 552216 216288 552244 216328
rect 545960 216260 549576 216288
rect 552216 216260 552888 216288
rect 545868 216056 548472 216084
rect 545776 215784 545896 215812
rect 545868 215472 545896 215784
rect 545868 215444 548288 215472
rect 548260 214996 548288 215444
rect 548444 215404 548472 216056
rect 549548 215676 549576 216260
rect 552860 215880 552888 216260
rect 553228 216016 553256 216396
rect 553780 216288 553808 216532
rect 553946 216384 553952 216436
rect 554004 216424 554010 216436
rect 559760 216424 559788 216668
rect 566182 216656 566188 216708
rect 566240 216696 566246 216708
rect 618346 216696 618352 216708
rect 566240 216668 618352 216696
rect 566240 216656 566246 216668
rect 618346 216656 618352 216668
rect 618404 216656 618410 216708
rect 670418 216656 670424 216708
rect 670476 216696 670482 216708
rect 675478 216696 675484 216708
rect 670476 216668 675484 216696
rect 670476 216656 670482 216668
rect 675478 216656 675484 216668
rect 675536 216656 675542 216708
rect 562502 216520 562508 216572
rect 562560 216560 562566 216572
rect 562560 216532 576854 216560
rect 562560 216520 562566 216532
rect 576826 216492 576854 216532
rect 600774 216492 600780 216504
rect 576826 216464 600780 216492
rect 600774 216452 600780 216464
rect 600832 216452 600838 216504
rect 600958 216452 600964 216504
rect 601016 216492 601022 216504
rect 606754 216492 606760 216504
rect 601016 216464 606760 216492
rect 601016 216452 601022 216464
rect 606754 216452 606760 216464
rect 606812 216452 606818 216504
rect 566182 216424 566188 216436
rect 554004 216396 558914 216424
rect 559760 216396 566188 216424
rect 554004 216384 554010 216396
rect 558886 216356 558914 216396
rect 566182 216384 566188 216396
rect 566240 216384 566246 216436
rect 567838 216384 567844 216436
rect 567896 216424 567902 216436
rect 573726 216424 573732 216436
rect 567896 216396 573732 216424
rect 567896 216384 567902 216396
rect 573726 216384 573732 216396
rect 573784 216384 573790 216436
rect 558886 216328 559604 216356
rect 559576 216288 559604 216328
rect 574002 216316 574008 216368
rect 574060 216356 574066 216368
rect 627178 216356 627184 216368
rect 574060 216328 627184 216356
rect 574060 216316 574066 216328
rect 627178 216316 627184 216328
rect 627236 216316 627242 216368
rect 553780 216260 554774 216288
rect 559576 216260 559696 216288
rect 554746 216152 554774 216260
rect 559668 216220 559696 216260
rect 600958 216220 600964 216232
rect 559668 216192 600964 216220
rect 600958 216180 600964 216192
rect 601016 216180 601022 216232
rect 616690 216220 616696 216232
rect 601160 216192 616696 216220
rect 554746 216124 558914 216152
rect 558886 216084 558914 216124
rect 576578 216084 576584 216096
rect 558886 216056 576584 216084
rect 576578 216044 576584 216056
rect 576636 216044 576642 216096
rect 576762 216044 576768 216096
rect 576820 216084 576826 216096
rect 576820 216044 576854 216084
rect 600774 216044 600780 216096
rect 600832 216084 600838 216096
rect 601160 216084 601188 216192
rect 616690 216180 616696 216192
rect 616748 216180 616754 216232
rect 600832 216056 601188 216084
rect 600832 216044 600838 216056
rect 602890 216044 602896 216096
rect 602948 216084 602954 216096
rect 626074 216084 626080 216096
rect 602948 216056 626080 216084
rect 602948 216044 602954 216056
rect 626074 216044 626080 216056
rect 626132 216044 626138 216096
rect 576826 216016 576854 216044
rect 553228 215988 554774 216016
rect 576826 215988 600636 216016
rect 554746 215948 554774 215988
rect 600608 215948 600636 215988
rect 601234 215948 601240 215960
rect 554746 215920 558914 215948
rect 558886 215880 558914 215920
rect 560266 215920 575474 215948
rect 600608 215920 601240 215948
rect 560266 215880 560294 215920
rect 552860 215852 553394 215880
rect 558886 215852 560294 215880
rect 575446 215880 575474 215920
rect 601234 215908 601240 215920
rect 601292 215908 601298 215960
rect 601510 215908 601516 215960
rect 601568 215948 601574 215960
rect 623774 215948 623780 215960
rect 601568 215920 623780 215948
rect 601568 215908 601574 215920
rect 623774 215908 623780 215920
rect 623832 215908 623838 215960
rect 599578 215880 599584 215892
rect 575446 215852 599584 215880
rect 553366 215812 553394 215852
rect 599578 215840 599584 215852
rect 599636 215840 599642 215892
rect 553366 215784 555740 215812
rect 555712 215744 555740 215784
rect 563026 215784 569954 215812
rect 555712 215716 561674 215744
rect 549548 215648 553394 215676
rect 553366 215608 553394 215648
rect 553366 215580 554774 215608
rect 554746 215540 554774 215580
rect 556126 215580 560294 215608
rect 556126 215540 556154 215580
rect 554746 215512 556154 215540
rect 560266 215404 560294 215580
rect 561646 215540 561674 215716
rect 563026 215540 563054 215784
rect 561646 215512 563054 215540
rect 569926 215472 569954 215784
rect 576808 215704 576814 215756
rect 576866 215744 576872 215756
rect 596266 215744 596272 215756
rect 576866 215716 596272 215744
rect 576866 215704 576872 215716
rect 596266 215704 596272 215716
rect 596324 215704 596330 215756
rect 596450 215704 596456 215756
rect 596508 215744 596514 215756
rect 600682 215744 600688 215756
rect 596508 215716 600688 215744
rect 596508 215704 596514 215716
rect 600682 215704 600688 215716
rect 600740 215704 600746 215756
rect 573910 215568 573916 215620
rect 573968 215608 573974 215620
rect 573968 215580 596312 215608
rect 573968 215568 573974 215580
rect 586468 215472 586474 215484
rect 564406 215444 568574 215472
rect 569926 215444 586474 215472
rect 564406 215404 564434 215444
rect 548444 215376 549208 215404
rect 560266 215376 564434 215404
rect 549180 215200 549208 215376
rect 568546 215268 568574 215444
rect 586468 215432 586474 215444
rect 586526 215432 586532 215484
rect 586698 215432 586704 215484
rect 586756 215472 586762 215484
rect 595990 215472 595996 215484
rect 586756 215444 595996 215472
rect 586756 215432 586762 215444
rect 595990 215432 595996 215444
rect 596048 215432 596054 215484
rect 596284 215472 596312 215580
rect 596634 215568 596640 215620
rect 596692 215608 596698 215620
rect 614114 215608 614120 215620
rect 596692 215580 614120 215608
rect 596692 215568 596698 215580
rect 614114 215568 614120 215580
rect 614172 215568 614178 215620
rect 600314 215472 600320 215484
rect 596284 215444 600320 215472
rect 600314 215432 600320 215444
rect 600372 215432 600378 215484
rect 600498 215432 600504 215484
rect 600556 215472 600562 215484
rect 603994 215472 604000 215484
rect 600556 215444 604000 215472
rect 600556 215432 600562 215444
rect 603994 215432 604000 215444
rect 604052 215432 604058 215484
rect 673914 215432 673920 215484
rect 673972 215472 673978 215484
rect 675478 215472 675484 215484
rect 673972 215444 675484 215472
rect 673972 215432 673978 215444
rect 675478 215432 675484 215444
rect 675536 215432 675542 215484
rect 573726 215296 573732 215348
rect 573784 215336 573790 215348
rect 576578 215336 576584 215348
rect 573784 215308 576584 215336
rect 573784 215296 573790 215308
rect 576578 215296 576584 215308
rect 576636 215296 576642 215348
rect 664162 215336 664168 215348
rect 579586 215308 664168 215336
rect 568546 215240 569954 215268
rect 549180 215172 554774 215200
rect 554746 215132 554774 215172
rect 556126 215172 557534 215200
rect 556126 215132 556154 215172
rect 554746 215104 556154 215132
rect 557506 215132 557534 215172
rect 569926 215132 569954 215240
rect 579586 215200 579614 215308
rect 664162 215296 664168 215308
rect 664220 215296 664226 215348
rect 675294 215336 675300 215348
rect 673748 215308 675300 215336
rect 673748 215212 673776 215308
rect 675294 215296 675300 215308
rect 675352 215296 675358 215348
rect 571306 215172 574094 215200
rect 571306 215132 571334 215172
rect 557506 215104 560294 215132
rect 560266 215064 560294 215104
rect 561646 215104 564434 215132
rect 569926 215104 571334 215132
rect 574066 215132 574094 215172
rect 575446 215172 579614 215200
rect 575446 215132 575474 215172
rect 673730 215160 673736 215212
rect 673788 215160 673794 215212
rect 574066 215104 575474 215132
rect 561646 215064 561674 215104
rect 560266 215036 561674 215064
rect 564406 215064 564434 215104
rect 581638 215092 581644 215144
rect 581696 215132 581702 215144
rect 616874 215132 616880 215144
rect 581696 215104 616880 215132
rect 581696 215092 581702 215104
rect 616874 215092 616880 215104
rect 616932 215092 616938 215144
rect 564406 215036 568574 215064
rect 568546 214996 568574 215036
rect 576026 214996 576032 215008
rect 548260 214968 556154 214996
rect 568546 214968 569954 214996
rect 556126 214928 556154 214968
rect 569926 214928 569954 214968
rect 571306 214968 574094 214996
rect 571306 214928 571334 214968
rect 556126 214900 560294 214928
rect 560266 214860 560294 214900
rect 561646 214900 563054 214928
rect 561646 214860 561674 214900
rect 560266 214832 561674 214860
rect 563026 214860 563054 214900
rect 564406 214900 565032 214928
rect 569926 214900 571334 214928
rect 564406 214860 564434 214900
rect 563026 214832 564434 214860
rect 565004 214792 565032 214900
rect 574066 214860 574094 214968
rect 575446 214968 576032 214996
rect 575446 214860 575474 214968
rect 576026 214956 576032 214968
rect 576084 214956 576090 215008
rect 581454 214956 581460 215008
rect 581512 214996 581518 215008
rect 618898 214996 618904 215008
rect 581512 214968 618904 214996
rect 581512 214956 581518 214968
rect 618898 214956 618904 214968
rect 618956 214956 618962 215008
rect 574066 214832 575474 214860
rect 575658 214820 575664 214872
rect 575716 214860 575722 214872
rect 620002 214860 620008 214872
rect 575716 214832 620008 214860
rect 575716 214820 575722 214832
rect 620002 214820 620008 214832
rect 620060 214820 620066 214872
rect 565004 214764 565814 214792
rect 565786 214724 565814 214764
rect 573910 214724 573916 214736
rect 565786 214696 573916 214724
rect 573910 214684 573916 214696
rect 573968 214684 573974 214736
rect 574738 214684 574744 214736
rect 574796 214684 574802 214736
rect 574922 214684 574928 214736
rect 574980 214724 574986 214736
rect 581454 214724 581460 214736
rect 574980 214696 581460 214724
rect 574980 214684 574986 214696
rect 581454 214684 581460 214696
rect 581512 214684 581518 214736
rect 619634 214724 619640 214736
rect 581656 214696 619640 214724
rect 573726 214588 573732 214600
rect 543016 214560 550634 214588
rect 539566 214492 542768 214520
rect 550606 214520 550634 214560
rect 560266 214560 573732 214588
rect 560266 214520 560294 214560
rect 573726 214548 573732 214560
rect 573784 214548 573790 214600
rect 574756 214588 574784 214684
rect 574664 214560 574784 214588
rect 550606 214492 560294 214520
rect 574664 214452 574692 214560
rect 575842 214548 575848 214600
rect 575900 214588 575906 214600
rect 581656 214588 581684 214696
rect 619634 214684 619640 214696
rect 619692 214684 619698 214736
rect 622394 214588 622400 214600
rect 575900 214560 581684 214588
rect 586486 214560 622400 214588
rect 575900 214548 575906 214560
rect 574830 214452 574836 214464
rect 574664 214424 574836 214452
rect 574830 214412 574836 214424
rect 574888 214412 574894 214464
rect 575290 214412 575296 214464
rect 575348 214452 575354 214464
rect 586486 214452 586514 214560
rect 622394 214548 622400 214560
rect 622452 214548 622458 214600
rect 655514 214548 655520 214600
rect 655572 214588 655578 214600
rect 656434 214588 656440 214600
rect 655572 214560 656440 214588
rect 655572 214548 655578 214560
rect 656434 214548 656440 214560
rect 656492 214548 656498 214600
rect 659654 214548 659660 214600
rect 659712 214588 659718 214600
rect 660298 214588 660304 214600
rect 659712 214560 660304 214588
rect 659712 214548 659718 214560
rect 660298 214548 660304 214560
rect 660356 214548 660362 214600
rect 661310 214548 661316 214600
rect 661368 214588 661374 214600
rect 661954 214588 661960 214600
rect 661368 214560 661960 214588
rect 661368 214548 661374 214560
rect 661954 214548 661960 214560
rect 662012 214548 662018 214600
rect 575348 214424 586514 214452
rect 575348 214412 575354 214424
rect 608778 214412 608784 214464
rect 608836 214452 608842 214464
rect 609514 214452 609520 214464
rect 608836 214424 609520 214452
rect 608836 214412 608842 214424
rect 609514 214412 609520 214424
rect 609572 214412 609578 214464
rect 575106 214276 575112 214328
rect 575164 214316 575170 214328
rect 581638 214316 581644 214328
rect 575164 214288 581644 214316
rect 575164 214276 575170 214288
rect 581638 214276 581644 214288
rect 581696 214276 581702 214328
rect 35802 214072 35808 214124
rect 35860 214112 35866 214124
rect 39942 214112 39948 214124
rect 35860 214084 39948 214112
rect 35860 214072 35866 214084
rect 39942 214072 39948 214084
rect 40000 214072 40006 214124
rect 673086 214072 673092 214124
rect 673144 214112 673150 214124
rect 675478 214112 675484 214124
rect 673144 214084 675484 214112
rect 673144 214072 673150 214084
rect 675478 214072 675484 214084
rect 675536 214072 675542 214124
rect 580350 213868 580356 213920
rect 580408 213908 580414 213920
rect 595714 213908 595720 213920
rect 580408 213880 595720 213908
rect 580408 213868 580414 213880
rect 595714 213868 595720 213880
rect 595772 213868 595778 213920
rect 596358 213908 596364 213920
rect 596146 213880 596364 213908
rect 574646 213732 574652 213784
rect 574704 213772 574710 213784
rect 595162 213772 595168 213784
rect 574704 213744 595168 213772
rect 574704 213732 574710 213744
rect 595162 213732 595168 213744
rect 595220 213732 595226 213784
rect 595346 213732 595352 213784
rect 595404 213772 595410 213784
rect 596146 213772 596174 213880
rect 596358 213868 596364 213880
rect 596416 213868 596422 213920
rect 603074 213868 603080 213920
rect 603132 213908 603138 213920
rect 605926 213908 605932 213920
rect 603132 213880 605932 213908
rect 603132 213868 603138 213880
rect 605926 213868 605932 213880
rect 605984 213868 605990 213920
rect 609238 213868 609244 213920
rect 609296 213908 609302 213920
rect 610618 213908 610624 213920
rect 609296 213880 610624 213908
rect 609296 213868 609302 213880
rect 610618 213868 610624 213880
rect 610676 213868 610682 213920
rect 624142 213868 624148 213920
rect 624200 213908 624206 213920
rect 625246 213908 625252 213920
rect 624200 213880 625252 213908
rect 624200 213868 624206 213880
rect 625246 213868 625252 213880
rect 625304 213868 625310 213920
rect 628558 213868 628564 213920
rect 628616 213908 628622 213920
rect 633802 213908 633808 213920
rect 628616 213880 633808 213908
rect 628616 213868 628622 213880
rect 633802 213868 633808 213880
rect 633860 213868 633866 213920
rect 639966 213868 639972 213920
rect 640024 213908 640030 213920
rect 651374 213908 651380 213920
rect 640024 213880 651380 213908
rect 640024 213868 640030 213880
rect 651374 213868 651380 213880
rect 651432 213868 651438 213920
rect 595404 213744 596174 213772
rect 595404 213732 595410 213744
rect 602062 213732 602068 213784
rect 602120 213772 602126 213784
rect 605098 213772 605104 213784
rect 602120 213744 605104 213772
rect 602120 213732 602126 213744
rect 605098 213732 605104 213744
rect 605156 213732 605162 213784
rect 605282 213732 605288 213784
rect 605340 213772 605346 213784
rect 606202 213772 606208 213784
rect 605340 213744 606208 213772
rect 605340 213732 605346 213744
rect 606202 213732 606208 213744
rect 606260 213732 606266 213784
rect 638862 213732 638868 213784
rect 638920 213772 638926 213784
rect 649994 213772 650000 213784
rect 638920 213744 650000 213772
rect 638920 213732 638926 213744
rect 649994 213732 650000 213744
rect 650052 213732 650058 213784
rect 671798 213664 671804 213716
rect 671856 213704 671862 213716
rect 675478 213704 675484 213716
rect 671856 213676 675484 213704
rect 671856 213664 671862 213676
rect 675478 213664 675484 213676
rect 675536 213664 675542 213716
rect 574462 213596 574468 213648
rect 574520 213636 574526 213648
rect 603626 213636 603632 213648
rect 574520 213608 603632 213636
rect 574520 213596 574526 213608
rect 603626 213596 603632 213608
rect 603684 213596 603690 213648
rect 638310 213596 638316 213648
rect 638368 213636 638374 213648
rect 651742 213636 651748 213648
rect 638368 213608 651748 213636
rect 638368 213596 638374 213608
rect 651742 213596 651748 213608
rect 651800 213596 651806 213648
rect 574094 213460 574100 213512
rect 574152 213500 574158 213512
rect 604546 213500 604552 213512
rect 574152 213472 604552 213500
rect 574152 213460 574158 213472
rect 604546 213460 604552 213472
rect 604604 213460 604610 213512
rect 636654 213460 636660 213512
rect 636712 213500 636718 213512
rect 650178 213500 650184 213512
rect 636712 213472 650184 213500
rect 636712 213460 636718 213472
rect 650178 213460 650184 213472
rect 650236 213460 650242 213512
rect 575474 213324 575480 213376
rect 575532 213364 575538 213376
rect 629386 213364 629392 213376
rect 575532 213336 629392 213364
rect 575532 213324 575538 213336
rect 629386 213324 629392 213336
rect 629444 213324 629450 213376
rect 635550 213324 635556 213376
rect 635608 213364 635614 213376
rect 649074 213364 649080 213376
rect 635608 213336 649080 213364
rect 635608 213324 635614 213336
rect 649074 213324 649080 213336
rect 649132 213324 649138 213376
rect 672258 213256 672264 213308
rect 672316 213296 672322 213308
rect 675478 213296 675484 213308
rect 672316 213268 675484 213296
rect 672316 213256 672322 213268
rect 675478 213256 675484 213268
rect 675536 213256 675542 213308
rect 574830 213188 574836 213240
rect 574888 213228 574894 213240
rect 630674 213228 630680 213240
rect 574888 213200 630680 213228
rect 574888 213188 574894 213200
rect 630674 213188 630680 213200
rect 630732 213188 630738 213240
rect 637206 213188 637212 213240
rect 637264 213228 637270 213240
rect 650730 213228 650736 213240
rect 637264 213200 650736 213228
rect 637264 213188 637270 213200
rect 650730 213188 650736 213200
rect 650788 213188 650794 213240
rect 640242 213052 640248 213104
rect 640300 213092 640306 213104
rect 650914 213092 650920 213104
rect 640300 213064 650920 213092
rect 640300 213052 640306 213064
rect 650914 213052 650920 213064
rect 650972 213052 650978 213104
rect 616690 212984 616696 213036
rect 616748 213024 616754 213036
rect 623314 213024 623320 213036
rect 616748 212996 623320 213024
rect 616748 212984 616754 212996
rect 623314 212984 623320 212996
rect 623372 212984 623378 213036
rect 35802 212916 35808 212968
rect 35860 212956 35866 212968
rect 40310 212956 40316 212968
rect 35860 212928 40316 212956
rect 35860 212916 35866 212928
rect 40310 212916 40316 212928
rect 40368 212916 40374 212968
rect 641622 212916 641628 212968
rect 641680 212956 641686 212968
rect 650362 212956 650368 212968
rect 641680 212928 650368 212956
rect 641680 212916 641686 212928
rect 650362 212916 650368 212928
rect 650420 212916 650426 212968
rect 632698 212780 632704 212832
rect 632756 212820 632762 212832
rect 634354 212820 634360 212832
rect 632756 212792 634360 212820
rect 632756 212780 632762 212792
rect 634354 212780 634360 212792
rect 634412 212780 634418 212832
rect 35618 212644 35624 212696
rect 35676 212684 35682 212696
rect 40678 212684 40684 212696
rect 35676 212656 40684 212684
rect 35676 212644 35682 212656
rect 40678 212644 40684 212656
rect 40736 212644 40742 212696
rect 630030 212644 630036 212696
rect 630088 212684 630094 212696
rect 632698 212684 632704 212696
rect 630088 212656 632704 212684
rect 630088 212644 630094 212656
rect 632698 212644 632704 212656
rect 632756 212644 632762 212696
rect 35434 212508 35440 212560
rect 35492 212548 35498 212560
rect 39942 212548 39948 212560
rect 35492 212520 39948 212548
rect 35492 212508 35498 212520
rect 39942 212508 39948 212520
rect 40000 212508 40006 212560
rect 579246 211964 579252 212016
rect 579304 212004 579310 212016
rect 581914 212004 581920 212016
rect 579304 211976 581920 212004
rect 579304 211964 579310 211976
rect 581914 211964 581920 211976
rect 581972 211964 581978 212016
rect 675846 211760 675852 211812
rect 675904 211800 675910 211812
rect 683114 211800 683120 211812
rect 675904 211772 683120 211800
rect 675904 211760 675910 211772
rect 683114 211760 683120 211772
rect 683172 211760 683178 211812
rect 35802 211556 35808 211608
rect 35860 211596 35866 211608
rect 40954 211596 40960 211608
rect 35860 211568 40960 211596
rect 35860 211556 35866 211568
rect 40954 211556 40960 211568
rect 41012 211556 41018 211608
rect 39666 211392 39672 211404
rect 36004 211364 39672 211392
rect 35802 211284 35808 211336
rect 35860 211324 35866 211336
rect 36004 211324 36032 211364
rect 39666 211352 39672 211364
rect 39724 211352 39730 211404
rect 35860 211296 36032 211324
rect 35860 211284 35866 211296
rect 578510 211284 578516 211336
rect 578568 211324 578574 211336
rect 583294 211324 583300 211336
rect 578568 211296 583300 211324
rect 578568 211284 578574 211296
rect 583294 211284 583300 211296
rect 583352 211284 583358 211336
rect 35618 211148 35624 211200
rect 35676 211188 35682 211200
rect 41506 211188 41512 211200
rect 35676 211160 41512 211188
rect 35676 211148 35682 211160
rect 41506 211148 41512 211160
rect 41564 211148 41570 211200
rect 42334 211148 42340 211200
rect 42392 211188 42398 211200
rect 51718 211188 51724 211200
rect 42392 211160 51724 211188
rect 42392 211148 42398 211160
rect 51718 211148 51724 211160
rect 51776 211148 51782 211200
rect 578878 211148 578884 211200
rect 578936 211188 578942 211200
rect 580902 211188 580908 211200
rect 578936 211160 580908 211188
rect 578936 211148 578942 211160
rect 580902 211148 580908 211160
rect 580960 211148 580966 211200
rect 664806 211080 664812 211132
rect 664864 211120 664870 211132
rect 667566 211120 667572 211132
rect 664864 211092 667572 211120
rect 664864 211080 664870 211092
rect 667566 211080 667572 211092
rect 667624 211080 667630 211132
rect 644474 211012 644480 211064
rect 644532 211052 644538 211064
rect 644842 211052 644848 211064
rect 644532 211024 644848 211052
rect 644532 211012 644538 211024
rect 644842 211012 644848 211024
rect 644900 211012 644906 211064
rect 652018 210400 652024 210452
rect 652076 210440 652082 210452
rect 652076 210412 669314 210440
rect 652076 210400 652082 210412
rect 669286 210304 669314 210412
rect 670970 210304 670976 210316
rect 669286 210276 670976 210304
rect 670970 210264 670976 210276
rect 671028 210264 671034 210316
rect 608594 210060 608600 210112
rect 608652 210100 608658 210112
rect 608962 210100 608968 210112
rect 608652 210072 608968 210100
rect 608652 210060 608658 210072
rect 608962 210060 608968 210072
rect 609020 210060 609026 210112
rect 35802 209924 35808 209976
rect 35860 209964 35866 209976
rect 40034 209964 40040 209976
rect 35860 209936 40040 209964
rect 35860 209924 35866 209936
rect 40034 209924 40040 209936
rect 40092 209924 40098 209976
rect 35618 209788 35624 209840
rect 35676 209828 35682 209840
rect 41690 209828 41696 209840
rect 35676 209800 41696 209828
rect 35676 209788 35682 209800
rect 41690 209788 41696 209800
rect 41748 209788 41754 209840
rect 579246 209788 579252 209840
rect 579304 209828 579310 209840
rect 581638 209828 581644 209840
rect 579304 209800 581644 209828
rect 579304 209788 579310 209800
rect 581638 209788 581644 209800
rect 581696 209788 581702 209840
rect 591298 209788 591304 209840
rect 591356 209828 591362 209840
rect 632146 209828 632152 209840
rect 591356 209800 632152 209828
rect 591356 209788 591362 209800
rect 632146 209788 632152 209800
rect 632204 209788 632210 209840
rect 652202 209516 652208 209568
rect 652260 209556 652266 209568
rect 652260 209528 654134 209556
rect 652260 209516 652266 209528
rect 654106 209080 654134 209528
rect 669406 209080 669412 209092
rect 654106 209052 669412 209080
rect 669406 209040 669412 209052
rect 669464 209040 669470 209092
rect 35802 208700 35808 208752
rect 35860 208740 35866 208752
rect 35860 208700 35894 208740
rect 35866 208672 35894 208700
rect 39942 208672 39948 208684
rect 35866 208644 39948 208672
rect 39942 208632 39948 208644
rect 40000 208632 40006 208684
rect 35802 208360 35808 208412
rect 35860 208400 35866 208412
rect 41690 208400 41696 208412
rect 35860 208372 41696 208400
rect 35860 208360 35866 208372
rect 41690 208360 41696 208372
rect 41748 208360 41754 208412
rect 42058 208360 42064 208412
rect 42116 208400 42122 208412
rect 43070 208400 43076 208412
rect 42116 208372 43076 208400
rect 42116 208360 42122 208372
rect 43070 208360 43076 208372
rect 43128 208360 43134 208412
rect 578694 208292 578700 208344
rect 578752 208332 578758 208344
rect 589458 208332 589464 208344
rect 578752 208304 589464 208332
rect 578752 208292 578758 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 669590 208088 669596 208140
rect 669648 208128 669654 208140
rect 675478 208128 675484 208140
rect 669648 208100 675484 208128
rect 669648 208088 669654 208100
rect 675478 208088 675484 208100
rect 675536 208088 675542 208140
rect 578418 208020 578424 208072
rect 578476 208060 578482 208072
rect 580626 208060 580632 208072
rect 578476 208032 580632 208060
rect 578476 208020 578482 208032
rect 580626 208020 580632 208032
rect 580684 208020 580690 208072
rect 35802 207272 35808 207324
rect 35860 207312 35866 207324
rect 40126 207312 40132 207324
rect 35860 207284 40132 207312
rect 35860 207272 35866 207284
rect 40126 207272 40132 207284
rect 40184 207272 40190 207324
rect 35526 207000 35532 207052
rect 35584 207040 35590 207052
rect 40954 207040 40960 207052
rect 35584 207012 40960 207040
rect 35584 207000 35590 207012
rect 40954 207000 40960 207012
rect 41012 207000 41018 207052
rect 581914 206932 581920 206984
rect 581972 206972 581978 206984
rect 589458 206972 589464 206984
rect 581972 206944 589464 206972
rect 581972 206932 581978 206944
rect 589458 206932 589464 206944
rect 589516 206932 589522 206984
rect 35802 205912 35808 205964
rect 35860 205952 35866 205964
rect 39758 205952 39764 205964
rect 35860 205924 39764 205952
rect 35860 205912 35866 205924
rect 39758 205912 39764 205924
rect 39816 205912 39822 205964
rect 674834 205708 674840 205760
rect 674892 205748 674898 205760
rect 675386 205748 675392 205760
rect 674892 205720 675392 205748
rect 674892 205708 674898 205720
rect 675386 205708 675392 205720
rect 675444 205708 675450 205760
rect 35802 205640 35808 205692
rect 35860 205680 35866 205692
rect 41690 205680 41696 205692
rect 35860 205652 41696 205680
rect 35860 205640 35866 205652
rect 41690 205640 41696 205652
rect 41748 205640 41754 205692
rect 42058 205640 42064 205692
rect 42116 205680 42122 205692
rect 43438 205680 43444 205692
rect 42116 205652 43444 205680
rect 42116 205640 42122 205652
rect 43438 205640 43444 205652
rect 43496 205640 43502 205692
rect 578694 205640 578700 205692
rect 578752 205680 578758 205692
rect 581822 205680 581828 205692
rect 578752 205652 581828 205680
rect 578752 205640 578758 205652
rect 581822 205640 581828 205652
rect 581880 205640 581886 205692
rect 583294 205572 583300 205624
rect 583352 205612 583358 205624
rect 589458 205612 589464 205624
rect 583352 205584 589464 205612
rect 583352 205572 583358 205584
rect 589458 205572 589464 205584
rect 589516 205572 589522 205624
rect 579062 205232 579068 205284
rect 579120 205272 579126 205284
rect 584398 205272 584404 205284
rect 579120 205244 584404 205272
rect 579120 205232 579126 205244
rect 584398 205232 584404 205244
rect 584456 205232 584462 205284
rect 35802 204892 35808 204944
rect 35860 204932 35866 204944
rect 40770 204932 40776 204944
rect 35860 204904 40776 204932
rect 35860 204892 35866 204904
rect 40770 204892 40776 204904
rect 40828 204892 40834 204944
rect 41690 204728 41696 204740
rect 41386 204700 41696 204728
rect 35618 204620 35624 204672
rect 35676 204660 35682 204672
rect 41386 204660 41414 204700
rect 41690 204688 41696 204700
rect 41748 204688 41754 204740
rect 42058 204688 42064 204740
rect 42116 204728 42122 204740
rect 44358 204728 44364 204740
rect 42116 204700 44364 204728
rect 42116 204688 42122 204700
rect 44358 204688 44364 204700
rect 44416 204688 44422 204740
rect 35676 204632 41414 204660
rect 35676 204620 35682 204632
rect 42058 204552 42064 204604
rect 42116 204592 42122 204604
rect 50338 204592 50344 204604
rect 42116 204564 50344 204592
rect 42116 204552 42122 204564
rect 50338 204552 50344 204564
rect 50396 204552 50402 204604
rect 35802 204484 35808 204536
rect 35860 204524 35866 204536
rect 41690 204524 41696 204536
rect 35860 204496 41696 204524
rect 35860 204484 35866 204496
rect 41690 204484 41696 204496
rect 41748 204484 41754 204536
rect 35526 204280 35532 204332
rect 35584 204320 35590 204332
rect 41690 204320 41696 204332
rect 35584 204292 41696 204320
rect 35584 204280 35590 204292
rect 41690 204280 41696 204292
rect 41748 204280 41754 204332
rect 42058 204280 42064 204332
rect 42116 204320 42122 204332
rect 48958 204320 48964 204332
rect 42116 204292 48964 204320
rect 42116 204280 42122 204292
rect 48958 204280 48964 204292
rect 49016 204280 49022 204332
rect 580902 204144 580908 204196
rect 580960 204184 580966 204196
rect 589458 204184 589464 204196
rect 580960 204156 589464 204184
rect 580960 204144 580966 204156
rect 589458 204144 589464 204156
rect 589516 204144 589522 204196
rect 35618 203124 35624 203176
rect 35676 203164 35682 203176
rect 41598 203164 41604 203176
rect 35676 203136 41604 203164
rect 35676 203124 35682 203136
rect 41598 203124 41604 203136
rect 41656 203124 41662 203176
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 40034 202892 40040 202904
rect 35860 202864 40040 202892
rect 35860 202852 35866 202864
rect 40034 202852 40040 202864
rect 40092 202852 40098 202904
rect 578694 202852 578700 202904
rect 578752 202892 578758 202904
rect 583202 202892 583208 202904
rect 578752 202864 583208 202892
rect 578752 202852 578758 202864
rect 583202 202852 583208 202864
rect 583260 202852 583266 202904
rect 581638 202716 581644 202768
rect 581696 202756 581702 202768
rect 589366 202756 589372 202768
rect 581696 202728 589372 202756
rect 581696 202716 581702 202728
rect 589366 202716 589372 202728
rect 589424 202716 589430 202768
rect 578234 201628 578240 201680
rect 578292 201668 578298 201680
rect 580902 201668 580908 201680
rect 578292 201640 580908 201668
rect 578292 201628 578298 201640
rect 580902 201628 580908 201640
rect 580960 201628 580966 201680
rect 673914 201424 673920 201476
rect 673972 201464 673978 201476
rect 675386 201464 675392 201476
rect 673972 201436 675392 201464
rect 673972 201424 673978 201436
rect 675386 201424 675392 201436
rect 675444 201424 675450 201476
rect 671798 201220 671804 201272
rect 671856 201260 671862 201272
rect 675110 201260 675116 201272
rect 671856 201232 675116 201260
rect 671856 201220 671862 201232
rect 675110 201220 675116 201232
rect 675168 201220 675174 201272
rect 581822 200744 581828 200796
rect 581880 200784 581886 200796
rect 590378 200784 590384 200796
rect 581880 200756 590384 200784
rect 581880 200744 581886 200756
rect 590378 200744 590384 200756
rect 590436 200744 590442 200796
rect 673730 200744 673736 200796
rect 673788 200784 673794 200796
rect 674926 200784 674932 200796
rect 673788 200756 674932 200784
rect 673788 200744 673794 200756
rect 674926 200744 674932 200756
rect 674984 200744 674990 200796
rect 578510 200404 578516 200456
rect 578568 200444 578574 200456
rect 581730 200444 581736 200456
rect 578568 200416 581736 200444
rect 578568 200404 578574 200416
rect 581730 200404 581736 200416
rect 581788 200404 581794 200456
rect 580626 199996 580632 200048
rect 580684 200036 580690 200048
rect 589458 200036 589464 200048
rect 580684 200008 589464 200036
rect 580684 199996 580690 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 578878 198704 578884 198756
rect 578936 198744 578942 198756
rect 583018 198744 583024 198756
rect 578936 198716 583024 198744
rect 578936 198704 578942 198716
rect 583018 198704 583024 198716
rect 583076 198704 583082 198756
rect 671982 198636 671988 198688
rect 672040 198676 672046 198688
rect 675294 198676 675300 198688
rect 672040 198648 675300 198676
rect 672040 198636 672046 198648
rect 675294 198636 675300 198648
rect 675352 198636 675358 198688
rect 673086 197752 673092 197804
rect 673144 197792 673150 197804
rect 675294 197792 675300 197804
rect 673144 197764 675300 197792
rect 673144 197752 673150 197764
rect 675294 197752 675300 197764
rect 675352 197752 675358 197804
rect 578326 197412 578332 197464
rect 578384 197452 578390 197464
rect 580258 197452 580264 197464
rect 578384 197424 580264 197452
rect 578384 197412 578390 197424
rect 580258 197412 580264 197424
rect 580316 197412 580322 197464
rect 668026 197344 668032 197396
rect 668084 197384 668090 197396
rect 670142 197384 670148 197396
rect 668084 197356 670148 197384
rect 668084 197344 668090 197356
rect 670142 197344 670148 197356
rect 670200 197344 670206 197396
rect 584398 197276 584404 197328
rect 584456 197316 584462 197328
rect 589458 197316 589464 197328
rect 584456 197288 589464 197316
rect 584456 197276 584462 197288
rect 589458 197276 589464 197288
rect 589516 197276 589522 197328
rect 581730 196596 581736 196648
rect 581788 196636 581794 196648
rect 589642 196636 589648 196648
rect 581788 196608 589648 196636
rect 581788 196596 581794 196608
rect 589642 196596 589648 196608
rect 589700 196596 589706 196648
rect 579246 196120 579252 196172
rect 579304 196160 579310 196172
rect 581638 196160 581644 196172
rect 579304 196132 581644 196160
rect 579304 196120 579310 196132
rect 581638 196120 581644 196132
rect 581696 196120 581702 196172
rect 583202 195916 583208 195968
rect 583260 195956 583266 195968
rect 589458 195956 589464 195968
rect 583260 195928 589464 195956
rect 583260 195916 583266 195928
rect 589458 195916 589464 195928
rect 589516 195916 589522 195968
rect 42426 195644 42432 195696
rect 42484 195684 42490 195696
rect 43622 195684 43628 195696
rect 42484 195656 43628 195684
rect 42484 195644 42490 195656
rect 43622 195644 43628 195656
rect 43680 195644 43686 195696
rect 580902 194488 580908 194540
rect 580960 194528 580966 194540
rect 589458 194528 589464 194540
rect 580960 194500 589464 194528
rect 580960 194488 580966 194500
rect 589458 194488 589464 194500
rect 589516 194488 589522 194540
rect 578510 193400 578516 193452
rect 578568 193440 578574 193452
rect 583754 193440 583760 193452
rect 578568 193412 583760 193440
rect 578568 193400 578574 193412
rect 583754 193400 583760 193412
rect 583812 193400 583818 193452
rect 42426 193128 42432 193180
rect 42484 193168 42490 193180
rect 43806 193168 43812 193180
rect 42484 193140 43812 193168
rect 42484 193128 42490 193140
rect 43806 193128 43812 193140
rect 43864 193128 43870 193180
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 588538 191876 588544 191888
rect 579580 191848 588544 191876
rect 579580 191836 579586 191848
rect 588538 191836 588544 191848
rect 588596 191836 588602 191888
rect 42426 191768 42432 191820
rect 42484 191808 42490 191820
rect 44542 191808 44548 191820
rect 42484 191780 44548 191808
rect 42484 191768 42490 191780
rect 44542 191768 44548 191780
rect 44600 191768 44606 191820
rect 42426 191632 42432 191684
rect 42484 191672 42490 191684
rect 44358 191672 44364 191684
rect 42484 191644 44364 191672
rect 42484 191632 42490 191644
rect 44358 191632 44364 191644
rect 44416 191632 44422 191684
rect 583754 191088 583760 191140
rect 583812 191128 583818 191140
rect 590378 191128 590384 191140
rect 583812 191100 590384 191128
rect 583812 191088 583818 191100
rect 590378 191088 590384 191100
rect 590436 191088 590442 191140
rect 583018 190408 583024 190460
rect 583076 190448 583082 190460
rect 589458 190448 589464 190460
rect 583076 190420 589464 190448
rect 583076 190408 583082 190420
rect 589458 190408 589464 190420
rect 589516 190408 589522 190460
rect 42426 190340 42432 190392
rect 42484 190380 42490 190392
rect 42978 190380 42984 190392
rect 42484 190352 42984 190380
rect 42484 190340 42490 190352
rect 42978 190340 42984 190352
rect 43036 190340 43042 190392
rect 669268 190272 669274 190324
rect 669326 190312 669332 190324
rect 675294 190312 675300 190324
rect 669326 190284 675300 190312
rect 669326 190272 669332 190284
rect 675294 190272 675300 190284
rect 675352 190272 675358 190324
rect 578234 189048 578240 189100
rect 578292 189088 578298 189100
rect 585962 189088 585968 189100
rect 578292 189060 585968 189088
rect 578292 189048 578298 189060
rect 585962 189048 585968 189060
rect 586020 189048 586026 189100
rect 581638 188912 581644 188964
rect 581696 188952 581702 188964
rect 589458 188952 589464 188964
rect 581696 188924 589464 188952
rect 581696 188912 581702 188924
rect 589458 188912 589464 188924
rect 589516 188912 589522 188964
rect 579246 188776 579252 188828
rect 579304 188816 579310 188828
rect 581822 188816 581828 188828
rect 579304 188788 581828 188816
rect 579304 188776 579310 188788
rect 581822 188776 581828 188788
rect 581880 188776 581886 188828
rect 42426 187620 42432 187672
rect 42484 187660 42490 187672
rect 43438 187660 43444 187672
rect 42484 187632 43444 187660
rect 42484 187620 42490 187632
rect 43438 187620 43444 187632
rect 43496 187620 43502 187672
rect 580258 187552 580264 187604
rect 580316 187592 580322 187604
rect 589366 187592 589372 187604
rect 580316 187564 589372 187592
rect 580316 187552 580322 187564
rect 589366 187552 589372 187564
rect 589424 187552 589430 187604
rect 578510 187144 578516 187196
rect 578568 187184 578574 187196
rect 584582 187184 584588 187196
rect 578568 187156 584588 187184
rect 578568 187144 578574 187156
rect 584582 187144 584588 187156
rect 584640 187144 584646 187196
rect 578878 186192 578884 186244
rect 578936 186232 578942 186244
rect 589458 186232 589464 186244
rect 578936 186204 589464 186232
rect 578936 186192 578942 186204
rect 589458 186192 589464 186204
rect 589516 186192 589522 186244
rect 578326 185240 578332 185292
rect 578384 185280 578390 185292
rect 580442 185280 580448 185292
rect 578384 185252 580448 185280
rect 578384 185240 578390 185252
rect 580442 185240 580448 185252
rect 580500 185240 580506 185292
rect 668210 184832 668216 184884
rect 668268 184872 668274 184884
rect 672534 184872 672540 184884
rect 668268 184844 672540 184872
rect 668268 184832 668274 184844
rect 672534 184832 672540 184844
rect 672592 184832 672598 184884
rect 579522 183540 579528 183592
rect 579580 183580 579586 183592
rect 587158 183580 587164 183592
rect 579580 183552 587164 183580
rect 579580 183540 579586 183552
rect 587158 183540 587164 183552
rect 587216 183540 587222 183592
rect 42426 183472 42432 183524
rect 42484 183512 42490 183524
rect 44174 183512 44180 183524
rect 42484 183484 44180 183512
rect 42484 183472 42490 183484
rect 44174 183472 44180 183484
rect 44232 183472 44238 183524
rect 578878 182180 578884 182232
rect 578936 182220 578942 182232
rect 583018 182220 583024 182232
rect 578936 182192 583024 182220
rect 578936 182180 578942 182192
rect 583018 182180 583024 182192
rect 583076 182180 583082 182232
rect 578510 181296 578516 181348
rect 578568 181336 578574 181348
rect 581638 181336 581644 181348
rect 578568 181308 581644 181336
rect 578568 181296 578574 181308
rect 581638 181296 581644 181308
rect 581696 181296 581702 181348
rect 585962 180752 585968 180804
rect 586020 180792 586026 180804
rect 589458 180792 589464 180804
rect 586020 180764 589464 180792
rect 586020 180752 586026 180764
rect 589458 180752 589464 180764
rect 589516 180752 589522 180804
rect 578970 179664 578976 179716
rect 579028 179704 579034 179716
rect 585778 179704 585784 179716
rect 579028 179676 585784 179704
rect 579028 179664 579034 179676
rect 585778 179664 585784 179676
rect 585836 179664 585842 179716
rect 581822 179256 581828 179308
rect 581880 179296 581886 179308
rect 589550 179296 589556 179308
rect 581880 179268 589556 179296
rect 581880 179256 581886 179268
rect 589550 179256 589556 179268
rect 589608 179256 589614 179308
rect 578602 178304 578608 178356
rect 578660 178344 578666 178356
rect 580258 178344 580264 178356
rect 578660 178316 580264 178344
rect 578660 178304 578666 178316
rect 580258 178304 580264 178316
rect 580316 178304 580322 178356
rect 667382 178236 667388 178288
rect 667440 178276 667446 178288
rect 675478 178276 675484 178288
rect 667440 178248 675484 178276
rect 667440 178236 667446 178248
rect 675478 178236 675484 178248
rect 675536 178236 675542 178288
rect 670970 178100 670976 178152
rect 671028 178140 671034 178152
rect 675478 178140 675484 178152
rect 671028 178112 675484 178140
rect 671028 178100 671034 178112
rect 675478 178100 675484 178112
rect 675536 178100 675542 178152
rect 584582 177964 584588 178016
rect 584640 178004 584646 178016
rect 589458 178004 589464 178016
rect 584640 177976 589464 178004
rect 584640 177964 584646 177976
rect 589458 177964 589464 177976
rect 589516 177964 589522 178016
rect 668578 177964 668584 178016
rect 668636 178004 668642 178016
rect 672534 178004 672540 178016
rect 668636 177976 672540 178004
rect 668636 177964 668642 177976
rect 672534 177964 672540 177976
rect 672592 177964 672598 178016
rect 673546 177692 673552 177744
rect 673604 177732 673610 177744
rect 675478 177732 675484 177744
rect 673604 177704 675484 177732
rect 673604 177692 673610 177704
rect 675478 177692 675484 177704
rect 675536 177692 675542 177744
rect 579522 176808 579528 176860
rect 579580 176848 579586 176860
rect 584398 176848 584404 176860
rect 579580 176820 584404 176848
rect 579580 176808 579586 176820
rect 584398 176808 584404 176820
rect 584456 176808 584462 176860
rect 673914 176808 673920 176860
rect 673972 176848 673978 176860
rect 675478 176848 675484 176860
rect 673972 176820 675484 176848
rect 673972 176808 673978 176820
rect 675478 176808 675484 176820
rect 675536 176808 675542 176860
rect 580442 176536 580448 176588
rect 580500 176576 580506 176588
rect 589458 176576 589464 176588
rect 580500 176548 589464 176576
rect 580500 176536 580506 176548
rect 589458 176536 589464 176548
rect 589516 176536 589522 176588
rect 667842 175380 667848 175432
rect 667900 175420 667906 175432
rect 675478 175420 675484 175432
rect 667900 175392 675484 175420
rect 667900 175380 667906 175392
rect 675478 175380 675484 175392
rect 675536 175380 675542 175432
rect 673362 175176 673368 175228
rect 673420 175216 673426 175228
rect 675478 175216 675484 175228
rect 673420 175188 675484 175216
rect 673420 175176 673426 175188
rect 675478 175176 675484 175188
rect 675536 175176 675542 175228
rect 579614 174496 579620 174548
rect 579672 174536 579678 174548
rect 589918 174536 589924 174548
rect 579672 174508 589924 174536
rect 579672 174496 579678 174508
rect 589918 174496 589924 174508
rect 589976 174496 589982 174548
rect 672994 174360 673000 174412
rect 673052 174400 673058 174412
rect 675478 174400 675484 174412
rect 673052 174372 675484 174400
rect 673052 174360 673058 174372
rect 675478 174360 675484 174372
rect 675536 174360 675542 174412
rect 587158 173816 587164 173868
rect 587216 173856 587222 173868
rect 589274 173856 589280 173868
rect 587216 173828 589280 173856
rect 587216 173816 587222 173828
rect 589274 173816 589280 173828
rect 589332 173816 589338 173868
rect 578326 172524 578332 172576
rect 578384 172564 578390 172576
rect 583202 172564 583208 172576
rect 578384 172536 583208 172564
rect 578384 172524 578390 172536
rect 583202 172524 583208 172536
rect 583260 172524 583266 172576
rect 583018 172388 583024 172440
rect 583076 172428 583082 172440
rect 589366 172428 589372 172440
rect 583076 172400 589372 172428
rect 583076 172388 583082 172400
rect 589366 172388 589372 172400
rect 589424 172388 589430 172440
rect 579062 171640 579068 171692
rect 579120 171680 579126 171692
rect 581822 171680 581828 171692
rect 579120 171652 581828 171680
rect 579120 171640 579126 171652
rect 581822 171640 581828 171652
rect 581880 171640 581886 171692
rect 670418 171096 670424 171148
rect 670476 171136 670482 171148
rect 675478 171136 675484 171148
rect 670476 171108 675484 171136
rect 670476 171096 670482 171108
rect 675478 171096 675484 171108
rect 675536 171096 675542 171148
rect 581638 170960 581644 171012
rect 581696 171000 581702 171012
rect 589458 171000 589464 171012
rect 581696 170972 589464 171000
rect 581696 170960 581702 170972
rect 589458 170960 589464 170972
rect 589516 170960 589522 171012
rect 579522 169736 579528 169788
rect 579580 169776 579586 169788
rect 588722 169776 588728 169788
rect 579580 169748 588728 169776
rect 579580 169736 579586 169748
rect 588722 169736 588728 169748
rect 588780 169736 588786 169788
rect 585778 169600 585784 169652
rect 585836 169640 585842 169652
rect 589458 169640 589464 169652
rect 585836 169612 589464 169640
rect 585836 169600 585842 169612
rect 589458 169600 589464 169612
rect 589516 169600 589522 169652
rect 671798 169464 671804 169516
rect 671856 169504 671862 169516
rect 675478 169504 675484 169516
rect 671856 169476 675484 169504
rect 671856 169464 671862 169476
rect 675478 169464 675484 169476
rect 675536 169464 675542 169516
rect 670602 169056 670608 169108
rect 670660 169096 670666 169108
rect 675478 169096 675484 169108
rect 670660 169068 675484 169096
rect 670660 169056 670666 169068
rect 675478 169056 675484 169068
rect 675536 169056 675542 169108
rect 673178 168648 673184 168700
rect 673236 168688 673242 168700
rect 675478 168688 675484 168700
rect 673236 168660 675484 168688
rect 673236 168648 673242 168660
rect 675478 168648 675484 168660
rect 675536 168648 675542 168700
rect 578234 168376 578240 168428
rect 578292 168416 578298 168428
rect 580442 168416 580448 168428
rect 578292 168388 580448 168416
rect 578292 168376 578298 168388
rect 580442 168376 580448 168388
rect 580500 168376 580506 168428
rect 580258 168240 580264 168292
rect 580316 168280 580322 168292
rect 589458 168280 589464 168292
rect 580316 168252 589464 168280
rect 580316 168240 580322 168252
rect 589458 168240 589464 168252
rect 589516 168240 589522 168292
rect 672626 167016 672632 167068
rect 672684 167056 672690 167068
rect 675478 167056 675484 167068
rect 672684 167028 675484 167056
rect 672684 167016 672690 167028
rect 675478 167016 675484 167028
rect 675536 167016 675542 167068
rect 669958 166812 669964 166864
rect 670016 166852 670022 166864
rect 675478 166852 675484 166864
rect 670016 166824 675484 166852
rect 670016 166812 670022 166824
rect 675478 166812 675484 166824
rect 675536 166812 675542 166864
rect 579614 166268 579620 166320
rect 579672 166308 579678 166320
rect 590378 166308 590384 166320
rect 579672 166280 590384 166308
rect 579672 166268 579678 166280
rect 590378 166268 590384 166280
rect 590436 166268 590442 166320
rect 579062 165588 579068 165640
rect 579120 165628 579126 165640
rect 584582 165628 584588 165640
rect 579120 165600 584588 165628
rect 579120 165588 579126 165600
rect 584582 165588 584588 165600
rect 584640 165588 584646 165640
rect 589458 165560 589464 165572
rect 586486 165532 589464 165560
rect 584398 165452 584404 165504
rect 584456 165492 584462 165504
rect 586486 165492 586514 165532
rect 589458 165520 589464 165532
rect 589516 165520 589522 165572
rect 584456 165464 586514 165492
rect 584456 165452 584462 165464
rect 579522 164296 579528 164348
rect 579580 164336 579586 164348
rect 583018 164336 583024 164348
rect 579580 164308 583024 164336
rect 579580 164296 579586 164308
rect 583018 164296 583024 164308
rect 583076 164296 583082 164348
rect 578694 162868 578700 162920
rect 578752 162908 578758 162920
rect 581638 162908 581644 162920
rect 578752 162880 581644 162908
rect 578752 162868 578758 162880
rect 581638 162868 581644 162880
rect 581696 162868 581702 162920
rect 583202 162800 583208 162852
rect 583260 162840 583266 162852
rect 589458 162840 589464 162852
rect 583260 162812 589464 162840
rect 583260 162800 583266 162812
rect 589458 162800 589464 162812
rect 589516 162800 589522 162852
rect 671798 162052 671804 162104
rect 671856 162092 671862 162104
rect 673546 162092 673552 162104
rect 671856 162064 673552 162092
rect 671856 162052 671862 162064
rect 673546 162052 673552 162064
rect 673604 162052 673610 162104
rect 581822 161372 581828 161424
rect 581880 161412 581886 161424
rect 589458 161412 589464 161424
rect 581880 161384 589464 161412
rect 581880 161372 581886 161384
rect 589458 161372 589464 161384
rect 589516 161372 589522 161424
rect 578510 160216 578516 160268
rect 578568 160256 578574 160268
rect 580258 160256 580264 160268
rect 578568 160228 580264 160256
rect 578568 160216 578574 160228
rect 580258 160216 580264 160228
rect 580316 160216 580322 160268
rect 579522 158720 579528 158772
rect 579580 158760 579586 158772
rect 588538 158760 588544 158772
rect 579580 158732 588544 158760
rect 579580 158720 579586 158732
rect 588538 158720 588544 158732
rect 588596 158720 588602 158772
rect 580442 158584 580448 158636
rect 580500 158624 580506 158636
rect 589458 158624 589464 158636
rect 580500 158596 589464 158624
rect 580500 158584 580506 158596
rect 589458 158584 589464 158596
rect 589516 158584 589522 158636
rect 579614 156612 579620 156664
rect 579672 156652 579678 156664
rect 589918 156652 589924 156664
rect 579672 156624 589924 156652
rect 579672 156612 579678 156624
rect 589918 156612 589924 156624
rect 589976 156612 589982 156664
rect 673546 155796 673552 155848
rect 673604 155836 673610 155848
rect 675386 155836 675392 155848
rect 673604 155808 675392 155836
rect 673604 155796 673610 155808
rect 675386 155796 675392 155808
rect 675444 155796 675450 155848
rect 670418 154912 670424 154964
rect 670476 154952 670482 154964
rect 675110 154952 675116 154964
rect 670476 154924 675116 154952
rect 670476 154912 670482 154924
rect 675110 154912 675116 154924
rect 675168 154912 675174 154964
rect 579246 154572 579252 154624
rect 579304 154612 579310 154624
rect 587342 154612 587348 154624
rect 579304 154584 587348 154612
rect 579304 154572 579310 154584
rect 587342 154572 587348 154584
rect 587400 154572 587406 154624
rect 584582 154436 584588 154488
rect 584640 154476 584646 154488
rect 589366 154476 589372 154488
rect 584640 154448 589372 154476
rect 584640 154436 584646 154448
rect 589366 154436 589372 154448
rect 589424 154436 589430 154488
rect 579246 153280 579252 153332
rect 579304 153320 579310 153332
rect 585778 153320 585784 153332
rect 579304 153292 585784 153320
rect 579304 153280 579310 153292
rect 585778 153280 585784 153292
rect 585836 153280 585842 153332
rect 583018 153076 583024 153128
rect 583076 153116 583082 153128
rect 589458 153116 589464 153128
rect 583076 153088 589464 153116
rect 583076 153076 583082 153088
rect 589458 153076 589464 153088
rect 589516 153076 589522 153128
rect 578694 152260 578700 152312
rect 578752 152300 578758 152312
rect 584398 152300 584404 152312
rect 578752 152272 584404 152300
rect 578752 152260 578758 152272
rect 584398 152260 584404 152272
rect 584456 152260 584462 152312
rect 673178 151716 673184 151768
rect 673236 151756 673242 151768
rect 675110 151756 675116 151768
rect 673236 151728 675116 151756
rect 673236 151716 673242 151728
rect 675110 151716 675116 151728
rect 675168 151716 675174 151768
rect 581638 151648 581644 151700
rect 581696 151688 581702 151700
rect 589458 151688 589464 151700
rect 581696 151660 589464 151688
rect 581696 151648 581702 151660
rect 589458 151648 589464 151660
rect 589516 151648 589522 151700
rect 579154 150424 579160 150476
rect 579212 150464 579218 150476
rect 583202 150464 583208 150476
rect 579212 150436 583208 150464
rect 579212 150424 579218 150436
rect 583202 150424 583208 150436
rect 583260 150424 583266 150476
rect 670602 150356 670608 150408
rect 670660 150396 670666 150408
rect 674926 150396 674932 150408
rect 670660 150368 674932 150396
rect 670660 150356 670666 150368
rect 674926 150356 674932 150368
rect 674984 150356 674990 150408
rect 578878 150288 578884 150340
rect 578936 150328 578942 150340
rect 589458 150328 589464 150340
rect 578936 150300 589464 150328
rect 578936 150288 578942 150300
rect 589458 150288 589464 150300
rect 589516 150288 589522 150340
rect 578878 149064 578884 149116
rect 578936 149104 578942 149116
rect 581638 149104 581644 149116
rect 578936 149076 581644 149104
rect 578936 149064 578942 149076
rect 581638 149064 581644 149076
rect 581696 149064 581702 149116
rect 674466 148928 674472 148980
rect 674524 148968 674530 148980
rect 675294 148968 675300 148980
rect 674524 148940 675300 148968
rect 674524 148928 674530 148940
rect 675294 148928 675300 148940
rect 675352 148928 675358 148980
rect 668762 148180 668768 148232
rect 668820 148220 668826 148232
rect 674098 148220 674104 148232
rect 668820 148192 674104 148220
rect 668820 148180 668826 148192
rect 674098 148180 674104 148192
rect 674156 148180 674162 148232
rect 579522 147636 579528 147688
rect 579580 147676 579586 147688
rect 588722 147676 588728 147688
rect 579580 147648 588728 147676
rect 579580 147636 579586 147648
rect 588722 147636 588728 147648
rect 588780 147636 588786 147688
rect 579246 147500 579252 147552
rect 579304 147540 579310 147552
rect 591298 147540 591304 147552
rect 579304 147512 591304 147540
rect 579304 147500 579310 147512
rect 591298 147500 591304 147512
rect 591356 147500 591362 147552
rect 580258 147364 580264 147416
rect 580316 147404 580322 147416
rect 589458 147404 589464 147416
rect 580316 147376 589464 147404
rect 580316 147364 580322 147376
rect 589458 147364 589464 147376
rect 589516 147364 589522 147416
rect 668762 146208 668768 146260
rect 668820 146248 668826 146260
rect 671430 146248 671436 146260
rect 668820 146220 671436 146248
rect 668820 146208 668826 146220
rect 671430 146208 671436 146220
rect 671488 146208 671494 146260
rect 579614 144168 579620 144220
rect 579672 144208 579678 144220
rect 590378 144208 590384 144220
rect 579672 144180 590384 144208
rect 579672 144168 579678 144180
rect 590378 144168 590384 144180
rect 590436 144168 590442 144220
rect 668762 144168 668768 144220
rect 668820 144208 668826 144220
rect 674282 144208 674288 144220
rect 668820 144180 674288 144208
rect 668820 144168 668826 144180
rect 674282 144168 674288 144180
rect 674340 144168 674346 144220
rect 578510 143624 578516 143676
rect 578568 143664 578574 143676
rect 580258 143664 580264 143676
rect 578568 143636 580264 143664
rect 578568 143624 578574 143636
rect 580258 143624 580264 143636
rect 580316 143624 580322 143676
rect 587342 143488 587348 143540
rect 587400 143528 587406 143540
rect 590010 143528 590016 143540
rect 587400 143500 590016 143528
rect 587400 143488 587406 143500
rect 590010 143488 590016 143500
rect 590068 143488 590074 143540
rect 579522 142128 579528 142180
rect 579580 142168 579586 142180
rect 587158 142168 587164 142180
rect 579580 142140 587164 142168
rect 579580 142128 579586 142140
rect 587158 142128 587164 142140
rect 587216 142128 587222 142180
rect 585778 141992 585784 142044
rect 585836 142032 585842 142044
rect 589458 142032 589464 142044
rect 585836 142004 589464 142032
rect 585836 141992 585842 142004
rect 589458 141992 589464 142004
rect 589516 141992 589522 142044
rect 584398 140700 584404 140752
rect 584456 140740 584462 140752
rect 589458 140740 589464 140752
rect 584456 140712 589464 140740
rect 584456 140700 584462 140712
rect 589458 140700 589464 140712
rect 589516 140700 589522 140752
rect 668762 140700 668768 140752
rect 668820 140740 668826 140752
rect 671614 140740 671620 140752
rect 668820 140712 671620 140740
rect 668820 140700 668826 140712
rect 671614 140700 671620 140712
rect 671672 140700 671678 140752
rect 579522 139408 579528 139460
rect 579580 139448 579586 139460
rect 584582 139448 584588 139460
rect 579580 139420 584588 139448
rect 579580 139408 579586 139420
rect 584582 139408 584588 139420
rect 584640 139408 584646 139460
rect 668762 139340 668768 139392
rect 668820 139380 668826 139392
rect 671154 139380 671160 139392
rect 668820 139352 671160 139380
rect 668820 139340 668826 139352
rect 671154 139340 671160 139352
rect 671212 139340 671218 139392
rect 668026 137980 668032 138032
rect 668084 138020 668090 138032
rect 672166 138020 672172 138032
rect 668084 137992 672172 138020
rect 668084 137980 668090 137992
rect 672166 137980 672172 137992
rect 672224 137980 672230 138032
rect 579246 137912 579252 137964
rect 579304 137952 579310 137964
rect 583018 137952 583024 137964
rect 579304 137924 583024 137952
rect 579304 137912 579310 137924
rect 583018 137912 583024 137924
rect 583076 137912 583082 137964
rect 583202 137912 583208 137964
rect 583260 137952 583266 137964
rect 589458 137952 589464 137964
rect 583260 137924 589464 137952
rect 583260 137912 583266 137924
rect 589458 137912 589464 137924
rect 589516 137912 589522 137964
rect 668578 137300 668584 137352
rect 668636 137340 668642 137352
rect 669130 137340 669136 137352
rect 668636 137312 669136 137340
rect 668636 137300 668642 137312
rect 669130 137300 669136 137312
rect 669188 137300 669194 137352
rect 581638 136484 581644 136536
rect 581696 136524 581702 136536
rect 589366 136524 589372 136536
rect 581696 136496 589372 136524
rect 581696 136484 581702 136496
rect 589366 136484 589372 136496
rect 589424 136484 589430 136536
rect 579062 135328 579068 135380
rect 579120 135368 579126 135380
rect 581086 135368 581092 135380
rect 579120 135340 581092 135368
rect 579120 135328 579126 135340
rect 581086 135328 581092 135340
rect 581144 135328 581150 135380
rect 578234 134512 578240 134564
rect 578292 134552 578298 134564
rect 585962 134552 585968 134564
rect 578292 134524 585968 134552
rect 578292 134512 578298 134524
rect 585962 134512 585968 134524
rect 586020 134512 586026 134564
rect 669222 133764 669228 133816
rect 669280 133804 669286 133816
rect 672810 133804 672816 133816
rect 669280 133776 672816 133804
rect 669280 133764 669286 133776
rect 672810 133764 672816 133776
rect 672868 133764 672874 133816
rect 669406 133356 669412 133408
rect 669464 133396 669470 133408
rect 675478 133396 675484 133408
rect 669464 133368 675484 133396
rect 669464 133356 669470 133368
rect 675478 133356 675484 133368
rect 675536 133356 675542 133408
rect 581086 133152 581092 133204
rect 581144 133192 581150 133204
rect 589918 133192 589924 133204
rect 581144 133164 589924 133192
rect 581144 133152 581150 133164
rect 589918 133152 589924 133164
rect 589976 133152 589982 133204
rect 578510 132880 578516 132932
rect 578568 132920 578574 132932
rect 581638 132920 581644 132932
rect 578568 132892 581644 132920
rect 578568 132880 578574 132892
rect 581638 132880 581644 132892
rect 581696 132880 581702 132932
rect 667198 132880 667204 132932
rect 667256 132920 667262 132932
rect 675478 132920 675484 132932
rect 667256 132892 675484 132920
rect 667256 132880 667262 132892
rect 675478 132880 675484 132892
rect 675536 132880 675542 132932
rect 667566 132744 667572 132796
rect 667624 132784 667630 132796
rect 675478 132784 675484 132796
rect 667624 132756 675484 132784
rect 667624 132744 667630 132756
rect 675478 132744 675484 132756
rect 675536 132744 675542 132796
rect 580258 132336 580264 132388
rect 580316 132376 580322 132388
rect 589458 132376 589464 132388
rect 580316 132348 589464 132376
rect 580316 132336 580322 132348
rect 589458 132336 589464 132348
rect 589516 132336 589522 132388
rect 673914 132132 673920 132184
rect 673972 132172 673978 132184
rect 675478 132172 675484 132184
rect 673972 132144 675484 132172
rect 673972 132132 673978 132144
rect 675478 132132 675484 132144
rect 675536 132132 675542 132184
rect 668394 131180 668400 131232
rect 668452 131220 668458 131232
rect 668762 131220 668768 131232
rect 668452 131192 668768 131220
rect 668452 131180 668458 131192
rect 668762 131180 668768 131192
rect 668820 131220 668826 131232
rect 675478 131220 675484 131232
rect 668820 131192 675484 131220
rect 668820 131180 668826 131192
rect 675478 131180 675484 131192
rect 675536 131180 675542 131232
rect 668302 131044 668308 131096
rect 668360 131084 668366 131096
rect 670234 131084 670240 131096
rect 668360 131056 670240 131084
rect 668360 131044 668366 131056
rect 670234 131044 670240 131056
rect 670292 131044 670298 131096
rect 671338 130840 671344 130892
rect 671396 130880 671402 130892
rect 675478 130880 675484 130892
rect 671396 130852 675484 130880
rect 671396 130840 671402 130852
rect 675478 130840 675484 130852
rect 675536 130840 675542 130892
rect 673362 130500 673368 130552
rect 673420 130540 673426 130552
rect 675478 130540 675484 130552
rect 673420 130512 675484 130540
rect 673420 130500 673426 130512
rect 675478 130500 675484 130512
rect 675536 130500 675542 130552
rect 578418 130364 578424 130416
rect 578476 130404 578482 130416
rect 588538 130404 588544 130416
rect 578476 130376 588544 130404
rect 578476 130364 578482 130376
rect 588538 130364 588544 130376
rect 588596 130364 588602 130416
rect 578602 129888 578608 129940
rect 578660 129928 578666 129940
rect 580442 129928 580448 129940
rect 578660 129900 580448 129928
rect 578660 129888 578666 129900
rect 580442 129888 580448 129900
rect 580500 129888 580506 129940
rect 668578 129888 668584 129940
rect 668636 129928 668642 129940
rect 675478 129928 675484 129940
rect 668636 129900 675484 129928
rect 668636 129888 668642 129900
rect 675478 129888 675484 129900
rect 675536 129888 675542 129940
rect 584582 129684 584588 129736
rect 584640 129724 584646 129736
rect 589458 129724 589464 129736
rect 584640 129696 589464 129724
rect 584640 129684 584646 129696
rect 589458 129684 589464 129696
rect 589516 129684 589522 129736
rect 672994 129684 673000 129736
rect 673052 129724 673058 129736
rect 675478 129724 675484 129736
rect 673052 129696 675484 129724
rect 673052 129684 673058 129696
rect 675478 129684 675484 129696
rect 675536 129684 675542 129736
rect 669222 129616 669228 129668
rect 669280 129656 669286 129668
rect 672350 129656 672356 129668
rect 669280 129628 672356 129656
rect 669280 129616 669286 129628
rect 672350 129616 672356 129628
rect 672408 129616 672414 129668
rect 668210 129208 668216 129260
rect 668268 129248 668274 129260
rect 669774 129248 669780 129260
rect 668268 129220 669780 129248
rect 668268 129208 668274 129220
rect 669774 129208 669780 129220
rect 669832 129208 669838 129260
rect 578878 128324 578884 128376
rect 578936 128364 578942 128376
rect 578936 128336 583800 128364
rect 578936 128324 578942 128336
rect 583772 128296 583800 128336
rect 668946 128324 668952 128376
rect 669004 128364 669010 128376
rect 675478 128364 675484 128376
rect 669004 128336 675484 128364
rect 669004 128324 669010 128336
rect 675478 128324 675484 128336
rect 675536 128324 675542 128376
rect 583772 128268 586514 128296
rect 586486 128228 586514 128268
rect 589458 128228 589464 128240
rect 586486 128200 589464 128228
rect 589458 128188 589464 128200
rect 589516 128188 589522 128240
rect 578326 126964 578332 127016
rect 578384 127004 578390 127016
rect 580258 127004 580264 127016
rect 578384 126976 580264 127004
rect 578384 126964 578390 126976
rect 580258 126964 580264 126976
rect 580316 126964 580322 127016
rect 587158 126896 587164 126948
rect 587216 126936 587222 126948
rect 589734 126936 589740 126948
rect 587216 126908 589740 126936
rect 587216 126896 587222 126908
rect 589734 126896 589740 126908
rect 589792 126896 589798 126948
rect 579430 126216 579436 126268
rect 579488 126256 579494 126268
rect 587342 126256 587348 126268
rect 579488 126228 587348 126256
rect 579488 126216 579494 126228
rect 587342 126216 587348 126228
rect 587400 126216 587406 126268
rect 675018 126148 675024 126200
rect 675076 126188 675082 126200
rect 675478 126188 675484 126200
rect 675076 126160 675484 126188
rect 675076 126148 675082 126160
rect 675478 126148 675484 126160
rect 675536 126148 675542 126200
rect 675846 126148 675852 126200
rect 675904 126188 675910 126200
rect 676398 126188 676404 126200
rect 675904 126160 676404 126188
rect 675904 126148 675910 126160
rect 676398 126148 676404 126160
rect 676456 126148 676462 126200
rect 673178 125944 673184 125996
rect 673236 125984 673242 125996
rect 675478 125984 675484 125996
rect 673236 125956 675484 125984
rect 673236 125944 673242 125956
rect 675478 125944 675484 125956
rect 675536 125944 675542 125996
rect 578510 125808 578516 125860
rect 578568 125848 578574 125860
rect 584398 125848 584404 125860
rect 578568 125820 584404 125848
rect 578568 125808 578574 125820
rect 584398 125808 584404 125820
rect 584456 125808 584462 125860
rect 672994 125740 673000 125792
rect 673052 125780 673058 125792
rect 675478 125780 675484 125792
rect 673052 125752 675484 125780
rect 673052 125740 673058 125752
rect 675478 125740 675484 125752
rect 675536 125740 675542 125792
rect 585962 124856 585968 124908
rect 586020 124896 586026 124908
rect 590378 124896 590384 124908
rect 586020 124868 590384 124896
rect 586020 124856 586026 124868
rect 590378 124856 590384 124868
rect 590436 124856 590442 124908
rect 578878 124176 578884 124228
rect 578936 124216 578942 124228
rect 585778 124216 585784 124228
rect 578936 124188 585784 124216
rect 578936 124176 578942 124188
rect 585778 124176 585784 124188
rect 585836 124176 585842 124228
rect 583018 124040 583024 124092
rect 583076 124080 583082 124092
rect 589458 124080 589464 124092
rect 583076 124052 589464 124080
rect 583076 124040 583082 124052
rect 589458 124040 589464 124052
rect 589516 124040 589522 124092
rect 673362 123904 673368 123956
rect 673420 123944 673426 123956
rect 675478 123944 675484 123956
rect 673420 123916 675484 123944
rect 673420 123904 673426 123916
rect 675478 123904 675484 123916
rect 675536 123904 675542 123956
rect 674006 123088 674012 123140
rect 674064 123128 674070 123140
rect 675478 123128 675484 123140
rect 674064 123100 675484 123128
rect 674064 123088 674070 123100
rect 675478 123088 675484 123100
rect 675536 123088 675542 123140
rect 670142 122408 670148 122460
rect 670200 122448 670206 122460
rect 675478 122448 675484 122460
rect 670200 122420 675484 122448
rect 670200 122408 670206 122420
rect 675478 122408 675484 122420
rect 675536 122408 675542 122460
rect 579522 121456 579528 121508
rect 579580 121496 579586 121508
rect 583018 121496 583024 121508
rect 579580 121468 583024 121496
rect 579580 121456 579586 121468
rect 583018 121456 583024 121468
rect 583076 121456 583082 121508
rect 671522 121388 671528 121440
rect 671580 121428 671586 121440
rect 675478 121428 675484 121440
rect 671580 121400 675484 121428
rect 671580 121388 671586 121400
rect 675478 121388 675484 121400
rect 675536 121388 675542 121440
rect 580258 120708 580264 120760
rect 580316 120748 580322 120760
rect 589918 120748 589924 120760
rect 580316 120720 589924 120748
rect 580316 120708 580322 120720
rect 589918 120708 589924 120720
rect 589976 120708 589982 120760
rect 581638 120028 581644 120080
rect 581696 120068 581702 120080
rect 589458 120068 589464 120080
rect 581696 120040 589464 120068
rect 581696 120028 581702 120040
rect 589458 120028 589464 120040
rect 589516 120028 589522 120080
rect 669222 120028 669228 120080
rect 669280 120068 669286 120080
rect 671798 120068 671804 120080
rect 669280 120040 671804 120068
rect 669280 120028 669286 120040
rect 671798 120028 671804 120040
rect 671856 120028 671862 120080
rect 579246 118668 579252 118720
rect 579304 118708 579310 118720
rect 587158 118708 587164 118720
rect 579304 118680 587164 118708
rect 579304 118668 579310 118680
rect 587158 118668 587164 118680
rect 587216 118668 587222 118720
rect 579062 117308 579068 117360
rect 579120 117348 579126 117360
rect 581638 117348 581644 117360
rect 579120 117320 581644 117348
rect 579120 117308 579126 117320
rect 581638 117308 581644 117320
rect 581696 117308 581702 117360
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 679618 117280 679624 117292
rect 675904 117252 679624 117280
rect 675904 117240 675910 117252
rect 679618 117240 679624 117252
rect 679676 117240 679682 117292
rect 580442 117172 580448 117224
rect 580500 117212 580506 117224
rect 589458 117212 589464 117224
rect 580500 117184 589464 117212
rect 580500 117172 580506 117184
rect 589458 117172 589464 117184
rect 589516 117172 589522 117224
rect 578326 116968 578332 117020
rect 578384 117008 578390 117020
rect 580258 117008 580264 117020
rect 578384 116980 580264 117008
rect 578384 116968 578390 116980
rect 580258 116968 580264 116980
rect 580316 116968 580322 117020
rect 587342 115880 587348 115932
rect 587400 115920 587406 115932
rect 589274 115920 589280 115932
rect 587400 115892 589280 115920
rect 587400 115880 587406 115892
rect 589274 115880 589280 115892
rect 589332 115880 589338 115932
rect 669222 115812 669228 115864
rect 669280 115852 669286 115864
rect 672626 115852 672632 115864
rect 669280 115824 672632 115852
rect 669280 115812 669286 115824
rect 672626 115812 672632 115824
rect 672684 115812 672690 115864
rect 675018 115472 675024 115524
rect 675076 115512 675082 115524
rect 675386 115512 675392 115524
rect 675076 115484 675392 115512
rect 675076 115472 675082 115484
rect 675386 115472 675392 115484
rect 675444 115472 675450 115524
rect 585778 114452 585784 114504
rect 585836 114492 585842 114504
rect 589458 114492 589464 114504
rect 585836 114464 589464 114492
rect 585836 114452 585842 114464
rect 589458 114452 589464 114464
rect 589516 114452 589522 114504
rect 669222 114112 669228 114164
rect 669280 114152 669286 114164
rect 674006 114152 674012 114164
rect 669280 114124 674012 114152
rect 669280 114112 669286 114124
rect 674006 114112 674012 114124
rect 674064 114112 674070 114164
rect 668302 112820 668308 112872
rect 668360 112860 668366 112872
rect 670142 112860 670148 112872
rect 668360 112832 670148 112860
rect 668360 112820 668366 112832
rect 670142 112820 670148 112832
rect 670200 112820 670206 112872
rect 584398 111732 584404 111784
rect 584456 111772 584462 111784
rect 589458 111772 589464 111784
rect 584456 111744 589464 111772
rect 584456 111732 584462 111744
rect 589458 111732 589464 111744
rect 589516 111732 589522 111784
rect 669038 111732 669044 111784
rect 669096 111772 669102 111784
rect 671522 111772 671528 111784
rect 669096 111744 671528 111772
rect 669096 111732 669102 111744
rect 671522 111732 671528 111744
rect 671580 111732 671586 111784
rect 673178 111732 673184 111784
rect 673236 111772 673242 111784
rect 675110 111772 675116 111784
rect 673236 111744 675116 111772
rect 673236 111732 673242 111744
rect 675110 111732 675116 111744
rect 675168 111732 675174 111784
rect 672994 111120 673000 111172
rect 673052 111160 673058 111172
rect 675386 111160 675392 111172
rect 673052 111132 675392 111160
rect 673052 111120 673058 111132
rect 675386 111120 675392 111132
rect 675444 111120 675450 111172
rect 578878 108944 578884 108996
rect 578936 108984 578942 108996
rect 589458 108984 589464 108996
rect 578936 108956 589464 108984
rect 578936 108944 578942 108956
rect 589458 108944 589464 108956
rect 589516 108944 589522 108996
rect 669130 108944 669136 108996
rect 669188 108984 669194 108996
rect 671338 108984 671344 108996
rect 669188 108956 671344 108984
rect 669188 108944 669194 108956
rect 671338 108944 671344 108956
rect 671396 108944 671402 108996
rect 583018 107584 583024 107636
rect 583076 107624 583082 107636
rect 589366 107624 589372 107636
rect 583076 107596 589372 107624
rect 583076 107584 583082 107596
rect 589366 107584 589372 107596
rect 589424 107584 589430 107636
rect 674190 106972 674196 107024
rect 674248 107012 674254 107024
rect 675294 107012 675300 107024
rect 674248 106984 675300 107012
rect 674248 106972 674254 106984
rect 675294 106972 675300 106984
rect 675352 106972 675358 107024
rect 673362 106496 673368 106548
rect 673420 106536 673426 106548
rect 675110 106536 675116 106548
rect 673420 106508 675116 106536
rect 673420 106496 673426 106508
rect 675110 106496 675116 106508
rect 675168 106496 675174 106548
rect 587158 106224 587164 106276
rect 587216 106264 587222 106276
rect 589274 106264 589280 106276
rect 587216 106236 589280 106264
rect 587216 106224 587222 106236
rect 589274 106224 589280 106236
rect 589332 106224 589338 106276
rect 581638 104796 581644 104848
rect 581696 104836 581702 104848
rect 589366 104836 589372 104848
rect 581696 104808 589372 104836
rect 581696 104796 581702 104808
rect 589366 104796 589372 104808
rect 589424 104796 589430 104848
rect 580258 102076 580264 102128
rect 580316 102116 580322 102128
rect 589458 102116 589464 102128
rect 580316 102088 589464 102116
rect 580316 102076 580322 102088
rect 589458 102076 589464 102088
rect 589516 102076 589522 102128
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 632146 99192 632152 99204
rect 623740 99164 632152 99192
rect 623740 99152 623746 99164
rect 632146 99152 632152 99164
rect 632204 99152 632210 99204
rect 625062 99016 625068 99068
rect 625120 99056 625126 99068
rect 634446 99056 634452 99068
rect 625120 99028 634452 99056
rect 625120 99016 625126 99028
rect 634446 99016 634452 99028
rect 634504 99016 634510 99068
rect 629754 98880 629760 98932
rect 629812 98920 629818 98932
rect 640978 98920 640984 98932
rect 629812 98892 640984 98920
rect 629812 98880 629818 98892
rect 640978 98880 640984 98892
rect 641036 98880 641042 98932
rect 621658 98744 621664 98796
rect 621716 98784 621722 98796
rect 628374 98784 628380 98796
rect 621716 98756 628380 98784
rect 621716 98744 621722 98756
rect 628374 98744 628380 98756
rect 628432 98744 628438 98796
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 639874 98784 639880 98796
rect 629076 98756 639880 98784
rect 629076 98744 629082 98756
rect 639874 98744 639880 98756
rect 639932 98744 639938 98796
rect 622302 98608 622308 98660
rect 622360 98648 622366 98660
rect 629478 98648 629484 98660
rect 622360 98620 629484 98648
rect 622360 98608 622366 98620
rect 629478 98608 629484 98620
rect 629536 98608 629542 98660
rect 630490 98608 630496 98660
rect 630548 98648 630554 98660
rect 642082 98648 642088 98660
rect 630548 98620 642088 98648
rect 630548 98608 630554 98620
rect 642082 98608 642088 98620
rect 642140 98608 642146 98660
rect 577498 97928 577504 97980
rect 577556 97968 577562 97980
rect 577556 97940 586514 97968
rect 577556 97928 577562 97940
rect 586486 97832 586514 97940
rect 594058 97928 594064 97980
rect 594116 97968 594122 97980
rect 596174 97968 596180 97980
rect 594116 97940 596180 97968
rect 594116 97928 594122 97940
rect 596174 97928 596180 97940
rect 596232 97928 596238 97980
rect 624602 97928 624608 97980
rect 624660 97968 624666 97980
rect 632974 97968 632980 97980
rect 624660 97940 632980 97968
rect 624660 97928 624666 97940
rect 632974 97928 632980 97940
rect 633032 97928 633038 97980
rect 634170 97928 634176 97980
rect 634228 97968 634234 97980
rect 643370 97968 643376 97980
rect 634228 97940 643376 97968
rect 634228 97928 634234 97940
rect 643370 97928 643376 97940
rect 643428 97928 643434 97980
rect 659746 97968 659752 97980
rect 649966 97940 659752 97968
rect 595254 97832 595260 97844
rect 586486 97804 595260 97832
rect 595254 97792 595260 97804
rect 595312 97832 595318 97844
rect 595622 97832 595628 97844
rect 595312 97804 595628 97832
rect 595312 97792 595318 97804
rect 595622 97792 595628 97804
rect 595680 97792 595686 97844
rect 626074 97792 626080 97844
rect 626132 97832 626138 97844
rect 635274 97832 635280 97844
rect 626132 97804 635280 97832
rect 626132 97792 626138 97804
rect 635274 97792 635280 97804
rect 635332 97792 635338 97844
rect 643554 97832 643560 97844
rect 639156 97804 643560 97832
rect 592678 97656 592684 97708
rect 592736 97696 592742 97708
rect 597554 97696 597560 97708
rect 592736 97668 597560 97696
rect 592736 97656 592742 97668
rect 597554 97656 597560 97668
rect 597612 97656 597618 97708
rect 620186 97656 620192 97708
rect 620244 97696 620250 97708
rect 626074 97696 626080 97708
rect 620244 97668 626080 97696
rect 620244 97656 620250 97668
rect 626074 97656 626080 97668
rect 626132 97656 626138 97708
rect 633342 97656 633348 97708
rect 633400 97696 633406 97708
rect 639156 97696 639184 97804
rect 643554 97792 643560 97804
rect 643612 97792 643618 97844
rect 633400 97668 639184 97696
rect 633400 97656 633406 97668
rect 639322 97656 639328 97708
rect 639380 97696 639386 97708
rect 639380 97668 641760 97696
rect 639380 97656 639386 97668
rect 595438 97520 595444 97572
rect 595496 97560 595502 97572
rect 600406 97560 600412 97572
rect 595496 97532 600412 97560
rect 595496 97520 595502 97532
rect 600406 97520 600412 97532
rect 600464 97520 600470 97572
rect 623130 97520 623136 97572
rect 623188 97560 623194 97572
rect 630674 97560 630680 97572
rect 623188 97532 630680 97560
rect 623188 97520 623194 97532
rect 630674 97520 630680 97532
rect 630732 97520 630738 97572
rect 632698 97520 632704 97572
rect 632756 97560 632762 97572
rect 632756 97532 639644 97560
rect 632756 97520 632762 97532
rect 618714 97384 618720 97436
rect 618772 97424 618778 97436
rect 626258 97424 626264 97436
rect 618772 97396 626264 97424
rect 618772 97384 618778 97396
rect 626258 97384 626264 97396
rect 626316 97384 626322 97436
rect 627546 97384 627552 97436
rect 627604 97424 627610 97436
rect 637574 97424 637580 97436
rect 627604 97396 637580 97424
rect 627604 97384 627610 97396
rect 637574 97384 637580 97396
rect 637632 97384 637638 97436
rect 578878 97248 578884 97300
rect 578936 97288 578942 97300
rect 598934 97288 598940 97300
rect 578936 97260 598940 97288
rect 578936 97248 578942 97260
rect 598934 97248 598940 97260
rect 598992 97248 598998 97300
rect 605466 97248 605472 97300
rect 605524 97288 605530 97300
rect 611906 97288 611912 97300
rect 605524 97260 611912 97288
rect 605524 97248 605530 97260
rect 611906 97248 611912 97260
rect 611964 97248 611970 97300
rect 628190 97248 628196 97300
rect 628248 97288 628254 97300
rect 639046 97288 639052 97300
rect 628248 97260 639052 97288
rect 628248 97248 628254 97260
rect 639046 97248 639052 97260
rect 639104 97248 639110 97300
rect 639616 97288 639644 97532
rect 641732 97424 641760 97668
rect 647142 97656 647148 97708
rect 647200 97696 647206 97708
rect 649966 97696 649994 97940
rect 659746 97928 659752 97940
rect 659804 97928 659810 97980
rect 659930 97928 659936 97980
rect 659988 97968 659994 97980
rect 665174 97968 665180 97980
rect 659988 97940 665180 97968
rect 659988 97928 659994 97940
rect 665174 97928 665180 97940
rect 665232 97928 665238 97980
rect 655422 97792 655428 97844
rect 655480 97832 655486 97844
rect 662506 97832 662512 97844
rect 655480 97804 662512 97832
rect 655480 97792 655486 97804
rect 662506 97792 662512 97804
rect 662564 97792 662570 97844
rect 647200 97668 649994 97696
rect 647200 97656 647206 97668
rect 651834 97656 651840 97708
rect 651892 97696 651898 97708
rect 659562 97696 659568 97708
rect 651892 97668 659568 97696
rect 651892 97656 651898 97668
rect 659562 97656 659568 97668
rect 659620 97656 659626 97708
rect 659746 97656 659752 97708
rect 659804 97696 659810 97708
rect 661954 97696 661960 97708
rect 659804 97668 661960 97696
rect 659804 97656 659810 97668
rect 661954 97656 661960 97668
rect 662012 97656 662018 97708
rect 644290 97520 644296 97572
rect 644348 97560 644354 97572
rect 658826 97560 658832 97572
rect 644348 97532 649304 97560
rect 644348 97520 644354 97532
rect 646498 97424 646504 97436
rect 641732 97396 646504 97424
rect 646498 97384 646504 97396
rect 646556 97384 646562 97436
rect 649276 97424 649304 97532
rect 649966 97532 658832 97560
rect 649966 97424 649994 97532
rect 658826 97520 658832 97532
rect 658884 97520 658890 97572
rect 649276 97396 649994 97424
rect 658182 97384 658188 97436
rect 658240 97424 658246 97436
rect 663058 97424 663064 97436
rect 658240 97396 663064 97424
rect 658240 97384 658246 97396
rect 663058 97384 663064 97396
rect 663116 97384 663122 97436
rect 644750 97288 644756 97300
rect 639616 97260 644756 97288
rect 644750 97248 644756 97260
rect 644808 97248 644814 97300
rect 656802 97248 656808 97300
rect 656860 97288 656866 97300
rect 661402 97288 661408 97300
rect 656860 97260 661408 97288
rect 656860 97248 656866 97260
rect 661402 97248 661408 97260
rect 661460 97248 661466 97300
rect 651098 97180 651104 97232
rect 651156 97220 651162 97232
rect 654318 97220 654324 97232
rect 651156 97192 654324 97220
rect 651156 97180 651162 97192
rect 654318 97180 654324 97192
rect 654376 97180 654382 97232
rect 626810 97112 626816 97164
rect 626868 97152 626874 97164
rect 636378 97152 636384 97164
rect 626868 97124 636384 97152
rect 626868 97112 626874 97124
rect 636378 97112 636384 97124
rect 636436 97112 636442 97164
rect 650362 96976 650368 97028
rect 650420 97016 650426 97028
rect 658274 97016 658280 97028
rect 650420 96988 658280 97016
rect 650420 96976 650426 96988
rect 658274 96976 658280 96988
rect 658332 96976 658338 97028
rect 601050 96908 601056 96960
rect 601108 96948 601114 96960
rect 601878 96948 601884 96960
rect 601108 96920 601884 96948
rect 601108 96908 601114 96920
rect 601878 96908 601884 96920
rect 601936 96908 601942 96960
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 606938 96948 606944 96960
rect 606260 96920 606944 96948
rect 606260 96908 606266 96920
rect 606938 96908 606944 96920
rect 606996 96908 607002 96960
rect 612642 96908 612648 96960
rect 612700 96948 612706 96960
rect 613378 96948 613384 96960
rect 612700 96920 613384 96948
rect 612700 96908 612706 96920
rect 613378 96908 613384 96920
rect 613436 96908 613442 96960
rect 614022 96908 614028 96960
rect 614080 96948 614086 96960
rect 614758 96948 614764 96960
rect 614080 96920 614764 96948
rect 614080 96908 614086 96920
rect 614758 96908 614764 96920
rect 614816 96908 614822 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 645210 96908 645216 96960
rect 645268 96948 645274 96960
rect 645762 96948 645768 96960
rect 645268 96920 645768 96948
rect 645268 96908 645274 96920
rect 645762 96908 645768 96920
rect 645820 96908 645826 96960
rect 660114 96948 660120 96960
rect 659626 96920 660120 96948
rect 609146 96840 609152 96892
rect 609204 96880 609210 96892
rect 609698 96880 609704 96892
rect 609204 96852 609704 96880
rect 609204 96840 609210 96852
rect 609698 96840 609704 96852
rect 609756 96840 609762 96892
rect 646682 96840 646688 96892
rect 646740 96880 646746 96892
rect 647142 96880 647148 96892
rect 646740 96852 647148 96880
rect 646740 96840 646746 96852
rect 647142 96840 647148 96852
rect 647200 96840 647206 96892
rect 654778 96840 654784 96892
rect 654836 96880 654842 96892
rect 655238 96880 655244 96892
rect 654836 96852 655244 96880
rect 654836 96840 654842 96852
rect 655238 96840 655244 96852
rect 655296 96840 655302 96892
rect 656710 96840 656716 96892
rect 656768 96880 656774 96892
rect 659626 96880 659654 96920
rect 660114 96908 660120 96920
rect 660172 96908 660178 96960
rect 656768 96852 659654 96880
rect 656768 96840 656774 96852
rect 613562 96772 613568 96824
rect 613620 96812 613626 96824
rect 614022 96812 614028 96824
rect 613620 96784 614028 96812
rect 613620 96772 613626 96784
rect 614022 96772 614028 96784
rect 614080 96772 614086 96824
rect 641530 96772 641536 96824
rect 641588 96812 641594 96824
rect 642818 96812 642824 96824
rect 641588 96784 642824 96812
rect 641588 96772 641594 96784
rect 642818 96772 642824 96784
rect 642876 96772 642882 96824
rect 612090 96704 612096 96756
rect 612148 96744 612154 96756
rect 612550 96744 612556 96756
rect 612148 96716 612556 96744
rect 612148 96704 612154 96716
rect 612550 96704 612556 96716
rect 612608 96704 612614 96756
rect 617242 96704 617248 96756
rect 617300 96744 617306 96756
rect 618070 96744 618076 96756
rect 617300 96716 618076 96744
rect 617300 96704 617306 96716
rect 618070 96704 618076 96716
rect 618128 96704 618134 96756
rect 643002 96704 643008 96756
rect 643060 96744 643066 96756
rect 660114 96744 660120 96756
rect 643060 96716 660120 96744
rect 643060 96704 643066 96716
rect 660114 96704 660120 96716
rect 660172 96704 660178 96756
rect 642266 96568 642272 96620
rect 642324 96608 642330 96620
rect 644106 96608 644112 96620
rect 642324 96580 644112 96608
rect 642324 96568 642330 96580
rect 644106 96568 644112 96580
rect 644164 96568 644170 96620
rect 651282 96608 651288 96620
rect 644308 96580 651288 96608
rect 638586 96432 638592 96484
rect 638644 96472 638650 96484
rect 644308 96472 644336 96580
rect 651282 96568 651288 96580
rect 651340 96568 651346 96620
rect 652570 96568 652576 96620
rect 652628 96608 652634 96620
rect 654962 96608 654968 96620
rect 652628 96580 654968 96608
rect 652628 96568 652634 96580
rect 654962 96568 654968 96580
rect 655020 96568 655026 96620
rect 638644 96444 644336 96472
rect 638644 96432 638650 96444
rect 653306 96432 653312 96484
rect 653364 96472 653370 96484
rect 663978 96472 663984 96484
rect 653364 96444 663984 96472
rect 653364 96432 653370 96444
rect 663978 96432 663984 96444
rect 664036 96432 664042 96484
rect 631226 96296 631232 96348
rect 631284 96336 631290 96348
rect 642634 96336 642640 96348
rect 631284 96308 642640 96336
rect 631284 96296 631290 96308
rect 642634 96296 642640 96308
rect 642692 96296 642698 96348
rect 642818 96296 642824 96348
rect 642876 96336 642882 96348
rect 648798 96336 648804 96348
rect 642876 96308 648804 96336
rect 642876 96296 642882 96308
rect 648798 96296 648804 96308
rect 648856 96296 648862 96348
rect 648982 96296 648988 96348
rect 649040 96336 649046 96348
rect 649040 96308 654824 96336
rect 649040 96296 649046 96308
rect 620922 96228 620928 96280
rect 620980 96268 620986 96280
rect 626442 96268 626448 96280
rect 620980 96240 626448 96268
rect 620980 96228 620986 96240
rect 626442 96228 626448 96240
rect 626500 96228 626506 96280
rect 631870 96160 631876 96212
rect 631928 96200 631934 96212
rect 644474 96200 644480 96212
rect 631928 96172 644480 96200
rect 631928 96160 631934 96172
rect 644474 96160 644480 96172
rect 644532 96160 644538 96212
rect 652018 96200 652024 96212
rect 648264 96172 652024 96200
rect 610618 96024 610624 96076
rect 610676 96064 610682 96076
rect 621658 96064 621664 96076
rect 610676 96036 621664 96064
rect 610676 96024 610682 96036
rect 621658 96024 621664 96036
rect 621716 96024 621722 96076
rect 635642 96024 635648 96076
rect 635700 96064 635706 96076
rect 635700 96036 639920 96064
rect 635700 96024 635706 96036
rect 608410 95888 608416 95940
rect 608468 95928 608474 95940
rect 620278 95928 620284 95940
rect 608468 95900 620284 95928
rect 608468 95888 608474 95900
rect 620278 95888 620284 95900
rect 620336 95888 620342 95940
rect 637758 95888 637764 95940
rect 637816 95888 637822 95940
rect 634722 95548 634728 95600
rect 634780 95588 634786 95600
rect 634780 95548 634814 95588
rect 634786 95384 634814 95548
rect 637776 95520 637804 95888
rect 639892 95792 639920 96036
rect 640058 96024 640064 96076
rect 640116 96064 640122 96076
rect 648264 96064 648292 96172
rect 652018 96160 652024 96172
rect 652076 96160 652082 96212
rect 654796 96200 654824 96308
rect 654962 96296 654968 96348
rect 655020 96336 655026 96348
rect 665542 96336 665548 96348
rect 655020 96308 665548 96336
rect 655020 96296 655026 96308
rect 665542 96296 665548 96308
rect 665600 96296 665606 96348
rect 663794 96200 663800 96212
rect 654796 96172 663800 96200
rect 663794 96160 663800 96172
rect 663852 96160 663858 96212
rect 640116 96036 648292 96064
rect 640116 96024 640122 96036
rect 649258 96024 649264 96076
rect 649316 96064 649322 96076
rect 660666 96064 660672 96076
rect 649316 96036 660672 96064
rect 649316 96024 649322 96036
rect 660666 96024 660672 96036
rect 660724 96024 660730 96076
rect 640794 95888 640800 95940
rect 640852 95928 640858 95940
rect 665358 95928 665364 95940
rect 640852 95900 665364 95928
rect 640852 95888 640858 95900
rect 665358 95888 665364 95900
rect 665416 95888 665422 95940
rect 642818 95792 642824 95804
rect 639892 95764 642824 95792
rect 642818 95752 642824 95764
rect 642876 95752 642882 95804
rect 645578 95616 645584 95668
rect 645636 95656 645642 95668
rect 656158 95656 656164 95668
rect 645636 95628 656164 95656
rect 645636 95616 645642 95628
rect 656158 95616 656164 95628
rect 656216 95616 656222 95668
rect 659194 95616 659200 95668
rect 659252 95656 659258 95668
rect 664162 95656 664168 95668
rect 659252 95628 664168 95656
rect 659252 95616 659258 95628
rect 664162 95616 664168 95628
rect 664220 95616 664226 95668
rect 649258 95520 649264 95532
rect 637776 95492 649264 95520
rect 649258 95480 649264 95492
rect 649316 95480 649322 95532
rect 643094 95384 643100 95396
rect 634786 95356 643100 95384
rect 643094 95344 643100 95356
rect 643152 95344 643158 95396
rect 616506 95140 616512 95192
rect 616564 95180 616570 95192
rect 623038 95180 623044 95192
rect 616564 95152 623044 95180
rect 616564 95140 616570 95152
rect 623038 95140 623044 95152
rect 623096 95140 623102 95192
rect 649626 95140 649632 95192
rect 649684 95180 649690 95192
rect 650638 95180 650644 95192
rect 649684 95152 650644 95180
rect 649684 95140 649690 95152
rect 650638 95140 650644 95152
rect 650696 95140 650702 95192
rect 643738 94596 643744 94648
rect 643796 94636 643802 94648
rect 653398 94636 653404 94648
rect 643796 94608 653404 94636
rect 643796 94596 643802 94608
rect 653398 94596 653404 94608
rect 653456 94596 653462 94648
rect 607674 94460 607680 94512
rect 607732 94500 607738 94512
rect 624970 94500 624976 94512
rect 607732 94472 624976 94500
rect 607732 94460 607738 94472
rect 624970 94460 624976 94472
rect 625028 94460 625034 94512
rect 642910 94460 642916 94512
rect 642968 94500 642974 94512
rect 663242 94500 663248 94512
rect 642968 94472 663248 94500
rect 642968 94460 642974 94472
rect 663242 94460 663248 94472
rect 663300 94460 663306 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 644106 93780 644112 93832
rect 644164 93820 644170 93832
rect 644164 93792 644474 93820
rect 644164 93780 644170 93792
rect 644446 93752 644474 93792
rect 654134 93752 654140 93764
rect 644446 93724 654140 93752
rect 654134 93712 654140 93724
rect 654192 93712 654198 93764
rect 609698 93100 609704 93152
rect 609756 93140 609762 93152
rect 618898 93140 618904 93152
rect 609756 93112 618904 93140
rect 609756 93100 609762 93112
rect 618898 93100 618904 93112
rect 618956 93100 618962 93152
rect 617886 92420 617892 92472
rect 617944 92460 617950 92472
rect 625430 92460 625436 92472
rect 617944 92432 625436 92460
rect 617944 92420 617950 92432
rect 625430 92420 625436 92432
rect 625488 92420 625494 92472
rect 651282 92420 651288 92472
rect 651340 92460 651346 92472
rect 654318 92460 654324 92472
rect 651340 92432 654324 92460
rect 651340 92420 651346 92432
rect 654318 92420 654324 92432
rect 654376 92420 654382 92472
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 617334 91032 617340 91044
rect 611320 91004 617340 91032
rect 611320 90992 611326 91004
rect 617334 90992 617340 91004
rect 617392 90992 617398 91044
rect 618070 90992 618076 91044
rect 618128 91032 618134 91044
rect 626442 91032 626448 91044
rect 618128 91004 626448 91032
rect 618128 90992 618134 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 646498 90992 646504 91044
rect 646556 91032 646562 91044
rect 654134 91032 654140 91044
rect 646556 91004 654140 91032
rect 646556 90992 646562 91004
rect 654134 90992 654140 91004
rect 654192 90992 654198 91044
rect 623038 89632 623044 89684
rect 623096 89672 623102 89684
rect 626442 89672 626448 89684
rect 623096 89644 626448 89672
rect 623096 89632 623102 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 647142 88952 647148 89004
rect 647200 88992 647206 89004
rect 656894 88992 656900 89004
rect 647200 88964 656900 88992
rect 647200 88952 647206 88964
rect 656894 88952 656900 88964
rect 656952 88952 656958 89004
rect 656158 88748 656164 88800
rect 656216 88788 656222 88800
rect 657446 88788 657452 88800
rect 656216 88760 657452 88788
rect 656216 88748 656222 88760
rect 657446 88748 657452 88760
rect 657504 88748 657510 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 664162 88788 664168 88800
rect 662380 88760 664168 88788
rect 662380 88748 662386 88760
rect 664162 88748 664168 88760
rect 664220 88748 664226 88800
rect 656710 88612 656716 88664
rect 656768 88652 656774 88664
rect 659286 88652 659292 88664
rect 656768 88624 659292 88652
rect 656768 88612 656774 88624
rect 659286 88612 659292 88624
rect 659344 88612 659350 88664
rect 607306 88272 607312 88324
rect 607364 88312 607370 88324
rect 626442 88312 626448 88324
rect 607364 88284 626448 88312
rect 607364 88272 607370 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 617334 88136 617340 88188
rect 617392 88176 617398 88188
rect 625614 88176 625620 88188
rect 617392 88148 625620 88176
rect 617392 88136 617398 88148
rect 625614 88136 625620 88148
rect 625672 88136 625678 88188
rect 648154 87116 648160 87168
rect 648212 87156 648218 87168
rect 662506 87156 662512 87168
rect 648212 87128 662512 87156
rect 648212 87116 648218 87128
rect 662506 87116 662512 87128
rect 662564 87116 662570 87168
rect 645762 86980 645768 87032
rect 645820 87020 645826 87032
rect 660666 87020 660672 87032
rect 645820 86992 660672 87020
rect 645820 86980 645826 86992
rect 660666 86980 660672 86992
rect 660724 86980 660730 87032
rect 652018 86708 652024 86760
rect 652076 86748 652082 86760
rect 660114 86748 660120 86760
rect 652076 86720 660120 86748
rect 652076 86708 652082 86720
rect 660114 86708 660120 86720
rect 660172 86708 660178 86760
rect 653398 86572 653404 86624
rect 653456 86612 653462 86624
rect 661402 86612 661408 86624
rect 653456 86584 661408 86612
rect 653456 86572 653462 86584
rect 661402 86572 661408 86584
rect 661460 86572 661466 86624
rect 650638 86436 650644 86488
rect 650696 86476 650702 86488
rect 658826 86476 658832 86488
rect 650696 86448 658832 86476
rect 650696 86436 650702 86448
rect 658826 86436 658832 86448
rect 658884 86436 658890 86488
rect 621658 86232 621664 86284
rect 621716 86272 621722 86284
rect 626442 86272 626448 86284
rect 621716 86244 626448 86272
rect 621716 86232 621722 86244
rect 626442 86232 626448 86244
rect 626500 86232 626506 86284
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 620278 84124 620284 84176
rect 620336 84164 620342 84176
rect 626258 84164 626264 84176
rect 620336 84136 626264 84164
rect 620336 84124 620342 84136
rect 626258 84124 626264 84136
rect 626316 84124 626322 84176
rect 618898 83988 618904 84040
rect 618956 84028 618962 84040
rect 618956 84000 625154 84028
rect 618956 83988 618962 84000
rect 625126 83960 625154 84000
rect 626442 83960 626448 83972
rect 625126 83932 626448 83960
rect 626442 83920 626448 83932
rect 626500 83920 626506 83972
rect 628558 80928 628564 80980
rect 628616 80968 628622 80980
rect 642450 80968 642456 80980
rect 628616 80940 642456 80968
rect 628616 80928 628622 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 612550 80792 612556 80844
rect 612608 80832 612614 80844
rect 645854 80832 645860 80844
rect 612608 80804 645860 80832
rect 612608 80792 612614 80804
rect 645854 80792 645860 80804
rect 645912 80792 645918 80844
rect 595622 80656 595628 80708
rect 595680 80696 595686 80708
rect 636102 80696 636108 80708
rect 595680 80668 636108 80696
rect 595680 80656 595686 80668
rect 636102 80656 636108 80668
rect 636160 80656 636166 80708
rect 629202 79432 629208 79484
rect 629260 79472 629266 79484
rect 637482 79472 637488 79484
rect 629260 79444 637488 79472
rect 629260 79432 629266 79444
rect 637482 79432 637488 79444
rect 637540 79432 637546 79484
rect 616782 79296 616788 79348
rect 616840 79336 616846 79348
rect 647418 79336 647424 79348
rect 616840 79308 647424 79336
rect 616840 79296 616846 79308
rect 647418 79296 647424 79308
rect 647476 79296 647482 79348
rect 637482 78208 637488 78260
rect 637540 78248 637546 78260
rect 645302 78248 645308 78260
rect 637540 78220 645308 78248
rect 637540 78208 637546 78220
rect 645302 78208 645308 78220
rect 645360 78208 645366 78260
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 638954 78112 638960 78124
rect 631100 78084 638960 78112
rect 631100 78072 631106 78084
rect 638954 78072 638960 78084
rect 639012 78072 639018 78124
rect 614022 77936 614028 77988
rect 614080 77976 614086 77988
rect 647602 77976 647608 77988
rect 614080 77948 647608 77976
rect 614080 77936 614086 77948
rect 647602 77936 647608 77948
rect 647660 77936 647666 77988
rect 631042 77704 631048 77716
rect 625126 77676 631048 77704
rect 591298 77392 591304 77444
rect 591356 77432 591362 77444
rect 625126 77432 625154 77676
rect 631042 77664 631048 77676
rect 631100 77664 631106 77716
rect 628282 77528 628288 77580
rect 628340 77568 628346 77580
rect 631502 77568 631508 77580
rect 628340 77540 631508 77568
rect 628340 77528 628346 77540
rect 631502 77528 631508 77540
rect 631560 77528 631566 77580
rect 591356 77404 625154 77432
rect 591356 77392 591362 77404
rect 625798 77392 625804 77444
rect 625856 77432 625862 77444
rect 633894 77432 633900 77444
rect 625856 77404 633900 77432
rect 625856 77392 625862 77404
rect 633894 77392 633900 77404
rect 633952 77392 633958 77444
rect 577498 77256 577504 77308
rect 577556 77296 577562 77308
rect 637114 77296 637120 77308
rect 577556 77268 637120 77296
rect 577556 77256 577562 77268
rect 637114 77256 637120 77268
rect 637172 77296 637178 77308
rect 639598 77296 639604 77308
rect 637172 77268 639604 77296
rect 637172 77256 637178 77268
rect 639598 77256 639604 77268
rect 639656 77256 639662 77308
rect 614758 76644 614764 76696
rect 614816 76684 614822 76696
rect 646314 76684 646320 76696
rect 614816 76656 646320 76684
rect 614816 76644 614822 76656
rect 646314 76644 646320 76656
rect 646372 76644 646378 76696
rect 613378 76508 613384 76560
rect 613436 76548 613442 76560
rect 649166 76548 649172 76560
rect 613436 76520 649172 76548
rect 613436 76508 613442 76520
rect 649166 76508 649172 76520
rect 649224 76508 649230 76560
rect 580258 75896 580264 75948
rect 580316 75936 580322 75948
rect 628282 75936 628288 75948
rect 580316 75908 628288 75936
rect 580316 75896 580322 75908
rect 628282 75896 628288 75908
rect 628340 75896 628346 75948
rect 615402 75284 615408 75336
rect 615460 75324 615466 75336
rect 646130 75324 646136 75336
rect 615460 75296 646136 75324
rect 615460 75284 615466 75296
rect 646130 75284 646136 75296
rect 646188 75284 646194 75336
rect 607122 75148 607128 75200
rect 607180 75188 607186 75200
rect 646866 75188 646872 75200
rect 607180 75160 646872 75188
rect 607180 75148 607186 75160
rect 646866 75148 646872 75160
rect 646924 75148 646930 75200
rect 611998 57196 612004 57248
rect 612056 57236 612062 57248
rect 662414 57236 662420 57248
rect 612056 57208 662420 57236
rect 612056 57196 612062 57208
rect 662414 57196 662420 57208
rect 662472 57196 662478 57248
rect 580258 53088 580264 53100
rect 151786 53060 580264 53088
rect 145374 52912 145380 52964
rect 145432 52952 145438 52964
rect 151786 52952 151814 53060
rect 580258 53048 580264 53060
rect 580316 53048 580322 53100
rect 145432 52924 151814 52952
rect 145432 52912 145438 52924
rect 288158 52368 288164 52420
rect 288216 52408 288222 52420
rect 625798 52408 625804 52420
rect 288216 52380 625804 52408
rect 288216 52368 288222 52380
rect 625798 52368 625804 52380
rect 625856 52368 625862 52420
rect 391934 52232 391940 52284
rect 391992 52272 391998 52284
rect 392578 52272 392584 52284
rect 391992 52244 392584 52272
rect 391992 52232 391998 52244
rect 392578 52232 392584 52244
rect 392636 52272 392642 52284
rect 577498 52272 577504 52284
rect 392636 52244 577504 52272
rect 392636 52232 392642 52244
rect 577498 52232 577504 52244
rect 577556 52232 577562 52284
rect 235810 51008 235816 51060
rect 235868 51048 235874 51060
rect 288158 51048 288164 51060
rect 235868 51020 288164 51048
rect 235868 51008 235874 51020
rect 288158 51008 288164 51020
rect 288216 51008 288222 51060
rect 340506 51008 340512 51060
rect 340564 51048 340570 51060
rect 391934 51048 391940 51060
rect 340564 51020 391940 51048
rect 340564 51008 340570 51020
rect 391934 51008 391940 51020
rect 391992 51008 391998 51060
rect 405090 50464 405096 50516
rect 405148 50504 405154 50516
rect 578878 50504 578884 50516
rect 405148 50476 578884 50504
rect 405148 50464 405154 50476
rect 578878 50464 578884 50476
rect 578936 50464 578942 50516
rect 183462 50328 183468 50380
rect 183520 50368 183526 50380
rect 406378 50368 406384 50380
rect 183520 50340 406384 50368
rect 183520 50328 183526 50340
rect 406378 50328 406384 50340
rect 406436 50328 406442 50380
rect 461026 47200 461032 47252
rect 461084 47240 461090 47252
rect 465902 47240 465908 47252
rect 461084 47212 465908 47240
rect 461084 47200 461090 47212
rect 465902 47200 465908 47212
rect 465960 47200 465966 47252
rect 194042 44820 194048 44872
rect 194100 44860 194106 44872
rect 661586 44860 661592 44872
rect 194100 44832 661592 44860
rect 194100 44820 194106 44832
rect 661586 44820 661592 44832
rect 661644 44820 661650 44872
rect 315942 43392 315948 43444
rect 316000 43432 316006 43444
rect 661126 43432 661132 43444
rect 316000 43404 661132 43432
rect 316000 43392 316006 43404
rect 661126 43392 661132 43404
rect 661184 43392 661190 43444
rect 464890 42328 464896 42380
rect 464948 42328 464954 42380
rect 315942 42173 315948 42225
rect 316000 42173 316006 42225
<< via1 >>
rect 366180 1027828 366232 1027880
rect 366548 1027828 366600 1027880
rect 366180 1024360 366232 1024412
rect 366548 1024360 366600 1024412
rect 505008 1007156 505060 1007208
rect 513840 1007156 513892 1007208
rect 357716 1007088 357768 1007140
rect 368940 1007088 368992 1007140
rect 505376 1007020 505428 1007072
rect 515588 1007020 515640 1007072
rect 357716 1006884 357768 1006936
rect 373264 1006952 373316 1007004
rect 425520 1006952 425572 1007004
rect 439688 1006952 439740 1007004
rect 503352 1006884 503404 1006936
rect 520924 1006952 520976 1007004
rect 551100 1006952 551152 1007004
rect 569224 1006952 569276 1007004
rect 427544 1006816 427596 1006868
rect 438124 1006816 438176 1006868
rect 554136 1006816 554188 1006868
rect 559656 1006816 559708 1006868
rect 358544 1006748 358596 1006800
rect 369124 1006748 369176 1006800
rect 400864 1006680 400916 1006732
rect 430856 1006680 430908 1006732
rect 555976 1006680 556028 1006732
rect 566464 1006680 566516 1006732
rect 506204 1006612 506256 1006664
rect 514024 1006612 514076 1006664
rect 94688 1006544 94740 1006596
rect 103152 1006544 103204 1006596
rect 145564 1006544 145616 1006596
rect 153752 1006544 153804 1006596
rect 298836 1006544 298888 1006596
rect 306932 1006544 306984 1006596
rect 429200 1006544 429252 1006596
rect 471244 1006544 471296 1006596
rect 505376 1006476 505428 1006528
rect 516784 1006476 516836 1006528
rect 102784 1006408 102836 1006460
rect 103980 1006408 104032 1006460
rect 145748 1006408 145800 1006460
rect 152924 1006408 152976 1006460
rect 300308 1006408 300360 1006460
rect 307760 1006408 307812 1006460
rect 360200 1006408 360252 1006460
rect 376024 1006408 376076 1006460
rect 553124 1006408 553176 1006460
rect 210424 1006340 210476 1006392
rect 228364 1006340 228416 1006392
rect 93124 1006272 93176 1006324
rect 100300 1006272 100352 1006324
rect 144276 1006272 144328 1006324
rect 152096 1006272 152148 1006324
rect 158260 1006272 158312 1006324
rect 175924 1006272 175976 1006324
rect 249064 1006272 249116 1006324
rect 256148 1006272 256200 1006324
rect 299296 1006272 299348 1006324
rect 311808 1006272 311860 1006324
rect 314660 1006272 314712 1006324
rect 319444 1006272 319496 1006324
rect 360568 1006272 360620 1006324
rect 208400 1006204 208452 1006256
rect 94504 1006136 94556 1006188
rect 101956 1006136 102008 1006188
rect 106832 1006136 106884 1006188
rect 124864 1006136 124916 1006188
rect 144460 1006136 144512 1006188
rect 159456 1006136 159508 1006188
rect 160284 1006136 160336 1006188
rect 164884 1006136 164936 1006188
rect 247040 1006136 247092 1006188
rect 252468 1006136 252520 1006188
rect 262680 1006136 262732 1006188
rect 278044 1006136 278096 1006188
rect 300124 1006136 300176 1006188
rect 306104 1006136 306156 1006188
rect 93308 1006000 93360 1006052
rect 98276 1006000 98328 1006052
rect 101404 1006000 101456 1006052
rect 103980 1006000 104032 1006052
rect 107660 1006000 107712 1006052
rect 126244 1006000 126296 1006052
rect 148876 1006000 148928 1006052
rect 150072 1006000 150124 1006052
rect 152648 1006000 152700 1006052
rect 155776 1006000 155828 1006052
rect 158628 1006000 158680 1006052
rect 177304 1006000 177356 1006052
rect 198648 1006000 198700 1006052
rect 201040 1006000 201092 1006052
rect 229744 1006000 229796 1006052
rect 249800 1006000 249852 1006052
rect 254124 1006000 254176 1006052
rect 261852 1006000 261904 1006052
rect 280804 1006000 280856 1006052
rect 302148 1006000 302200 1006052
rect 304080 1006000 304132 1006052
rect 314660 1006000 314712 1006052
rect 323584 1006000 323636 1006052
rect 354588 1006000 354640 1006052
rect 354864 1006000 354916 1006052
rect 355692 1006000 355744 1006052
rect 359556 1006000 359608 1006052
rect 361396 1006000 361448 1006052
rect 365260 1006136 365312 1006188
rect 369124 1006272 369176 1006324
rect 374644 1006272 374696 1006324
rect 425152 1006272 425204 1006324
rect 443644 1006272 443696 1006324
rect 502156 1006272 502208 1006324
rect 518164 1006272 518216 1006324
rect 556804 1006272 556856 1006324
rect 560208 1006272 560260 1006324
rect 571984 1006272 572036 1006324
rect 371884 1006136 371936 1006188
rect 422024 1006136 422076 1006188
rect 423496 1006136 423548 1006188
rect 508228 1006136 508280 1006188
rect 522304 1006136 522356 1006188
rect 557172 1006136 557224 1006188
rect 365076 1006000 365128 1006052
rect 367744 1006000 367796 1006052
rect 368940 1006000 368992 1006052
rect 378140 1006000 378192 1006052
rect 422668 1006000 422720 1006052
rect 429844 1006000 429896 1006052
rect 430028 1006000 430080 1006052
rect 471428 1006000 471480 1006052
rect 497924 1006000 497976 1006052
rect 498844 1006000 498896 1006052
rect 501328 1006000 501380 1006052
rect 506480 1006000 506532 1006052
rect 509056 1006000 509108 1006052
rect 514024 1006000 514076 1006052
rect 522488 1006000 522540 1006052
rect 574744 1006000 574796 1006052
rect 515404 1005864 515456 1005916
rect 432052 1005796 432104 1005848
rect 433524 1005796 433576 1005848
rect 423496 1005660 423548 1005712
rect 446404 1005660 446456 1005712
rect 560852 1005660 560904 1005712
rect 570604 1005660 570656 1005712
rect 428372 1005524 428424 1005576
rect 460204 1005524 460256 1005576
rect 555148 1005524 555200 1005576
rect 567844 1005524 567896 1005576
rect 436928 1005388 436980 1005440
rect 465724 1005388 465776 1005440
rect 553952 1005388 554004 1005440
rect 573364 1005388 573416 1005440
rect 149888 1005320 149940 1005372
rect 152924 1005320 152976 1005372
rect 427176 1005320 427228 1005372
rect 195704 1005252 195756 1005304
rect 202696 1005252 202748 1005304
rect 263048 1005252 263100 1005304
rect 279424 1005252 279476 1005304
rect 360568 1005252 360620 1005304
rect 377404 1005252 377456 1005304
rect 456064 1005252 456116 1005304
rect 552296 1005252 552348 1005304
rect 570788 1005252 570840 1005304
rect 430856 1005184 430908 1005236
rect 431914 1005184 431966 1005236
rect 507032 1005184 507084 1005236
rect 509976 1005184 510028 1005236
rect 432052 1005116 432104 1005168
rect 436928 1005116 436980 1005168
rect 209228 1005048 209280 1005100
rect 211804 1005048 211856 1005100
rect 363420 1005048 363472 1005100
rect 366364 1005048 366416 1005100
rect 508228 1005048 508280 1005100
rect 510896 1005048 510948 1005100
rect 432420 1004980 432472 1005032
rect 434168 1004980 434220 1005032
rect 151084 1004912 151136 1004964
rect 153752 1004912 153804 1004964
rect 154396 1004912 154448 1004964
rect 160652 1004912 160704 1004964
rect 207572 1004912 207624 1004964
rect 209872 1004912 209924 1004964
rect 365076 1004912 365128 1004964
rect 370504 1004912 370556 1004964
rect 429200 1004912 429252 1004964
rect 432236 1004912 432288 1004964
rect 507860 1004912 507912 1004964
rect 509700 1004912 509752 1004964
rect 151268 1004776 151320 1004828
rect 154120 1004776 154172 1004828
rect 159456 1004776 159508 1004828
rect 162124 1004776 162176 1004828
rect 313832 1004776 313884 1004828
rect 316040 1004776 316092 1004828
rect 352840 1004776 352892 1004828
rect 355692 1004776 355744 1004828
rect 362592 1004776 362644 1004828
rect 364984 1004776 365036 1004828
rect 431684 1004776 431736 1004828
rect 106188 1004640 106240 1004692
rect 108488 1004640 108540 1004692
rect 149704 1004640 149756 1004692
rect 151728 1004640 151780 1004692
rect 160652 1004640 160704 1004692
rect 162860 1004640 162912 1004692
rect 209228 1004640 209280 1004692
rect 211160 1004640 211212 1004692
rect 212540 1004640 212592 1004692
rect 217324 1004640 217376 1004692
rect 250444 1004640 250496 1004692
rect 256516 1004640 256568 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 364248 1004640 364300 1004692
rect 366548 1004640 366600 1004692
rect 430028 1004640 430080 1004692
rect 431868 1004640 431920 1004692
rect 498108 1004776 498160 1004828
rect 499672 1004776 499724 1004828
rect 507400 1004776 507452 1004828
rect 509240 1004776 509292 1004828
rect 555976 1004776 556028 1004828
rect 558184 1004776 558236 1004828
rect 433984 1004640 434036 1004692
rect 499488 1004640 499540 1004692
rect 500500 1004640 500552 1004692
rect 509056 1004640 509108 1004692
rect 510712 1004640 510764 1004692
rect 557632 1004640 557684 1004692
rect 559564 1004640 559616 1004692
rect 504548 1004436 504600 1004488
rect 510160 1004436 510212 1004488
rect 356520 1003892 356572 1003944
rect 381452 1003892 381504 1003944
rect 422024 1003892 422076 1003944
rect 469864 1003892 469916 1003944
rect 298652 1003280 298704 1003332
rect 331128 1003280 331180 1003332
rect 354588 1002804 354640 1002856
rect 355140 1002804 355192 1002856
rect 456064 1002804 456116 1002856
rect 462320 1002804 462372 1002856
rect 98644 1002736 98696 1002788
rect 101956 1002736 102008 1002788
rect 252008 1002736 252060 1002788
rect 255320 1002736 255372 1002788
rect 424692 1002668 424744 1002720
rect 449164 1002668 449216 1002720
rect 97264 1002600 97316 1002652
rect 100300 1002600 100352 1002652
rect 157432 1002600 157484 1002652
rect 159364 1002600 159416 1002652
rect 560208 1002600 560260 1002652
rect 567200 1002600 567252 1002652
rect 246764 1002532 246816 1002584
rect 255320 1002532 255372 1002584
rect 426348 1002532 426400 1002584
rect 458088 1002532 458140 1002584
rect 98828 1002464 98880 1002516
rect 101128 1002464 101180 1002516
rect 106004 1002464 106056 1002516
rect 109500 1002464 109552 1002516
rect 158628 1002464 158680 1002516
rect 160192 1002464 160244 1002516
rect 261024 1002464 261076 1002516
rect 264244 1002464 264296 1002516
rect 501696 1002464 501748 1002516
rect 504364 1002464 504416 1002516
rect 558828 1002464 558880 1002516
rect 562324 1002464 562376 1002516
rect 96528 1002328 96580 1002380
rect 99104 1002328 99156 1002380
rect 105636 1002328 105688 1002380
rect 107752 1002328 107804 1002380
rect 108028 1002328 108080 1002380
rect 110420 1002328 110472 1002380
rect 144736 1002328 144788 1002380
rect 150900 1002328 150952 1002380
rect 156604 1002328 156656 1002380
rect 158720 1002328 158772 1002380
rect 211252 1002328 211304 1002380
rect 215944 1002328 215996 1002380
rect 500224 1002328 500276 1002380
rect 502156 1002328 502208 1002380
rect 558000 1002328 558052 1002380
rect 560300 1002328 560352 1002380
rect 560484 1002328 560536 1002380
rect 563060 1002328 563112 1002380
rect 99012 1002192 99064 1002244
rect 101128 1002192 101180 1002244
rect 104808 1002192 104860 1002244
rect 106464 1002192 106516 1002244
rect 108488 1002192 108540 1002244
rect 111064 1002192 111116 1002244
rect 148324 1002192 148376 1002244
rect 151728 1002192 151780 1002244
rect 155776 1002192 155828 1002244
rect 157340 1002192 157392 1002244
rect 203340 1002192 203392 1002244
rect 206376 1002192 206428 1002244
rect 210056 1002192 210108 1002244
rect 212540 1002192 212592 1002244
rect 251824 1002192 251876 1002244
rect 254492 1002192 254544 1002244
rect 428004 1002192 428056 1002244
rect 431132 1002192 431184 1002244
rect 500500 1002192 500552 1002244
rect 502984 1002192 503036 1002244
rect 509884 1002192 509936 1002244
rect 512644 1002192 512696 1002244
rect 553124 1002192 553176 1002244
rect 554320 1002192 554372 1002244
rect 560024 1002192 560076 1002244
rect 562508 1002192 562560 1002244
rect 97448 1002056 97500 1002108
rect 99472 1002056 99524 1002108
rect 100024 1002056 100076 1002108
rect 103152 1002056 103204 1002108
rect 106832 1002056 106884 1002108
rect 109040 1002056 109092 1002108
rect 109684 1002056 109736 1002108
rect 111892 1002056 111944 1002108
rect 148968 1002056 149020 1002108
rect 150900 1002056 150952 1002108
rect 155224 1002056 155276 1002108
rect 156604 1002056 156656 1002108
rect 203708 1002056 203760 1002108
rect 205548 1002056 205600 1002108
rect 211252 1002056 211304 1002108
rect 213184 1002056 213236 1002108
rect 253480 1002056 253532 1002108
rect 256148 1002056 256200 1002108
rect 263508 1002056 263560 1002108
rect 265624 1002056 265676 1002108
rect 310980 1002056 311032 1002108
rect 313280 1002056 313332 1002108
rect 355784 1002056 355836 1002108
rect 358544 1002056 358596 1002108
rect 359740 1002056 359792 1002108
rect 362224 1002056 362276 1002108
rect 423588 1002056 423640 1002108
rect 425152 1002056 425204 1002108
rect 428372 1002056 428424 1002108
rect 431316 1002056 431368 1002108
rect 433340 1002056 433392 1002108
rect 435364 1002056 435416 1002108
rect 500684 1002056 500736 1002108
rect 502524 1002056 502576 1002108
rect 510344 1002056 510396 1002108
rect 512828 1002056 512880 1002108
rect 555148 1002056 555200 1002108
rect 556804 1002056 556856 1002108
rect 558000 1002056 558052 1002108
rect 560668 1002056 560720 1002108
rect 560852 1002056 560904 1002108
rect 563704 1002056 563756 1002108
rect 152464 1001988 152516 1002040
rect 154580 1001988 154632 1002040
rect 96344 1001920 96396 1001972
rect 98276 1001920 98328 1001972
rect 100208 1001920 100260 1001972
rect 102324 1001920 102376 1001972
rect 106004 1001920 106056 1001972
rect 108120 1001920 108172 1001972
rect 108856 1001920 108908 1001972
rect 112076 1001920 112128 1001972
rect 147588 1001920 147640 1001972
rect 149244 1001920 149296 1001972
rect 154948 1001920 155000 1001972
rect 155960 1001920 156012 1001972
rect 157800 1001920 157852 1001972
rect 160376 1001920 160428 1001972
rect 195152 1001920 195204 1001972
rect 198648 1001920 198700 1001972
rect 204904 1001920 204956 1001972
rect 206744 1001920 206796 1001972
rect 212080 1001920 212132 1001972
rect 213920 1001920 213972 1001972
rect 261024 1001920 261076 1001972
rect 263600 1001920 263652 1001972
rect 263876 1001920 263928 1001972
rect 267004 1001920 267056 1001972
rect 310152 1001920 310204 1001972
rect 311900 1001920 311952 1001972
rect 312636 1001920 312688 1001972
rect 314660 1001920 314712 1001972
rect 351828 1001920 351880 1001972
rect 354036 1001920 354088 1001972
rect 356060 1001920 356112 1001972
rect 356520 1001920 356572 1001972
rect 357348 1001920 357400 1001972
rect 360844 1001920 360896 1001972
rect 361396 1001920 361448 1001972
rect 363604 1001920 363656 1001972
rect 365904 1001920 365956 1001972
rect 369124 1001920 369176 1001972
rect 419448 1001920 419500 1001972
rect 421472 1001920 421524 1001972
rect 424324 1001920 424376 1001972
rect 425060 1001920 425112 1001972
rect 426348 1001920 426400 1001972
rect 428464 1001920 428516 1001972
rect 432880 1001920 432932 1001972
rect 436744 1001920 436796 1001972
rect 496728 1001920 496780 1001972
rect 498476 1001920 498528 1001972
rect 502248 1001920 502300 1001972
rect 503352 1001920 503404 1001972
rect 504180 1001920 504232 1001972
rect 505744 1001920 505796 1001972
rect 506204 1001920 506256 1001972
rect 507860 1001920 507912 1001972
rect 554320 1001920 554372 1001972
rect 555424 1001920 555476 1001972
rect 558828 1001920 558880 1001972
rect 560208 1001920 560260 1001972
rect 561680 1001920 561732 1001972
rect 565084 1001920 565136 1001972
rect 512828 1001376 512880 1001428
rect 519544 1001376 519596 1001428
rect 246580 1001172 246632 1001224
rect 256976 1001172 257028 1001224
rect 355784 1001172 355836 1001224
rect 378784 1001172 378836 1001224
rect 510160 1000900 510212 1000952
rect 517244 1000900 517296 1000952
rect 92664 999744 92716 999796
rect 99012 999744 99064 999796
rect 195520 999744 195572 999796
rect 209872 999744 209924 999796
rect 591304 999268 591356 999320
rect 616788 999268 616840 999320
rect 298928 999132 298980 999184
rect 305276 999132 305328 999184
rect 378140 999132 378192 999184
rect 383292 999132 383344 999184
rect 458088 999132 458140 999184
rect 373264 999064 373316 999116
rect 375564 999064 375616 999116
rect 446404 999064 446456 999116
rect 452292 999064 452344 999116
rect 591120 999132 591172 999184
rect 625620 999132 625672 999184
rect 516784 999064 516836 999116
rect 523316 999064 523368 999116
rect 472624 998928 472676 998980
rect 513840 998928 513892 998980
rect 523684 998928 523736 998980
rect 428464 998792 428516 998844
rect 466460 998792 466512 998844
rect 504364 998792 504416 998844
rect 516692 998792 516744 998844
rect 196624 998656 196676 998708
rect 204352 998656 204404 998708
rect 199384 998520 199436 998572
rect 203524 998520 203576 998572
rect 303252 998520 303304 998572
rect 308956 998520 309008 998572
rect 355140 998520 355192 998572
rect 378600 998724 378652 998776
rect 431316 998656 431368 998708
rect 472440 998656 472492 998708
rect 499488 998656 499540 998708
rect 510068 998656 510120 998708
rect 377404 998588 377456 998640
rect 383568 998588 383620 998640
rect 425060 998520 425112 998572
rect 472072 998520 472124 998572
rect 506480 998520 506532 998572
rect 524052 998520 524104 998572
rect 200856 998384 200908 998436
rect 203892 998384 203944 998436
rect 247868 998384 247920 998436
rect 259000 998384 259052 998436
rect 304448 998384 304500 998436
rect 307300 998384 307352 998436
rect 356060 998384 356112 998436
rect 383476 998384 383528 998436
rect 423588 998384 423640 998436
rect 472256 998384 472308 998436
rect 500224 998384 500276 998436
rect 523132 998384 523184 998436
rect 616788 998384 616840 998436
rect 625436 998384 625488 998436
rect 196808 998248 196860 998300
rect 202696 998248 202748 998300
rect 302884 998248 302936 998300
rect 306104 998248 306156 998300
rect 443644 998248 443696 998300
rect 446864 998248 446916 998300
rect 510068 998248 510120 998300
rect 520556 998248 520608 998300
rect 254584 998180 254636 998232
rect 257344 998180 257396 998232
rect 198648 998112 198700 998164
rect 200672 998112 200724 998164
rect 202144 998112 202196 998164
rect 204076 998112 204128 998164
rect 247684 998112 247736 998164
rect 253664 998112 253716 998164
rect 305644 998112 305696 998164
rect 308128 998112 308180 998164
rect 143724 998044 143776 998096
rect 146944 998044 146996 998096
rect 255964 998044 256016 998096
rect 258172 998044 258224 998096
rect 260196 998044 260248 998096
rect 262864 998044 262916 998096
rect 92296 997976 92348 998028
rect 94688 997976 94740 998028
rect 200028 997976 200080 998028
rect 201868 997976 201920 998028
rect 250996 997976 251048 998028
rect 253296 997976 253348 998028
rect 304264 997976 304316 998028
rect 306932 997976 306984 998028
rect 308404 997976 308456 998028
rect 310612 997976 310664 998028
rect 549168 997976 549220 998028
rect 551100 997976 551152 998028
rect 202328 997908 202380 997960
rect 204720 997908 204772 997960
rect 257344 997908 257396 997960
rect 259000 997908 259052 997960
rect 259828 997908 259880 997960
rect 262220 997908 262272 997960
rect 143908 997840 143960 997892
rect 151268 997840 151320 997892
rect 249708 997840 249760 997892
rect 252468 997840 252520 997892
rect 303528 997840 303580 997892
rect 304908 997840 304960 997892
rect 307024 997840 307076 997892
rect 308956 997840 309008 997892
rect 547788 997840 547840 997892
rect 550272 997840 550324 997892
rect 550548 997840 550600 997892
rect 553308 997840 553360 997892
rect 200948 997772 201000 997824
rect 203524 997772 203576 997824
rect 258172 997772 258224 997824
rect 259460 997772 259512 997824
rect 260196 997772 260248 997824
rect 260932 997772 260984 997824
rect 378784 997772 378836 997824
rect 383108 997772 383160 997824
rect 488908 997772 488960 997824
rect 493508 997772 493560 997824
rect 520924 997772 520976 997824
rect 523868 997772 523920 997824
rect 592040 997772 592092 997824
rect 625804 997772 625856 997824
rect 144828 997704 144880 997756
rect 152648 997704 152700 997756
rect 247224 997704 247276 997756
rect 254584 997704 254636 997756
rect 299112 997704 299164 997756
rect 310428 997704 310480 997756
rect 363604 997704 363656 997756
rect 372344 997704 372396 997756
rect 431132 997704 431184 997756
rect 439688 997704 439740 997756
rect 515588 997704 515640 997756
rect 516876 997704 516928 997756
rect 164884 997636 164936 997688
rect 170312 997636 170364 997688
rect 566464 997636 566516 997688
rect 623688 997636 623740 997688
rect 438124 997568 438176 997620
rect 439872 997568 439924 997620
rect 573364 997500 573416 997552
rect 553124 997364 553176 997416
rect 581276 997364 581328 997416
rect 581828 997500 581880 997552
rect 591304 997500 591356 997552
rect 590384 997364 590436 997416
rect 319444 997296 319496 997348
rect 332600 997296 332652 997348
rect 97080 997228 97132 997280
rect 98828 997228 98880 997280
rect 331128 997160 331180 997212
rect 357348 997160 357400 997212
rect 569224 997160 569276 997212
rect 620284 997160 620336 997212
rect 318064 997024 318116 997076
rect 349160 997024 349212 997076
rect 360844 997024 360896 997076
rect 380900 997024 380952 997076
rect 558184 997024 558236 997076
rect 617340 997024 617392 997076
rect 106924 996888 106976 996940
rect 111892 996888 111944 996940
rect 570788 996888 570840 996940
rect 581460 996888 581512 996940
rect 574744 996752 574796 996804
rect 592040 996888 592092 996940
rect 581276 996616 581328 996668
rect 590568 996616 590620 996668
rect 200212 996412 200264 996464
rect 203708 996412 203760 996464
rect 421012 996412 421064 996464
rect 426440 996412 426492 996464
rect 92480 996344 92532 996396
rect 121736 996344 121788 996396
rect 555424 996276 555476 996328
rect 591120 996276 591172 996328
rect 551928 996208 551980 996260
rect 554320 996208 554372 996260
rect 109500 996072 109552 996124
rect 158720 996072 158772 996124
rect 159364 996072 159416 996124
rect 208400 996072 208452 996124
rect 229744 996072 229796 996124
rect 262220 996072 262272 996124
rect 278044 996072 278096 996124
rect 316040 996072 316092 996124
rect 366548 996072 366600 996124
rect 433524 996072 433576 996124
rect 433984 996072 434036 996124
rect 510712 996072 510764 996124
rect 522488 996072 522540 996124
rect 560576 996072 560628 996124
rect 111064 995936 111116 995988
rect 144460 995936 144512 995988
rect 162124 995936 162176 995988
rect 210240 995936 210292 995988
rect 228364 995936 228416 995988
rect 263600 995936 263652 995988
rect 264244 995936 264296 995988
rect 299296 995936 299348 995988
rect 365260 995936 365312 995988
rect 432236 995936 432288 995988
rect 434168 995936 434220 995988
rect 510896 995936 510948 995988
rect 522304 995936 522356 995988
rect 563060 995936 563112 995988
rect 124864 995800 124916 995852
rect 160376 995800 160428 995852
rect 175924 995800 175976 995852
rect 211160 995800 211212 995852
rect 213184 995800 213236 995852
rect 261116 995800 261168 995852
rect 280804 995800 280856 995852
rect 314660 995800 314712 995852
rect 364984 995800 365036 995852
rect 432052 995800 432104 995852
rect 471244 995800 471296 995852
rect 507860 995800 507912 995852
rect 509700 995800 509752 995852
rect 554136 995800 554188 995852
rect 554320 995800 554372 995852
rect 625436 995800 625488 995852
rect 195060 995528 195112 995580
rect 200948 995528 201000 995580
rect 246212 995528 246264 995580
rect 252008 995528 252060 995580
rect 298468 995528 298520 995580
rect 304448 995528 304500 995580
rect 323584 995528 323636 995580
rect 364984 995528 365036 995580
rect 366364 995528 366416 995580
rect 177304 995460 177356 995512
rect 126244 995392 126296 995444
rect 160192 995392 160244 995444
rect 212540 995392 212592 995444
rect 262864 995392 262916 995444
rect 313280 995392 313332 995444
rect 88984 995324 89036 995376
rect 92480 995324 92532 995376
rect 472624 995528 472676 995580
rect 474004 995528 474056 995580
rect 493508 995528 493560 995580
rect 511080 995528 511132 995580
rect 523868 995528 523920 995580
rect 525340 995528 525392 995580
rect 625804 995528 625856 995580
rect 627920 995528 627972 995580
rect 475936 995460 475988 995512
rect 478788 995460 478840 995512
rect 472440 995392 472492 995444
rect 474740 995392 474792 995444
rect 400864 995324 400916 995376
rect 142804 995256 142856 995308
rect 149888 995256 149940 995308
rect 194324 995256 194376 995308
rect 195244 995256 195296 995308
rect 211804 995256 211856 995308
rect 77668 995120 77720 995172
rect 100208 995120 100260 995172
rect 137928 995120 137980 995172
rect 144644 995120 144696 995172
rect 77024 994984 77076 995036
rect 102784 994984 102836 995036
rect 128452 994916 128504 994968
rect 157340 994916 157392 994968
rect 180800 995188 180852 995240
rect 244372 995256 244424 995308
rect 260932 995256 260984 995308
rect 291108 995256 291160 995308
rect 302884 995256 302936 995308
rect 244096 995188 244148 995240
rect 194692 995120 194744 995172
rect 199384 995120 199436 995172
rect 293592 995120 293644 995172
rect 298836 995120 298888 995172
rect 78312 994848 78364 994900
rect 104164 994848 104216 994900
rect 132132 994780 132184 994832
rect 145564 994780 145616 994832
rect 80152 994712 80204 994764
rect 101404 994712 101456 994764
rect 132408 994644 132460 994696
rect 149704 994644 149756 994696
rect 81348 994576 81400 994628
rect 98644 994576 98696 994628
rect 131580 994508 131632 994560
rect 155960 994780 156012 994832
rect 183284 994916 183336 994968
rect 205640 994916 205692 994968
rect 229192 994916 229244 994968
rect 234712 995052 234764 995104
rect 358728 994984 358780 995036
rect 398840 995052 398892 995104
rect 234528 994916 234580 994968
rect 259460 994916 259512 994968
rect 286508 994916 286560 994968
rect 300308 994916 300360 994968
rect 397000 994916 397052 994968
rect 402980 995324 403032 995376
rect 471428 995256 471480 995308
rect 509240 995392 509292 995444
rect 509884 995392 509936 995444
rect 560300 995392 560352 995444
rect 620284 995392 620336 995444
rect 639512 995324 639564 995376
rect 505744 995256 505796 995308
rect 532148 995256 532200 995308
rect 567200 995256 567252 995308
rect 630588 995256 630640 995308
rect 489736 995188 489788 995240
rect 472256 995120 472308 995172
rect 477684 995120 477736 995172
rect 429844 994916 429896 994968
rect 523316 995120 523368 995172
rect 526076 995120 526128 995172
rect 526260 995120 526312 995172
rect 529020 995120 529072 995172
rect 556804 995120 556856 995172
rect 640708 995120 640760 995172
rect 500684 994984 500736 995036
rect 528744 994984 528796 995036
rect 359556 994848 359608 994900
rect 393964 994848 394016 994900
rect 520556 994848 520608 994900
rect 534080 995052 534132 995104
rect 550640 994984 550692 995036
rect 635832 994984 635884 995036
rect 533068 994916 533120 994968
rect 537852 994916 537904 994968
rect 550364 994848 550416 994900
rect 625804 994848 625856 994900
rect 630772 994848 630824 994900
rect 638684 994984 638736 995036
rect 638500 994848 638552 994900
rect 640800 994916 640852 994968
rect 180616 994780 180668 994832
rect 192852 994780 192904 994832
rect 195244 994780 195296 994832
rect 207020 994780 207072 994832
rect 231584 994780 231636 994832
rect 255964 994780 256016 994832
rect 180616 994644 180668 994696
rect 204904 994644 204956 994696
rect 232872 994644 232924 994696
rect 257344 994644 257396 994696
rect 285956 994644 286008 994696
rect 289452 994644 289504 994696
rect 195244 994508 195296 994560
rect 229008 994508 229060 994560
rect 239404 994508 239456 994560
rect 283472 994508 283524 994560
rect 305644 994780 305696 994832
rect 460204 994780 460256 994832
rect 485964 994780 486016 994832
rect 486608 994780 486660 994832
rect 489736 994780 489788 994832
rect 371884 994712 371936 994764
rect 388076 994712 388128 994764
rect 388260 994712 388312 994764
rect 393320 994712 393372 994764
rect 502984 994712 503036 994764
rect 538220 994712 538272 994764
rect 571984 994712 572036 994764
rect 635188 994712 635240 994764
rect 81992 994440 82044 994492
rect 93124 994440 93176 994492
rect 192852 994372 192904 994424
rect 202144 994372 202196 994424
rect 207020 994372 207072 994424
rect 213920 994372 213972 994424
rect 232228 994372 232280 994424
rect 250444 994372 250496 994424
rect 282828 994372 282880 994424
rect 311900 994644 311952 994696
rect 469864 994644 469916 994696
rect 481364 994644 481416 994696
rect 362224 994576 362276 994628
rect 393504 994576 393556 994628
rect 502248 994576 502300 994628
rect 539232 994576 539284 994628
rect 625804 994576 625856 994628
rect 637028 994576 637080 994628
rect 140136 994236 140188 994288
rect 186504 994236 186556 994288
rect 191840 994236 191892 994288
rect 251456 994236 251508 994288
rect 284116 994236 284168 994288
rect 301504 994508 301556 994560
rect 309784 994508 309836 994560
rect 563704 994508 563756 994560
rect 624608 994508 624660 994560
rect 380900 994440 380952 994492
rect 388260 994440 388312 994492
rect 308404 994372 308456 994424
rect 397644 994440 397696 994492
rect 402980 994440 403032 994492
rect 497924 994440 497976 994492
rect 538036 994440 538088 994492
rect 357348 994236 357400 994288
rect 381176 994236 381228 994288
rect 184480 994100 184532 994152
rect 196624 994100 196676 994152
rect 239404 994100 239456 994152
rect 249064 994100 249116 994152
rect 265624 994100 265676 994152
rect 267740 994100 267792 994152
rect 289452 994100 289504 994152
rect 301504 994100 301556 994152
rect 378600 994100 378652 994152
rect 388076 994168 388128 994220
rect 549168 994372 549220 994424
rect 667112 994372 667164 994424
rect 426440 994236 426492 994288
rect 446128 994236 446180 994288
rect 547788 994236 547840 994288
rect 666560 994236 666612 994288
rect 240048 993964 240100 994016
rect 246212 993964 246264 994016
rect 496728 993284 496780 993336
rect 666928 993284 666980 993336
rect 280712 993148 280764 993200
rect 316408 993148 316460 993200
rect 351828 993148 351880 993200
rect 665180 993148 665232 993200
rect 51724 993012 51776 993064
rect 107752 993012 107804 993064
rect 147588 993012 147640 993064
rect 650000 993012 650052 993064
rect 46204 992876 46256 992928
rect 108120 992876 108172 992928
rect 148968 992876 149020 992928
rect 651380 992876 651432 992928
rect 512644 991856 512696 991908
rect 527640 991856 527692 991908
rect 267004 991720 267056 991772
rect 284300 991720 284352 991772
rect 367744 991720 367796 991772
rect 415032 991720 415084 991772
rect 419448 991720 419500 991772
rect 668032 991720 668084 991772
rect 73436 991584 73488 991636
rect 112076 991584 112128 991636
rect 200028 991584 200080 991636
rect 651748 991584 651800 991636
rect 50344 991448 50396 991500
rect 110420 991448 110472 991500
rect 138296 991448 138348 991500
rect 162860 991448 162912 991500
rect 198648 991448 198700 991500
rect 650736 991448 650788 991500
rect 562508 990496 562560 990548
rect 672724 990496 672776 990548
rect 435364 990360 435416 990412
rect 463608 990360 463660 990412
rect 498108 990360 498160 990412
rect 666744 990360 666796 990412
rect 303528 990224 303580 990276
rect 665456 990224 665508 990276
rect 48964 990088 49016 990140
rect 109040 990088 109092 990140
rect 249708 990088 249760 990140
rect 648896 990088 648948 990140
rect 422208 988864 422260 988916
rect 668216 988864 668268 988916
rect 250996 988728 251048 988780
rect 650184 988728 650236 988780
rect 559564 987640 559616 987692
rect 669964 987640 670016 987692
rect 352840 987504 352892 987556
rect 668400 987504 668452 987556
rect 96344 987368 96396 987420
rect 650920 987368 650972 987420
rect 203156 986620 203208 986672
rect 207020 986620 207072 986672
rect 217324 986620 217376 986672
rect 219440 986620 219492 986672
rect 570604 986212 570656 986264
rect 592500 986212 592552 986264
rect 370504 986076 370556 986128
rect 397828 986076 397880 986128
rect 463608 986076 463660 986128
rect 478972 986076 479024 986128
rect 519544 986076 519596 986128
rect 543832 986076 543884 986128
rect 565084 986076 565136 986128
rect 608784 986076 608836 986128
rect 89628 985940 89680 985992
rect 106924 985940 106976 985992
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 279424 985940 279476 985992
rect 300492 985940 300544 985992
rect 369124 985940 369176 985992
rect 414112 985940 414164 985992
rect 415032 985940 415084 985992
rect 430304 985940 430356 985992
rect 436744 985940 436796 985992
rect 462780 985940 462832 985992
rect 465724 985940 465776 985992
rect 495164 985940 495216 985992
rect 515404 985940 515456 985992
rect 560116 985940 560168 985992
rect 562324 985940 562376 985992
rect 658924 985940 658976 985992
rect 560944 984852 560996 984904
rect 660304 984852 660356 984904
rect 302148 984716 302200 984768
rect 665640 984716 665692 984768
rect 96528 984580 96580 984632
rect 650368 984580 650420 984632
rect 55864 975672 55916 975724
rect 62120 975672 62172 975724
rect 651564 975672 651616 975724
rect 661684 975672 661736 975724
rect 42524 969416 42576 969468
rect 55864 969416 55916 969468
rect 42248 966832 42300 966884
rect 42708 966832 42760 966884
rect 673368 966152 673420 966204
rect 675116 966152 675168 966204
rect 42432 964656 42484 964708
rect 42892 964656 42944 964708
rect 42432 963840 42484 963892
rect 44180 963840 44232 963892
rect 42432 963432 42484 963484
rect 43076 963432 43128 963484
rect 42432 961868 42484 961920
rect 44456 961868 44508 961920
rect 47584 961868 47636 961920
rect 62120 961868 62172 961920
rect 651564 961868 651616 961920
rect 663064 961868 663116 961920
rect 674288 961868 674340 961920
rect 675116 961868 675168 961920
rect 42432 959080 42484 959132
rect 43260 959080 43312 959132
rect 42432 958264 42484 958316
rect 44640 958264 44692 958316
rect 674472 957856 674524 957908
rect 675116 957856 675168 957908
rect 660488 957720 660540 957772
rect 675300 957312 675352 957364
rect 673184 956360 673236 956412
rect 675116 956360 675168 956412
rect 35164 951464 35216 951516
rect 41696 951464 41748 951516
rect 675852 949424 675904 949476
rect 678244 949424 678296 949476
rect 675852 948744 675904 948796
rect 682384 948744 682436 948796
rect 651564 948064 651616 948116
rect 671344 948064 671396 948116
rect 43536 945956 43588 946008
rect 62120 945956 62172 946008
rect 663064 941808 663116 941860
rect 675484 941808 675536 941860
rect 41328 941468 41380 941520
rect 41696 941468 41748 941520
rect 43628 941332 43680 941384
rect 48964 941332 49016 941384
rect 43444 941196 43496 941248
rect 50344 941196 50396 941248
rect 40960 940108 41012 940160
rect 41696 940108 41748 940160
rect 43444 939768 43496 939820
rect 51724 939768 51776 939820
rect 672724 938680 672776 938732
rect 675484 938680 675536 938732
rect 40960 938544 41012 938596
rect 41512 938544 41564 938596
rect 671344 938544 671396 938596
rect 675300 938544 675352 938596
rect 41144 938408 41196 938460
rect 41512 938408 41564 938460
rect 661684 938408 661736 938460
rect 674932 938408 674984 938460
rect 671528 937524 671580 937576
rect 675484 937524 675536 937576
rect 660304 937320 660356 937372
rect 675484 937320 675536 937372
rect 658924 937184 658976 937236
rect 674932 937184 674984 937236
rect 671160 937048 671212 937100
rect 675300 937048 675352 937100
rect 44640 936980 44692 937032
rect 62120 936980 62172 937032
rect 651564 936980 651616 937032
rect 660488 936980 660540 937032
rect 669964 935892 670016 935944
rect 675484 935892 675536 935944
rect 672080 935756 672132 935808
rect 675484 935756 675536 935808
rect 672448 935620 672500 935672
rect 675300 935620 675352 935672
rect 673000 933308 673052 933360
rect 675484 933308 675536 933360
rect 673368 932968 673420 933020
rect 675484 932968 675536 933020
rect 43444 932900 43496 932952
rect 54484 932900 54536 932952
rect 42800 931540 42852 931592
rect 53104 931540 53156 931592
rect 673184 930112 673236 930164
rect 675484 930112 675536 930164
rect 678244 930044 678296 930096
rect 683120 930044 683172 930096
rect 669780 928752 669832 928804
rect 675484 928752 675536 928804
rect 670608 927392 670660 927444
rect 675484 927392 675536 927444
rect 47584 923244 47636 923296
rect 62120 923244 62172 923296
rect 651564 921816 651616 921868
rect 661684 921816 661736 921868
rect 50344 909440 50396 909492
rect 62120 909440 62172 909492
rect 651564 909440 651616 909492
rect 664444 909440 664496 909492
rect 46204 896996 46256 897048
rect 62120 896996 62172 897048
rect 651564 895636 651616 895688
rect 663064 895636 663116 895688
rect 42432 884688 42484 884740
rect 62120 884688 62172 884740
rect 652392 881832 652444 881884
rect 671344 881832 671396 881884
rect 669596 879044 669648 879096
rect 675300 879044 675352 879096
rect 43444 870816 43496 870868
rect 62120 870816 62172 870868
rect 651564 869388 651616 869440
rect 658924 869388 658976 869440
rect 673000 869388 673052 869440
rect 675116 869388 675168 869440
rect 671344 868980 671396 869032
rect 675024 868980 675076 869032
rect 674656 868028 674708 868080
rect 675116 868028 675168 868080
rect 670976 866804 671028 866856
rect 675116 866804 675168 866856
rect 669228 866668 669280 866720
rect 675024 866396 675076 866448
rect 674472 864628 674524 864680
rect 675300 864628 675352 864680
rect 673368 862860 673420 862912
rect 675116 862860 675168 862912
rect 51908 858372 51960 858424
rect 62120 858372 62172 858424
rect 651564 855584 651616 855636
rect 671344 855584 671396 855636
rect 44824 844568 44876 844620
rect 62120 844568 62172 844620
rect 651564 841780 651616 841832
rect 659108 841780 659160 841832
rect 55864 832124 55916 832176
rect 62120 832124 62172 832176
rect 651564 829404 651616 829456
rect 660304 829404 660356 829456
rect 51724 818320 51776 818372
rect 62120 818320 62172 818372
rect 35808 817096 35860 817148
rect 40684 817096 40736 817148
rect 35624 816960 35676 817012
rect 39948 816960 40000 817012
rect 35624 816008 35676 816060
rect 41696 816008 41748 816060
rect 35440 815872 35492 815924
rect 41696 815872 41748 815924
rect 35808 815736 35860 815788
rect 41328 815736 41380 815788
rect 35256 815600 35308 815652
rect 41696 815600 41748 815652
rect 42156 815600 42208 815652
rect 50344 815600 50396 815652
rect 651564 815600 651616 815652
rect 661868 815600 661920 815652
rect 35808 814648 35860 814700
rect 41696 814716 41748 814768
rect 35624 814376 35676 814428
rect 40316 814376 40368 814428
rect 35440 814240 35492 814292
rect 41696 814240 41748 814292
rect 42064 814240 42116 814292
rect 44180 814240 44232 814292
rect 41144 812948 41196 813000
rect 41512 812948 41564 813000
rect 41328 811588 41380 811640
rect 41696 811588 41748 811640
rect 43628 807440 43680 807492
rect 48964 807440 49016 807492
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 651564 803224 651616 803276
rect 663248 803224 663300 803276
rect 32404 802544 32456 802596
rect 41696 802544 41748 802596
rect 31668 802272 31720 802324
rect 39764 802272 39816 802324
rect 36544 801728 36596 801780
rect 39856 801728 39908 801780
rect 33784 800912 33836 800964
rect 40040 800912 40092 800964
rect 43628 799008 43680 799060
rect 47584 799008 47636 799060
rect 47768 793568 47820 793620
rect 62120 793568 62172 793620
rect 42248 792548 42300 792600
rect 43076 792548 43128 792600
rect 42708 790236 42760 790288
rect 42156 789964 42208 790016
rect 651564 789352 651616 789404
rect 662052 789352 662104 789404
rect 670240 789352 670292 789404
rect 675116 789352 675168 789404
rect 670792 787992 670844 788044
rect 675116 787992 675168 788044
rect 674288 784116 674340 784168
rect 675116 784116 675168 784168
rect 672264 782620 672316 782672
rect 675116 782620 675168 782672
rect 668768 782484 668820 782536
rect 675300 782484 675352 782536
rect 56232 780036 56284 780088
rect 62120 780036 62172 780088
rect 673644 779764 673696 779816
rect 675116 779764 675168 779816
rect 673828 779084 673880 779136
rect 675116 779084 675168 779136
rect 660304 778948 660356 779000
rect 675116 778948 675168 779000
rect 672816 778336 672868 778388
rect 675300 778336 675352 778388
rect 674196 776976 674248 777028
rect 675300 776976 675352 777028
rect 674840 775888 674892 775940
rect 675208 775888 675260 775940
rect 675024 775752 675076 775804
rect 651564 775548 651616 775600
rect 660488 775548 660540 775600
rect 674840 775548 674892 775600
rect 35808 774324 35860 774376
rect 39764 774324 39816 774376
rect 35532 773372 35584 773424
rect 40868 773372 40920 773424
rect 35808 773236 35860 773288
rect 35808 773100 35860 773152
rect 41696 773100 41748 773152
rect 42064 773100 42116 773152
rect 44456 773100 44508 773152
rect 41696 772964 41748 773016
rect 42064 772964 42116 773016
rect 55864 772964 55916 773016
rect 35348 772828 35400 772880
rect 51908 772828 51960 772880
rect 41696 772692 41748 772744
rect 42064 772692 42116 772744
rect 676036 772216 676088 772268
rect 683304 772216 683356 772268
rect 675852 772080 675904 772132
rect 684132 772080 684184 772132
rect 35532 771672 35584 771724
rect 39856 771672 39908 771724
rect 35808 771536 35860 771588
rect 41696 771536 41748 771588
rect 42064 771536 42116 771588
rect 42892 771536 42944 771588
rect 35348 771400 35400 771452
rect 41696 771400 41748 771452
rect 42064 771400 42116 771452
rect 44180 771400 44232 771452
rect 35808 770448 35860 770500
rect 39856 770448 39908 770500
rect 35624 770176 35676 770228
rect 41696 770244 41748 770296
rect 42064 770244 42116 770296
rect 43260 770244 43312 770296
rect 35808 770040 35860 770092
rect 41696 770040 41748 770092
rect 42064 770040 42116 770092
rect 44640 770040 44692 770092
rect 35808 768816 35860 768868
rect 39304 768816 39356 768868
rect 35624 768680 35676 768732
rect 41328 768680 41380 768732
rect 35808 767592 35860 767644
rect 40040 767592 40092 767644
rect 35624 767456 35676 767508
rect 36544 767456 36596 767508
rect 43628 767320 43680 767372
rect 62120 767320 62172 767372
rect 674932 766368 674984 766420
rect 675392 766368 675444 766420
rect 35808 766300 35860 766352
rect 39764 766164 39816 766216
rect 35808 765892 35860 765944
rect 41696 765960 41748 766012
rect 42064 765892 42116 765944
rect 44456 765892 44508 765944
rect 40040 765144 40092 765196
rect 41696 765144 41748 765196
rect 42064 765008 42116 765060
rect 42524 765008 42576 765060
rect 35808 764668 35860 764720
rect 39120 764668 39172 764720
rect 35808 763308 35860 763360
rect 37924 763308 37976 763360
rect 35624 763172 35676 763224
rect 41696 763240 41748 763292
rect 651564 763240 651616 763292
rect 660304 763172 660356 763224
rect 35808 761880 35860 761932
rect 40224 761880 40276 761932
rect 664444 760860 664496 760912
rect 675484 760860 675536 760912
rect 661684 760520 661736 760572
rect 675300 760520 675352 760572
rect 663064 760384 663116 760436
rect 675484 760384 675536 760436
rect 671528 760248 671580 760300
rect 675300 760248 675352 760300
rect 671528 759840 671580 759892
rect 675484 759840 675536 759892
rect 671160 759500 671212 759552
rect 675484 759500 675536 759552
rect 36544 759024 36596 759076
rect 39948 759024 40000 759076
rect 671160 759024 671212 759076
rect 675484 759024 675536 759076
rect 672080 758684 672132 758736
rect 675484 758684 675536 758736
rect 673184 758208 673236 758260
rect 675484 758208 675536 758260
rect 35164 758140 35216 758192
rect 41696 758140 41748 758192
rect 42432 758140 42484 758192
rect 37924 757732 37976 757784
rect 41604 757732 41656 757784
rect 672448 757868 672500 757920
rect 675484 757868 675536 757920
rect 42432 757596 42484 757648
rect 672080 757392 672132 757444
rect 675484 757392 675536 757444
rect 674012 756236 674064 756288
rect 675116 756236 675168 756288
rect 673368 755012 673420 755064
rect 675484 755012 675536 755064
rect 44456 754876 44508 754928
rect 669596 754604 669648 754656
rect 675484 754604 675536 754656
rect 42248 754264 42300 754316
rect 672632 754196 672684 754248
rect 675484 754196 675536 754248
rect 43444 753516 43496 753568
rect 45008 753516 45060 753568
rect 50712 753516 50764 753568
rect 62120 753516 62172 753568
rect 670976 753380 671028 753432
rect 675484 753380 675536 753432
rect 673000 752156 673052 752208
rect 675484 752156 675536 752208
rect 671804 751748 671856 751800
rect 675484 751748 675536 751800
rect 675852 750932 675904 750984
rect 683120 750932 683172 750984
rect 669596 750048 669648 750100
rect 675484 750048 675536 750100
rect 651564 749368 651616 749420
rect 664444 749368 664496 749420
rect 42432 749300 42484 749352
rect 43260 749300 43312 749352
rect 669228 743656 669280 743708
rect 675116 743656 675168 743708
rect 671896 742772 671948 742824
rect 675300 742772 675352 742824
rect 666376 742432 666428 742484
rect 675300 742432 675352 742484
rect 674840 741616 674892 741668
rect 675484 741616 675536 741668
rect 56048 741072 56100 741124
rect 62120 741072 62172 741124
rect 674472 739712 674524 739764
rect 675116 739712 675168 739764
rect 674012 738624 674064 738676
rect 675392 738624 675444 738676
rect 651564 735564 651616 735616
rect 663064 735564 663116 735616
rect 670792 734952 670844 735004
rect 675300 734952 675352 735004
rect 660488 734816 660540 734868
rect 675300 734816 675352 734868
rect 667664 732776 667716 732828
rect 675116 732776 675168 732828
rect 43444 731144 43496 731196
rect 50344 731144 50396 731196
rect 43260 730124 43312 730176
rect 56232 730056 56284 730108
rect 41328 728628 41380 728680
rect 41696 728628 41748 728680
rect 42064 728628 42116 728680
rect 45008 728628 45060 728680
rect 670424 728628 670476 728680
rect 675116 728628 675168 728680
rect 41052 727404 41104 727456
rect 41696 727404 41748 727456
rect 42064 727404 42116 727456
rect 43076 727404 43128 727456
rect 40868 727268 40920 727320
rect 41696 727268 41748 727320
rect 42064 727268 42116 727320
rect 44272 727268 44324 727320
rect 51908 727268 51960 727320
rect 62120 727268 62172 727320
rect 675852 726792 675904 726844
rect 684224 726792 684276 726844
rect 676036 726520 676088 726572
rect 683212 726520 683264 726572
rect 41328 726316 41380 726368
rect 41604 726316 41656 726368
rect 651564 723120 651616 723172
rect 659292 723120 659344 723172
rect 31760 720264 31812 720316
rect 40040 720264 40092 720316
rect 42340 719108 42392 719160
rect 55864 719108 55916 719160
rect 671344 716524 671396 716576
rect 675484 716524 675536 716576
rect 37924 716048 37976 716100
rect 40316 716048 40368 716100
rect 35164 715640 35216 715692
rect 41328 715640 41380 715692
rect 33784 715368 33836 715420
rect 41696 715368 41748 715420
rect 671528 715300 671580 715352
rect 675116 715300 675168 715352
rect 42064 715232 42116 715284
rect 42708 715232 42760 715284
rect 659108 715096 659160 715148
rect 675484 715096 675536 715148
rect 658924 714960 658976 715012
rect 675300 714960 675352 715012
rect 50528 714824 50580 714876
rect 62120 714824 62172 714876
rect 671528 714824 671580 714876
rect 675484 714824 675536 714876
rect 40040 714484 40092 714536
rect 41696 714484 41748 714536
rect 671160 714484 671212 714536
rect 675484 714484 675536 714536
rect 673000 714008 673052 714060
rect 675484 714008 675536 714060
rect 673184 713668 673236 713720
rect 675484 713668 675536 713720
rect 671160 713192 671212 713244
rect 675484 713192 675536 713244
rect 672080 712852 672132 712904
rect 675484 712852 675536 712904
rect 671344 712376 671396 712428
rect 675484 712376 675536 712428
rect 42892 712240 42944 712292
rect 51724 712240 51776 712292
rect 676220 712036 676272 712088
rect 677508 712036 677560 712088
rect 676036 711832 676088 711884
rect 676772 711832 676824 711884
rect 670976 711220 671028 711272
rect 675484 711220 675536 711272
rect 42248 710948 42300 711000
rect 42892 710948 42944 711000
rect 668584 709724 668636 709776
rect 675484 709724 675536 709776
rect 670240 709588 670292 709640
rect 675484 709588 675536 709640
rect 44180 709316 44232 709368
rect 651564 709316 651616 709368
rect 658924 709316 658976 709368
rect 668768 709316 668820 709368
rect 675300 709316 675352 709368
rect 42340 708364 42392 708416
rect 673828 707956 673880 708008
rect 675484 707956 675536 708008
rect 43076 707752 43128 707804
rect 43444 707752 43496 707804
rect 672356 707548 672408 707600
rect 675484 707548 675536 707600
rect 673644 707140 673696 707192
rect 675484 707140 675536 707192
rect 672816 706732 672868 706784
rect 675484 706732 675536 706784
rect 675852 705168 675904 705220
rect 683120 705168 683172 705220
rect 669964 705032 670016 705084
rect 675484 705032 675536 705084
rect 42248 702108 42300 702160
rect 42248 701836 42300 701888
rect 51724 701020 51776 701072
rect 62120 701020 62172 701072
rect 668768 699660 668820 699712
rect 675116 699660 675168 699712
rect 651564 696940 651616 696992
rect 664628 696940 664680 696992
rect 673644 694152 673696 694204
rect 675116 694152 675168 694204
rect 673828 693336 673880 693388
rect 675116 693336 675168 693388
rect 674656 692996 674708 693048
rect 675392 692996 675444 693048
rect 666100 692860 666152 692912
rect 675116 692860 675168 692912
rect 672816 690004 672868 690056
rect 675116 690004 675168 690056
rect 659292 689256 659344 689308
rect 674932 689256 674984 689308
rect 43812 688644 43864 688696
rect 62120 688644 62172 688696
rect 674196 687896 674248 687948
rect 675300 687896 675352 687948
rect 43444 687692 43496 687744
rect 50712 687692 50764 687744
rect 671252 687420 671304 687472
rect 675116 687420 675168 687472
rect 43260 687352 43312 687404
rect 51908 687352 51960 687404
rect 40960 687216 41012 687268
rect 41696 687216 41748 687268
rect 42064 687216 42116 687268
rect 56048 687216 56100 687268
rect 41144 685992 41196 686044
rect 41696 686060 41748 686112
rect 42064 686060 42116 686112
rect 44456 686060 44508 686112
rect 41328 685856 41380 685908
rect 41696 685856 41748 685908
rect 42064 685856 42116 685908
rect 45008 685856 45060 685908
rect 669412 685856 669464 685908
rect 675300 685516 675352 685568
rect 40868 684768 40920 684820
rect 41144 684632 41196 684684
rect 41696 684700 41748 684752
rect 42064 684700 42116 684752
rect 42892 684700 42944 684752
rect 41696 684496 41748 684548
rect 42064 684496 42116 684548
rect 44272 684496 44324 684548
rect 41328 683476 41380 683528
rect 41696 683476 41748 683528
rect 651564 683136 651616 683188
rect 659108 683136 659160 683188
rect 675852 682388 675904 682440
rect 683396 682388 683448 682440
rect 40776 679328 40828 679380
rect 41328 679328 41380 679380
rect 40592 679192 40644 679244
rect 41696 679192 41748 679244
rect 43996 676404 44048 676456
rect 50344 676404 50396 676456
rect 47768 674840 47820 674892
rect 62120 674840 62172 674892
rect 33784 672732 33836 672784
rect 39488 672732 39540 672784
rect 36544 672052 36596 672104
rect 41696 672052 41748 672104
rect 37924 671236 37976 671288
rect 40040 671236 40092 671288
rect 663248 670828 663300 670880
rect 675300 670828 675352 670880
rect 661868 670692 661920 670744
rect 675484 670692 675536 670744
rect 673000 669740 673052 669792
rect 674840 669740 674892 669792
rect 671528 669604 671580 669656
rect 675300 669604 675352 669656
rect 671620 669468 671672 669520
rect 675484 669468 675536 669520
rect 651564 669332 651616 669384
rect 661868 669332 661920 669384
rect 662052 669332 662104 669384
rect 675484 669332 675536 669384
rect 671068 668516 671120 668568
rect 675484 668516 675536 668568
rect 671068 668380 671120 668432
rect 675300 668380 675352 668432
rect 672356 668040 672408 668092
rect 675484 668040 675536 668092
rect 45192 667904 45244 667956
rect 42248 667768 42300 667820
rect 671436 667700 671488 667752
rect 675484 667700 675536 667752
rect 673276 667224 673328 667276
rect 675484 667224 675536 667276
rect 44640 666544 44692 666596
rect 671988 666068 672040 666120
rect 675484 666068 675536 666120
rect 42248 666000 42300 666052
rect 667664 665320 667716 665372
rect 675300 665320 675352 665372
rect 666376 665184 666428 665236
rect 675484 665184 675536 665236
rect 670424 664844 670476 664896
rect 675484 664844 675536 664896
rect 669228 663756 669280 663808
rect 675484 663756 675536 663808
rect 42524 663280 42576 663332
rect 42340 663212 42392 663264
rect 673460 663212 673512 663264
rect 675484 663212 675536 663264
rect 42708 663008 42760 663060
rect 43444 663008 43496 663060
rect 42524 662940 42576 662992
rect 672540 662804 672592 662856
rect 675484 662804 675536 662856
rect 42524 662668 42576 662720
rect 43444 662396 43496 662448
rect 62120 662396 62172 662448
rect 670792 661988 670844 662040
rect 675484 661988 675536 662040
rect 671804 661580 671856 661632
rect 675484 661580 675536 661632
rect 670792 661104 670844 661156
rect 675484 661104 675536 661156
rect 42156 660492 42208 660544
rect 42708 660492 42760 660544
rect 670976 659948 671028 660000
rect 675484 659948 675536 660000
rect 675852 659812 675904 659864
rect 683120 659812 683172 659864
rect 42064 657364 42116 657416
rect 42616 657364 42668 657416
rect 651564 656888 651616 656940
rect 661684 656888 661736 656940
rect 664996 654100 665048 654152
rect 675300 654100 675352 654152
rect 671896 651380 671948 651432
rect 675300 651380 675352 651432
rect 668952 649068 669004 649120
rect 674840 649136 674892 649188
rect 51908 647844 51960 647896
rect 62120 647844 62172 647896
rect 669228 647708 669280 647760
rect 675392 647708 675444 647760
rect 35808 644716 35860 644768
rect 39396 644716 39448 644768
rect 35532 644444 35584 644496
rect 39764 644444 39816 644496
rect 670240 644444 670292 644496
rect 674840 644444 674892 644496
rect 661868 643696 661920 643748
rect 675300 643628 675352 643680
rect 35808 643492 35860 643544
rect 39672 643492 39724 643544
rect 35532 643220 35584 643272
rect 41696 643288 41748 643340
rect 42064 643288 42116 643340
rect 44456 643288 44508 643340
rect 35348 643084 35400 643136
rect 41696 643084 41748 643136
rect 42064 643084 42116 643136
rect 51724 643084 51776 643136
rect 651564 643084 651616 643136
rect 663248 643084 663300 643136
rect 35808 642132 35860 642184
rect 38936 642200 38988 642252
rect 35440 641860 35492 641912
rect 39580 641996 39632 642048
rect 666284 641860 666336 641912
rect 674840 641860 674892 641912
rect 35624 641724 35676 641776
rect 41696 641724 41748 641776
rect 42064 641724 42116 641776
rect 44180 641724 44232 641776
rect 665916 641724 665968 641776
rect 670424 641724 670476 641776
rect 670424 641248 670476 641300
rect 675300 641248 675352 641300
rect 35808 640772 35860 640824
rect 39672 640704 39724 640756
rect 673644 640568 673696 640620
rect 673828 640568 673880 640620
rect 35624 640432 35676 640484
rect 39856 640432 39908 640484
rect 35808 640296 35860 640348
rect 41696 640296 41748 640348
rect 42064 640296 42116 640348
rect 43076 640296 43128 640348
rect 673644 640296 673696 640348
rect 673828 640296 673880 640348
rect 35808 639072 35860 639124
rect 40224 639072 40276 639124
rect 35532 638936 35584 638988
rect 40040 638936 40092 638988
rect 35348 638188 35400 638240
rect 41696 638188 41748 638240
rect 35532 637916 35584 637968
rect 40960 637916 41012 637968
rect 35808 637712 35860 637764
rect 41512 637712 41564 637764
rect 676036 637508 676088 637560
rect 682384 637508 682436 637560
rect 676036 636828 676088 636880
rect 683304 636828 683356 636880
rect 35808 636352 35860 636404
rect 40684 636352 40736 636404
rect 49148 636216 49200 636268
rect 62120 636216 62172 636268
rect 35808 635060 35860 635112
rect 39580 635060 39632 635112
rect 35624 634788 35676 634840
rect 40500 634788 40552 634840
rect 35808 633836 35860 633888
rect 41696 633700 41748 633752
rect 42064 633700 42116 633752
rect 53288 633700 53340 633752
rect 35808 633496 35860 633548
rect 41696 633496 41748 633548
rect 42064 633496 42116 633548
rect 51724 633564 51776 633616
rect 675852 633564 675904 633616
rect 682568 633564 682620 633616
rect 33784 630028 33836 630080
rect 41696 630028 41748 630080
rect 42064 629960 42116 630012
rect 42708 629960 42760 630012
rect 32404 629892 32456 629944
rect 41696 629892 41748 629944
rect 651564 629280 651616 629332
rect 661868 629280 661920 629332
rect 42892 626628 42944 626680
rect 50528 626628 50580 626680
rect 664444 625676 664496 625728
rect 675484 625676 675536 625728
rect 663064 625404 663116 625456
rect 42524 625336 42576 625388
rect 42248 625132 42300 625184
rect 675484 625268 675536 625320
rect 660304 625132 660356 625184
rect 675116 625132 675168 625184
rect 671528 624928 671580 624980
rect 675484 624928 675536 624980
rect 42340 624656 42392 624708
rect 43812 624656 43864 624708
rect 672908 624656 672960 624708
rect 675484 624656 675536 624708
rect 671160 624316 671212 624368
rect 675484 624316 675536 624368
rect 47768 623772 47820 623824
rect 62120 623772 62172 623824
rect 672356 623500 672408 623552
rect 675484 623500 675536 623552
rect 671528 623024 671580 623076
rect 675484 623024 675536 623076
rect 673460 622888 673512 622940
rect 673460 622684 673512 622736
rect 673644 622684 673696 622736
rect 675484 622684 675536 622736
rect 672080 622208 672132 622260
rect 675484 622208 675536 622260
rect 669412 619828 669464 619880
rect 675024 619828 675076 619880
rect 666100 619624 666152 619676
rect 675484 619624 675536 619676
rect 673092 619080 673144 619132
rect 674840 619080 674892 619132
rect 42616 618876 42668 618928
rect 43628 618876 43680 618928
rect 668768 618264 668820 618316
rect 675484 618264 675536 618316
rect 671344 618128 671396 618180
rect 675484 618128 675536 618180
rect 673276 616972 673328 617024
rect 675484 616972 675536 617024
rect 651564 616836 651616 616888
rect 660488 616836 660540 616888
rect 668584 616768 668636 616820
rect 669780 616768 669832 616820
rect 672724 616564 672776 616616
rect 675484 616564 675536 616616
rect 670424 616088 670476 616140
rect 675484 616088 675536 616140
rect 42248 615680 42300 615732
rect 675852 615612 675904 615664
rect 683120 615612 683172 615664
rect 42248 615476 42300 615528
rect 672172 614864 672224 614916
rect 675484 614864 675536 614916
rect 42156 613572 42208 613624
rect 44364 613572 44416 613624
rect 43628 609220 43680 609272
rect 62120 609220 62172 609272
rect 663524 608608 663576 608660
rect 675208 608812 675260 608864
rect 670332 607112 670384 607164
rect 670148 606840 670200 606892
rect 674288 604324 674340 604376
rect 675300 604324 675352 604376
rect 673644 603440 673696 603492
rect 675392 603440 675444 603492
rect 652576 603100 652628 603152
rect 660304 603100 660356 603152
rect 667848 603100 667900 603152
rect 674840 603100 674892 603152
rect 35808 601672 35860 601724
rect 41696 601672 41748 601724
rect 42064 601672 42116 601724
rect 49148 601672 49200 601724
rect 670424 601672 670476 601724
rect 675300 601672 675352 601724
rect 43812 600380 43864 600432
rect 51908 600312 51960 600364
rect 660488 599564 660540 599616
rect 675300 599564 675352 599616
rect 41328 598952 41380 599004
rect 41696 598952 41748 599004
rect 42064 598952 42116 599004
rect 44456 598952 44508 599004
rect 41052 597796 41104 597848
rect 41696 597864 41748 597916
rect 42064 597864 42116 597916
rect 42892 597864 42944 597916
rect 40868 597660 40920 597712
rect 41696 597728 41748 597780
rect 42064 597728 42116 597780
rect 43168 597728 43220 597780
rect 41328 597524 41380 597576
rect 41696 597524 41748 597576
rect 42064 597524 42116 597576
rect 43812 597524 43864 597576
rect 49148 597524 49200 597576
rect 62120 597524 62172 597576
rect 666100 596164 666152 596216
rect 674748 596164 674800 596216
rect 41144 595892 41196 595944
rect 41696 595892 41748 595944
rect 668768 595212 668820 595264
rect 675300 595212 675352 595264
rect 674748 595008 674800 595060
rect 675300 595008 675352 595060
rect 40776 592832 40828 592884
rect 41696 592832 41748 592884
rect 675852 592628 675904 592680
rect 683304 592628 683356 592680
rect 675852 592492 675904 592544
rect 678244 592492 678296 592544
rect 42064 591880 42116 591932
rect 42432 591880 42484 591932
rect 675852 591404 675904 591456
rect 683488 591404 683540 591456
rect 675852 591268 675904 591320
rect 684132 591268 684184 591320
rect 43260 590792 43312 590844
rect 50528 590792 50580 590844
rect 651564 590656 651616 590708
rect 664444 590656 664496 590708
rect 668768 589228 668820 589280
rect 669412 589228 669464 589280
rect 33048 587120 33100 587172
rect 39580 587120 39632 587172
rect 36544 586372 36596 586424
rect 39580 586372 39632 586424
rect 35164 585896 35216 585948
rect 40500 585896 40552 585948
rect 31024 585556 31076 585608
rect 39672 585556 39724 585608
rect 51908 583720 51960 583772
rect 62120 583720 62172 583772
rect 43168 581000 43220 581052
rect 44640 581000 44692 581052
rect 664628 581000 664680 581052
rect 675484 581000 675536 581052
rect 673000 579980 673052 580032
rect 675484 579980 675536 580032
rect 658924 579776 658976 579828
rect 674932 579776 674984 579828
rect 659108 579640 659160 579692
rect 675300 579640 675352 579692
rect 673276 578484 673328 578536
rect 675300 578484 675352 578536
rect 42248 578416 42300 578468
rect 673092 578348 673144 578400
rect 675484 578348 675536 578400
rect 672908 578212 672960 578264
rect 674932 578212 674984 578264
rect 42248 577804 42300 577856
rect 673460 577600 673512 577652
rect 675484 577600 675536 577652
rect 671344 577260 671396 577312
rect 675300 577260 675352 577312
rect 671988 577124 672040 577176
rect 675484 577124 675536 577176
rect 671528 576988 671580 577040
rect 673368 576988 673420 577040
rect 651564 576852 651616 576904
rect 659292 576852 659344 576904
rect 671160 576852 671212 576904
rect 675484 576920 675536 576972
rect 671896 575492 671948 575544
rect 675484 575492 675536 575544
rect 672540 574336 672592 574388
rect 675484 574336 675536 574388
rect 666284 574200 666336 574252
rect 675300 574200 675352 574252
rect 664996 574064 665048 574116
rect 675484 574064 675536 574116
rect 42156 573452 42208 573504
rect 42616 573452 42668 573504
rect 670240 572840 670292 572892
rect 675484 572840 675536 572892
rect 668860 572704 668912 572756
rect 675300 572704 675352 572756
rect 43444 571344 43496 571396
rect 62120 571344 62172 571396
rect 671712 571208 671764 571260
rect 675300 571208 675352 571260
rect 675852 570052 675904 570104
rect 683120 570052 683172 570104
rect 665916 569984 665968 570036
rect 675484 569984 675536 570036
rect 671344 569576 671396 569628
rect 675484 569576 675536 569628
rect 675852 565156 675904 565208
rect 676220 565156 676272 565208
rect 664996 564544 665048 564596
rect 675300 564544 675352 564596
rect 663708 564408 663760 564460
rect 675484 564408 675536 564460
rect 652392 563048 652444 563100
rect 658924 563048 658976 563100
rect 674656 558220 674708 558272
rect 675392 558220 675444 558272
rect 43444 557812 43496 557864
rect 49148 557812 49200 557864
rect 673276 557676 673328 557728
rect 675300 557676 675352 557728
rect 43260 557540 43312 557592
rect 51908 557540 51960 557592
rect 54852 557540 54904 557592
rect 62120 557540 62172 557592
rect 666376 557540 666428 557592
rect 675300 557540 675352 557592
rect 40868 554888 40920 554940
rect 41696 554888 41748 554940
rect 42064 554888 42116 554940
rect 42800 554888 42852 554940
rect 40592 554752 40644 554804
rect 41696 554752 41748 554804
rect 42064 554752 42116 554804
rect 44364 554752 44416 554804
rect 671804 554752 671856 554804
rect 675116 554752 675168 554804
rect 673460 554140 673512 554192
rect 675116 554140 675168 554192
rect 658924 554004 658976 554056
rect 675116 554004 675168 554056
rect 42064 550672 42116 550724
rect 43168 550672 43220 550724
rect 651564 550604 651616 550656
rect 658924 550604 658976 550656
rect 40040 550400 40092 550452
rect 41696 550400 41748 550452
rect 42064 550332 42116 550384
rect 42524 550332 42576 550384
rect 674472 549720 674524 549772
rect 675300 549720 675352 549772
rect 41144 548088 41196 548140
rect 41696 548088 41748 548140
rect 43444 547884 43496 547936
rect 56048 547884 56100 547936
rect 31760 547408 31812 547460
rect 38476 547408 38528 547460
rect 675944 546796 675996 546848
rect 681004 546796 681056 546848
rect 43444 546524 43496 546576
rect 49148 546524 49200 546576
rect 676128 545708 676180 545760
rect 683212 545708 683264 545760
rect 674472 545436 674524 545488
rect 675024 545436 675076 545488
rect 43444 545096 43496 545148
rect 62120 545096 62172 545148
rect 34428 544348 34480 544400
rect 39488 544348 39540 544400
rect 38476 542172 38528 542224
rect 39764 542172 39816 542224
rect 42708 540676 42760 540728
rect 43628 540676 43680 540728
rect 42432 537616 42484 537668
rect 44088 537616 44140 537668
rect 651564 536800 651616 536852
rect 663064 536800 663116 536852
rect 42708 536596 42760 536648
rect 45376 536596 45428 536648
rect 663248 535576 663300 535628
rect 675484 535644 675536 535696
rect 661684 535440 661736 535492
rect 675484 535440 675536 535492
rect 42340 535236 42392 535288
rect 43904 535236 43956 535288
rect 673092 534556 673144 534608
rect 674932 534556 674984 534608
rect 672908 534352 672960 534404
rect 675484 534420 675536 534472
rect 661868 534216 661920 534268
rect 674472 534216 674524 534268
rect 673000 534080 673052 534132
rect 675484 534080 675536 534132
rect 42432 533400 42484 533452
rect 43076 533400 43128 533452
rect 671528 533332 671580 533384
rect 675484 533332 675536 533384
rect 672540 532720 672592 532772
rect 675484 532720 675536 532772
rect 42708 532652 42760 532704
rect 45192 532652 45244 532704
rect 671160 532516 671212 532568
rect 675484 532516 675536 532568
rect 663524 531428 663576 531480
rect 675484 531360 675536 531412
rect 667848 530068 667900 530120
rect 675484 530068 675536 530120
rect 669044 529932 669096 529984
rect 674932 529932 674984 529984
rect 42524 529048 42576 529100
rect 43260 529048 43312 529100
rect 666100 528572 666152 528624
rect 675484 528572 675536 528624
rect 673644 528436 673696 528488
rect 675484 528436 675536 528488
rect 673828 528028 673880 528080
rect 675484 528028 675536 528080
rect 670424 526804 670476 526856
rect 675484 526804 675536 526856
rect 672724 526396 672776 526448
rect 675484 526396 675536 526448
rect 673736 525784 673788 525836
rect 675484 525784 675536 525836
rect 681004 525716 681056 525768
rect 683120 525716 683172 525768
rect 43260 523676 43312 523728
rect 62764 523676 62816 523728
rect 651564 522996 651616 523048
rect 661684 522996 661736 523048
rect 42064 518916 42116 518968
rect 62120 518916 62172 518968
rect 651564 510620 651616 510672
rect 660488 510620 660540 510672
rect 52092 506472 52144 506524
rect 62120 506472 62172 506524
rect 676036 503480 676088 503532
rect 679624 503480 679676 503532
rect 676036 498244 676088 498296
rect 679808 498244 679860 498296
rect 651564 496816 651616 496868
rect 659108 496816 659160 496868
rect 43628 491920 43680 491972
rect 62120 491920 62172 491972
rect 664444 491580 664496 491632
rect 675300 491580 675352 491632
rect 660304 491444 660356 491496
rect 675484 491444 675536 491496
rect 659292 491308 659344 491360
rect 675484 491308 675536 491360
rect 676220 490152 676272 490204
rect 677416 490152 677468 490204
rect 673000 490016 673052 490068
rect 675484 490016 675536 490068
rect 672540 488656 672592 488708
rect 675484 488656 675536 488708
rect 676220 488520 676272 488572
rect 677232 488520 677284 488572
rect 666376 485936 666428 485988
rect 675484 485936 675536 485988
rect 663708 485800 663760 485852
rect 675300 485800 675352 485852
rect 670240 485596 670292 485648
rect 675484 485596 675536 485648
rect 651564 484440 651616 484492
rect 664812 484372 664864 484424
rect 664996 484372 665048 484424
rect 675484 484372 675536 484424
rect 673460 483556 673512 483608
rect 675484 483556 675536 483608
rect 673276 483148 673328 483200
rect 675484 483148 675536 483200
rect 671804 482740 671856 482792
rect 675484 482740 675536 482792
rect 671988 482332 672040 482384
rect 675484 482332 675536 482384
rect 674104 481856 674156 481908
rect 675484 481856 675536 481908
rect 671528 480632 671580 480684
rect 675484 480632 675536 480684
rect 47952 480224 48004 480276
rect 62120 480224 62172 480276
rect 651564 470568 651616 470620
rect 661868 470568 661920 470620
rect 49332 466420 49384 466472
rect 62120 466420 62172 466472
rect 651564 456764 651616 456816
rect 663248 456764 663300 456816
rect 55036 454044 55088 454096
rect 62120 454044 62172 454096
rect 651564 444456 651616 444508
rect 660672 444388 660724 444440
rect 50712 440240 50764 440292
rect 62120 440240 62172 440292
rect 651564 430584 651616 430636
rect 660304 430584 660356 430636
rect 41328 429564 41380 429616
rect 41696 429564 41748 429616
rect 41328 429428 41380 429480
rect 41696 429428 41748 429480
rect 42064 429428 42116 429480
rect 43260 429428 43312 429480
rect 41144 429292 41196 429344
rect 41696 429292 41748 429344
rect 42064 429292 42116 429344
rect 43444 429292 43496 429344
rect 40960 429156 41012 429208
rect 41696 429156 41748 429208
rect 42064 429156 42116 429208
rect 44548 429156 44600 429208
rect 42064 428408 42116 428460
rect 42892 428408 42944 428460
rect 41696 428000 41748 428052
rect 41328 427932 41380 427984
rect 41144 427796 41196 427848
rect 41696 427796 41748 427848
rect 42064 427796 42116 427848
rect 44272 427796 44324 427848
rect 46572 427796 46624 427848
rect 62120 427796 62172 427848
rect 41144 426572 41196 426624
rect 41696 426640 41748 426692
rect 42064 426640 42116 426692
rect 43812 426640 43864 426692
rect 40960 426436 41012 426488
rect 41696 426436 41748 426488
rect 42064 426436 42116 426488
rect 44272 426436 44324 426488
rect 41328 424328 41380 424380
rect 41696 424328 41748 424380
rect 42432 419500 42484 419552
rect 51908 419500 51960 419552
rect 45744 418140 45796 418192
rect 54668 418140 54720 418192
rect 651564 416780 651616 416832
rect 664444 416780 664496 416832
rect 56232 415420 56284 415472
rect 62120 415420 62172 415472
rect 42248 409776 42300 409828
rect 43444 409776 43496 409828
rect 42432 408416 42484 408468
rect 54852 408416 54904 408468
rect 42432 408280 42484 408332
rect 45376 408280 45428 408332
rect 42432 407056 42484 407108
rect 43076 407056 43128 407108
rect 42340 405968 42392 406020
rect 45560 405968 45612 406020
rect 651564 404336 651616 404388
rect 659292 404336 659344 404388
rect 669320 403384 669372 403436
rect 675300 403384 675352 403436
rect 663064 403248 663116 403300
rect 675484 403248 675536 403300
rect 661684 403112 661736 403164
rect 675484 403044 675536 403096
rect 658924 402976 658976 403028
rect 42248 402908 42300 402960
rect 43812 402908 43864 402960
rect 669320 402908 669372 402960
rect 42432 402500 42484 402552
rect 45192 402500 45244 402552
rect 43444 401616 43496 401668
rect 62120 401616 62172 401668
rect 672816 400528 672868 400580
rect 675484 400528 675536 400580
rect 42432 400120 42484 400172
rect 43996 400120 44048 400172
rect 673184 399712 673236 399764
rect 675484 399712 675536 399764
rect 671160 397264 671212 397316
rect 675484 397264 675536 397316
rect 670424 396040 670476 396092
rect 675484 396040 675536 396092
rect 673920 395632 673972 395684
rect 675484 395632 675536 395684
rect 673368 394408 673420 394460
rect 675484 394408 675536 394460
rect 672540 394136 672592 394188
rect 672908 394136 672960 394188
rect 673000 394000 673052 394052
rect 675484 394000 675536 394052
rect 671620 392368 671672 392420
rect 675484 392368 675536 392420
rect 675852 392096 675904 392148
rect 683120 392096 683172 392148
rect 651564 390532 651616 390584
rect 661684 390532 661736 390584
rect 48136 389240 48188 389292
rect 62120 389240 62172 389292
rect 35808 387540 35860 387592
rect 41696 387540 41748 387592
rect 42064 387472 42116 387524
rect 49332 387472 49384 387524
rect 35624 386792 35676 386844
rect 39948 386792 40000 386844
rect 40132 386656 40184 386708
rect 35808 386520 35860 386572
rect 35440 386384 35492 386436
rect 41696 386452 41748 386504
rect 42064 386452 42116 386504
rect 47952 386452 48004 386504
rect 35808 385432 35860 385484
rect 40132 385432 40184 385484
rect 35532 385160 35584 385212
rect 41696 385228 41748 385280
rect 42064 385228 42116 385280
rect 42892 385228 42944 385280
rect 35348 385024 35400 385076
rect 41696 385024 41748 385076
rect 42064 385024 42116 385076
rect 45376 385024 45428 385076
rect 674932 384752 674984 384804
rect 675484 384752 675536 384804
rect 35808 384072 35860 384124
rect 39764 384072 39816 384124
rect 35624 383800 35676 383852
rect 39948 383868 40000 383920
rect 42064 383732 42116 383784
rect 44548 383732 44600 383784
rect 35808 383664 35860 383716
rect 41696 383664 41748 383716
rect 35808 382644 35860 382696
rect 41696 382644 41748 382696
rect 35624 382508 35676 382560
rect 40224 382508 40276 382560
rect 35440 382372 35492 382424
rect 40040 382372 40092 382424
rect 35256 382236 35308 382288
rect 39028 382236 39080 382288
rect 35808 381148 35860 381200
rect 41420 381148 41472 381200
rect 35624 381012 35676 381064
rect 40040 381012 40092 381064
rect 35808 379924 35860 379976
rect 41512 379924 41564 379976
rect 35624 379652 35676 379704
rect 39948 379652 40000 379704
rect 35808 379516 35860 379568
rect 39580 379516 39632 379568
rect 670424 379448 670476 379500
rect 675116 379448 675168 379500
rect 35808 378292 35860 378344
rect 41236 378292 41288 378344
rect 651564 378156 651616 378208
rect 663064 378156 663116 378208
rect 673368 377816 673420 377868
rect 675300 377816 675352 377868
rect 35624 377000 35676 377052
rect 41696 376932 41748 376984
rect 42064 376796 42116 376848
rect 35808 376728 35860 376780
rect 41696 376728 41748 376780
rect 53472 376728 53524 376780
rect 673000 376592 673052 376644
rect 675116 376592 675168 376644
rect 28816 375844 28868 375896
rect 33784 375844 33836 375896
rect 35808 375572 35860 375624
rect 41696 375572 41748 375624
rect 42064 375504 42116 375556
rect 52276 375504 52328 375556
rect 49332 375368 49384 375420
rect 62120 375368 62172 375420
rect 33784 373260 33836 373312
rect 41696 373260 41748 373312
rect 672816 372512 672868 372564
rect 675300 372512 675352 372564
rect 32404 371832 32456 371884
rect 41696 371832 41748 371884
rect 42064 371696 42116 371748
rect 42616 371696 42668 371748
rect 42248 365644 42300 365696
rect 45192 365644 45244 365696
rect 651564 364352 651616 364404
rect 664628 364352 664680 364404
rect 42340 364216 42392 364268
rect 52092 364216 52144 364268
rect 42340 364080 42392 364132
rect 43812 364080 43864 364132
rect 42432 360136 42484 360188
rect 44364 360136 44416 360188
rect 42156 359932 42208 359984
rect 43260 359932 43312 359984
rect 659108 357688 659160 357740
rect 675300 357824 675352 357876
rect 664812 357552 664864 357604
rect 675484 357552 675536 357604
rect 660488 357416 660540 357468
rect 675116 357416 675168 357468
rect 673920 357008 673972 357060
rect 675484 357008 675536 357060
rect 50896 356668 50948 356720
rect 62120 356668 62172 356720
rect 42432 355988 42484 356040
rect 42984 355988 43036 356040
rect 672448 355852 672500 355904
rect 675484 355852 675536 355904
rect 672448 355376 672500 355428
rect 675484 355376 675536 355428
rect 673184 355036 673236 355088
rect 675484 355036 675536 355088
rect 673184 354560 673236 354612
rect 675484 354560 675536 354612
rect 667848 353608 667900 353660
rect 675484 353608 675536 353660
rect 671804 353336 671856 353388
rect 675484 353336 675536 353388
rect 670424 352520 670476 352572
rect 675484 352520 675536 352572
rect 673368 350072 673420 350124
rect 675484 350072 675536 350124
rect 673552 349664 673604 349716
rect 675484 349664 675536 349716
rect 669780 349256 669832 349308
rect 675484 349256 675536 349308
rect 673000 348848 673052 348900
rect 675484 348848 675536 348900
rect 671160 348440 671212 348492
rect 675484 348440 675536 348492
rect 675852 347896 675904 347948
rect 676588 347896 676640 347948
rect 672356 347216 672408 347268
rect 675484 347216 675536 347268
rect 45192 347012 45244 347064
rect 62120 347012 62172 347064
rect 675852 346400 675904 346452
rect 683120 346400 683172 346452
rect 35808 344020 35860 344072
rect 39212 344020 39264 344072
rect 35808 343748 35860 343800
rect 41696 343816 41748 343868
rect 42064 343816 42116 343868
rect 50712 343816 50764 343868
rect 35624 343612 35676 343664
rect 41696 343612 41748 343664
rect 42064 343612 42116 343664
rect 56232 343612 56284 343664
rect 35808 342660 35860 342712
rect 40316 342660 40368 342712
rect 35624 342388 35676 342440
rect 40040 342388 40092 342440
rect 35624 342252 35676 342304
rect 41696 342252 41748 342304
rect 42064 342252 42116 342304
rect 44640 342252 44692 342304
rect 35808 341436 35860 341488
rect 41696 341436 41748 341488
rect 42064 341368 42116 341420
rect 42892 341368 42944 341420
rect 35348 341164 35400 341216
rect 41696 341232 41748 341284
rect 42064 341232 42116 341284
rect 42708 341232 42760 341284
rect 35808 341028 35860 341080
rect 41696 341028 41748 341080
rect 42064 341028 42116 341080
rect 43628 341028 43680 341080
rect 35624 340892 35676 340944
rect 41696 340892 41748 340944
rect 42064 340892 42116 340944
rect 44456 340892 44508 340944
rect 35808 339600 35860 339652
rect 41420 339600 41472 339652
rect 35808 338376 35860 338428
rect 41696 338376 41748 338428
rect 35624 338104 35676 338156
rect 41512 338104 41564 338156
rect 652208 338104 652260 338156
rect 667388 338104 667440 338156
rect 671804 338036 671856 338088
rect 675116 338036 675168 338088
rect 674472 337900 674524 337952
rect 675116 337900 675168 337952
rect 35808 337084 35860 337136
rect 39856 337084 39908 337136
rect 35808 336880 35860 336932
rect 40316 336880 40368 336932
rect 35532 336744 35584 336796
rect 41696 336744 41748 336796
rect 42064 336744 42116 336796
rect 43628 336744 43680 336796
rect 46572 336744 46624 336796
rect 62120 336744 62172 336796
rect 673368 335996 673420 336048
rect 674932 335996 674984 336048
rect 673552 335860 673604 335912
rect 675392 335860 675444 335912
rect 35808 335588 35860 335640
rect 40868 335588 40920 335640
rect 35624 335316 35676 335368
rect 40224 335316 40276 335368
rect 35624 334364 35676 334416
rect 40316 334364 40368 334416
rect 35440 334092 35492 334144
rect 40132 334092 40184 334144
rect 35808 333956 35860 334008
rect 41696 333956 41748 334008
rect 42064 333956 42116 334008
rect 50712 333956 50764 334008
rect 670424 333888 670476 333940
rect 675116 333888 675168 333940
rect 35808 333004 35860 333056
rect 39304 332868 39356 332920
rect 35808 332596 35860 332648
rect 41696 332596 41748 332648
rect 42064 332596 42116 332648
rect 56232 332596 56284 332648
rect 669780 332596 669832 332648
rect 675116 332596 675168 332648
rect 673000 331712 673052 331764
rect 675116 331712 675168 331764
rect 42432 327020 42484 327072
rect 45836 327020 45888 327072
rect 670240 325592 670292 325644
rect 675116 325592 675168 325644
rect 667848 325456 667900 325508
rect 674932 325456 674984 325508
rect 42432 325320 42484 325372
rect 44640 325320 44692 325372
rect 651564 324300 651616 324352
rect 673552 324300 673604 324352
rect 42432 321512 42484 321564
rect 55036 321512 55088 321564
rect 42432 321240 42484 321292
rect 43996 321240 44048 321292
rect 42248 319948 42300 320000
rect 45376 319948 45428 320000
rect 42432 319132 42484 319184
rect 46020 319132 46072 319184
rect 42616 318724 42668 318776
rect 46756 318724 46808 318776
rect 42432 317364 42484 317416
rect 43076 317364 43128 317416
rect 42432 316888 42484 316940
rect 43812 316888 43864 316940
rect 42432 315868 42484 315920
rect 43628 315868 43680 315920
rect 43812 313896 43864 313948
rect 62764 313896 62816 313948
rect 663248 313420 663300 313472
rect 675484 313420 675536 313472
rect 661868 313284 661920 313336
rect 675484 313284 675536 313336
rect 673920 312468 673972 312520
rect 675484 312468 675536 312520
rect 660672 311992 660724 312044
rect 675300 311992 675352 312044
rect 664260 311856 664312 311908
rect 675484 311856 675536 311908
rect 666376 310700 666428 310752
rect 675484 310700 675536 310752
rect 651564 310496 651616 310548
rect 667204 310496 667256 310548
rect 42432 310428 42484 310480
rect 45560 310428 45612 310480
rect 670424 310360 670476 310412
rect 675484 310360 675536 310412
rect 673184 310020 673236 310072
rect 675484 310020 675536 310072
rect 664996 309136 665048 309188
rect 675484 309136 675536 309188
rect 673276 305464 673328 305516
rect 675484 305464 675536 305516
rect 673092 303832 673144 303884
rect 675484 303832 675536 303884
rect 672816 303424 672868 303476
rect 675484 303424 675536 303476
rect 670240 302200 670292 302252
rect 675484 302200 675536 302252
rect 680360 302200 680412 302252
rect 683120 302200 683172 302252
rect 43628 301248 43680 301300
rect 50896 301248 50948 301300
rect 43076 300976 43128 301028
rect 49332 300976 49384 301028
rect 41144 299616 41196 299668
rect 41696 299684 41748 299736
rect 42064 299684 42116 299736
rect 43260 299684 43312 299736
rect 40960 299480 41012 299532
rect 41696 299480 41748 299532
rect 42064 299480 42116 299532
rect 48136 299480 48188 299532
rect 40960 298256 41012 298308
rect 41144 298256 41196 298308
rect 41696 298324 41748 298376
rect 42064 298324 42116 298376
rect 42892 298324 42944 298376
rect 42064 298188 42116 298240
rect 44456 298188 44508 298240
rect 41696 298120 41748 298172
rect 49332 298120 49384 298172
rect 62120 298120 62172 298172
rect 41144 296828 41196 296880
rect 41696 296896 41748 296948
rect 42064 296896 42116 296948
rect 44180 296896 44232 296948
rect 675852 296896 675904 296948
rect 681004 296896 681056 296948
rect 40960 296692 41012 296744
rect 41696 296692 41748 296744
rect 42064 296692 42116 296744
rect 44548 296692 44600 296744
rect 675484 296352 675536 296404
rect 675484 295876 675536 295928
rect 41328 293972 41380 294024
rect 41696 293972 41748 294024
rect 42064 293972 42116 294024
rect 47216 293972 47268 294024
rect 40500 292544 40552 292596
rect 41604 292544 41656 292596
rect 674472 292272 674524 292324
rect 675116 292272 675168 292324
rect 41144 291184 41196 291236
rect 41696 291184 41748 291236
rect 42064 291184 42116 291236
rect 43996 291184 44048 291236
rect 43628 290300 43680 290352
rect 49516 290300 49568 290352
rect 42064 290028 42116 290080
rect 60004 289960 60056 290012
rect 40960 289824 41012 289876
rect 41696 289824 41748 289876
rect 42064 289824 42116 289876
rect 64144 289824 64196 289876
rect 41144 289076 41196 289128
rect 41696 289076 41748 289128
rect 37924 284996 37976 285048
rect 41696 284996 41748 285048
rect 43628 284316 43680 284368
rect 62120 284316 62172 284368
rect 651564 284316 651616 284368
rect 664812 284316 664864 284368
rect 42432 281460 42484 281512
rect 43444 281460 43496 281512
rect 42432 280100 42484 280152
rect 42984 280100 43036 280152
rect 406936 278672 406988 278724
rect 499580 278672 499632 278724
rect 437204 278536 437256 278588
rect 546684 278536 546736 278588
rect 48964 278400 49016 278452
rect 644664 278400 644716 278452
rect 64144 278264 64196 278316
rect 661040 278264 661092 278316
rect 56232 278128 56284 278180
rect 658280 278128 658332 278180
rect 49516 277992 49568 278044
rect 659660 277992 659712 278044
rect 424692 277788 424744 277840
rect 527732 277788 527784 277840
rect 413744 277652 413796 277704
rect 510068 277652 510120 277704
rect 422208 277516 422260 277568
rect 524512 277516 524564 277568
rect 467656 277380 467708 277432
rect 570972 277380 571024 277432
rect 42340 277176 42392 277228
rect 44088 277176 44140 277228
rect 457444 277176 457496 277228
rect 563520 277176 563572 277228
rect 42340 277040 42392 277092
rect 43996 277040 44048 277092
rect 409420 277040 409472 277092
rect 499488 277040 499540 277092
rect 499764 277040 499816 277092
rect 509056 277040 509108 277092
rect 509240 277040 509292 277092
rect 601424 277040 601476 277092
rect 380716 276904 380768 276956
rect 457168 276904 457220 276956
rect 472992 276904 473044 276956
rect 606116 276904 606168 276956
rect 387340 276768 387392 276820
rect 467840 276768 467892 276820
rect 469036 276768 469088 276820
rect 599032 276768 599084 276820
rect 52276 276632 52328 276684
rect 655520 276632 655572 276684
rect 402428 276496 402480 276548
rect 492220 276496 492272 276548
rect 493324 276496 493376 276548
rect 499396 276496 499448 276548
rect 499534 276496 499586 276548
rect 616788 276496 616840 276548
rect 420368 276360 420420 276412
rect 521016 276360 521068 276412
rect 442908 276224 442960 276276
rect 557632 276224 557684 276276
rect 410892 276088 410944 276140
rect 110788 275952 110840 276004
rect 156696 275952 156748 276004
rect 171048 275952 171100 276004
rect 107200 275816 107252 275868
rect 153844 275816 153896 275868
rect 160468 275816 160520 275868
rect 174452 275816 174504 275868
rect 175832 275952 175884 276004
rect 177856 275952 177908 276004
rect 317144 275952 317196 276004
rect 319996 275952 320048 276004
rect 331220 275952 331272 276004
rect 340144 275952 340196 276004
rect 342260 275952 342312 276004
rect 350724 275952 350776 276004
rect 355324 275952 355376 276004
rect 369676 275952 369728 276004
rect 369952 275952 370004 276004
rect 407488 275952 407540 276004
rect 408224 275952 408276 276004
rect 436560 276088 436612 276140
rect 175924 275816 175976 275868
rect 305092 275816 305144 275868
rect 316500 275816 316552 275868
rect 317328 275816 317380 275868
rect 336556 275816 336608 275868
rect 343824 275816 343876 275868
rect 354312 275816 354364 275868
rect 356888 275816 356940 275868
rect 399208 275816 399260 275868
rect 400220 275816 400272 275868
rect 411076 275816 411128 275868
rect 421656 275952 421708 276004
rect 421840 275952 421892 276004
rect 425244 275952 425296 276004
rect 426072 275952 426124 276004
rect 436744 275952 436796 276004
rect 450728 276088 450780 276140
rect 531228 276088 531280 276140
rect 465724 275952 465776 276004
rect 465908 275952 465960 276004
rect 466644 275952 466696 276004
rect 467104 275952 467156 276004
rect 475568 275952 475620 276004
rect 475752 275952 475804 276004
rect 480168 275952 480220 276004
rect 480352 275952 480404 276004
rect 484308 275952 484360 276004
rect 485780 275952 485832 276004
rect 489736 275952 489788 276004
rect 489920 275952 489972 276004
rect 494980 275952 495032 276004
rect 495348 275952 495400 276004
rect 504364 275952 504416 276004
rect 504732 275952 504784 276004
rect 501788 275816 501840 275868
rect 501972 275816 502024 275868
rect 508688 275816 508740 275868
rect 509056 275952 509108 276004
rect 512000 275952 512052 276004
rect 512184 275952 512236 276004
rect 516232 275952 516284 276004
rect 523684 275952 523736 276004
rect 533344 275952 533396 276004
rect 616788 275952 616840 276004
rect 635648 275952 635700 276004
rect 574192 275816 574244 275868
rect 103704 275680 103756 275732
rect 160560 275680 160612 275732
rect 174636 275680 174688 275732
rect 197544 275680 197596 275732
rect 199476 275680 199528 275732
rect 210884 275680 210936 275732
rect 297272 275680 297324 275732
rect 311716 275680 311768 275732
rect 319996 275680 320048 275732
rect 343640 275680 343692 275732
rect 345388 275680 345440 275732
rect 370872 275680 370924 275732
rect 374184 275680 374236 275732
rect 393320 275680 393372 275732
rect 395436 275680 395488 275732
rect 399668 275680 399720 275732
rect 399852 275680 399904 275732
rect 400588 275680 400640 275732
rect 400772 275680 400824 275732
rect 480812 275680 480864 275732
rect 480996 275680 481048 275732
rect 487896 275680 487948 275732
rect 488080 275680 488132 275732
rect 489874 275680 489926 275732
rect 490012 275680 490064 275732
rect 604920 275680 604972 275732
rect 610072 275680 610124 275732
rect 614396 275680 614448 275732
rect 74080 275544 74132 275596
rect 77760 275544 77812 275596
rect 85948 275544 86000 275596
rect 149060 275544 149112 275596
rect 149796 275544 149848 275596
rect 179972 275544 180024 275596
rect 181720 275544 181772 275596
rect 207020 275544 207072 275596
rect 282920 275544 282972 275596
rect 285772 275544 285824 275596
rect 302516 275544 302568 275596
rect 318800 275544 318852 275596
rect 329196 275544 329248 275596
rect 374368 275544 374420 275596
rect 374644 275544 374696 275596
rect 379152 275544 379204 275596
rect 380900 275544 380952 275596
rect 386420 275544 386472 275596
rect 391572 275544 391624 275596
rect 473452 275544 473504 275596
rect 474004 275544 474056 275596
rect 475200 275544 475252 275596
rect 475384 275544 475436 275596
rect 68192 275408 68244 275460
rect 135260 275408 135312 275460
rect 136824 275408 136876 275460
rect 152740 275408 152792 275460
rect 153292 275408 153344 275460
rect 185584 275408 185636 275460
rect 188804 275408 188856 275460
rect 213920 275476 213972 275528
rect 236092 275408 236144 275460
rect 242256 275408 242308 275460
rect 285680 275408 285732 275460
rect 303436 275408 303488 275460
rect 311072 275408 311124 275460
rect 329472 275408 329524 275460
rect 333612 275408 333664 275460
rect 381544 275408 381596 275460
rect 382648 275408 382700 275460
rect 388628 275408 388680 275460
rect 210056 275340 210108 275392
rect 226432 275340 226484 275392
rect 70584 275272 70636 275324
rect 139308 275272 139360 275324
rect 152188 275272 152240 275324
rect 162584 275272 162636 275324
rect 167552 275272 167604 275324
rect 200028 275272 200080 275324
rect 227812 275272 227864 275324
rect 237380 275272 237432 275324
rect 238484 275272 238536 275324
rect 243728 275272 243780 275324
rect 265900 275272 265952 275324
rect 271512 275272 271564 275324
rect 278412 275272 278464 275324
rect 292856 275272 292908 275324
rect 295340 275272 295392 275324
rect 299940 275272 299992 275324
rect 301136 275272 301188 275324
rect 322388 275272 322440 275324
rect 322572 275272 322624 275324
rect 333060 275272 333112 275324
rect 340236 275272 340288 275324
rect 392124 275408 392176 275460
rect 396724 275408 396776 275460
rect 400404 275408 400456 275460
rect 400588 275408 400640 275460
rect 480168 275408 480220 275460
rect 480352 275408 480404 275460
rect 484860 275408 484912 275460
rect 485044 275408 485096 275460
rect 391940 275272 391992 275324
rect 396908 275272 396960 275324
rect 397460 275272 397512 275324
rect 211252 275204 211304 275256
rect 212448 275204 212500 275256
rect 113180 275136 113232 275188
rect 142988 275136 143040 275188
rect 156880 275136 156932 275188
rect 166172 275136 166224 275188
rect 245568 275136 245620 275188
rect 246304 275136 246356 275188
rect 350540 275136 350592 275188
rect 357900 275136 357952 275188
rect 365628 275136 365680 275188
rect 375564 275136 375616 275188
rect 386420 275136 386472 275188
rect 414388 275136 414440 275188
rect 415216 275272 415268 275324
rect 418344 275272 418396 275324
rect 418528 275272 418580 275324
rect 421840 275272 421892 275324
rect 422024 275272 422076 275324
rect 422944 275272 422996 275324
rect 465540 275272 465592 275324
rect 465724 275272 465776 275324
rect 475384 275272 475436 275324
rect 475568 275272 475620 275324
rect 423312 275136 423364 275188
rect 427084 275136 427136 275188
rect 427268 275136 427320 275188
rect 431132 275136 431184 275188
rect 431316 275136 431368 275188
rect 436560 275136 436612 275188
rect 436744 275136 436796 275188
rect 485044 275136 485096 275188
rect 485228 275136 485280 275188
rect 489874 275136 489926 275188
rect 494520 275136 494572 275188
rect 494980 275544 495032 275596
rect 612004 275544 612056 275596
rect 494980 275408 495032 275460
rect 498568 275408 498620 275460
rect 498752 275408 498804 275460
rect 501972 275272 502024 275324
rect 504364 275408 504416 275460
rect 640432 275408 640484 275460
rect 648528 275272 648580 275324
rect 523500 275136 523552 275188
rect 194692 275068 194744 275120
rect 195888 275068 195940 275120
rect 378784 275068 378836 275120
rect 386236 275068 386288 275120
rect 142712 275000 142764 275052
rect 169760 275000 169812 275052
rect 249064 275000 249116 275052
rect 250352 275000 250404 275052
rect 386420 275000 386472 275052
rect 414572 275000 414624 275052
rect 415492 275000 415544 275052
rect 501788 275000 501840 275052
rect 501972 275000 502024 275052
rect 537576 275136 537628 275188
rect 537760 275136 537812 275188
rect 552940 275136 552992 275188
rect 556160 275136 556212 275188
rect 565912 275136 565964 275188
rect 570972 275136 571024 275188
rect 596088 275136 596140 275188
rect 597468 275136 597520 275188
rect 610808 275136 610860 275188
rect 71780 274932 71832 274984
rect 73804 274932 73856 274984
rect 81256 274932 81308 274984
rect 86224 274932 86276 274984
rect 186412 274932 186464 274984
rect 188068 274932 188120 274984
rect 207756 274932 207808 274984
rect 208400 274932 208452 274984
rect 135628 274864 135680 274916
rect 158720 274864 158772 274916
rect 376116 274864 376168 274916
rect 403992 274864 404044 274916
rect 404176 274864 404228 274916
rect 412272 274864 412324 274916
rect 414388 274864 414440 274916
rect 418160 274864 418212 274916
rect 418344 274864 418396 274916
rect 421932 274864 421984 274916
rect 422300 274864 422352 274916
rect 214840 274796 214892 274848
rect 221740 274796 221792 274848
rect 338856 274728 338908 274780
rect 344836 274728 344888 274780
rect 353392 274728 353444 274780
rect 355508 274728 355560 274780
rect 358728 274728 358780 274780
rect 364984 274728 365036 274780
rect 365444 274728 365496 274780
rect 382648 274728 382700 274780
rect 382832 274728 382884 274780
rect 386420 274728 386472 274780
rect 388076 274728 388128 274780
rect 408684 274728 408736 274780
rect 411260 274728 411312 274780
rect 415768 274728 415820 274780
rect 417976 274728 418028 274780
rect 422668 274728 422720 274780
rect 423220 274864 423272 274916
rect 509194 274864 509246 274916
rect 509332 274864 509384 274916
rect 513932 274864 513984 274916
rect 514116 274864 514168 274916
rect 633348 275000 633400 275052
rect 531228 274864 531280 274916
rect 570696 274864 570748 274916
rect 619640 274796 619692 274848
rect 623872 274796 623924 274848
rect 523316 274728 523368 274780
rect 523500 274728 523552 274780
rect 530492 274728 530544 274780
rect 533344 274728 533396 274780
rect 549352 274728 549404 274780
rect 552848 274728 552900 274780
rect 556436 274728 556488 274780
rect 89536 274660 89588 274712
rect 92480 274660 92532 274712
rect 161572 274660 161624 274712
rect 163688 274660 163740 274712
rect 163964 274660 164016 274712
rect 167644 274660 167696 274712
rect 178132 274660 178184 274712
rect 179328 274660 179380 274712
rect 185216 274660 185268 274712
rect 186964 274660 187016 274712
rect 241980 274660 242032 274712
rect 246028 274660 246080 274712
rect 246764 274660 246816 274712
rect 248880 274660 248932 274712
rect 271144 274660 271196 274712
rect 276296 274660 276348 274712
rect 276664 274660 276716 274712
rect 278688 274660 278740 274712
rect 280712 274660 280764 274712
rect 283380 274660 283432 274712
rect 293224 274660 293276 274712
rect 294052 274660 294104 274712
rect 319628 274660 319680 274712
rect 327080 274660 327132 274712
rect 614764 274660 614816 274712
rect 616604 274660 616656 274712
rect 618904 274660 618956 274712
rect 620284 274660 620336 274712
rect 643744 274660 643796 274712
rect 645124 274660 645176 274712
rect 42248 274592 42300 274644
rect 47032 274592 47084 274644
rect 96620 274456 96672 274508
rect 119344 274592 119396 274644
rect 120264 274592 120316 274644
rect 161434 274592 161486 274644
rect 329656 274592 329708 274644
rect 365628 274592 365680 274644
rect 390284 274592 390336 274644
rect 470232 274592 470284 274644
rect 470416 274592 470468 274644
rect 475384 274592 475436 274644
rect 475568 274592 475620 274644
rect 479616 274592 479668 274644
rect 479800 274592 479852 274644
rect 597468 274592 597520 274644
rect 119068 274456 119120 274508
rect 168472 274456 168524 274508
rect 169760 274456 169812 274508
rect 185124 274456 185176 274508
rect 294604 274456 294656 274508
rect 307024 274456 307076 274508
rect 318708 274456 318760 274508
rect 350540 274456 350592 274508
rect 351828 274456 351880 274508
rect 400220 274456 400272 274508
rect 401324 274456 401376 274508
rect 489920 274456 489972 274508
rect 490104 274456 490156 274508
rect 494888 274456 494940 274508
rect 495072 274456 495124 274508
rect 497004 274456 497056 274508
rect 497188 274456 497240 274508
rect 617984 274456 618036 274508
rect 111984 274320 112036 274372
rect 164240 274320 164292 274372
rect 177856 274320 177908 274372
rect 204260 274320 204312 274372
rect 302884 274320 302936 274372
rect 317696 274320 317748 274372
rect 336556 274320 336608 274372
rect 378784 274320 378836 274372
rect 393228 274320 393280 274372
rect 476120 274320 476172 274372
rect 478604 274320 478656 274372
rect 610072 274320 610124 274372
rect 102508 274184 102560 274236
rect 157892 274184 157944 274236
rect 166356 274184 166408 274236
rect 198924 274184 198976 274236
rect 200580 274184 200632 274236
rect 213184 274184 213236 274236
rect 283932 274184 283984 274236
rect 302332 274184 302384 274236
rect 307576 274184 307628 274236
rect 331220 274184 331272 274236
rect 343548 274184 343600 274236
rect 391940 274184 391992 274236
rect 394332 274184 394384 274236
rect 475200 274184 475252 274236
rect 475384 274184 475436 274236
rect 485044 274184 485096 274236
rect 485228 274184 485280 274236
rect 489736 274184 489788 274236
rect 489920 274184 489972 274236
rect 621480 274184 621532 274236
rect 234896 274116 234948 274168
rect 239496 274116 239548 274168
rect 77576 274048 77628 274100
rect 143632 274048 143684 274100
rect 158076 274048 158128 274100
rect 193312 274048 193364 274100
rect 198280 274048 198332 274100
rect 218704 274048 218756 274100
rect 279884 274048 279936 274100
rect 295156 274048 295208 274100
rect 300124 274048 300176 274100
rect 325976 274048 326028 274100
rect 371884 274048 371936 274100
rect 395712 274048 395764 274100
rect 397276 274048 397328 274100
rect 483204 274048 483256 274100
rect 72976 273912 73028 273964
rect 140964 273912 141016 273964
rect 141516 273912 141568 273964
rect 183744 273912 183796 273964
rect 184112 273912 184164 273964
rect 206284 273912 206336 273964
rect 206560 273912 206612 273964
rect 223856 273912 223908 273964
rect 224224 273912 224276 273964
rect 234896 273912 234948 273964
rect 274364 273912 274416 273964
rect 286876 273912 286928 273964
rect 288072 273912 288124 273964
rect 309416 273912 309468 273964
rect 314476 273912 314528 273964
rect 342260 273912 342312 273964
rect 344652 273912 344704 273964
rect 396724 273912 396776 273964
rect 398748 273912 398800 273964
rect 486700 274048 486752 274100
rect 487068 274048 487120 274100
rect 485044 273912 485096 273964
rect 494520 273912 494572 273964
rect 494888 274048 494940 274100
rect 625068 274048 625120 274100
rect 628564 273912 628616 273964
rect 632704 273912 632756 273964
rect 643928 273912 643980 273964
rect 130844 273776 130896 273828
rect 176752 273776 176804 273828
rect 322756 273776 322808 273828
rect 358728 273776 358780 273828
rect 367008 273776 367060 273828
rect 435916 273776 435968 273828
rect 124956 273640 125008 273692
rect 149704 273640 149756 273692
rect 161480 273640 161532 273692
rect 169944 273640 169996 273692
rect 374368 273640 374420 273692
rect 420552 273640 420604 273692
rect 422668 273640 422720 273692
rect 446496 273776 446548 273828
rect 448152 273776 448204 273828
rect 446404 273640 446456 273692
rect 460756 273640 460808 273692
rect 461032 273776 461084 273828
rect 569500 273776 569552 273828
rect 556160 273640 556212 273692
rect 358084 273504 358136 273556
rect 389732 273504 389784 273556
rect 394792 273504 394844 273556
rect 397460 273504 397512 273556
rect 405188 273504 405240 273556
rect 494336 273504 494388 273556
rect 494520 273504 494572 273556
rect 529296 273504 529348 273556
rect 332508 273368 332560 273420
rect 374644 273368 374696 273420
rect 378968 273368 379020 273420
rect 409880 273368 409932 273420
rect 416412 273368 416464 273420
rect 515128 273368 515180 273420
rect 414664 273300 414716 273352
rect 353944 273232 353996 273284
rect 382372 273232 382424 273284
rect 385960 273232 386012 273284
rect 394792 273232 394844 273284
rect 42432 273164 42484 273216
rect 45376 273164 45428 273216
rect 127348 273164 127400 273216
rect 174636 273164 174688 273216
rect 326988 273164 327040 273216
rect 345388 273164 345440 273216
rect 394976 273164 395028 273216
rect 415676 273164 415728 273216
rect 432052 273232 432104 273284
rect 446404 273232 446456 273284
rect 431868 273164 431920 273216
rect 451004 273164 451056 273216
rect 568304 273164 568356 273216
rect 121368 273028 121420 273080
rect 171600 273028 171652 273080
rect 174452 273028 174504 273080
rect 196164 273028 196216 273080
rect 317512 273028 317564 273080
rect 343824 273028 343876 273080
rect 345480 273028 345532 273080
rect 372068 273028 372120 273080
rect 372436 273028 372488 273080
rect 443828 273028 443880 273080
rect 444012 273028 444064 273080
rect 450544 273028 450596 273080
rect 109592 272892 109644 272944
rect 163412 272892 163464 272944
rect 180800 272892 180852 272944
rect 207480 272892 207532 272944
rect 295064 272892 295116 272944
rect 302516 272892 302568 272944
rect 310060 272892 310112 272944
rect 319996 272892 320048 272944
rect 321468 272892 321520 272944
rect 361396 272892 361448 272944
rect 376576 272892 376628 272944
rect 451280 273028 451332 273080
rect 454040 273028 454092 273080
rect 458180 273028 458232 273080
rect 461400 273028 461452 273080
rect 571800 273028 571852 273080
rect 571984 273028 572036 273080
rect 608508 273028 608560 273080
rect 451096 272892 451148 272944
rect 97724 272756 97776 272808
rect 155408 272756 155460 272808
rect 168656 272756 168708 272808
rect 198740 272756 198792 272808
rect 298744 272756 298796 272808
rect 310520 272756 310572 272808
rect 324044 272756 324096 272808
rect 366088 272756 366140 272808
rect 371792 272756 371844 272808
rect 377956 272756 378008 272808
rect 378140 272756 378192 272808
rect 437388 272756 437440 272808
rect 437572 272756 437624 272808
rect 441620 272756 441672 272808
rect 442264 272756 442316 272808
rect 454040 272756 454092 272808
rect 454684 272892 454736 272944
rect 575388 272892 575440 272944
rect 564716 272756 564768 272808
rect 578884 272756 578936 272808
rect 636844 272756 636896 272808
rect 91836 272620 91888 272672
rect 152372 272620 152424 272672
rect 159272 272620 159324 272672
rect 194784 272620 194836 272672
rect 195704 272620 195756 272672
rect 217232 272620 217284 272672
rect 217416 272620 217468 272672
rect 230664 272620 230716 272672
rect 286876 272620 286928 272672
rect 305828 272620 305880 272672
rect 306288 272620 306340 272672
rect 317328 272620 317380 272672
rect 325516 272620 325568 272672
rect 368480 272620 368532 272672
rect 369768 272620 369820 272672
rect 436928 272620 436980 272672
rect 437112 272620 437164 272672
rect 455972 272620 456024 272672
rect 239680 272552 239732 272604
rect 244556 272552 244608 272604
rect 77760 272484 77812 272536
rect 142160 272484 142212 272536
rect 154488 272484 154540 272536
rect 190736 272484 190788 272536
rect 197084 272484 197136 272536
rect 218060 272484 218112 272536
rect 218336 272484 218388 272536
rect 231216 272484 231268 272536
rect 231400 272484 231452 272536
rect 239312 272484 239364 272536
rect 271696 272484 271748 272536
rect 280988 272484 281040 272536
rect 282184 272484 282236 272536
rect 297548 272484 297600 272536
rect 303436 272484 303488 272536
rect 322572 272484 322624 272536
rect 333244 272484 333296 272536
rect 371792 272484 371844 272536
rect 371976 272484 372028 272536
rect 374184 272484 374236 272536
rect 375012 272484 375064 272536
rect 378140 272484 378192 272536
rect 384304 272484 384356 272536
rect 388260 272484 388312 272536
rect 388444 272484 388496 272536
rect 454224 272484 454276 272536
rect 454408 272484 454460 272536
rect 461400 272620 461452 272672
rect 456524 272484 456576 272536
rect 578516 272620 578568 272672
rect 461768 272484 461820 272536
rect 466276 272484 466328 272536
rect 466460 272484 466512 272536
rect 582472 272484 582524 272536
rect 585784 272484 585836 272536
rect 622676 272484 622728 272536
rect 93032 272348 93084 272400
rect 137560 272348 137612 272400
rect 137928 272348 137980 272400
rect 181168 272348 181220 272400
rect 364248 272348 364300 272400
rect 424508 272348 424560 272400
rect 116676 272212 116728 272264
rect 159640 272212 159692 272264
rect 362776 272212 362828 272264
rect 405372 272212 405424 272264
rect 442264 272348 442316 272400
rect 442448 272348 442500 272400
rect 444012 272348 444064 272400
rect 444196 272348 444248 272400
rect 475660 272348 475712 272400
rect 476028 272348 476080 272400
rect 480076 272348 480128 272400
rect 480214 272348 480266 272400
rect 487620 272348 487672 272400
rect 490656 272348 490708 272400
rect 499028 272348 499080 272400
rect 499396 272348 499448 272400
rect 551560 272348 551612 272400
rect 552664 272348 552716 272400
rect 586060 272348 586112 272400
rect 340696 272076 340748 272128
rect 371976 272076 372028 272128
rect 355876 271940 355928 271992
rect 380900 272076 380952 272128
rect 382188 272076 382240 272128
rect 427084 272212 427136 272264
rect 437388 272212 437440 272264
rect 437572 272212 437624 272264
rect 447692 272212 447744 272264
rect 447876 272212 447928 272264
rect 489736 272212 489788 272264
rect 490196 272212 490248 272264
rect 561220 272212 561272 272264
rect 411904 272076 411956 272128
rect 487804 272076 487856 272128
rect 499028 272076 499080 272128
rect 499672 272076 499724 272128
rect 500224 272076 500276 272128
rect 552664 272076 552716 272128
rect 490012 272008 490064 272060
rect 498844 272008 498896 272060
rect 378784 271940 378836 271992
rect 388444 271940 388496 271992
rect 388628 271940 388680 271992
rect 394976 271940 395028 271992
rect 405372 271940 405424 271992
rect 415216 271940 415268 271992
rect 415676 271940 415728 271992
rect 427084 271940 427136 271992
rect 427728 271940 427780 271992
rect 489874 271940 489926 271992
rect 499534 271940 499586 271992
rect 532792 271940 532844 271992
rect 551560 271940 551612 271992
rect 555240 271940 555292 271992
rect 101312 271804 101364 271856
rect 157616 271804 157668 271856
rect 179144 271804 179196 271856
rect 204904 271804 204956 271856
rect 232504 271804 232556 271856
rect 233884 271804 233936 271856
rect 304908 271804 304960 271856
rect 334164 271804 334216 271856
rect 334624 271804 334676 271856
rect 349620 271804 349672 271856
rect 361304 271804 361356 271856
rect 426440 271804 426492 271856
rect 427544 271804 427596 271856
rect 531596 271804 531648 271856
rect 263416 271736 263468 271788
rect 269212 271736 269264 271788
rect 88616 271668 88668 271720
rect 145656 271668 145708 271720
rect 170128 271668 170180 271720
rect 201040 271668 201092 271720
rect 296628 271668 296680 271720
rect 301136 271668 301188 271720
rect 309048 271668 309100 271720
rect 342444 271668 342496 271720
rect 347780 271668 347832 271720
rect 363604 271668 363656 271720
rect 363788 271668 363840 271720
rect 429752 271668 429804 271720
rect 98920 271532 98972 271584
rect 156512 271532 156564 271584
rect 165160 271532 165212 271584
rect 197360 271532 197412 271584
rect 213644 271532 213696 271584
rect 228272 271532 228324 271584
rect 289636 271532 289688 271584
rect 297272 271532 297324 271584
rect 301504 271532 301556 271584
rect 314108 271532 314160 271584
rect 315948 271532 316000 271584
rect 345664 271532 345716 271584
rect 346584 271532 346636 271584
rect 352196 271600 352248 271652
rect 359464 271532 359516 271584
rect 365444 271532 365496 271584
rect 383200 271532 383252 271584
rect 388628 271532 388680 271584
rect 388812 271532 388864 271584
rect 391756 271532 391808 271584
rect 391940 271532 391992 271584
rect 435180 271668 435232 271720
rect 435364 271668 435416 271720
rect 538772 271804 538824 271856
rect 533528 271668 533580 271720
rect 551744 271668 551796 271720
rect 554044 271668 554096 271720
rect 615684 271668 615736 271720
rect 430212 271532 430264 271584
rect 440608 271532 440660 271584
rect 440976 271532 441028 271584
rect 447094 271532 447146 271584
rect 451234 271532 451286 271584
rect 451372 271532 451424 271584
rect 480260 271532 480312 271584
rect 480536 271532 480588 271584
rect 489276 271532 489328 271584
rect 489644 271532 489696 271584
rect 562416 271532 562468 271584
rect 625804 271532 625856 271584
rect 629760 271532 629812 271584
rect 92480 271396 92532 271448
rect 150440 271396 150492 271448
rect 150992 271396 151044 271448
rect 188252 271396 188304 271448
rect 201776 271396 201828 271448
rect 221004 271396 221056 271448
rect 229008 271396 229060 271448
rect 237840 271396 237892 271448
rect 268844 271396 268896 271448
rect 277492 271396 277544 271448
rect 286324 271396 286376 271448
rect 296352 271396 296404 271448
rect 300676 271396 300728 271448
rect 311072 271396 311124 271448
rect 311716 271396 311768 271448
rect 346768 271396 346820 271448
rect 350080 271396 350132 271448
rect 388076 271396 388128 271448
rect 84752 271260 84804 271312
rect 147680 271260 147732 271312
rect 155684 271260 155736 271312
rect 192208 271260 192260 271312
rect 193496 271260 193548 271312
rect 215760 271260 215812 271312
rect 221924 271260 221976 271312
rect 232504 271260 232556 271312
rect 273076 271260 273128 271312
rect 284576 271260 284628 271312
rect 285312 271260 285364 271312
rect 304632 271260 304684 271312
rect 319996 271260 320048 271312
rect 360200 271260 360252 271312
rect 370320 271260 370372 271312
rect 413468 271396 413520 271448
rect 413928 271396 413980 271448
rect 427084 271396 427136 271448
rect 430028 271396 430080 271448
rect 433432 271396 433484 271448
rect 433616 271396 433668 271448
rect 435364 271396 435416 271448
rect 439136 271396 439188 271448
rect 446680 271396 446732 271448
rect 553860 271396 553912 271448
rect 388628 271260 388680 271312
rect 461584 271260 461636 271312
rect 461768 271260 461820 271312
rect 465172 271260 465224 271312
rect 465356 271260 465408 271312
rect 480720 271260 480772 271312
rect 487620 271260 487672 271312
rect 580080 271260 580132 271312
rect 65892 271124 65944 271176
rect 136640 271124 136692 271176
rect 139124 271124 139176 271176
rect 140504 271124 140556 271176
rect 145012 271124 145064 271176
rect 184940 271124 184992 271176
rect 185584 271124 185636 271176
rect 191840 271124 191892 271176
rect 192392 271124 192444 271176
rect 215300 271124 215352 271176
rect 215944 271124 215996 271176
rect 229744 271124 229796 271176
rect 233700 271124 233752 271176
rect 240784 271124 240836 271176
rect 277308 271124 277360 271176
rect 291660 271124 291712 271176
rect 292396 271124 292448 271176
rect 315304 271124 315356 271176
rect 321284 271124 321336 271176
rect 362592 271124 362644 271176
rect 365628 271124 365680 271176
rect 424508 271124 424560 271176
rect 114284 270988 114336 271040
rect 167184 270988 167236 271040
rect 337752 270988 337804 271040
rect 359464 270988 359516 271040
rect 360108 270988 360160 271040
rect 413284 270988 413336 271040
rect 413468 270988 413520 271040
rect 430212 271124 430264 271176
rect 427084 270988 427136 271040
rect 456754 271124 456806 271176
rect 456892 271124 456944 271176
rect 466414 271124 466466 271176
rect 466552 271124 466604 271176
rect 480260 271124 480312 271176
rect 489920 271124 489972 271176
rect 594340 271124 594392 271176
rect 431776 270988 431828 271040
rect 539876 270988 539928 271040
rect 123760 270852 123812 270904
rect 172704 270852 172756 270904
rect 344192 270852 344244 270904
rect 356888 270852 356940 270904
rect 357164 270852 357216 270904
rect 417700 270852 417752 270904
rect 418160 270852 418212 270904
rect 418988 270852 419040 270904
rect 419448 270852 419500 270904
rect 509194 270852 509246 270904
rect 509424 270852 509476 270904
rect 533528 270852 533580 270904
rect 538864 270852 538916 270904
rect 597836 270852 597888 270904
rect 134432 270716 134484 270768
rect 178960 270716 179012 270768
rect 345664 270716 345716 270768
rect 353116 270716 353168 270768
rect 354588 270716 354640 270768
rect 402888 270716 402940 270768
rect 403072 270716 403124 270768
rect 403992 270716 404044 270768
rect 412916 270716 412968 270768
rect 413284 270716 413336 270768
rect 422484 270716 422536 270768
rect 424508 270716 424560 270768
rect 430028 270716 430080 270768
rect 430304 270716 430356 270768
rect 431316 270716 431368 270768
rect 432420 270716 432472 270768
rect 436100 270716 436152 270768
rect 436284 270716 436336 270768
rect 535184 270716 535236 270768
rect 142988 270580 143040 270632
rect 165712 270580 165764 270632
rect 343364 270580 343416 270632
rect 348148 270580 348200 270632
rect 353208 270580 353260 270632
rect 402796 270580 402848 270632
rect 402934 270580 402986 270632
rect 405924 270580 405976 270632
rect 489920 270580 489972 270632
rect 490104 270580 490156 270632
rect 499488 270580 499540 270632
rect 499672 270580 499724 270632
rect 639236 270580 639288 270632
rect 108948 270444 109000 270496
rect 162400 270444 162452 270496
rect 176936 270444 176988 270496
rect 78864 270308 78916 270360
rect 132592 270308 132644 270360
rect 133788 270308 133840 270360
rect 177580 270308 177632 270360
rect 179144 270444 179196 270496
rect 202144 270444 202196 270496
rect 207020 270444 207072 270496
rect 209504 270444 209556 270496
rect 221740 270444 221792 270496
rect 229376 270444 229428 270496
rect 244372 270444 244424 270496
rect 247776 270444 247828 270496
rect 250168 270444 250220 270496
rect 251456 270444 251508 270496
rect 258816 270444 258868 270496
rect 261300 270444 261352 270496
rect 292672 270444 292724 270496
rect 305092 270444 305144 270496
rect 325792 270444 325844 270496
rect 355324 270444 355376 270496
rect 367744 270444 367796 270496
rect 432420 270444 432472 270496
rect 432604 270444 432656 270496
rect 442264 270444 442316 270496
rect 442448 270444 442500 270496
rect 444932 270444 444984 270496
rect 445116 270444 445168 270496
rect 549536 270444 549588 270496
rect 205824 270308 205876 270360
rect 208400 270308 208452 270360
rect 224960 270308 225012 270360
rect 243176 270308 243228 270360
rect 247040 270308 247092 270360
rect 261024 270308 261076 270360
rect 264980 270308 265032 270360
rect 274824 270308 274876 270360
rect 278964 270308 279016 270360
rect 301964 270308 302016 270360
rect 320180 270308 320232 270360
rect 332324 270308 332376 270360
rect 379152 270308 379204 270360
rect 379336 270308 379388 270360
rect 383384 270308 383436 270360
rect 383568 270308 383620 270360
rect 388444 270308 388496 270360
rect 388628 270308 388680 270360
rect 459836 270308 459888 270360
rect 94228 270172 94280 270224
rect 153568 270172 153620 270224
rect 163688 270172 163740 270224
rect 166448 270172 166500 270224
rect 172428 270172 172480 270224
rect 179144 270172 179196 270224
rect 179512 270172 179564 270224
rect 203616 270172 203668 270224
rect 205548 270172 205600 270224
rect 223488 270172 223540 270224
rect 278872 270172 278924 270224
rect 288440 270172 288492 270224
rect 290464 270172 290516 270224
rect 311900 270172 311952 270224
rect 312820 270172 312872 270224
rect 331404 270172 331456 270224
rect 351644 270172 351696 270224
rect 359648 270172 359700 270224
rect 359832 270172 359884 270224
rect 67548 270036 67600 270088
rect 78588 270036 78640 270088
rect 80060 270036 80112 270088
rect 144460 270036 144512 270088
rect 152740 270036 152792 270088
rect 179788 270036 179840 270088
rect 183468 270036 183520 270088
rect 194508 270036 194560 270088
rect 202972 270036 203024 270088
rect 222016 270036 222068 270088
rect 226616 270036 226668 270088
rect 236736 270036 236788 270088
rect 266176 270036 266228 270088
rect 273260 270036 273312 270088
rect 276480 270036 276532 270088
rect 289820 270036 289872 270088
rect 297824 270036 297876 270088
rect 324320 270036 324372 270088
rect 334992 270036 335044 270088
rect 374460 270036 374512 270088
rect 374828 270172 374880 270224
rect 376760 270172 376812 270224
rect 376944 270172 376996 270224
rect 405740 270172 405792 270224
rect 405924 270172 405976 270224
rect 406752 270172 406804 270224
rect 407396 270172 407448 270224
rect 393688 270036 393740 270088
rect 75828 269900 75880 269952
rect 141792 269900 141844 269952
rect 143908 269900 143960 269952
rect 184480 269900 184532 269952
rect 191656 269900 191708 269952
rect 211160 269900 211212 269952
rect 212264 269900 212316 269952
rect 219440 269900 219492 269952
rect 219624 269900 219676 269952
rect 227720 269900 227772 269952
rect 230388 269900 230440 269952
rect 238944 269900 238996 269952
rect 266912 269900 266964 269952
rect 274640 269900 274692 269952
rect 275008 269900 275060 269952
rect 287060 269900 287112 269952
rect 287520 269900 287572 269952
rect 307760 269900 307812 269952
rect 310336 269900 310388 269952
rect 338856 269900 338908 269952
rect 339040 269900 339092 269952
rect 359464 269900 359516 269952
rect 359648 269900 359700 269952
rect 397644 270036 397696 270088
rect 398288 270036 398340 270088
rect 408040 270172 408092 270224
rect 408500 270172 408552 270224
rect 408776 270172 408828 270224
rect 442080 270172 442132 270224
rect 442264 270172 442316 270224
rect 469772 270308 469824 270360
rect 469956 270308 470008 270360
rect 474740 270308 474792 270360
rect 474924 270308 474976 270360
rect 599308 270308 599360 270360
rect 461768 270172 461820 270224
rect 582748 270172 582800 270224
rect 395896 269900 395948 269952
rect 407580 269900 407632 269952
rect 408592 270036 408644 270088
rect 408960 270036 409012 270088
rect 499396 270036 499448 270088
rect 499534 270036 499586 270088
rect 620284 270172 620336 270224
rect 69388 269764 69440 269816
rect 138848 269764 138900 269816
rect 140688 269764 140740 269816
rect 173532 269764 173584 269816
rect 122748 269628 122800 269680
rect 84108 269492 84160 269544
rect 126704 269492 126756 269544
rect 126888 269492 126940 269544
rect 166080 269492 166132 269544
rect 166448 269628 166500 269680
rect 195520 269764 195572 269816
rect 195888 269764 195940 269816
rect 216864 269764 216916 269816
rect 223304 269764 223356 269816
rect 234528 269764 234580 269816
rect 237196 269764 237248 269816
rect 243360 269764 243412 269816
rect 261760 269764 261812 269816
rect 263600 269764 263652 269816
rect 265440 269764 265492 269816
rect 271880 269764 271932 269816
rect 283104 269764 283156 269816
rect 300860 269764 300912 269816
rect 306104 269764 306156 269816
rect 335360 269764 335412 269816
rect 337200 269764 337252 269816
rect 383568 269764 383620 269816
rect 383752 269764 383804 269816
rect 173900 269628 173952 269680
rect 179512 269628 179564 269680
rect 179972 269628 180024 269680
rect 189632 269628 189684 269680
rect 197544 269628 197596 269680
rect 205088 269628 205140 269680
rect 271880 269628 271932 269680
rect 281540 269628 281592 269680
rect 313924 269628 313976 269680
rect 338120 269628 338172 269680
rect 341248 269628 341300 269680
rect 359280 269628 359332 269680
rect 359464 269628 359516 269680
rect 373724 269628 373776 269680
rect 171232 269492 171284 269544
rect 173532 269492 173584 269544
rect 182272 269492 182324 269544
rect 310796 269492 310848 269544
rect 327540 269492 327592 269544
rect 330208 269492 330260 269544
rect 372988 269492 373040 269544
rect 373448 269492 373500 269544
rect 397920 269628 397972 269680
rect 398472 269764 398524 269816
rect 476028 269764 476080 269816
rect 477040 269764 477092 269816
rect 480076 269764 480128 269816
rect 480536 269900 480588 269952
rect 488172 269900 488224 269952
rect 488356 269900 488408 269952
rect 494520 269900 494572 269952
rect 626540 270036 626592 270088
rect 484492 269764 484544 269816
rect 486240 269764 486292 269816
rect 620284 269900 620336 269952
rect 630680 269900 630732 269952
rect 494888 269764 494940 269816
rect 499304 269764 499356 269816
rect 499580 269764 499632 269816
rect 619640 269764 619692 269816
rect 636200 269764 636252 269816
rect 647240 269764 647292 269816
rect 407396 269628 407448 269680
rect 407580 269628 407632 269680
rect 413468 269628 413520 269680
rect 414112 269628 414164 269680
rect 509056 269628 509108 269680
rect 509240 269628 509292 269680
rect 633624 269628 633676 269680
rect 375196 269492 375248 269544
rect 384120 269492 384172 269544
rect 384488 269492 384540 269544
rect 388628 269492 388680 269544
rect 388996 269492 389048 269544
rect 390560 269492 390612 269544
rect 391296 269492 391348 269544
rect 469588 269492 469640 269544
rect 469772 269492 469824 269544
rect 481640 269492 481692 269544
rect 484308 269492 484360 269544
rect 489736 269492 489788 269544
rect 489920 269492 489972 269544
rect 590660 269492 590712 269544
rect 259736 269424 259788 269476
rect 260840 269424 260892 269476
rect 129372 269356 129424 269408
rect 175648 269356 175700 269408
rect 354772 269356 354824 269408
rect 393688 269356 393740 269408
rect 393872 269356 393924 269408
rect 398472 269356 398524 269408
rect 398932 269356 398984 269408
rect 401784 269356 401836 269408
rect 401968 269356 402020 269408
rect 264704 269288 264756 269340
rect 265900 269288 265952 269340
rect 128544 269220 128596 269272
rect 163596 269220 163648 269272
rect 166080 269220 166132 269272
rect 173440 269220 173492 269272
rect 328000 269220 328052 269272
rect 372620 269220 372672 269272
rect 372988 269220 373040 269272
rect 374276 269220 374328 269272
rect 374460 269152 374512 269204
rect 383936 269220 383988 269272
rect 388444 269220 388496 269272
rect 408454 269220 408506 269272
rect 408684 269220 408736 269272
rect 412640 269220 412692 269272
rect 413468 269356 413520 269408
rect 432604 269356 432656 269408
rect 432788 269356 432840 269408
rect 535460 269356 535512 269408
rect 423680 269220 423732 269272
rect 423864 269220 423916 269272
rect 521660 269220 521712 269272
rect 384120 269152 384172 269204
rect 384488 269152 384540 269204
rect 248328 269084 248380 269136
rect 249984 269084 250036 269136
rect 42432 269016 42484 269068
rect 45560 269016 45612 269068
rect 118608 269016 118660 269068
rect 169760 269016 169812 269068
rect 225420 269016 225472 269068
rect 226340 269016 226392 269068
rect 324320 269016 324372 269068
rect 336740 269016 336792 269068
rect 339408 269016 339460 269068
rect 358912 269016 358964 269068
rect 375840 269016 375892 269068
rect 407764 269016 407816 269068
rect 407948 269016 408000 269068
rect 104900 268880 104952 268932
rect 160192 268880 160244 268932
rect 203892 268880 203944 268932
rect 269120 268880 269172 268932
rect 276664 268880 276716 268932
rect 299296 268880 299348 268932
rect 319628 268880 319680 268932
rect 319812 268880 319864 268932
rect 345204 268880 345256 268932
rect 349344 268880 349396 268932
rect 209872 268812 209924 268864
rect 77208 268744 77260 268796
rect 104900 268744 104952 268796
rect 106280 268744 106332 268796
rect 161664 268744 161716 268796
rect 187608 268744 187660 268796
rect 208492 268744 208544 268796
rect 316960 268744 317012 268796
rect 353392 268744 353444 268796
rect 358544 268880 358596 268932
rect 369308 268880 369360 268932
rect 369492 268880 369544 268932
rect 432788 269016 432840 269068
rect 449900 269016 449952 269068
rect 453120 269016 453172 269068
rect 95424 268608 95476 268660
rect 155040 268608 155092 268660
rect 162584 268608 162636 268660
rect 190092 268608 190144 268660
rect 190368 268608 190420 268660
rect 203340 268608 203392 268660
rect 273536 268608 273588 268660
rect 282920 268608 282972 268660
rect 294880 268608 294932 268660
rect 317144 268608 317196 268660
rect 329472 268608 329524 268660
rect 340880 268608 340932 268660
rect 353760 268608 353812 268660
rect 364800 268744 364852 268796
rect 432236 268744 432288 268796
rect 441344 268880 441396 268932
rect 437020 268744 437072 268796
rect 437388 268744 437440 268796
rect 447048 268880 447100 268932
rect 452384 268880 452436 268932
rect 455604 268880 455656 268932
rect 456800 268880 456852 268932
rect 460020 268880 460072 268932
rect 461400 268880 461452 268932
rect 87144 268472 87196 268524
rect 149888 268472 149940 268524
rect 162768 268472 162820 268524
rect 196992 268472 197044 268524
rect 208860 268472 208912 268524
rect 225696 268472 225748 268524
rect 282368 268472 282420 268524
rect 295340 268472 295392 268524
rect 297088 268472 297140 268524
rect 322940 268472 322992 268524
rect 324688 268472 324740 268524
rect 359280 268472 359332 268524
rect 369952 268608 370004 268660
rect 374644 268608 374696 268660
rect 385040 268608 385092 268660
rect 388352 268608 388404 268660
rect 452660 268744 452712 268796
rect 461768 269016 461820 269068
rect 572720 269016 572772 269068
rect 461860 268880 461912 268932
rect 576860 268880 576912 268932
rect 442080 268608 442132 268660
rect 455604 268608 455656 268660
rect 461400 268608 461452 268660
rect 462136 268744 462188 268796
rect 466414 268744 466466 268796
rect 467012 268744 467064 268796
rect 583852 268744 583904 268796
rect 466276 268608 466328 268660
rect 466828 268608 466880 268660
rect 499396 268608 499448 268660
rect 499534 268608 499586 268660
rect 581000 268608 581052 268660
rect 82728 268336 82780 268388
rect 146944 268336 146996 268388
rect 148876 268336 148928 268388
rect 187884 268336 187936 268388
rect 188068 268336 188120 268388
rect 115848 268200 115900 268252
rect 166816 268200 166868 268252
rect 210884 268336 210936 268388
rect 219808 268336 219860 268388
rect 220728 268336 220780 268388
rect 233056 268336 233108 268388
rect 281632 268336 281684 268388
rect 298100 268336 298152 268388
rect 304172 268336 304224 268388
rect 329840 268336 329892 268388
rect 342168 268336 342220 268388
rect 374644 268336 374696 268388
rect 382464 268472 382516 268524
rect 455144 268472 455196 268524
rect 455328 268472 455380 268524
rect 461768 268472 461820 268524
rect 461952 268472 462004 268524
rect 480076 268472 480128 268524
rect 382832 268336 382884 268388
rect 387616 268336 387668 268388
rect 462136 268336 462188 268388
rect 462320 268336 462372 268388
rect 466552 268336 466604 268388
rect 466736 268336 466788 268388
rect 594800 268472 594852 268524
rect 601608 268472 601660 268524
rect 645860 268472 645912 268524
rect 480352 268336 480404 268388
rect 608876 268336 608928 268388
rect 210976 268200 211028 268252
rect 317696 268200 317748 268252
rect 356060 268200 356112 268252
rect 359280 268200 359332 268252
rect 367192 268200 367244 268252
rect 135260 268064 135312 268116
rect 138112 268064 138164 268116
rect 147496 268064 147548 268116
rect 186688 268064 186740 268116
rect 360384 268064 360436 268116
rect 413100 268200 413152 268252
rect 369308 268064 369360 268116
rect 407304 268064 407356 268116
rect 407764 268064 407816 268116
rect 432420 268200 432472 268252
rect 432604 268200 432656 268252
rect 442080 268200 442132 268252
rect 413468 268064 413520 268116
rect 416688 268064 416740 268116
rect 416872 268064 416924 268116
rect 437020 268064 437072 268116
rect 437204 268064 437256 268116
rect 547880 268200 547932 268252
rect 664444 268132 664496 268184
rect 675300 268132 675352 268184
rect 442448 268064 442500 268116
rect 541256 268064 541308 268116
rect 659292 267996 659344 268048
rect 668952 267996 669004 268048
rect 158720 267928 158772 267980
rect 180800 267928 180852 267980
rect 365812 267928 365864 267980
rect 347136 267792 347188 267844
rect 376116 267792 376168 267844
rect 378048 267792 378100 267844
rect 388352 267792 388404 267844
rect 390100 267792 390152 267844
rect 391940 267792 391992 267844
rect 396172 267928 396224 267980
rect 407948 267928 408000 267980
rect 411168 267928 411220 267980
rect 412916 267928 412968 267980
rect 413100 267928 413152 267980
rect 418528 267928 418580 267980
rect 422944 267928 422996 267980
rect 424876 267928 424928 267980
rect 428464 267928 428516 267980
rect 524696 267928 524748 267980
rect 404360 267792 404412 267844
rect 407304 267792 407356 267844
rect 410892 267792 410944 267844
rect 412640 267792 412692 267844
rect 415492 267792 415544 267844
rect 415676 267792 415728 267844
rect 263968 267724 264020 267776
rect 269580 267724 269632 267776
rect 42616 267656 42668 267708
rect 47216 267656 47268 267708
rect 132408 267656 132460 267708
rect 178592 267656 178644 267708
rect 213184 267656 213236 267708
rect 220544 267656 220596 267708
rect 305920 267656 305972 267708
rect 324320 267656 324372 267708
rect 333888 267656 333940 267708
rect 353944 267656 353996 267708
rect 357440 267656 357492 267708
rect 365996 267656 366048 267708
rect 100668 267520 100720 267572
rect 158720 267520 158772 267572
rect 166264 267520 166316 267572
rect 194048 267520 194100 267572
rect 203340 267520 203392 267572
rect 213184 267520 213236 267572
rect 286692 267520 286744 267572
rect 294604 267520 294656 267572
rect 295616 267520 295668 267572
rect 301964 267520 302016 267572
rect 308128 267520 308180 267572
rect 329472 267520 329524 267572
rect 342720 267520 342772 267572
rect 343548 267520 343600 267572
rect 346400 267520 346452 267572
rect 373448 267656 373500 267708
rect 373632 267656 373684 267708
rect 417700 267656 417752 267708
rect 418068 267792 418120 267844
rect 660304 267860 660356 267912
rect 675484 267996 675536 268048
rect 506480 267792 506532 267844
rect 668952 267724 669004 267776
rect 427084 267656 427136 267708
rect 432788 267656 432840 267708
rect 436008 267656 436060 267708
rect 437388 267656 437440 267708
rect 132592 267384 132644 267436
rect 145472 267384 145524 267436
rect 145656 267384 145708 267436
rect 149520 267384 149572 267436
rect 149704 267384 149756 267436
rect 174176 267384 174228 267436
rect 179328 267384 179380 267436
rect 207296 267384 207348 267436
rect 233884 267384 233936 267436
rect 240416 267384 240468 267436
rect 293408 267384 293460 267436
rect 302884 267384 302936 267436
rect 313280 267384 313332 267436
rect 334624 267384 334676 267436
rect 335360 267384 335412 267436
rect 342168 267384 342220 267436
rect 371608 267520 371660 267572
rect 371792 267520 371844 267572
rect 377128 267520 377180 267572
rect 377312 267520 377364 267572
rect 379336 267520 379388 267572
rect 379520 267520 379572 267572
rect 86224 267248 86276 267300
rect 145932 267248 145984 267300
rect 146208 267248 146260 267300
rect 187424 267248 187476 267300
rect 194508 267248 194560 267300
rect 208768 267248 208820 267300
rect 257344 267248 257396 267300
rect 259460 267248 259512 267300
rect 322112 267248 322164 267300
rect 341800 267248 341852 267300
rect 341984 267248 342036 267300
rect 355232 267248 355284 267300
rect 380532 267384 380584 267436
rect 381360 267520 381412 267572
rect 384304 267520 384356 267572
rect 384488 267520 384540 267572
rect 388168 267520 388220 267572
rect 388352 267520 388404 267572
rect 392584 267520 392636 267572
rect 392768 267520 392820 267572
rect 427360 267520 427412 267572
rect 428004 267520 428056 267572
rect 471060 267520 471112 267572
rect 471428 267656 471480 267708
rect 538864 267656 538916 267708
rect 675484 267792 675536 267844
rect 490472 267520 490524 267572
rect 490656 267520 490708 267572
rect 494152 267520 494204 267572
rect 494520 267520 494572 267572
rect 585784 267520 585836 267572
rect 391756 267384 391808 267436
rect 392032 267384 392084 267436
rect 393228 267384 393280 267436
rect 393412 267384 393464 267436
rect 464712 267384 464764 267436
rect 466828 267384 466880 267436
rect 480168 267384 480220 267436
rect 480352 267384 480404 267436
rect 483112 267384 483164 267436
rect 483296 267384 483348 267436
rect 489736 267384 489788 267436
rect 490196 267384 490248 267436
rect 625804 267384 625856 267436
rect 370504 267248 370556 267300
rect 390100 267248 390152 267300
rect 390468 267248 390520 267300
rect 398472 267248 398524 267300
rect 401968 267248 402020 267300
rect 402980 267248 403032 267300
rect 91008 267112 91060 267164
rect 146760 267112 146812 267164
rect 149520 267112 149572 267164
rect 151360 267112 151412 267164
rect 167644 267112 167696 267164
rect 198464 267112 198516 267164
rect 209872 267112 209924 267164
rect 222752 267112 222804 267164
rect 227720 267112 227772 267164
rect 232320 267112 232372 267164
rect 267648 267112 267700 267164
rect 271144 267112 271196 267164
rect 272064 267112 272116 267164
rect 280712 267112 280764 267164
rect 291200 267112 291252 267164
rect 301504 267112 301556 267164
rect 302240 267112 302292 267164
rect 312820 267112 312872 267164
rect 313004 267112 313056 267164
rect 343364 267112 343416 267164
rect 350816 267112 350868 267164
rect 73804 266976 73856 267028
rect 140320 266976 140372 267028
rect 140504 266976 140556 267028
rect 183008 266976 183060 267028
rect 186964 266976 187016 267028
rect 211712 266976 211764 267028
rect 212448 266976 212500 267028
rect 104900 266840 104952 266892
rect 143264 266840 143316 266892
rect 146760 266840 146812 266892
rect 152096 266840 152148 266892
rect 153844 266840 153896 266892
rect 163136 266840 163188 266892
rect 163688 266840 163740 266892
rect 176384 266840 176436 266892
rect 119344 266704 119396 266756
rect 156236 266704 156288 266756
rect 156788 266704 156840 266756
rect 165344 266704 165396 266756
rect 175924 266704 175976 266756
rect 202880 266840 202932 266892
rect 226340 266976 226392 267028
rect 236000 266976 236052 267028
rect 278688 266976 278740 267028
rect 293224 266976 293276 267028
rect 300400 266976 300452 267028
rect 310796 266976 310848 267028
rect 314752 266976 314804 267028
rect 340052 266976 340104 267028
rect 227168 266840 227220 266892
rect 256516 266840 256568 266892
rect 258080 266840 258132 266892
rect 262864 266840 262916 266892
rect 267924 266840 267976 266892
rect 275744 266840 275796 266892
rect 278872 266840 278924 266892
rect 288992 266840 289044 266892
rect 298744 266840 298796 266892
rect 311072 266840 311124 266892
rect 319812 266840 319864 266892
rect 327264 266840 327316 266892
rect 333428 266840 333480 266892
rect 338304 266840 338356 266892
rect 341800 266976 341852 267028
rect 347780 266976 347832 267028
rect 348608 266976 348660 267028
rect 358084 266840 358136 266892
rect 359648 266840 359700 266892
rect 362960 266840 363012 266892
rect 365996 266976 366048 267028
rect 371424 267112 371476 267164
rect 396172 267112 396224 267164
rect 369124 266840 369176 266892
rect 378968 266976 379020 267028
rect 379704 266976 379756 267028
rect 413008 266976 413060 267028
rect 319168 266704 319220 266756
rect 339408 266704 339460 266756
rect 340052 266704 340104 266756
rect 206284 266636 206336 266688
rect 210240 266636 210292 266688
rect 126704 266568 126756 266620
rect 148416 266568 148468 266620
rect 159640 266568 159692 266620
rect 168288 266568 168340 266620
rect 246304 266568 246356 266620
rect 248512 266568 248564 266620
rect 333428 266568 333480 266620
rect 343456 266704 343508 266756
rect 351644 266704 351696 266756
rect 353024 266704 353076 266756
rect 369308 266704 369360 266756
rect 370688 266840 370740 266892
rect 412824 266840 412876 266892
rect 417056 267248 417108 267300
rect 417884 267248 417936 267300
rect 418068 267248 418120 267300
rect 413468 267180 413520 267232
rect 416872 267180 416924 267232
rect 466184 267112 466236 267164
rect 417240 266976 417292 267028
rect 421748 266976 421800 267028
rect 426900 266976 426952 267028
rect 427084 266976 427136 267028
rect 466184 266976 466236 267028
rect 469680 267248 469732 267300
rect 470508 267248 470560 267300
rect 471060 267248 471112 267300
rect 476304 267248 476356 267300
rect 476488 267248 476540 267300
rect 543740 267248 543792 267300
rect 467012 267112 467064 267164
rect 487804 267112 487856 267164
rect 489920 267112 489972 267164
rect 491208 267112 491260 267164
rect 491392 267112 491444 267164
rect 494704 267112 494756 267164
rect 494888 267112 494940 267164
rect 497648 267112 497700 267164
rect 499534 267112 499586 267164
rect 632704 267112 632756 267164
rect 479524 266976 479576 267028
rect 479708 266976 479760 267028
rect 554044 266976 554096 267028
rect 422392 266840 422444 266892
rect 514024 266840 514076 266892
rect 514208 266840 514260 266892
rect 525892 266840 525944 266892
rect 374092 266704 374144 266756
rect 375104 266704 375156 266756
rect 379704 266704 379756 266756
rect 380992 266704 381044 266756
rect 382188 266704 382240 266756
rect 385408 266704 385460 266756
rect 388812 266704 388864 266756
rect 390560 266704 390612 266756
rect 391572 266704 391624 266756
rect 391756 266704 391808 266756
rect 424968 266704 425020 266756
rect 425152 266704 425204 266756
rect 426256 266704 426308 266756
rect 426624 266704 426676 266756
rect 427544 266704 427596 266756
rect 427912 266704 427964 266756
rect 432788 266704 432840 266756
rect 433248 266704 433300 266756
rect 437388 266704 437440 266756
rect 437664 266704 437716 266756
rect 476488 266704 476540 266756
rect 478880 266704 478932 266756
rect 479708 266704 479760 266756
rect 479892 266704 479944 266756
rect 571984 266704 572036 266756
rect 666376 266636 666428 266688
rect 675484 266636 675536 266688
rect 211160 266500 211212 266552
rect 214656 266500 214708 266552
rect 241336 266500 241388 266552
rect 245568 266500 245620 266552
rect 259552 266500 259604 266552
rect 262588 266500 262640 266552
rect 269856 266500 269908 266552
rect 274824 266500 274876 266552
rect 280160 266500 280212 266552
rect 286324 266500 286376 266552
rect 301504 266500 301556 266552
rect 304172 266500 304224 266552
rect 304448 266500 304500 266552
rect 306104 266500 306156 266552
rect 330944 266500 330996 266552
rect 333244 266500 333296 266552
rect 78588 266432 78640 266484
rect 137376 266432 137428 266484
rect 137560 266432 137612 266484
rect 154304 266432 154356 266484
rect 346584 266568 346636 266620
rect 347872 266568 347924 266620
rect 365812 266568 365864 266620
rect 372896 266568 372948 266620
rect 405924 266568 405976 266620
rect 406384 266500 406436 266552
rect 417608 266500 417660 266552
rect 345480 266432 345532 266484
rect 362960 266432 363012 266484
rect 396264 266432 396316 266484
rect 157892 266364 157944 266416
rect 159456 266364 159508 266416
rect 204904 266364 204956 266416
rect 206560 266364 206612 266416
rect 208492 266364 208544 266416
rect 212448 266364 212500 266416
rect 219440 266364 219492 266416
rect 227904 266364 227956 266416
rect 232504 266364 232556 266416
rect 233792 266364 233844 266416
rect 239496 266364 239548 266416
rect 241888 266364 241940 266416
rect 251180 266364 251232 266416
rect 252192 266364 252244 266416
rect 255872 266364 255924 266416
rect 256700 266364 256752 266416
rect 258080 266364 258132 266416
rect 259736 266364 259788 266416
rect 260288 266364 260340 266416
rect 261760 266364 261812 266416
rect 262128 266364 262180 266416
rect 266360 266364 266412 266416
rect 270592 266364 270644 266416
rect 271604 266364 271656 266416
rect 280896 266364 280948 266416
rect 282184 266364 282236 266416
rect 284576 266364 284628 266416
rect 285496 266364 285548 266416
rect 286048 266364 286100 266416
rect 286876 266364 286928 266416
rect 294144 266364 294196 266416
rect 295064 266364 295116 266416
rect 298560 266364 298612 266416
rect 300124 266364 300176 266416
rect 303712 266364 303764 266416
rect 304908 266364 304960 266416
rect 305184 266364 305236 266416
rect 306288 266364 306340 266416
rect 306656 266364 306708 266416
rect 313924 266364 313976 266416
rect 316224 266364 316276 266416
rect 317328 266364 317380 266416
rect 320640 266364 320692 266416
rect 321468 266364 321520 266416
rect 331680 266364 331732 266416
rect 332508 266364 332560 266416
rect 345664 266364 345716 266416
rect 352288 266364 352340 266416
rect 353208 266364 353260 266416
rect 354772 266364 354824 266416
rect 358912 266364 358964 266416
rect 360108 266364 360160 266416
rect 361856 266364 361908 266416
rect 362776 266364 362828 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 397184 266228 397236 266280
rect 401600 266364 401652 266416
rect 402888 266364 402940 266416
rect 403072 266364 403124 266416
rect 404176 266364 404228 266416
rect 414848 266364 414900 266416
rect 417240 266364 417292 266416
rect 417424 266364 417476 266416
rect 490104 266568 490156 266620
rect 421932 266432 421984 266484
rect 465816 266432 465868 266484
rect 466920 266432 466972 266484
rect 493324 266568 493376 266620
rect 494704 266568 494756 266620
rect 513840 266568 513892 266620
rect 514024 266568 514076 266620
rect 518900 266568 518952 266620
rect 664260 266500 664312 266552
rect 675116 266500 675168 266552
rect 492864 266432 492916 266484
rect 493692 266432 493744 266484
rect 494336 266432 494388 266484
rect 495348 266432 495400 266484
rect 495808 266432 495860 266484
rect 496728 266432 496780 266484
rect 498660 266432 498712 266484
rect 499212 266432 499264 266484
rect 499396 266432 499448 266484
rect 601608 266432 601660 266484
rect 418528 266364 418580 266416
rect 419448 266364 419500 266416
rect 415676 266228 415728 266280
rect 419448 266228 419500 266280
rect 664444 266364 664496 266416
rect 675300 266364 675352 266416
rect 422392 266296 422444 266348
rect 424048 266296 424100 266348
rect 427912 266296 427964 266348
rect 435088 266296 435140 266348
rect 437664 266296 437716 266348
rect 448704 266296 448756 266348
rect 566096 266296 566148 266348
rect 382096 266160 382148 266212
rect 384120 266160 384172 266212
rect 421840 266160 421892 266212
rect 422208 266160 422260 266212
rect 442080 266160 442132 266212
rect 448888 266160 448940 266212
rect 449072 266160 449124 266212
rect 456754 266160 456806 266212
rect 456892 266160 456944 266212
rect 575664 266160 575716 266212
rect 362592 266024 362644 266076
rect 428280 266024 428332 266076
rect 447600 266024 447652 266076
rect 448336 266024 448388 266076
rect 448520 266024 448572 266076
rect 184940 265888 184992 265940
rect 185676 265888 185728 265940
rect 198740 265888 198792 265940
rect 199660 265888 199712 265940
rect 384672 265888 384724 265940
rect 461032 265888 461084 265940
rect 461768 266024 461820 266076
rect 463976 266024 464028 266076
rect 464160 266024 464212 266076
rect 591028 266024 591080 266076
rect 467380 265888 467432 265940
rect 470784 265888 470836 265940
rect 601792 265888 601844 265940
rect 670424 265820 670476 265872
rect 675300 265820 675352 265872
rect 368480 265752 368532 265804
rect 369768 265752 369820 265804
rect 389088 265752 389140 265804
rect 470600 265752 470652 265804
rect 477408 265752 477460 265804
rect 612740 265752 612792 265804
rect 404544 265616 404596 265668
rect 495624 265616 495676 265668
rect 497280 265616 497332 265668
rect 643744 265616 643796 265668
rect 669320 265548 669372 265600
rect 675484 265548 675536 265600
rect 403808 265480 403860 265532
rect 448520 265480 448572 265532
rect 444288 265344 444340 265396
rect 559288 265480 559340 265532
rect 448888 265344 448940 265396
rect 552848 265344 552900 265396
rect 417792 265208 417844 265260
rect 516416 265208 516468 265260
rect 666008 265208 666060 265260
rect 675484 265208 675536 265260
rect 439872 265072 439924 265124
rect 537760 265072 537812 265124
rect 664996 265072 665048 265124
rect 675484 265004 675536 265056
rect 437664 264936 437716 264988
rect 523684 264936 523736 264988
rect 664260 264936 664312 264988
rect 669320 264868 669372 264920
rect 435456 264732 435508 264784
rect 545120 264732 545172 264784
rect 461216 264596 461268 264648
rect 586520 264596 586572 264648
rect 471888 264460 471940 264512
rect 603080 264460 603132 264512
rect 482192 264324 482244 264376
rect 618904 264324 618956 264376
rect 51908 264188 51960 264240
rect 655704 264188 655756 264240
rect 665088 263576 665140 263628
rect 675484 263576 675536 263628
rect 673276 262896 673328 262948
rect 675484 262896 675536 262948
rect 511540 261468 511592 261520
rect 568580 261468 568632 261520
rect 671804 261264 671856 261316
rect 675484 261264 675536 261316
rect 511356 259972 511408 260024
rect 514024 259972 514076 260024
rect 669228 259700 669280 259752
rect 675484 259700 675536 259752
rect 666376 259564 666428 259616
rect 675484 259564 675536 259616
rect 666192 259428 666244 259480
rect 675300 259428 675352 259480
rect 670424 259224 670476 259276
rect 675484 259224 675536 259276
rect 672356 258408 672408 258460
rect 675484 258408 675536 258460
rect 35808 258204 35860 258256
rect 39948 258204 40000 258256
rect 35808 257116 35860 257168
rect 39580 257116 39632 257168
rect 42064 256980 42116 257032
rect 43812 256980 43864 257032
rect 35624 256844 35676 256896
rect 41696 256912 41748 256964
rect 35440 256708 35492 256760
rect 41696 256708 41748 256760
rect 42064 256708 42116 256760
rect 45192 256708 45244 256760
rect 511448 256708 511500 256760
rect 519544 256708 519596 256760
rect 675944 256708 675996 256760
rect 683120 256708 683172 256760
rect 669780 256572 669832 256624
rect 675484 256572 675536 256624
rect 35808 255688 35860 255740
rect 40408 255688 40460 255740
rect 35624 255416 35676 255468
rect 41696 255484 41748 255536
rect 42064 255484 42116 255536
rect 42800 255484 42852 255536
rect 35440 255280 35492 255332
rect 41696 255280 41748 255332
rect 42064 255280 42116 255332
rect 45008 255280 45060 255332
rect 35808 254532 35860 254584
rect 39764 254532 39816 254584
rect 35808 254260 35860 254312
rect 40040 254260 40092 254312
rect 35624 254124 35676 254176
rect 41236 254056 41288 254108
rect 35440 253920 35492 253972
rect 41696 253920 41748 253972
rect 42064 253920 42116 253972
rect 44548 253920 44600 253972
rect 35808 252696 35860 252748
rect 41696 252696 41748 252748
rect 35532 252560 35584 252612
rect 40040 252560 40092 252612
rect 511908 252560 511960 252612
rect 562324 252560 562376 252612
rect 35808 251472 35860 251524
rect 41512 251472 41564 251524
rect 35532 251200 35584 251252
rect 41696 251200 41748 251252
rect 35808 250180 35860 250232
rect 39396 250180 39448 250232
rect 35440 249908 35492 249960
rect 39856 249908 39908 249960
rect 35624 249772 35676 249824
rect 41696 249772 41748 249824
rect 42064 249772 42116 249824
rect 47216 249772 47268 249824
rect 510620 249772 510672 249824
rect 513288 249772 513340 249824
rect 40040 249500 40092 249552
rect 41696 249500 41748 249552
rect 42064 249432 42116 249484
rect 42616 249432 42668 249484
rect 511172 249024 511224 249076
rect 571340 249024 571392 249076
rect 35808 248820 35860 248872
rect 40132 248820 40184 248872
rect 35440 248548 35492 248600
rect 39120 248548 39172 248600
rect 35624 248412 35676 248464
rect 41696 248412 41748 248464
rect 42064 248412 42116 248464
rect 44364 248412 44416 248464
rect 35808 247460 35860 247512
rect 40408 247460 40460 247512
rect 35624 247188 35676 247240
rect 41696 247188 41748 247240
rect 42064 247188 42116 247240
rect 129004 247188 129056 247240
rect 35808 247052 35860 247104
rect 41696 247052 41748 247104
rect 42064 247052 42116 247104
rect 128820 247052 128872 247104
rect 674472 246984 674524 247036
rect 674840 246984 674892 247036
rect 513288 246304 513340 246356
rect 569960 246304 570012 246356
rect 669412 245148 669464 245200
rect 675392 245148 675444 245200
rect 666192 242836 666244 242888
rect 669412 242836 669464 242888
rect 670424 242836 670476 242888
rect 675116 242836 675168 242888
rect 511264 242292 511316 242344
rect 628564 242292 628616 242344
rect 31024 242156 31076 242208
rect 41696 242156 41748 242208
rect 512000 242156 512052 242208
rect 633440 242156 633492 242208
rect 669228 241680 669280 241732
rect 675116 241680 675168 241732
rect 674656 241408 674708 241460
rect 675116 241408 675168 241460
rect 519544 240728 519596 240780
rect 567200 240728 567252 240780
rect 44180 239912 44232 239964
rect 44640 239912 44692 239964
rect 514024 238144 514076 238196
rect 568764 238144 568816 238196
rect 511264 238008 511316 238060
rect 632704 238008 632756 238060
rect 666376 237328 666428 237380
rect 675300 237328 675352 237380
rect 42432 235900 42484 235952
rect 44640 235900 44692 235952
rect 42432 234540 42484 234592
rect 43812 234540 43864 234592
rect 42432 234200 42484 234252
rect 42984 234200 43036 234252
rect 510896 233996 510948 234048
rect 577504 233996 577556 234048
rect 510712 233860 510764 233912
rect 629944 233860 629996 233912
rect 42432 231820 42484 231872
rect 47032 231820 47084 231872
rect 55864 231752 55916 231804
rect 646044 231752 646096 231804
rect 42432 231684 42484 231736
rect 44364 231684 44416 231736
rect 46204 231616 46256 231668
rect 643100 231616 643152 231668
rect 51724 231480 51776 231532
rect 650552 231480 650604 231532
rect 47584 231344 47636 231396
rect 645860 231344 645912 231396
rect 44824 231208 44876 231260
rect 644480 231208 644532 231260
rect 50528 231072 50580 231124
rect 652760 231072 652812 231124
rect 53104 230936 53156 230988
rect 641812 230936 641864 230988
rect 132592 230800 132644 230852
rect 661316 230800 661368 230852
rect 108948 230732 109000 230784
rect 117044 230732 117096 230784
rect 117228 230732 117280 230784
rect 132408 230732 132460 230784
rect 181260 230664 181312 230716
rect 183100 230664 183152 230716
rect 474648 230664 474700 230716
rect 478052 230664 478104 230716
rect 481272 230664 481324 230716
rect 507492 230664 507544 230716
rect 89628 230596 89680 230648
rect 171232 230596 171284 230648
rect 79968 230460 80020 230512
rect 116860 230460 116912 230512
rect 117044 230460 117096 230512
rect 184480 230528 184532 230580
rect 42156 230392 42208 230444
rect 43168 230392 43220 230444
rect 176844 230392 176896 230444
rect 181260 230392 181312 230444
rect 181444 230392 181496 230444
rect 189172 230528 189224 230580
rect 191748 230528 191800 230580
rect 193588 230528 193640 230580
rect 204720 230528 204772 230580
rect 187424 230392 187476 230444
rect 190276 230392 190328 230444
rect 190460 230392 190512 230444
rect 107568 230256 107620 230308
rect 182824 230256 182876 230308
rect 183468 230256 183520 230308
rect 203248 230256 203300 230308
rect 82912 230120 82964 230172
rect 153752 230120 153804 230172
rect 153936 230120 153988 230172
rect 156328 230120 156380 230172
rect 88248 229984 88300 230036
rect 166816 230120 166868 230172
rect 167000 230120 167052 230172
rect 204720 230120 204772 230172
rect 205456 230392 205508 230444
rect 206008 230392 206060 230444
rect 244648 230392 244700 230444
rect 256332 230392 256384 230444
rect 279976 230392 280028 230444
rect 290464 230392 290516 230444
rect 295432 230392 295484 230444
rect 388168 230392 388220 230444
rect 390744 230392 390796 230444
rect 284944 230324 284996 230376
rect 286600 230324 286652 230376
rect 296720 230324 296772 230376
rect 299296 230324 299348 230376
rect 300492 230324 300544 230376
rect 301504 230324 301556 230376
rect 319444 230324 319496 230376
rect 320272 230324 320324 230376
rect 331864 230324 331916 230376
rect 333060 230324 333112 230376
rect 333520 230324 333572 230376
rect 334532 230324 334584 230376
rect 339592 230324 339644 230376
rect 340972 230324 341024 230376
rect 353392 230324 353444 230376
rect 354588 230324 354640 230376
rect 355048 230324 355100 230376
rect 356704 230324 356756 230376
rect 359464 230324 359516 230376
rect 361488 230324 361540 230376
rect 364432 230324 364484 230376
rect 365628 230324 365680 230376
rect 371608 230324 371660 230376
rect 373632 230324 373684 230376
rect 376576 230324 376628 230376
rect 377864 230324 377916 230376
rect 378232 230324 378284 230376
rect 379152 230324 379204 230376
rect 391480 230324 391532 230376
rect 392584 230324 392636 230376
rect 395896 230324 395948 230376
rect 396724 230324 396776 230376
rect 205088 230256 205140 230308
rect 240232 230256 240284 230308
rect 247776 230256 247828 230308
rect 275560 230256 275612 230308
rect 380992 230256 381044 230308
rect 389088 230256 389140 230308
rect 338028 230188 338080 230240
rect 341432 230188 341484 230240
rect 341800 230188 341852 230240
rect 343732 230188 343784 230240
rect 345664 230188 345716 230240
rect 349712 230188 349764 230240
rect 357256 230188 357308 230240
rect 359740 230188 359792 230240
rect 369400 230188 369452 230240
rect 371884 230188 371936 230240
rect 235816 230120 235868 230172
rect 236000 230120 236052 230172
rect 238576 230120 238628 230172
rect 240968 230120 241020 230172
rect 271144 230120 271196 230172
rect 279884 230120 279936 230172
rect 297640 230120 297692 230172
rect 335728 230120 335780 230172
rect 337292 230120 337344 230172
rect 361120 230120 361172 230172
rect 363972 230120 364024 230172
rect 374920 230120 374972 230172
rect 381176 230120 381228 230172
rect 298744 230052 298796 230104
rect 299848 230052 299900 230104
rect 338488 230052 338540 230104
rect 342720 230052 342772 230104
rect 383200 230052 383252 230104
rect 390008 230052 390060 230104
rect 390376 230052 390428 230104
rect 394056 230188 394108 230240
rect 394240 230188 394292 230240
rect 397184 230188 397236 230240
rect 159732 229984 159784 230036
rect 168840 229984 168892 230036
rect 169024 229984 169076 230036
rect 170128 229984 170180 230036
rect 171140 229984 171192 230036
rect 174544 229984 174596 230036
rect 175004 229984 175056 230036
rect 191748 229984 191800 230036
rect 192116 229984 192168 230036
rect 193312 229984 193364 230036
rect 195244 229984 195296 230036
rect 231400 229984 231452 230036
rect 243544 229984 243596 230036
rect 266728 229984 266780 230036
rect 275652 229984 275704 230036
rect 293224 229984 293276 230036
rect 305644 229984 305696 230036
rect 313096 229984 313148 230036
rect 344008 229984 344060 230036
rect 348240 229984 348292 230036
rect 349528 229984 349580 230036
rect 356336 229984 356388 230036
rect 363328 229984 363380 230036
rect 368388 229984 368440 230036
rect 372712 229984 372764 230036
rect 382280 229984 382332 230036
rect 339040 229916 339092 229968
rect 340144 229916 340196 229968
rect 390744 229916 390796 229968
rect 397920 229984 397972 230036
rect 69664 229848 69716 229900
rect 153936 229848 153988 229900
rect 154120 229848 154172 229900
rect 66904 229712 66956 229764
rect 144644 229712 144696 229764
rect 144828 229712 144880 229764
rect 150256 229712 150308 229764
rect 150440 229712 150492 229764
rect 159732 229712 159784 229764
rect 160744 229848 160796 229900
rect 214104 229848 214156 229900
rect 214472 229848 214524 229900
rect 216496 229848 216548 229900
rect 220452 229848 220504 229900
rect 257896 229848 257948 229900
rect 267004 229848 267056 229900
rect 288808 229848 288860 229900
rect 297364 229848 297416 229900
rect 308680 229848 308732 229900
rect 308864 229848 308916 229900
rect 317512 229848 317564 229900
rect 341248 229848 341300 229900
rect 344100 229848 344152 229900
rect 358912 229848 358964 229900
rect 362408 229848 362460 229900
rect 365812 229848 365864 229900
rect 378048 229848 378100 229900
rect 389272 229848 389324 229900
rect 390468 229848 390520 229900
rect 395160 229848 395212 229900
rect 403256 230392 403308 230444
rect 408776 230392 408828 230444
rect 416044 230392 416096 230444
rect 421288 230392 421340 230444
rect 422208 230392 422260 230444
rect 422392 230392 422444 230444
rect 438032 230528 438084 230580
rect 472624 230528 472676 230580
rect 544384 230460 544436 230512
rect 403624 230324 403676 230376
rect 405004 230324 405056 230376
rect 406384 230324 406436 230376
rect 408408 230324 408460 230376
rect 414112 230256 414164 230308
rect 427728 230256 427780 230308
rect 429568 230256 429620 230308
rect 432144 230256 432196 230308
rect 432328 230256 432380 230308
rect 442264 230392 442316 230444
rect 443920 230392 443972 230444
rect 445944 230392 445996 230444
rect 447232 230392 447284 230444
rect 448060 230392 448112 230444
rect 453304 230392 453356 230444
rect 454500 230392 454552 230444
rect 456616 230392 456668 230444
rect 465816 230392 465868 230444
rect 466552 230392 466604 230444
rect 467748 230392 467800 230444
rect 476488 230392 476540 230444
rect 477408 230392 477460 230444
rect 478052 230392 478104 230444
rect 480076 230392 480128 230444
rect 480904 230324 480956 230376
rect 483296 230324 483348 230376
rect 437848 230256 437900 230308
rect 480536 230256 480588 230308
rect 483756 230256 483808 230308
rect 488080 230256 488132 230308
rect 398748 230120 398800 230172
rect 413192 230120 413244 230172
rect 420736 230120 420788 230172
rect 451464 230120 451516 230172
rect 454960 230120 455012 230172
rect 459560 230120 459612 230172
rect 463240 230120 463292 230172
rect 399208 229984 399260 230036
rect 406660 229984 406712 230036
rect 409788 229984 409840 230036
rect 427544 229984 427596 230036
rect 431868 229984 431920 230036
rect 481824 229984 481876 230036
rect 482560 230120 482612 230172
rect 542452 230256 542504 230308
rect 488448 230120 488500 230172
rect 542084 230120 542136 230172
rect 483296 229984 483348 230036
rect 484216 229984 484268 230036
rect 549904 229984 549956 230036
rect 400864 229848 400916 229900
rect 336280 229780 336332 229832
rect 339776 229780 339828 229832
rect 392216 229780 392268 229832
rect 394700 229780 394752 229832
rect 213368 229712 213420 229764
rect 213552 229712 213604 229764
rect 253480 229712 253532 229764
rect 259092 229712 259144 229764
rect 284392 229712 284444 229764
rect 293868 229712 293920 229764
rect 304264 229712 304316 229764
rect 340512 229712 340564 229764
rect 343916 229712 343968 229764
rect 361672 229712 361724 229764
rect 369584 229712 369636 229764
rect 377128 229712 377180 229764
rect 321836 229644 321888 229696
rect 323584 229644 323636 229696
rect 396448 229712 396500 229764
rect 401692 229712 401744 229764
rect 405832 229712 405884 229764
rect 409788 229712 409840 229764
rect 417240 229848 417292 229900
rect 424232 229848 424284 229900
rect 427360 229848 427412 229900
rect 432604 229848 432656 229900
rect 432880 229848 432932 229900
rect 437848 229848 437900 229900
rect 438032 229848 438084 229900
rect 441896 229848 441948 229900
rect 442264 229848 442316 229900
rect 484860 229848 484912 229900
rect 485872 229848 485924 229900
rect 558184 229848 558236 229900
rect 420920 229712 420972 229764
rect 395160 229644 395212 229696
rect 117228 229576 117280 229628
rect 181444 229576 181496 229628
rect 182088 229576 182140 229628
rect 126888 229440 126940 229492
rect 190920 229440 190972 229492
rect 191564 229576 191616 229628
rect 192760 229576 192812 229628
rect 194232 229576 194284 229628
rect 195244 229440 195296 229492
rect 195888 229576 195940 229628
rect 202788 229576 202840 229628
rect 205088 229576 205140 229628
rect 205456 229576 205508 229628
rect 209320 229576 209372 229628
rect 211712 229576 211764 229628
rect 249064 229576 249116 229628
rect 342352 229576 342404 229628
rect 343548 229576 343600 229628
rect 349068 229576 349120 229628
rect 353024 229576 353076 229628
rect 356152 229576 356204 229628
rect 363144 229576 363196 229628
rect 387708 229576 387760 229628
rect 391756 229576 391808 229628
rect 404728 229576 404780 229628
rect 408776 229576 408828 229628
rect 416872 229576 416924 229628
rect 425520 229712 425572 229764
rect 429016 229712 429068 229764
rect 430028 229712 430080 229764
rect 430212 229712 430264 229764
rect 433616 229712 433668 229764
rect 433800 229712 433852 229764
rect 436192 229712 436244 229764
rect 438032 229712 438084 229764
rect 487344 229712 487396 229764
rect 487528 229712 487580 229764
rect 565084 229712 565136 229764
rect 421840 229576 421892 229628
rect 438584 229576 438636 229628
rect 438952 229576 439004 229628
rect 287704 229508 287756 229560
rect 291016 229508 291068 229560
rect 343732 229508 343784 229560
rect 345388 229508 345440 229560
rect 394056 229508 394108 229560
rect 399484 229508 399536 229560
rect 203524 229440 203576 229492
rect 222568 229440 222620 229492
rect 227352 229440 227404 229492
rect 262312 229440 262364 229492
rect 317512 229440 317564 229492
rect 319720 229440 319772 229492
rect 384856 229440 384908 229492
rect 388444 229440 388496 229492
rect 343364 229372 343416 229424
rect 346676 229372 346728 229424
rect 378784 229372 378836 229424
rect 383936 229372 383988 229424
rect 133788 229304 133840 229356
rect 200488 229304 200540 229356
rect 140688 229168 140740 229220
rect 202604 229304 202656 229356
rect 202788 229304 202840 229356
rect 205272 229304 205324 229356
rect 205548 229304 205600 229356
rect 214288 229304 214340 229356
rect 214656 229304 214708 229356
rect 218152 229304 218204 229356
rect 200856 229168 200908 229220
rect 206008 229168 206060 229220
rect 211160 229168 211212 229220
rect 220912 229304 220964 229356
rect 222200 229304 222252 229356
rect 227536 229304 227588 229356
rect 229192 229304 229244 229356
rect 250168 229304 250220 229356
rect 320088 229304 320140 229356
rect 321376 229304 321428 229356
rect 385960 229304 386012 229356
rect 392216 229440 392268 229492
rect 403072 229440 403124 229492
rect 417240 229440 417292 229492
rect 419080 229440 419132 229492
rect 429844 229440 429896 229492
rect 430028 229440 430080 229492
rect 432420 229440 432472 229492
rect 392032 229304 392084 229356
rect 394056 229304 394108 229356
rect 413560 229304 413612 229356
rect 418804 229304 418856 229356
rect 426808 229304 426860 229356
rect 440792 229440 440844 229492
rect 441160 229576 441212 229628
rect 490380 229576 490432 229628
rect 490564 229576 490616 229628
rect 510620 229576 510672 229628
rect 494704 229440 494756 229492
rect 250444 229236 250496 229288
rect 255688 229236 255740 229288
rect 334072 229236 334124 229288
rect 335544 229236 335596 229288
rect 350632 229236 350684 229288
rect 355324 229236 355376 229288
rect 367744 229236 367796 229288
rect 220820 229168 220872 229220
rect 225328 229168 225380 229220
rect 233884 229168 233936 229220
rect 243544 229168 243596 229220
rect 109776 229032 109828 229084
rect 176844 229032 176896 229084
rect 222200 229032 222252 229084
rect 229744 229100 229796 229152
rect 321376 229100 321428 229152
rect 325792 229100 325844 229152
rect 373816 229100 373868 229152
rect 374644 229100 374696 229152
rect 99840 228896 99892 228948
rect 96528 228760 96580 228812
rect 171140 228760 171192 228812
rect 176476 228896 176528 228948
rect 233700 229032 233752 229084
rect 261760 229032 261812 229084
rect 389824 229168 389876 229220
rect 392860 229168 392912 229220
rect 410248 229168 410300 229220
rect 412732 229168 412784 229220
rect 418528 229168 418580 229220
rect 422944 229236 422996 229288
rect 424600 229168 424652 229220
rect 430212 229168 430264 229220
rect 430672 229168 430724 229220
rect 431592 229168 431644 229220
rect 432420 229168 432472 229220
rect 433800 229304 433852 229356
rect 434536 229304 434588 229356
rect 438032 229304 438084 229356
rect 438584 229304 438636 229356
rect 439596 229304 439648 229356
rect 440608 229304 440660 229356
rect 441436 229304 441488 229356
rect 444472 229304 444524 229356
rect 445668 229304 445720 229356
rect 433432 229168 433484 229220
rect 434352 229168 434404 229220
rect 435088 229168 435140 229220
rect 436008 229168 436060 229220
rect 436744 229168 436796 229220
rect 488908 229304 488960 229356
rect 490380 229304 490432 229356
rect 497464 229304 497516 229356
rect 466000 229168 466052 229220
rect 474648 229168 474700 229220
rect 474832 229168 474884 229220
rect 477224 229168 477276 229220
rect 479248 229168 479300 229220
rect 522580 229168 522632 229220
rect 382464 229032 382516 229084
rect 384304 229032 384356 229084
rect 410432 229032 410484 229084
rect 419632 228964 419684 229016
rect 442264 229032 442316 229084
rect 451280 229032 451332 229084
rect 453948 229032 454000 229084
rect 458824 229032 458876 229084
rect 524052 229032 524104 229084
rect 229008 228896 229060 228948
rect 262864 228896 262916 228948
rect 275376 228896 275428 228948
rect 293500 228896 293552 228948
rect 390928 228896 390980 228948
rect 419448 228896 419500 228948
rect 424048 228896 424100 228948
rect 457076 228896 457128 228948
rect 458272 228896 458324 228948
rect 523132 228896 523184 228948
rect 176614 228760 176666 228812
rect 179236 228760 179288 228812
rect 182364 228760 182416 228812
rect 220820 228760 220872 228812
rect 222108 228760 222160 228812
rect 258448 228760 258500 228812
rect 265440 228760 265492 228812
rect 287152 228760 287204 228812
rect 291936 228760 291988 228812
rect 304816 228760 304868 228812
rect 360568 228760 360620 228812
rect 375656 228760 375708 228812
rect 382280 228760 382332 228812
rect 390744 228760 390796 228812
rect 401968 228760 402020 228812
rect 434720 228760 434772 228812
rect 442264 228760 442316 228812
rect 451280 228760 451332 228812
rect 451648 228760 451700 228812
rect 456248 228760 456300 228812
rect 464896 228760 464948 228812
rect 532700 228760 532752 228812
rect 93216 228624 93268 228676
rect 150440 228624 150492 228676
rect 150624 228624 150676 228676
rect 178960 228624 179012 228676
rect 182180 228624 182232 228676
rect 233056 228624 233108 228676
rect 245476 228624 245528 228676
rect 273904 228624 273956 228676
rect 276296 228624 276348 228676
rect 294880 228624 294932 228676
rect 295248 228624 295300 228676
rect 307024 228624 307076 228676
rect 360016 228624 360068 228676
rect 374184 228624 374236 228676
rect 377680 228624 377732 228676
rect 400496 228624 400548 228676
rect 404176 228624 404228 228676
rect 440424 228624 440476 228676
rect 441896 228624 441948 228676
rect 468392 228624 468444 228676
rect 471888 228624 471940 228676
rect 75828 228488 75880 228540
rect 162400 228488 162452 228540
rect 166264 228488 166316 228540
rect 211160 228488 211212 228540
rect 212264 228488 212316 228540
rect 251824 228488 251876 228540
rect 253756 228488 253808 228540
rect 278872 228488 278924 228540
rect 286968 228488 287020 228540
rect 300952 228488 301004 228540
rect 347320 228488 347372 228540
rect 356152 228488 356204 228540
rect 369952 228488 370004 228540
rect 386604 228488 386656 228540
rect 393228 228488 393280 228540
rect 423956 228488 424008 228540
rect 432604 228488 432656 228540
rect 472808 228488 472860 228540
rect 473728 228488 473780 228540
rect 540336 228488 540388 228540
rect 542452 228624 542504 228676
rect 559472 228624 559524 228676
rect 542820 228488 542872 228540
rect 68928 228352 68980 228404
rect 157984 228352 158036 228404
rect 159732 228352 159784 228404
rect 214472 228352 214524 228404
rect 214932 228352 214984 228404
rect 255136 228352 255188 228404
rect 256516 228352 256568 228404
rect 281632 228352 281684 228404
rect 282000 228352 282052 228404
rect 298192 228352 298244 228404
rect 304356 228352 304408 228404
rect 314752 228352 314804 228404
rect 351184 228352 351236 228404
rect 360752 228352 360804 228404
rect 363972 228352 364024 228404
rect 373080 228352 373132 228404
rect 373264 228352 373316 228404
rect 393320 228352 393372 228404
rect 397552 228352 397604 228404
rect 430580 228352 430632 228404
rect 433616 228352 433668 228404
rect 118792 228216 118844 228268
rect 150624 228216 150676 228268
rect 150808 228216 150860 228268
rect 195888 228216 195940 228268
rect 149520 228080 149572 228132
rect 209688 228080 209740 228132
rect 65984 227944 66036 227996
rect 155776 227944 155828 227996
rect 155960 227944 156012 227996
rect 205548 227944 205600 227996
rect 208952 227944 209004 227996
rect 249340 228216 249392 228268
rect 226616 228080 226668 228132
rect 233700 228080 233752 228132
rect 248880 228080 248932 228132
rect 276112 228216 276164 228268
rect 428464 228216 428516 228268
rect 455696 228216 455748 228268
rect 440792 228080 440844 228132
rect 463332 228216 463384 228268
rect 463884 228352 463936 228404
rect 474924 228352 474976 228404
rect 477592 228352 477644 228404
rect 552296 228352 552348 228404
rect 471980 228216 472032 228268
rect 474648 228216 474700 228268
rect 534724 228216 534776 228268
rect 540336 228216 540388 228268
rect 546500 228216 546552 228268
rect 456248 228080 456300 228132
rect 513196 228080 513248 228132
rect 356336 227944 356388 227996
rect 359096 227944 359148 227996
rect 454500 227944 454552 227996
rect 514760 227944 514812 227996
rect 127072 227808 127124 227860
rect 181720 227808 181772 227860
rect 204536 227808 204588 227860
rect 211528 227808 211580 227860
rect 455696 227808 455748 227860
rect 262128 227740 262180 227792
rect 268936 227740 268988 227792
rect 308496 227740 308548 227792
rect 315856 227740 315908 227792
rect 42524 227672 42576 227724
rect 47216 227672 47268 227724
rect 118608 227672 118660 227724
rect 127808 227672 127860 227724
rect 137100 227672 137152 227724
rect 137284 227672 137336 227724
rect 197728 227672 197780 227724
rect 199384 227672 199436 227724
rect 242992 227672 243044 227724
rect 272524 227672 272576 227724
rect 285496 227672 285548 227724
rect 97356 227400 97408 227452
rect 127256 227536 127308 227588
rect 315856 227604 315908 227656
rect 316960 227740 317012 227792
rect 317328 227740 317380 227792
rect 321836 227740 321888 227792
rect 408408 227672 408460 227724
rect 443552 227672 443604 227724
rect 459560 227808 459612 227860
rect 518072 227808 518124 227860
rect 459744 227672 459796 227724
rect 461032 227672 461084 227724
rect 527824 227672 527876 227724
rect 191104 227536 191156 227588
rect 192668 227536 192720 227588
rect 236000 227536 236052 227588
rect 249708 227536 249760 227588
rect 277216 227536 277268 227588
rect 383936 227536 383988 227588
rect 398840 227536 398892 227588
rect 415216 227536 415268 227588
rect 452568 227536 452620 227588
rect 468208 227536 468260 227588
rect 538220 227536 538272 227588
rect 115664 227400 115716 227452
rect 188896 227400 188948 227452
rect 189080 227400 189132 227452
rect 236368 227400 236420 227452
rect 242256 227400 242308 227452
rect 271696 227400 271748 227452
rect 372160 227400 372212 227452
rect 389732 227400 389784 227452
rect 395344 227400 395396 227452
rect 426440 227400 426492 227452
rect 432144 227400 432196 227452
rect 476212 227400 476264 227452
rect 477224 227400 477276 227452
rect 547972 227400 548024 227452
rect 82544 227264 82596 227316
rect 157432 227264 157484 227316
rect 157708 227196 157760 227248
rect 175832 227264 175884 227316
rect 179052 227264 179104 227316
rect 192116 227264 192168 227316
rect 72516 227128 72568 227180
rect 156604 227128 156656 227180
rect 165160 227128 165212 227180
rect 187240 227128 187292 227180
rect 234160 227264 234212 227316
rect 236000 227264 236052 227316
rect 266176 227264 266228 227316
rect 267556 227264 267608 227316
rect 287428 227264 287480 227316
rect 367192 227264 367244 227316
rect 385592 227264 385644 227316
rect 415768 227264 415820 227316
rect 458456 227264 458508 227316
rect 63592 226992 63644 227044
rect 142114 226992 142166 227044
rect 142252 226992 142304 227044
rect 157524 226992 157576 227044
rect 157800 226992 157852 227044
rect 122196 226856 122248 226908
rect 179052 226856 179104 226908
rect 182824 226992 182876 227044
rect 185952 226992 186004 227044
rect 186136 226992 186188 227044
rect 197452 227128 197504 227180
rect 204904 227128 204956 227180
rect 205088 227128 205140 227180
rect 212632 227128 212684 227180
rect 235724 227128 235776 227180
rect 267188 227128 267240 227180
rect 267372 227128 267424 227180
rect 290188 227128 290240 227180
rect 293684 227128 293736 227180
rect 305368 227128 305420 227180
rect 361488 227128 361540 227180
rect 371516 227128 371568 227180
rect 382096 227128 382148 227180
rect 407304 227128 407356 227180
rect 420184 227128 420236 227180
rect 465264 227264 465316 227316
rect 475384 227264 475436 227316
rect 548708 227264 548760 227316
rect 464988 227128 465040 227180
rect 478328 227128 478380 227180
rect 479800 227128 479852 227180
rect 554780 227128 554832 227180
rect 187976 226992 188028 227044
rect 231952 226992 232004 227044
rect 237288 226992 237340 227044
rect 128820 226720 128872 226772
rect 137284 226720 137336 226772
rect 137468 226720 137520 226772
rect 142114 226720 142166 226772
rect 142252 226720 142304 226772
rect 204904 226856 204956 226908
rect 240784 226856 240836 226908
rect 263416 226992 263468 227044
rect 272524 226992 272576 227044
rect 283656 226992 283708 227044
rect 298468 226992 298520 227044
rect 299388 226992 299440 227044
rect 310336 226992 310388 227044
rect 311072 226992 311124 227044
rect 319168 226992 319220 227044
rect 353944 226992 353996 227044
rect 365812 226992 365864 227044
rect 366824 226992 366876 227044
rect 383936 226992 383988 227044
rect 388720 226992 388772 227044
rect 417056 226992 417108 227044
rect 426256 226992 426308 227044
rect 473544 226992 473596 227044
rect 480536 226992 480588 227044
rect 484676 226992 484728 227044
rect 485320 226992 485372 227044
rect 563888 226992 563940 227044
rect 267832 226856 267884 226908
rect 399760 226856 399812 226908
rect 433616 226856 433668 226908
rect 436192 226856 436244 226908
rect 464988 226856 465040 226908
rect 465724 226856 465776 226908
rect 519176 226856 519228 226908
rect 132224 226584 132276 226636
rect 199660 226584 199712 226636
rect 205088 226720 205140 226772
rect 205640 226720 205692 226772
rect 248512 226788 248564 226840
rect 427728 226720 427780 226772
rect 452752 226720 452804 226772
rect 513380 226720 513432 226772
rect 206560 226584 206612 226636
rect 141884 226448 141936 226500
rect 142160 226448 142212 226500
rect 142344 226448 142396 226500
rect 204352 226448 204404 226500
rect 138756 226380 138808 226432
rect 141700 226380 141752 226432
rect 241888 226584 241940 226636
rect 452752 226584 452804 226636
rect 456064 226584 456116 226636
rect 465724 226584 465776 226636
rect 465908 226584 465960 226636
rect 520556 226584 520608 226636
rect 450544 226448 450596 226500
rect 489874 226448 489926 226500
rect 490932 226448 490984 226500
rect 495532 226448 495584 226500
rect 201960 226312 202012 226364
rect 243360 226380 243412 226432
rect 246856 226380 246908 226432
rect 289544 226312 289596 226364
rect 293868 226312 293920 226364
rect 97908 226244 97960 226296
rect 167000 226244 167052 226296
rect 167184 226244 167236 226296
rect 173440 226244 173492 226296
rect 173624 226244 173676 226296
rect 175648 226244 175700 226296
rect 175832 226244 175884 226296
rect 42432 226176 42484 226228
rect 45560 226176 45612 226228
rect 84936 226108 84988 226160
rect 92388 225972 92440 226024
rect 162400 226108 162452 226160
rect 88064 225836 88116 225888
rect 165988 225972 166040 226024
rect 166448 225972 166500 226024
rect 167368 225972 167420 226024
rect 78404 225700 78456 225752
rect 161848 225700 161900 225752
rect 167184 225836 167236 225888
rect 168472 225972 168524 226024
rect 173256 226108 173308 226160
rect 176476 226108 176528 226160
rect 176752 226244 176804 226296
rect 190276 226244 190328 226296
rect 190414 226244 190466 226296
rect 195060 226244 195112 226296
rect 195244 226244 195296 226296
rect 201776 226244 201828 226296
rect 205456 226244 205508 226296
rect 247408 226244 247460 226296
rect 413008 226244 413060 226296
rect 449072 226244 449124 226296
rect 469312 226244 469364 226296
rect 540336 226244 540388 226296
rect 181352 226108 181404 226160
rect 224224 226108 224276 226160
rect 225696 226108 225748 226160
rect 260656 226108 260708 226160
rect 273720 226108 273772 226160
rect 292120 226108 292172 226160
rect 379888 226108 379940 226160
rect 402980 226108 403032 226160
rect 408592 226108 408644 226160
rect 447048 226108 447100 226160
rect 478696 226108 478748 226160
rect 553676 226108 553728 226160
rect 168288 225836 168340 225888
rect 180800 225836 180852 225888
rect 226432 225972 226484 226024
rect 255228 225972 255280 226024
rect 280528 225972 280580 226024
rect 381176 225972 381228 226024
rect 394884 225972 394936 226024
rect 400680 225972 400732 226024
rect 219808 225836 219860 225888
rect 224224 225836 224276 225888
rect 230848 225836 230900 225888
rect 252744 225836 252796 225888
rect 279424 225836 279476 225888
rect 382648 225836 382700 225888
rect 408776 225836 408828 225888
rect 425152 225972 425204 226024
rect 469312 225972 469364 226024
rect 475108 225972 475160 226024
rect 483572 225972 483624 226024
rect 484032 225972 484084 226024
rect 489552 225972 489604 226024
rect 489736 225972 489788 226024
rect 556160 225972 556212 226024
rect 425796 225836 425848 225888
rect 427912 225836 427964 225888
rect 474188 225836 474240 225888
rect 482008 225836 482060 225888
rect 558920 225836 558972 225888
rect 167828 225700 167880 225752
rect 214380 225700 214432 225752
rect 214564 225700 214616 225752
rect 226984 225700 227036 225752
rect 227168 225700 227220 225752
rect 259552 225700 259604 225752
rect 260564 225700 260616 225752
rect 283288 225700 283340 225752
rect 290280 225700 290332 225752
rect 303160 225700 303212 225752
rect 303344 225700 303396 225752
rect 310888 225700 310940 225752
rect 312728 225700 312780 225752
rect 317512 225700 317564 225752
rect 352288 225700 352340 225752
rect 357624 225700 357676 225752
rect 362776 225700 362828 225752
rect 378968 225700 379020 225752
rect 386880 225700 386932 225752
rect 414020 225700 414072 225752
rect 438216 225700 438268 225752
rect 489874 225700 489926 225752
rect 490012 225700 490064 225752
rect 561220 225700 561272 225752
rect 62120 225564 62172 225616
rect 149704 225564 149756 225616
rect 151176 225564 151228 225616
rect 213184 225564 213236 225616
rect 214196 225564 214248 225616
rect 224224 225564 224276 225616
rect 246764 225564 246816 225616
rect 274180 225564 274232 225616
rect 279608 225564 279660 225616
rect 297088 225564 297140 225616
rect 298008 225564 298060 225616
rect 308128 225564 308180 225616
rect 357072 225564 357124 225616
rect 365260 225564 365312 225616
rect 365444 225564 365496 225616
rect 382648 225564 382700 225616
rect 393688 225564 393740 225616
rect 423036 225564 423088 225616
rect 433984 225564 434036 225616
rect 475108 225564 475160 225616
rect 480352 225564 480404 225616
rect 486792 225564 486844 225616
rect 486976 225564 487028 225616
rect 566096 225564 566148 225616
rect 81348 225428 81400 225480
rect 158444 225428 158496 225480
rect 158628 225428 158680 225480
rect 212356 225428 212408 225480
rect 212540 225428 212592 225480
rect 215392 225428 215444 225480
rect 215576 225428 215628 225480
rect 104808 225292 104860 225344
rect 178132 225292 178184 225344
rect 178500 225292 178552 225344
rect 214196 225292 214248 225344
rect 214748 225292 214800 225344
rect 217600 225292 217652 225344
rect 219164 225428 219216 225480
rect 255964 225428 256016 225480
rect 410800 225428 410852 225480
rect 437480 225428 437532 225480
rect 448888 225428 448940 225480
rect 509516 225428 509568 225480
rect 252928 225292 252980 225344
rect 417424 225292 417476 225344
rect 436744 225292 436796 225344
rect 442632 225292 442684 225344
rect 489874 225292 489926 225344
rect 490012 225292 490064 225344
rect 492588 225292 492640 225344
rect 492772 225292 492824 225344
rect 499028 225292 499080 225344
rect 134984 225156 135036 225208
rect 195244 225156 195296 225208
rect 195428 225156 195480 225208
rect 214564 225156 214616 225208
rect 215760 225156 215812 225208
rect 254032 225156 254084 225208
rect 407488 225156 407540 225208
rect 421104 225156 421156 225208
rect 440056 225156 440108 225208
rect 495716 225156 495768 225208
rect 120080 225020 120132 225072
rect 151636 225020 151688 225072
rect 151774 225020 151826 225072
rect 161296 225020 161348 225072
rect 161480 225020 161532 225072
rect 212540 225020 212592 225072
rect 214380 225020 214432 225072
rect 221464 225020 221516 225072
rect 222292 225020 222344 225072
rect 227168 225020 227220 225072
rect 231676 225020 231728 225072
rect 238024 225020 238076 225072
rect 445944 225020 445996 225072
rect 501512 225020 501564 225072
rect 378048 224952 378100 225004
rect 379796 224952 379848 225004
rect 42616 224884 42668 224936
rect 45744 224884 45796 224936
rect 121368 224884 121420 224936
rect 77024 224748 77076 224800
rect 151452 224748 151504 224800
rect 151728 224748 151780 224800
rect 159364 224748 159416 224800
rect 159732 224748 159784 224800
rect 180616 224748 180668 224800
rect 180800 224748 180852 224800
rect 181904 224748 181956 224800
rect 184848 224884 184900 224936
rect 194416 224884 194468 224936
rect 194876 224884 194928 224936
rect 198280 224884 198332 224936
rect 198464 224884 198516 224936
rect 243728 224884 243780 224936
rect 244556 224884 244608 224936
rect 272800 224884 272852 224936
rect 370504 224884 370556 224936
rect 376116 224884 376168 224936
rect 409788 224884 409840 224936
rect 441068 224884 441120 224936
rect 442816 224884 442868 224936
rect 187056 224748 187108 224800
rect 187240 224748 187292 224800
rect 234712 224748 234764 224800
rect 240600 224748 240652 224800
rect 270040 224748 270092 224800
rect 347872 224748 347924 224800
rect 353484 224748 353536 224800
rect 394700 224748 394752 224800
rect 411260 224748 411312 224800
rect 412456 224748 412508 224800
rect 451280 224748 451332 224800
rect 451464 224748 451516 224800
rect 462964 224748 463016 224800
rect 464344 224884 464396 224936
rect 471796 224884 471848 224936
rect 472256 224884 472308 224936
rect 534172 224884 534224 224936
rect 465080 224748 465132 224800
rect 467104 224748 467156 224800
rect 536380 224748 536432 224800
rect 99104 224612 99156 224664
rect 177856 224612 177908 224664
rect 178040 224612 178092 224664
rect 194876 224612 194928 224664
rect 197268 224612 197320 224664
rect 204536 224612 204588 224664
rect 204720 224612 204772 224664
rect 210700 224612 210752 224664
rect 210884 224612 210936 224664
rect 229192 224612 229244 224664
rect 231860 224612 231912 224664
rect 236920 224612 236972 224664
rect 238576 224612 238628 224664
rect 269488 224612 269540 224664
rect 281264 224612 281316 224664
rect 296720 224612 296772 224664
rect 375840 224612 375892 224664
rect 397552 224612 397604 224664
rect 397920 224612 397972 224664
rect 414572 224612 414624 224664
rect 414756 224612 414808 224664
rect 454316 224612 454368 224664
rect 460480 224612 460532 224664
rect 524236 224612 524288 224664
rect 524374 224612 524426 224664
rect 533344 224612 533396 224664
rect 75000 224476 75052 224528
rect 151728 224476 151780 224528
rect 152096 224476 152148 224528
rect 155040 224476 155092 224528
rect 155408 224476 155460 224528
rect 157294 224476 157346 224528
rect 157432 224476 157484 224528
rect 159732 224476 159784 224528
rect 159916 224476 159968 224528
rect 162952 224476 163004 224528
rect 163136 224476 163188 224528
rect 218704 224476 218756 224528
rect 232320 224476 232372 224528
rect 265072 224476 265124 224528
rect 270224 224476 270276 224528
rect 288256 224476 288308 224528
rect 305000 224476 305052 224528
rect 312544 224476 312596 224528
rect 368388 224476 368440 224528
rect 376760 224476 376812 224528
rect 384120 224476 384172 224528
rect 407948 224476 408000 224528
rect 423404 224476 423456 224528
rect 445300 224476 445352 224528
rect 446128 224476 446180 224528
rect 461584 224476 461636 224528
rect 465448 224476 465500 224528
rect 472256 224476 472308 224528
rect 61844 224340 61896 224392
rect 146024 224340 146076 224392
rect 146208 224340 146260 224392
rect 206836 224340 206888 224392
rect 207020 224340 207072 224392
rect 207940 224340 207992 224392
rect 210424 224340 210476 224392
rect 212080 224340 212132 224392
rect 214564 224340 214616 224392
rect 250720 224340 250772 224392
rect 271604 224340 271656 224392
rect 291568 224340 291620 224392
rect 296628 224340 296680 224392
rect 307576 224340 307628 224392
rect 359740 224340 359792 224392
rect 368480 224340 368532 224392
rect 376392 224340 376444 224392
rect 399024 224340 399076 224392
rect 423680 224340 423732 224392
rect 467932 224340 467984 224392
rect 470416 224340 470468 224392
rect 475384 224476 475436 224528
rect 475568 224476 475620 224528
rect 543924 224476 543976 224528
rect 472624 224340 472676 224392
rect 533160 224340 533212 224392
rect 533344 224340 533396 224392
rect 541348 224340 541400 224392
rect 542084 224340 542136 224392
rect 557356 224340 557408 224392
rect 68468 224204 68520 224256
rect 155224 224204 155276 224256
rect 155592 224204 155644 224256
rect 204720 224204 204772 224256
rect 204904 224204 204956 224256
rect 124680 224068 124732 224120
rect 190368 224068 190420 224120
rect 191748 224068 191800 224120
rect 231860 224068 231912 224120
rect 234620 224204 234672 224256
rect 268384 224204 268436 224256
rect 270408 224204 270460 224256
rect 289912 224204 289964 224256
rect 291200 224204 291252 224256
rect 305920 224204 305972 224256
rect 307484 224204 307536 224256
rect 315028 224204 315080 224256
rect 358360 224204 358412 224256
rect 372712 224204 372764 224256
rect 380440 224204 380492 224256
rect 405740 224204 405792 224256
rect 406660 224204 406712 224256
rect 431132 224204 431184 224256
rect 435640 224204 435692 224256
rect 485228 224204 485280 224256
rect 499488 224204 499540 224256
rect 505192 224204 505244 224256
rect 547420 224204 547472 224256
rect 562324 224204 562376 224256
rect 571340 224204 571392 224256
rect 234988 224068 235040 224120
rect 399484 224068 399536 224120
rect 418160 224068 418212 224120
rect 429844 224068 429896 224120
rect 461032 224068 461084 224120
rect 461584 224068 461636 224120
rect 466460 224068 466512 224120
rect 468760 224068 468812 224120
rect 472624 224068 472676 224120
rect 475384 224068 475436 224120
rect 480904 224068 480956 224120
rect 481088 224068 481140 224120
rect 499672 224136 499724 224188
rect 504916 224136 504968 224188
rect 485780 224068 485832 224120
rect 499488 224068 499540 224120
rect 509884 224068 509936 224120
rect 551284 224068 551336 224120
rect 131028 223932 131080 223984
rect 134708 223796 134760 223848
rect 193496 223796 193548 223848
rect 194416 223932 194468 223984
rect 204904 223932 204956 223984
rect 196900 223796 196952 223848
rect 200856 223796 200908 223848
rect 141240 223660 141292 223712
rect 203800 223660 203852 223712
rect 204536 223796 204588 223848
rect 241152 223932 241204 223984
rect 272984 223932 273036 223984
rect 275652 223932 275704 223984
rect 403256 223932 403308 223984
rect 424692 223932 424744 223984
rect 425520 223932 425572 223984
rect 457720 223932 457772 223984
rect 462136 223932 462188 223984
rect 528836 223932 528888 223984
rect 533160 223932 533212 223984
rect 538864 223932 538916 223984
rect 243176 223796 243228 223848
rect 412732 223796 412784 223848
rect 447692 223796 447744 223848
rect 454776 223796 454828 223848
rect 208400 223660 208452 223712
rect 214564 223660 214616 223712
rect 416320 223660 416372 223712
rect 429200 223660 429252 223712
rect 472440 223660 472492 223712
rect 475568 223660 475620 223712
rect 477040 223660 477092 223712
rect 242900 223592 242952 223644
rect 245200 223592 245252 223644
rect 94964 223524 95016 223576
rect 91560 223388 91612 223440
rect 161940 223388 161992 223440
rect 86684 223252 86736 223304
rect 167644 223388 167696 223440
rect 173808 223524 173860 223576
rect 172612 223388 172664 223440
rect 173532 223388 173584 223440
rect 177028 223388 177080 223440
rect 180708 223524 180760 223576
rect 230296 223524 230348 223576
rect 250536 223524 250588 223576
rect 276480 223524 276532 223576
rect 277124 223524 277176 223576
rect 294328 223524 294380 223576
rect 313096 223524 313148 223576
rect 318616 223524 318668 223576
rect 350172 223524 350224 223576
rect 355692 223524 355744 223576
rect 369584 223524 369636 223576
rect 374000 223524 374052 223576
rect 223120 223388 223172 223440
rect 226064 223388 226116 223440
rect 227352 223388 227404 223440
rect 227628 223388 227680 223440
rect 258632 223388 258684 223440
rect 258816 223388 258868 223440
rect 282460 223388 282512 223440
rect 310612 223388 310664 223440
rect 314200 223388 314252 223440
rect 345112 223388 345164 223440
rect 352472 223388 352524 223440
rect 368848 223388 368900 223440
rect 387248 223524 387300 223576
rect 392860 223524 392912 223576
rect 416228 223524 416280 223576
rect 424232 223524 424284 223576
rect 436192 223524 436244 223576
rect 443736 223524 443788 223576
rect 444196 223524 444248 223576
rect 480904 223660 480956 223712
rect 499304 223660 499356 223712
rect 499948 223796 500000 223848
rect 509884 223796 509936 223848
rect 510068 223796 510120 223848
rect 514576 223796 514628 223848
rect 516784 223796 516836 223848
rect 524236 223796 524288 223848
rect 524374 223796 524426 223848
rect 617708 223796 617760 223848
rect 504732 223660 504784 223712
rect 499534 223592 499586 223644
rect 485228 223524 485280 223576
rect 485872 223524 485924 223576
rect 499304 223524 499356 223576
rect 629852 223592 629904 223644
rect 505376 223456 505428 223508
rect 516784 223456 516836 223508
rect 379336 223388 379388 223440
rect 393504 223388 393556 223440
rect 401692 223388 401744 223440
rect 426624 223388 426676 223440
rect 436560 223388 436612 223440
rect 449900 223388 449952 223440
rect 452200 223388 452252 223440
rect 505192 223388 505244 223440
rect 522580 223388 522632 223440
rect 554964 223388 555016 223440
rect 74264 223116 74316 223168
rect 82912 223116 82964 223168
rect 83280 223116 83332 223168
rect 157294 223116 157346 223168
rect 157432 223116 157484 223168
rect 161112 223116 161164 223168
rect 161940 223116 161992 223168
rect 170680 223252 170732 223304
rect 170864 223252 170916 223304
rect 223672 223252 223724 223304
rect 227444 223252 227496 223304
rect 261116 223252 261168 223304
rect 261300 223252 261352 223304
rect 286048 223252 286100 223304
rect 293960 223252 294012 223304
rect 302056 223252 302108 223304
rect 362408 223252 362460 223304
rect 165252 223116 165304 223168
rect 173072 223116 173124 223168
rect 79784 222980 79836 223032
rect 163504 222980 163556 223032
rect 164148 222980 164200 223032
rect 185584 223116 185636 223168
rect 185768 223116 185820 223168
rect 174084 222980 174136 223032
rect 214564 222980 214616 223032
rect 214748 222980 214800 223032
rect 218980 222980 219032 223032
rect 224224 223116 224276 223168
rect 227628 223116 227680 223168
rect 228640 223116 228692 223168
rect 252284 223116 252336 223168
rect 278320 223116 278372 223168
rect 288348 223116 288400 223168
rect 302608 223116 302660 223168
rect 353024 223116 353076 223168
rect 357440 223116 357492 223168
rect 363144 223116 363196 223168
rect 377864 223252 377916 223304
rect 396356 223252 396408 223304
rect 397184 223252 397236 223304
rect 422852 223252 422904 223304
rect 427544 223252 427596 223304
rect 446036 223252 446088 223304
rect 447876 223252 447928 223304
rect 455696 223252 455748 223304
rect 455880 223252 455932 223304
rect 518992 223252 519044 223304
rect 519544 223252 519596 223304
rect 531320 223252 531372 223304
rect 228180 222980 228232 223032
rect 263968 222980 264020 223032
rect 278688 222980 278740 223032
rect 295984 222980 296036 223032
rect 302240 222980 302292 223032
rect 311440 222980 311492 223032
rect 354404 222980 354456 223032
rect 363236 222980 363288 223032
rect 369860 223116 369912 223168
rect 374368 223116 374420 223168
rect 379336 223116 379388 223168
rect 385776 223116 385828 223168
rect 409972 223116 410024 223168
rect 411904 223116 411956 223168
rect 444012 223116 444064 223168
rect 444196 223116 444248 223168
rect 485734 223116 485786 223168
rect 485872 223116 485924 223168
rect 560392 223116 560444 223168
rect 369032 222980 369084 223032
rect 373632 222980 373684 223032
rect 392216 222980 392268 223032
rect 394056 222980 394108 223032
rect 419724 222980 419776 223032
rect 426072 222980 426124 223032
rect 463884 222980 463936 223032
rect 464160 222980 464212 223032
rect 60372 222844 60424 222896
rect 142114 222844 142166 222896
rect 142436 222844 142488 222896
rect 152464 222844 152516 222896
rect 152648 222844 152700 222896
rect 157156 222844 157208 222896
rect 157340 222844 157392 222896
rect 158168 222844 158220 222896
rect 158352 222844 158404 222896
rect 165528 222844 165580 222896
rect 165712 222844 165764 222896
rect 215208 222844 215260 222896
rect 218060 222844 218112 222896
rect 257344 222844 257396 222896
rect 257988 222844 258040 222896
rect 283840 222844 283892 222896
rect 284024 222844 284076 222896
rect 300492 222844 300544 222896
rect 303528 222844 303580 222896
rect 311992 222844 312044 222896
rect 314384 222844 314436 222896
rect 320088 222844 320140 222896
rect 342904 222844 342956 222896
rect 349252 222844 349304 222896
rect 355968 222844 356020 222896
rect 367376 222844 367428 222896
rect 371056 222844 371108 222896
rect 390928 222844 390980 222896
rect 405280 222844 405332 222896
rect 439412 222844 439464 222896
rect 439872 222844 439924 222896
rect 485872 222844 485924 222896
rect 488908 222776 488960 222828
rect 490932 222776 490984 222828
rect 114468 222708 114520 222760
rect 185032 222708 185084 222760
rect 102140 222572 102192 222624
rect 152280 222572 152332 222624
rect 152464 222572 152516 222624
rect 173532 222572 173584 222624
rect 175188 222572 175240 222624
rect 185768 222708 185820 222760
rect 191564 222708 191616 222760
rect 239680 222708 239732 222760
rect 391756 222708 391808 222760
rect 412916 222708 412968 222760
rect 413192 222708 413244 222760
rect 429476 222708 429528 222760
rect 442080 222708 442132 222760
rect 486424 222708 486476 222760
rect 491392 222980 491444 223032
rect 563612 222980 563664 223032
rect 491576 222844 491628 222896
rect 565728 222844 565780 222896
rect 519544 222708 519596 222760
rect 185584 222572 185636 222624
rect 213368 222572 213420 222624
rect 213736 222572 213788 222624
rect 252100 222572 252152 222624
rect 299756 222572 299808 222624
rect 306472 222572 306524 222624
rect 390008 222572 390060 222624
rect 406292 222572 406344 222624
rect 406936 222572 406988 222624
rect 423772 222572 423824 222624
rect 448336 222572 448388 222624
rect 499488 222572 499540 222624
rect 499672 222572 499724 222624
rect 500868 222572 500920 222624
rect 501052 222572 501104 222624
rect 503444 222572 503496 222624
rect 505192 222572 505244 222624
rect 514024 222572 514076 222624
rect 554780 222572 554832 222624
rect 555424 222572 555476 222624
rect 557356 222572 557408 222624
rect 565728 222572 565780 222624
rect 611360 222572 611412 222624
rect 626540 222572 626592 222624
rect 661684 222572 661736 222624
rect 668400 222708 668452 222760
rect 675116 222640 675168 222692
rect 101496 222436 101548 222488
rect 125324 222436 125376 222488
rect 142114 222300 142166 222352
rect 142620 222300 142672 222352
rect 194600 222300 194652 222352
rect 194968 222436 195020 222488
rect 195612 222300 195664 222352
rect 207204 222436 207256 222488
rect 215944 222436 215996 222488
rect 220636 222436 220688 222488
rect 256792 222436 256844 222488
rect 389088 222436 389140 222488
rect 403164 222436 403216 222488
rect 411720 222436 411772 222488
rect 428096 222436 428148 222488
rect 450084 222436 450136 222488
rect 505008 222436 505060 222488
rect 505192 222436 505244 222488
rect 510712 222436 510764 222488
rect 555424 222436 555476 222488
rect 608600 222436 608652 222488
rect 663064 222436 663116 222488
rect 668400 222436 668452 222488
rect 675484 222504 675536 222556
rect 438400 222368 438452 222420
rect 442908 222368 442960 222420
rect 523132 222368 523184 222420
rect 523684 222368 523736 222420
rect 207388 222300 207440 222352
rect 214564 222300 214616 222352
rect 221740 222300 221792 222352
rect 420920 222300 420972 222352
rect 432788 222300 432840 222352
rect 444840 222300 444892 222352
rect 503168 222300 503220 222352
rect 503444 222300 503496 222352
rect 508504 222300 508556 222352
rect 119712 222096 119764 222148
rect 181168 222164 181220 222216
rect 181444 222096 181496 222148
rect 183468 222096 183520 222148
rect 184296 222096 184348 222148
rect 116400 221960 116452 222012
rect 181996 221960 182048 222012
rect 182180 221960 182232 222012
rect 185768 221960 185820 222012
rect 188988 222096 189040 222148
rect 192484 221960 192536 222012
rect 80796 221824 80848 221876
rect 111064 221824 111116 221876
rect 111432 221824 111484 221876
rect 183836 221824 183888 221876
rect 185584 221824 185636 221876
rect 191932 221824 191984 221876
rect 195152 222096 195204 222148
rect 201592 222232 201644 222284
rect 201224 222096 201276 222148
rect 245936 222096 245988 222148
rect 248144 222096 248196 222148
rect 251272 222096 251324 222148
rect 261668 222096 261720 222148
rect 265256 222096 265308 222148
rect 266268 222096 266320 222148
rect 267004 222096 267056 222148
rect 267188 222096 267240 222148
rect 284576 222096 284628 222148
rect 347136 222096 347188 222148
rect 354220 222096 354272 222148
rect 381912 222096 381964 222148
rect 388444 222096 388496 222148
rect 402704 222096 402756 222148
rect 438860 222096 438912 222148
rect 446864 222096 446916 222148
rect 499580 222096 499632 222148
rect 499764 222096 499816 222148
rect 519728 222232 519780 222284
rect 547420 222300 547472 222352
rect 623964 222300 624016 222352
rect 664628 222300 664680 222352
rect 675300 222368 675352 222420
rect 601700 222164 601752 222216
rect 664444 222164 664496 222216
rect 519544 222096 519596 222148
rect 530768 222096 530820 222148
rect 675484 222232 675536 222284
rect 192852 222028 192904 222080
rect 194232 222028 194284 222080
rect 246396 222028 246448 222080
rect 247776 222028 247828 222080
rect 194416 221960 194468 222012
rect 238944 221960 238996 222012
rect 247960 221960 248012 222012
rect 274732 221960 274784 222012
rect 237472 221824 237524 221876
rect 243912 221824 243964 221876
rect 272064 221824 272116 221876
rect 97724 221688 97776 221740
rect 171048 221688 171100 221740
rect 171232 221688 171284 221740
rect 181260 221688 181312 221740
rect 181444 221688 181496 221740
rect 225512 221688 225564 221740
rect 231860 221688 231912 221740
rect 233424 221688 233476 221740
rect 233700 221688 233752 221740
rect 261668 221688 261720 221740
rect 261944 221688 261996 221740
rect 267188 221688 267240 221740
rect 59820 221552 59872 221604
rect 144368 221552 144420 221604
rect 144552 221552 144604 221604
rect 200074 221552 200126 221604
rect 200304 221552 200356 221604
rect 202328 221552 202380 221604
rect 204720 221552 204772 221604
rect 227904 221552 227956 221604
rect 230388 221552 230440 221604
rect 263140 221552 263192 221604
rect 268752 221552 268804 221604
rect 288992 221960 289044 222012
rect 388628 221960 388680 222012
rect 412180 221960 412232 222012
rect 417792 221960 417844 222012
rect 461860 221960 461912 222012
rect 473176 221960 473228 222012
rect 545764 221960 545816 222012
rect 549904 221960 549956 222012
rect 560576 221960 560628 222012
rect 285312 221824 285364 221876
rect 300124 221824 300176 221876
rect 362592 221824 362644 221876
rect 377404 221824 377456 221876
rect 379152 221824 379204 221876
rect 402244 221824 402296 221876
rect 409604 221824 409656 221876
rect 448612 221824 448664 221876
rect 477408 221824 477460 221876
rect 550640 221824 550692 221876
rect 558184 221824 558236 221876
rect 564716 221824 564768 221876
rect 280068 221688 280120 221740
rect 296168 221688 296220 221740
rect 300124 221688 300176 221740
rect 309508 221688 309560 221740
rect 310060 221688 310112 221740
rect 316132 221688 316184 221740
rect 343548 221688 343600 221740
rect 347872 221688 347924 221740
rect 351736 221688 351788 221740
rect 362500 221688 362552 221740
rect 371884 221688 371936 221740
rect 389180 221688 389232 221740
rect 390468 221688 390520 221740
rect 418804 221688 418856 221740
rect 422208 221688 422260 221740
rect 464344 221688 464396 221740
rect 475936 221688 475988 221740
rect 549996 221688 550048 221740
rect 565084 221688 565136 221740
rect 567384 221688 567436 221740
rect 288624 221552 288676 221604
rect 303712 221552 303764 221604
rect 315120 221552 315172 221604
rect 319444 221552 319496 221604
rect 344836 221552 344888 221604
rect 350908 221552 350960 221604
rect 354588 221552 354640 221604
rect 364340 221552 364392 221604
rect 365628 221552 365680 221604
rect 380900 221552 380952 221604
rect 387524 221552 387576 221604
rect 415584 221552 415636 221604
rect 445668 221552 445720 221604
rect 475384 221552 475436 221604
rect 477868 221552 477920 221604
rect 70032 221416 70084 221468
rect 151636 221416 151688 221468
rect 151820 221416 151872 221468
rect 159824 221416 159876 221468
rect 160008 221416 160060 221468
rect 160744 221416 160796 221468
rect 160928 221416 160980 221468
rect 166816 221416 166868 221468
rect 166954 221416 167006 221468
rect 213276 221416 213328 221468
rect 122564 221280 122616 221332
rect 185584 221280 185636 221332
rect 185768 221280 185820 221332
rect 204720 221280 204772 221332
rect 232136 221416 232188 221468
rect 240048 221416 240100 221468
rect 270592 221416 270644 221468
rect 271236 221416 271288 221468
rect 292672 221416 292724 221468
rect 298560 221416 298612 221468
rect 309232 221416 309284 221468
rect 316040 221416 316092 221468
rect 321652 221416 321704 221468
rect 358176 221416 358228 221468
rect 370780 221416 370832 221468
rect 374644 221416 374696 221468
rect 395620 221416 395672 221468
rect 398564 221416 398616 221468
rect 432052 221416 432104 221468
rect 436008 221416 436060 221468
rect 485734 221416 485786 221468
rect 485872 221416 485924 221468
rect 495256 221416 495308 221468
rect 495394 221416 495446 221468
rect 519544 221416 519596 221468
rect 519728 221416 519780 221468
rect 129464 221144 129516 221196
rect 192300 221144 192352 221196
rect 192484 221144 192536 221196
rect 214748 221280 214800 221332
rect 245752 221280 245804 221332
rect 257160 221280 257212 221332
rect 280712 221280 280764 221332
rect 392584 221280 392636 221332
rect 422300 221280 422352 221332
rect 423220 221280 423272 221332
rect 459560 221280 459612 221332
rect 470232 221280 470284 221332
rect 540520 221280 540572 221332
rect 207480 221144 207532 221196
rect 247592 221144 247644 221196
rect 396724 221144 396776 221196
rect 428740 221144 428792 221196
rect 439596 221144 439648 221196
rect 466828 221144 466880 221196
rect 467748 221144 467800 221196
rect 535552 221144 535604 221196
rect 564716 221552 564768 221604
rect 596732 221688 596784 221740
rect 603448 221688 603500 221740
rect 568580 221416 568632 221468
rect 569500 221416 569552 221468
rect 553308 221280 553360 221332
rect 558000 221144 558052 221196
rect 558368 221280 558420 221332
rect 597100 221280 597152 221332
rect 620284 221416 620336 221468
rect 628196 221280 628248 221332
rect 608968 221144 609020 221196
rect 620284 221144 620336 221196
rect 628012 221144 628064 221196
rect 664260 221076 664312 221128
rect 675484 221076 675536 221128
rect 139124 221008 139176 221060
rect 171048 221008 171100 221060
rect 171232 221008 171284 221060
rect 210148 221008 210200 221060
rect 213276 221008 213328 221060
rect 216864 221008 216916 221060
rect 217416 221008 217468 221060
rect 254308 221008 254360 221060
rect 416044 221008 416096 221060
rect 441988 221008 442040 221060
rect 459928 221008 459980 221060
rect 526168 221008 526220 221060
rect 126152 220872 126204 220924
rect 127072 220872 127124 220924
rect 137928 220872 137980 220924
rect 195152 220872 195204 220924
rect 195336 220872 195388 220924
rect 199476 220872 199528 220924
rect 204168 220872 204220 220924
rect 214748 220872 214800 220924
rect 63960 220804 64012 220856
rect 66904 220804 66956 220856
rect 199844 220804 199896 220856
rect 201040 220804 201092 220856
rect 57612 220736 57664 220788
rect 62120 220736 62172 220788
rect 67364 220736 67416 220788
rect 69664 220736 69716 220788
rect 79140 220736 79192 220788
rect 79968 220736 80020 220788
rect 80152 220736 80204 220788
rect 102140 220736 102192 220788
rect 108120 220736 108172 220788
rect 63408 220600 63460 220652
rect 120080 220600 120132 220652
rect 123852 220736 123904 220788
rect 127808 220736 127860 220788
rect 127992 220736 128044 220788
rect 136548 220736 136600 220788
rect 136916 220736 136968 220788
rect 152464 220736 152516 220788
rect 153660 220736 153712 220788
rect 154120 220736 154172 220788
rect 154488 220736 154540 220788
rect 194968 220736 195020 220788
rect 195152 220736 195204 220788
rect 199660 220736 199712 220788
rect 203432 220736 203484 220788
rect 126152 220600 126204 220652
rect 126336 220600 126388 220652
rect 192484 220600 192536 220652
rect 193036 220600 193088 220652
rect 205272 220736 205324 220788
rect 239588 220736 239640 220788
rect 239772 220736 239824 220788
rect 240968 220736 241020 220788
rect 241244 220736 241296 220788
rect 244556 220736 244608 220788
rect 251088 220736 251140 220788
rect 252744 220736 252796 220788
rect 253020 220736 253072 220788
rect 256332 220736 256384 220788
rect 267096 220736 267148 220788
rect 267556 220736 267608 220788
rect 244740 220668 244792 220720
rect 247960 220668 248012 220720
rect 55956 220464 56008 220516
rect 56876 220464 56928 220516
rect 76656 220464 76708 220516
rect 80152 220464 80204 220516
rect 87420 220464 87472 220516
rect 88248 220464 88300 220516
rect 89076 220464 89128 220516
rect 89628 220464 89680 220516
rect 95700 220464 95752 220516
rect 97908 220464 97960 220516
rect 120540 220464 120592 220516
rect 127624 220464 127676 220516
rect 127808 220464 127860 220516
rect 161756 220464 161808 220516
rect 161940 220464 161992 220516
rect 162400 220464 162452 220516
rect 162584 220464 162636 220516
rect 165068 220464 165120 220516
rect 165620 220464 165672 220516
rect 166448 220464 166500 220516
rect 166632 220464 166684 220516
rect 203616 220464 203668 220516
rect 214564 220600 214616 220652
rect 216312 220600 216364 220652
rect 219716 220600 219768 220652
rect 219900 220600 219952 220652
rect 220452 220600 220504 220652
rect 221556 220600 221608 220652
rect 222292 220600 222344 220652
rect 222476 220600 222528 220652
rect 223856 220600 223908 220652
rect 224040 220600 224092 220652
rect 224500 220600 224552 220652
rect 232688 220600 232740 220652
rect 232872 220600 232924 220652
rect 233884 220600 233936 220652
rect 236460 220600 236512 220652
rect 243728 220600 243780 220652
rect 249524 220600 249576 220652
rect 277584 220872 277636 220924
rect 418988 220872 419040 220924
rect 455420 220872 455472 220924
rect 597100 221008 597152 221060
rect 608784 221008 608836 221060
rect 673276 220940 673328 220992
rect 675116 220940 675168 220992
rect 602252 220872 602304 220924
rect 296076 220804 296128 220856
rect 297364 220804 297416 220856
rect 275652 220736 275704 220788
rect 290464 220736 290516 220788
rect 302700 220736 302752 220788
rect 305644 220736 305696 220788
rect 277860 220600 277912 220652
rect 279608 220600 279660 220652
rect 304632 220600 304684 220652
rect 313464 220804 313516 220856
rect 461216 220804 461268 220856
rect 528376 220804 528428 220856
rect 596732 220804 596784 220856
rect 667848 220804 667900 220856
rect 675300 220804 675352 220856
rect 316776 220736 316828 220788
rect 320548 220736 320600 220788
rect 320916 220736 320968 220788
rect 321376 220736 321428 220788
rect 323400 220736 323452 220788
rect 324964 220736 325016 220788
rect 326712 220736 326764 220788
rect 327356 220736 327408 220788
rect 328184 220736 328236 220788
rect 328920 220736 328972 220788
rect 329104 220736 329156 220788
rect 330484 220736 330536 220788
rect 330852 220736 330904 220788
rect 332140 220736 332192 220788
rect 333888 220736 333940 220788
rect 334348 220736 334400 220788
rect 346216 220736 346268 220788
rect 351920 220736 351972 220788
rect 355324 220736 355376 220788
rect 358360 220736 358412 220788
rect 365260 220736 365312 220788
rect 366640 220736 366692 220788
rect 395160 220736 395212 220788
rect 398104 220736 398156 220788
rect 423036 220736 423088 220788
rect 425428 220736 425480 220788
rect 429200 220736 429252 220788
rect 456064 220736 456116 220788
rect 591304 220668 591356 220720
rect 321192 220600 321244 220652
rect 324688 220600 324740 220652
rect 327540 220600 327592 220652
rect 330208 220600 330260 220652
rect 355692 220600 355744 220652
rect 356704 220600 356756 220652
rect 357624 220600 357676 220652
rect 360200 220600 360252 220652
rect 393044 220600 393096 220652
rect 421288 220600 421340 220652
rect 425796 220600 425848 220652
rect 435548 220600 435600 220652
rect 444012 220600 444064 220652
rect 449440 220600 449492 220652
rect 449716 220600 449768 220652
rect 60648 220396 60700 220448
rect 61384 220396 61436 220448
rect 89444 220328 89496 220380
rect 165988 220328 166040 220380
rect 62580 220192 62632 220244
rect 63592 220192 63644 220244
rect 77208 220192 77260 220244
rect 156880 220192 156932 220244
rect 161296 220192 161348 220244
rect 161756 220192 161808 220244
rect 170036 220328 170088 220380
rect 170220 220328 170272 220380
rect 219532 220328 219584 220380
rect 219716 220328 219768 220380
rect 224040 220328 224092 220380
rect 250352 220464 250404 220516
rect 252836 220464 252888 220516
rect 253572 220464 253624 220516
rect 256332 220464 256384 220516
rect 281816 220464 281868 220516
rect 297732 220464 297784 220516
rect 299388 220464 299440 220516
rect 306840 220464 306892 220516
rect 310612 220464 310664 220516
rect 320088 220464 320140 220516
rect 323216 220464 323268 220516
rect 376116 220464 376168 220516
rect 388168 220464 388220 220516
rect 397368 220464 397420 220516
rect 427912 220464 427964 220516
rect 434720 220464 434772 220516
rect 437020 220464 437072 220516
rect 445300 220464 445352 220516
rect 445668 220464 445720 220516
rect 452568 220600 452620 220652
rect 456984 220600 457036 220652
rect 457168 220600 457220 220652
rect 470140 220600 470192 220652
rect 480352 220600 480404 220652
rect 471796 220464 471848 220516
rect 475200 220464 475252 220516
rect 475384 220464 475436 220516
rect 502340 220600 502392 220652
rect 504364 220600 504416 220652
rect 506020 220600 506072 220652
rect 506204 220600 506256 220652
rect 528560 220600 528612 220652
rect 548340 220600 548392 220652
rect 562508 220600 562560 220652
rect 562968 220600 563020 220652
rect 596272 220600 596324 220652
rect 481088 220464 481140 220516
rect 229468 220328 229520 220380
rect 231492 220328 231544 220380
rect 236000 220328 236052 220380
rect 239588 220328 239640 220380
rect 166954 220192 167006 220244
rect 171048 220192 171100 220244
rect 171876 220192 171928 220244
rect 173440 220192 173492 220244
rect 173624 220192 173676 220244
rect 181076 220192 181128 220244
rect 186872 220192 186924 220244
rect 187424 220192 187476 220244
rect 187608 220192 187660 220244
rect 58440 220056 58492 220108
rect 60372 220056 60424 220108
rect 64788 220056 64840 220108
rect 77024 220056 77076 220108
rect 103980 220056 104032 220108
rect 147634 220056 147686 220108
rect 147772 220056 147824 220108
rect 148968 220056 149020 220108
rect 149152 220056 149204 220108
rect 150164 220056 150216 220108
rect 151084 220056 151136 220108
rect 151820 220056 151872 220108
rect 152464 220056 152516 220108
rect 157340 220056 157392 220108
rect 204628 220056 204680 220108
rect 205088 220192 205140 220244
rect 242072 220192 242124 220244
rect 242624 220328 242676 220380
rect 273536 220328 273588 220380
rect 274364 220328 274416 220380
rect 276296 220328 276348 220380
rect 282552 220328 282604 220380
rect 298744 220328 298796 220380
rect 300768 220328 300820 220380
rect 305000 220328 305052 220380
rect 318432 220328 318484 220380
rect 322204 220328 322256 220380
rect 325608 220328 325660 220380
rect 328736 220328 328788 220380
rect 366456 220328 366508 220380
rect 381544 220328 381596 220380
rect 388444 220328 388496 220380
rect 404728 220328 404780 220380
rect 405004 220328 405056 220380
rect 437848 220328 437900 220380
rect 441436 220328 441488 220380
rect 495256 220328 495308 220380
rect 495394 220328 495446 220380
rect 504364 220328 504416 220380
rect 504548 220328 504600 220380
rect 511540 220328 511592 220380
rect 513380 220328 513432 220380
rect 515588 220328 515640 220380
rect 534724 220464 534776 220516
rect 542544 220464 542596 220516
rect 544568 220464 544620 220516
rect 548156 220464 548208 220516
rect 548524 220464 548576 220516
rect 572536 220464 572588 220516
rect 572674 220464 572726 220516
rect 590936 220464 590988 220516
rect 602896 220464 602948 220516
rect 532516 220328 532568 220380
rect 607220 220328 607272 220380
rect 307668 220260 307720 220312
rect 315856 220260 315908 220312
rect 242900 220192 242952 220244
rect 243544 220192 243596 220244
rect 252836 220192 252888 220244
rect 219348 220056 219400 220108
rect 219532 220056 219584 220108
rect 222476 220056 222528 220108
rect 223212 220056 223264 220108
rect 224500 220056 224552 220108
rect 224684 220056 224736 220108
rect 226616 220056 226668 220108
rect 101864 219920 101916 219972
rect 104808 219920 104860 219972
rect 113916 219920 113968 219972
rect 83924 219784 83976 219836
rect 88892 219784 88944 219836
rect 103152 219784 103204 219836
rect 118792 219784 118844 219836
rect 127624 219920 127676 219972
rect 166816 219920 166868 219972
rect 166954 219920 167006 219972
rect 187608 219920 187660 219972
rect 187792 219920 187844 219972
rect 231860 220056 231912 220108
rect 232688 220056 232740 220108
rect 259828 220192 259880 220244
rect 262956 220192 263008 220244
rect 284944 220192 284996 220244
rect 286140 220192 286192 220244
rect 293960 220192 294012 220244
rect 299204 220192 299256 220244
rect 303344 220192 303396 220244
rect 356888 220192 356940 220244
rect 365168 220192 365220 220244
rect 368112 220192 368164 220244
rect 385040 220192 385092 220244
rect 401416 220192 401468 220244
rect 434812 220192 434864 220244
rect 437480 220192 437532 220244
rect 450268 220192 450320 220244
rect 450912 220192 450964 220244
rect 512000 220192 512052 220244
rect 540336 220192 540388 220244
rect 622676 220192 622728 220244
rect 253572 220056 253624 220108
rect 264244 220056 264296 220108
rect 269580 220056 269632 220108
rect 287612 220056 287664 220108
rect 287796 220056 287848 220108
rect 288624 220056 288676 220108
rect 292304 220056 292356 220108
rect 299756 220056 299808 220108
rect 319260 220056 319312 220108
rect 323860 220056 323912 220108
rect 353208 220056 353260 220108
rect 361672 220056 361724 220108
rect 364156 220056 364208 220108
rect 378232 220056 378284 220108
rect 379520 220056 379572 220108
rect 401600 220056 401652 220108
rect 408132 220056 408184 220108
rect 444564 220056 444616 220108
rect 453948 220056 454000 220108
rect 463700 220056 463752 220108
rect 465080 220056 465132 220108
rect 475568 220056 475620 220108
rect 475752 220056 475804 220108
rect 480536 220056 480588 220108
rect 480720 220056 480772 220108
rect 481272 220056 481324 220108
rect 481456 220056 481508 220108
rect 542360 220056 542412 220108
rect 542544 219988 542596 220040
rect 548524 219988 548576 220040
rect 548892 219988 548944 220040
rect 601516 219988 601568 220040
rect 229836 219920 229888 219972
rect 243544 219920 243596 219972
rect 243728 219920 243780 219972
rect 262128 219920 262180 219972
rect 428096 219920 428148 219972
rect 451924 219920 451976 219972
rect 455696 219920 455748 219972
rect 507768 219920 507820 219972
rect 530400 219852 530452 219904
rect 562324 219852 562376 219904
rect 562508 219852 562560 219904
rect 562876 219852 562928 219904
rect 563060 219852 563112 219904
rect 567936 219852 567988 219904
rect 136916 219784 136968 219836
rect 137100 219784 137152 219836
rect 142068 219784 142120 219836
rect 142252 219784 142304 219836
rect 195336 219784 195388 219836
rect 195888 219784 195940 219836
rect 197452 219784 197504 219836
rect 201592 219784 201644 219836
rect 205088 219784 205140 219836
rect 206652 219784 206704 219836
rect 209688 219784 209740 219836
rect 209872 219784 209924 219836
rect 211436 219784 211488 219836
rect 211620 219784 211672 219836
rect 214380 219784 214432 219836
rect 214564 219784 214616 219836
rect 243360 219784 243412 219836
rect 322572 219716 322624 219768
rect 325976 219716 326028 219768
rect 70860 219648 70912 219700
rect 143080 219648 143132 219700
rect 143264 219648 143316 219700
rect 154488 219648 154540 219700
rect 154672 219648 154724 219700
rect 156788 219648 156840 219700
rect 156972 219648 157024 219700
rect 202328 219648 202380 219700
rect 202512 219648 202564 219700
rect 205272 219648 205324 219700
rect 205916 219648 205968 219700
rect 207204 219648 207256 219700
rect 209688 219648 209740 219700
rect 248144 219648 248196 219700
rect 254676 219648 254728 219700
rect 256516 219648 256568 219700
rect 421104 219648 421156 219700
rect 443000 219784 443052 219836
rect 436744 219648 436796 219700
rect 460204 219784 460256 219836
rect 463884 219784 463936 219836
rect 470968 219784 471020 219836
rect 471428 219784 471480 219836
rect 474464 219784 474516 219836
rect 264612 219580 264664 219632
rect 270224 219580 270276 219632
rect 311624 219580 311676 219632
rect 317788 219580 317840 219632
rect 324228 219580 324280 219632
rect 327724 219580 327776 219632
rect 88892 219512 88944 219564
rect 160928 219512 160980 219564
rect 161296 219512 161348 219564
rect 162584 219512 162636 219564
rect 163596 219512 163648 219564
rect 166908 219512 166960 219564
rect 169392 219512 169444 219564
rect 173808 219512 173860 219564
rect 174176 219512 174228 219564
rect 176568 219512 176620 219564
rect 177672 219512 177724 219564
rect 180524 219512 180576 219564
rect 181168 219512 181220 219564
rect 183284 219512 183336 219564
rect 183468 219512 183520 219564
rect 187792 219512 187844 219564
rect 187976 219512 188028 219564
rect 193036 219512 193088 219564
rect 118056 219376 118108 219428
rect 188160 219376 188212 219428
rect 190092 219376 190144 219428
rect 196716 219376 196768 219428
rect 201592 219376 201644 219428
rect 204628 219376 204680 219428
rect 210424 219376 210476 219428
rect 423772 219512 423824 219564
rect 445300 219512 445352 219564
rect 445668 219512 445720 219564
rect 466000 219648 466052 219700
rect 466460 219648 466512 219700
rect 505100 219784 505152 219836
rect 506572 219784 506624 219836
rect 509976 219784 510028 219836
rect 521660 219716 521712 219768
rect 522580 219716 522632 219768
rect 574928 219852 574980 219904
rect 575296 219852 575348 219904
rect 610348 219852 610400 219904
rect 568304 219716 568356 219768
rect 575664 219716 575716 219768
rect 575848 219716 575900 219768
rect 597560 219716 597612 219768
rect 666008 219716 666060 219768
rect 675300 219716 675352 219768
rect 475568 219648 475620 219700
rect 449072 219512 449124 219564
rect 453580 219512 453632 219564
rect 459744 219512 459796 219564
rect 231676 219444 231728 219496
rect 238116 219444 238168 219496
rect 240048 219444 240100 219496
rect 248052 219444 248104 219496
rect 249708 219444 249760 219496
rect 294420 219444 294472 219496
rect 298008 219444 298060 219496
rect 306012 219444 306064 219496
rect 307484 219444 307536 219496
rect 325056 219444 325108 219496
rect 326528 219444 326580 219496
rect 340696 219444 340748 219496
rect 345940 219444 345992 219496
rect 348884 219444 348936 219496
rect 355048 219444 355100 219496
rect 430396 219376 430448 219428
rect 475936 219376 475988 219428
rect 476580 219512 476632 219564
rect 481456 219512 481508 219564
rect 485872 219512 485924 219564
rect 495256 219512 495308 219564
rect 495532 219648 495584 219700
rect 504548 219648 504600 219700
rect 504732 219648 504784 219700
rect 506204 219580 506256 219632
rect 527824 219580 527876 219632
rect 563060 219580 563112 219632
rect 499948 219512 500000 219564
rect 476764 219376 476816 219428
rect 479892 219376 479944 219428
rect 490104 219376 490156 219428
rect 496820 219308 496872 219360
rect 535368 219444 535420 219496
rect 537484 219444 537536 219496
rect 548340 219444 548392 219496
rect 549996 219444 550048 219496
rect 112904 219240 112956 219292
rect 185400 219240 185452 219292
rect 431592 219240 431644 219292
rect 475752 219240 475804 219292
rect 483572 219240 483624 219292
rect 485780 219240 485832 219292
rect 515588 219240 515640 219292
rect 563060 219240 563112 219292
rect 563244 219240 563296 219292
rect 572168 219444 572220 219496
rect 575296 219444 575348 219496
rect 665088 219580 665140 219632
rect 675484 219580 675536 219632
rect 624148 219444 624200 219496
rect 564072 219308 564124 219360
rect 572996 219240 573048 219292
rect 609244 219240 609296 219292
rect 486424 219172 486476 219224
rect 498292 219172 498344 219224
rect 112260 219104 112312 219156
rect 186596 219104 186648 219156
rect 431776 219104 431828 219156
rect 476074 219104 476126 219156
rect 484676 219104 484728 219156
rect 485044 219104 485096 219156
rect 501052 219104 501104 219156
rect 596088 219104 596140 219156
rect 596272 219104 596324 219156
rect 627828 219104 627880 219156
rect 628012 219104 628064 219156
rect 628840 219104 628892 219156
rect 486148 219036 486200 219088
rect 494060 219036 494112 219088
rect 104808 218968 104860 219020
rect 176200 218968 176252 219020
rect 176568 218968 176620 219020
rect 181168 218968 181220 219020
rect 434352 218968 434404 219020
rect 485964 218968 486016 219020
rect 503168 218968 503220 219020
rect 503628 218968 503680 219020
rect 587900 218968 587952 219020
rect 591304 218968 591356 219020
rect 617248 218968 617300 219020
rect 106188 218832 106240 218884
rect 180984 218832 181036 218884
rect 448060 218832 448112 218884
rect 506572 218832 506624 218884
rect 539600 218832 539652 218884
rect 546132 218832 546184 218884
rect 546316 218832 546368 218884
rect 548524 218832 548576 218884
rect 552296 218832 552348 218884
rect 625528 218832 625580 218884
rect 105636 218696 105688 218748
rect 175832 218696 175884 218748
rect 176200 218696 176252 218748
rect 179696 218696 179748 218748
rect 445484 218696 445536 218748
rect 132960 218560 133012 218612
rect 199016 218560 199068 218612
rect 136272 218424 136324 218476
rect 200396 218424 200448 218476
rect 476396 218696 476448 218748
rect 481732 218696 481784 218748
rect 504364 218696 504416 218748
rect 528560 218696 528612 218748
rect 597376 218696 597428 218748
rect 597560 218696 597612 218748
rect 621664 218696 621716 218748
rect 508504 218560 508556 218612
rect 598480 218560 598532 218612
rect 498292 218424 498344 218476
rect 587532 218424 587584 218476
rect 146208 218288 146260 218340
rect 207756 218288 207808 218340
rect 494060 218288 494112 218340
rect 495256 218288 495308 218340
rect 571800 218288 571852 218340
rect 572444 218288 572496 218340
rect 580356 218288 580408 218340
rect 581644 218288 581696 218340
rect 591304 218424 591356 218476
rect 597376 218424 597428 218476
rect 597928 218424 597980 218476
rect 587900 218288 587952 218340
rect 597560 218288 597612 218340
rect 147588 218152 147640 218204
rect 207020 218152 207072 218204
rect 510712 218152 510764 218204
rect 599032 218152 599084 218204
rect 175832 218016 175884 218068
rect 182548 218016 182600 218068
rect 491668 218016 491720 218068
rect 563014 218016 563066 218068
rect 563152 218016 563204 218068
rect 573364 218016 573416 218068
rect 574468 218016 574520 218068
rect 581644 218016 581696 218068
rect 587532 218016 587584 218068
rect 595352 218016 595404 218068
rect 596180 218016 596232 218068
rect 596824 218016 596876 218068
rect 488540 217880 488592 217932
rect 594800 217880 594852 217932
rect 188436 217812 188488 217864
rect 188988 217812 189040 217864
rect 190920 217812 190972 217864
rect 191748 217812 191800 217864
rect 340972 217812 341024 217864
rect 341800 217812 341852 217864
rect 343916 217812 343968 217864
rect 344284 217812 344336 217864
rect 374000 217812 374052 217864
rect 374920 217812 374972 217864
rect 382464 217812 382516 217864
rect 383200 217812 383252 217864
rect 390744 217812 390796 217864
rect 391480 217812 391532 217864
rect 393320 217812 393372 217864
rect 393964 217812 394016 217864
rect 398840 217812 398892 217864
rect 399760 217812 399812 217864
rect 402980 217812 403032 217864
rect 403900 217812 403952 217864
rect 419540 217812 419592 217864
rect 420460 217812 420512 217864
rect 426440 217812 426492 217864
rect 427084 217812 427136 217864
rect 541716 217744 541768 217796
rect 542728 217744 542780 217796
rect 543096 217744 543148 217796
rect 544384 217744 544436 217796
rect 475936 217608 475988 217660
rect 477914 217608 477966 217660
rect 514760 217608 514812 217660
rect 516002 217608 516054 217660
rect 519176 217608 519228 217660
rect 520142 217608 520194 217660
rect 537668 217608 537720 217660
rect 546316 217744 546368 217796
rect 548524 217744 548576 217796
rect 553492 217744 553544 217796
rect 556804 217744 556856 217796
rect 607864 217744 607916 217796
rect 545580 217608 545632 217660
rect 570420 217608 570472 217660
rect 573364 217608 573416 217660
rect 609888 217608 609940 217660
rect 475752 217472 475804 217524
rect 481226 217472 481278 217524
rect 538680 217472 538732 217524
rect 541716 217472 541768 217524
rect 542176 217472 542228 217524
rect 543096 217472 543148 217524
rect 543326 217472 543378 217524
rect 42064 217268 42116 217320
rect 62764 217268 62816 217320
rect 33048 217200 33100 217252
rect 41512 217200 41564 217252
rect 110420 217200 110472 217252
rect 185216 217200 185268 217252
rect 545580 217336 545632 217388
rect 605288 217472 605340 217524
rect 548524 217336 548576 217388
rect 607404 217404 607456 217456
rect 610348 217404 610400 217456
rect 620560 217404 620612 217456
rect 607220 217268 607272 217320
rect 621112 217268 621164 217320
rect 100668 217064 100720 217116
rect 178040 217064 178092 217116
rect 510344 217064 510396 217116
rect 538220 217200 538272 217252
rect 602068 217200 602120 217252
rect 526444 217064 526496 217116
rect 531228 217064 531280 217116
rect 536196 217064 536248 217116
rect 567844 217064 567896 217116
rect 570420 217064 570472 217116
rect 616144 217064 616196 217116
rect 93860 216928 93912 216980
rect 174360 216928 174412 216980
rect 453396 216928 453448 216980
rect 516508 216928 516560 216980
rect 531228 216928 531280 216980
rect 573548 216928 573600 216980
rect 573732 216928 573784 216980
rect 575296 216928 575348 216980
rect 90732 216792 90784 216844
rect 171140 216792 171192 216844
rect 457536 216792 457588 216844
rect 521660 216792 521712 216844
rect 525432 216792 525484 216844
rect 531872 216792 531924 216844
rect 538036 216792 538088 216844
rect 539784 216792 539836 216844
rect 540980 216792 541032 216844
rect 603080 216792 603132 216844
rect 614028 216792 614080 216844
rect 614488 216792 614540 216844
rect 671988 216792 672040 216844
rect 675300 216792 675352 216844
rect 85580 216656 85632 216708
rect 168656 216656 168708 216708
rect 516140 216656 516192 216708
rect 518624 216656 518676 216708
rect 520280 216656 520332 216708
rect 525432 216520 525484 216572
rect 485504 216384 485556 216436
rect 500592 216384 500644 216436
rect 516140 216384 516192 216436
rect 516324 216384 516376 216436
rect 48964 215296 49016 215348
rect 35808 214820 35860 214872
rect 41512 214820 41564 214872
rect 43168 214752 43220 214804
rect 49332 214752 49384 214804
rect 518624 216384 518676 216436
rect 518808 216384 518860 216436
rect 520648 216384 520700 216436
rect 521200 216384 521252 216436
rect 526076 216384 526128 216436
rect 526444 216384 526496 216436
rect 531412 216520 531464 216572
rect 532700 216520 532752 216572
rect 533712 216520 533764 216572
rect 539600 216520 539652 216572
rect 539784 216520 539836 216572
rect 542176 216520 542228 216572
rect 542728 216452 542780 216504
rect 531228 216384 531280 216436
rect 531872 216384 531924 216436
rect 537392 216384 537444 216436
rect 537668 216384 537720 216436
rect 538036 216384 538088 216436
rect 538680 216384 538732 216436
rect 541164 216384 541216 216436
rect 541992 216384 542044 216436
rect 543004 216384 543056 216436
rect 543464 216384 543516 216436
rect 543648 216384 543700 216436
rect 545120 216384 545172 216436
rect 545488 216384 545540 216436
rect 545672 216384 545724 216436
rect 547972 216520 548024 216572
rect 546776 216384 546828 216436
rect 552664 216384 552716 216436
rect 553952 216384 554004 216436
rect 566188 216656 566240 216708
rect 618352 216656 618404 216708
rect 670424 216656 670476 216708
rect 675484 216656 675536 216708
rect 562508 216520 562560 216572
rect 600780 216452 600832 216504
rect 600964 216452 601016 216504
rect 606760 216452 606812 216504
rect 566188 216384 566240 216436
rect 567844 216384 567896 216436
rect 573732 216384 573784 216436
rect 574008 216316 574060 216368
rect 627184 216316 627236 216368
rect 600964 216180 601016 216232
rect 576584 216044 576636 216096
rect 576768 216044 576820 216096
rect 600780 216044 600832 216096
rect 616696 216180 616748 216232
rect 602896 216044 602948 216096
rect 626080 216044 626132 216096
rect 601240 215908 601292 215960
rect 601516 215908 601568 215960
rect 623780 215908 623832 215960
rect 599584 215840 599636 215892
rect 576814 215704 576866 215756
rect 596272 215704 596324 215756
rect 596456 215704 596508 215756
rect 600688 215704 600740 215756
rect 573916 215568 573968 215620
rect 586474 215432 586526 215484
rect 586704 215432 586756 215484
rect 595996 215432 596048 215484
rect 596640 215568 596692 215620
rect 614120 215568 614172 215620
rect 600320 215432 600372 215484
rect 600504 215432 600556 215484
rect 604000 215432 604052 215484
rect 673920 215432 673972 215484
rect 675484 215432 675536 215484
rect 573732 215296 573784 215348
rect 576584 215296 576636 215348
rect 664168 215296 664220 215348
rect 675300 215296 675352 215348
rect 673736 215160 673788 215212
rect 581644 215092 581696 215144
rect 616880 215092 616932 215144
rect 576032 214956 576084 215008
rect 581460 214956 581512 215008
rect 618904 214956 618956 215008
rect 575664 214820 575716 214872
rect 620008 214820 620060 214872
rect 573916 214684 573968 214736
rect 574744 214684 574796 214736
rect 574928 214684 574980 214736
rect 581460 214684 581512 214736
rect 573732 214548 573784 214600
rect 575848 214548 575900 214600
rect 619640 214684 619692 214736
rect 574836 214412 574888 214464
rect 575296 214412 575348 214464
rect 622400 214548 622452 214600
rect 655520 214548 655572 214600
rect 656440 214548 656492 214600
rect 659660 214548 659712 214600
rect 660304 214548 660356 214600
rect 661316 214548 661368 214600
rect 661960 214548 662012 214600
rect 608784 214412 608836 214464
rect 609520 214412 609572 214464
rect 575112 214276 575164 214328
rect 581644 214276 581696 214328
rect 35808 214072 35860 214124
rect 39948 214072 40000 214124
rect 673092 214072 673144 214124
rect 675484 214072 675536 214124
rect 580356 213868 580408 213920
rect 595720 213868 595772 213920
rect 574652 213732 574704 213784
rect 595168 213732 595220 213784
rect 595352 213732 595404 213784
rect 596364 213868 596416 213920
rect 603080 213868 603132 213920
rect 605932 213868 605984 213920
rect 609244 213868 609296 213920
rect 610624 213868 610676 213920
rect 624148 213868 624200 213920
rect 625252 213868 625304 213920
rect 628564 213868 628616 213920
rect 633808 213868 633860 213920
rect 639972 213868 640024 213920
rect 651380 213868 651432 213920
rect 602068 213732 602120 213784
rect 605104 213732 605156 213784
rect 605288 213732 605340 213784
rect 606208 213732 606260 213784
rect 638868 213732 638920 213784
rect 650000 213732 650052 213784
rect 671804 213664 671856 213716
rect 675484 213664 675536 213716
rect 574468 213596 574520 213648
rect 603632 213596 603684 213648
rect 638316 213596 638368 213648
rect 651748 213596 651800 213648
rect 574100 213460 574152 213512
rect 604552 213460 604604 213512
rect 636660 213460 636712 213512
rect 650184 213460 650236 213512
rect 575480 213324 575532 213376
rect 629392 213324 629444 213376
rect 635556 213324 635608 213376
rect 649080 213324 649132 213376
rect 672264 213256 672316 213308
rect 675484 213256 675536 213308
rect 574836 213188 574888 213240
rect 630680 213188 630732 213240
rect 637212 213188 637264 213240
rect 650736 213188 650788 213240
rect 640248 213052 640300 213104
rect 650920 213052 650972 213104
rect 616696 212984 616748 213036
rect 623320 212984 623372 213036
rect 35808 212916 35860 212968
rect 40316 212916 40368 212968
rect 641628 212916 641680 212968
rect 650368 212916 650420 212968
rect 632704 212780 632756 212832
rect 634360 212780 634412 212832
rect 35624 212644 35676 212696
rect 40684 212644 40736 212696
rect 630036 212644 630088 212696
rect 632704 212644 632756 212696
rect 35440 212508 35492 212560
rect 39948 212508 40000 212560
rect 579252 211964 579304 212016
rect 581920 211964 581972 212016
rect 675852 211760 675904 211812
rect 683120 211760 683172 211812
rect 35808 211556 35860 211608
rect 40960 211556 41012 211608
rect 35808 211284 35860 211336
rect 39672 211352 39724 211404
rect 578516 211284 578568 211336
rect 583300 211284 583352 211336
rect 35624 211148 35676 211200
rect 41512 211148 41564 211200
rect 42340 211148 42392 211200
rect 51724 211148 51776 211200
rect 578884 211148 578936 211200
rect 580908 211148 580960 211200
rect 664812 211080 664864 211132
rect 667572 211080 667624 211132
rect 644480 211012 644532 211064
rect 644848 211012 644900 211064
rect 652024 210400 652076 210452
rect 670976 210264 671028 210316
rect 608600 210060 608652 210112
rect 608968 210060 609020 210112
rect 35808 209924 35860 209976
rect 40040 209924 40092 209976
rect 35624 209788 35676 209840
rect 41696 209788 41748 209840
rect 579252 209788 579304 209840
rect 581644 209788 581696 209840
rect 591304 209788 591356 209840
rect 632152 209788 632204 209840
rect 652208 209516 652260 209568
rect 669412 209040 669464 209092
rect 35808 208700 35860 208752
rect 39948 208632 40000 208684
rect 35808 208360 35860 208412
rect 41696 208360 41748 208412
rect 42064 208360 42116 208412
rect 43076 208360 43128 208412
rect 578700 208292 578752 208344
rect 589464 208292 589516 208344
rect 669596 208088 669648 208140
rect 675484 208088 675536 208140
rect 578424 208020 578476 208072
rect 580632 208020 580684 208072
rect 35808 207272 35860 207324
rect 40132 207272 40184 207324
rect 35532 207000 35584 207052
rect 40960 207000 41012 207052
rect 581920 206932 581972 206984
rect 589464 206932 589516 206984
rect 35808 205912 35860 205964
rect 39764 205912 39816 205964
rect 674840 205708 674892 205760
rect 675392 205708 675444 205760
rect 35808 205640 35860 205692
rect 41696 205640 41748 205692
rect 42064 205640 42116 205692
rect 43444 205640 43496 205692
rect 578700 205640 578752 205692
rect 581828 205640 581880 205692
rect 583300 205572 583352 205624
rect 589464 205572 589516 205624
rect 579068 205232 579120 205284
rect 584404 205232 584456 205284
rect 35808 204892 35860 204944
rect 40776 204892 40828 204944
rect 35624 204620 35676 204672
rect 41696 204688 41748 204740
rect 42064 204688 42116 204740
rect 44364 204688 44416 204740
rect 42064 204552 42116 204604
rect 50344 204552 50396 204604
rect 35808 204484 35860 204536
rect 41696 204484 41748 204536
rect 35532 204280 35584 204332
rect 41696 204280 41748 204332
rect 42064 204280 42116 204332
rect 48964 204280 49016 204332
rect 580908 204144 580960 204196
rect 589464 204144 589516 204196
rect 35624 203124 35676 203176
rect 41604 203124 41656 203176
rect 35808 202852 35860 202904
rect 40040 202852 40092 202904
rect 578700 202852 578752 202904
rect 583208 202852 583260 202904
rect 581644 202716 581696 202768
rect 589372 202716 589424 202768
rect 578240 201628 578292 201680
rect 580908 201628 580960 201680
rect 673920 201424 673972 201476
rect 675392 201424 675444 201476
rect 671804 201220 671856 201272
rect 675116 201220 675168 201272
rect 581828 200744 581880 200796
rect 590384 200744 590436 200796
rect 673736 200744 673788 200796
rect 674932 200744 674984 200796
rect 578516 200404 578568 200456
rect 581736 200404 581788 200456
rect 580632 199996 580684 200048
rect 589464 199996 589516 200048
rect 578884 198704 578936 198756
rect 583024 198704 583076 198756
rect 671988 198636 672040 198688
rect 675300 198636 675352 198688
rect 673092 197752 673144 197804
rect 675300 197752 675352 197804
rect 578332 197412 578384 197464
rect 580264 197412 580316 197464
rect 668032 197344 668084 197396
rect 670148 197344 670200 197396
rect 584404 197276 584456 197328
rect 589464 197276 589516 197328
rect 581736 196596 581788 196648
rect 589648 196596 589700 196648
rect 579252 196120 579304 196172
rect 581644 196120 581696 196172
rect 583208 195916 583260 195968
rect 589464 195916 589516 195968
rect 42432 195644 42484 195696
rect 43628 195644 43680 195696
rect 580908 194488 580960 194540
rect 589464 194488 589516 194540
rect 578516 193400 578568 193452
rect 583760 193400 583812 193452
rect 42432 193128 42484 193180
rect 43812 193128 43864 193180
rect 579528 191836 579580 191888
rect 588544 191836 588596 191888
rect 42432 191768 42484 191820
rect 44548 191768 44600 191820
rect 42432 191632 42484 191684
rect 44364 191632 44416 191684
rect 583760 191088 583812 191140
rect 590384 191088 590436 191140
rect 583024 190408 583076 190460
rect 589464 190408 589516 190460
rect 42432 190340 42484 190392
rect 42984 190340 43036 190392
rect 669274 190272 669326 190324
rect 675300 190272 675352 190324
rect 578240 189048 578292 189100
rect 585968 189048 586020 189100
rect 581644 188912 581696 188964
rect 589464 188912 589516 188964
rect 579252 188776 579304 188828
rect 581828 188776 581880 188828
rect 42432 187620 42484 187672
rect 43444 187620 43496 187672
rect 580264 187552 580316 187604
rect 589372 187552 589424 187604
rect 578516 187144 578568 187196
rect 584588 187144 584640 187196
rect 578884 186192 578936 186244
rect 589464 186192 589516 186244
rect 578332 185240 578384 185292
rect 580448 185240 580500 185292
rect 668216 184832 668268 184884
rect 672540 184832 672592 184884
rect 579528 183540 579580 183592
rect 587164 183540 587216 183592
rect 42432 183472 42484 183524
rect 44180 183472 44232 183524
rect 578884 182180 578936 182232
rect 583024 182180 583076 182232
rect 578516 181296 578568 181348
rect 581644 181296 581696 181348
rect 585968 180752 586020 180804
rect 589464 180752 589516 180804
rect 578976 179664 579028 179716
rect 585784 179664 585836 179716
rect 581828 179256 581880 179308
rect 589556 179256 589608 179308
rect 578608 178304 578660 178356
rect 580264 178304 580316 178356
rect 667388 178236 667440 178288
rect 675484 178236 675536 178288
rect 670976 178100 671028 178152
rect 675484 178100 675536 178152
rect 584588 177964 584640 178016
rect 589464 177964 589516 178016
rect 668584 177964 668636 178016
rect 672540 177964 672592 178016
rect 673552 177692 673604 177744
rect 675484 177692 675536 177744
rect 579528 176808 579580 176860
rect 584404 176808 584456 176860
rect 673920 176808 673972 176860
rect 675484 176808 675536 176860
rect 580448 176536 580500 176588
rect 589464 176536 589516 176588
rect 667848 175380 667900 175432
rect 675484 175380 675536 175432
rect 673368 175176 673420 175228
rect 675484 175176 675536 175228
rect 579620 174496 579672 174548
rect 589924 174496 589976 174548
rect 673000 174360 673052 174412
rect 675484 174360 675536 174412
rect 587164 173816 587216 173868
rect 589280 173816 589332 173868
rect 578332 172524 578384 172576
rect 583208 172524 583260 172576
rect 583024 172388 583076 172440
rect 589372 172388 589424 172440
rect 579068 171640 579120 171692
rect 581828 171640 581880 171692
rect 670424 171096 670476 171148
rect 675484 171096 675536 171148
rect 581644 170960 581696 171012
rect 589464 170960 589516 171012
rect 579528 169736 579580 169788
rect 588728 169736 588780 169788
rect 585784 169600 585836 169652
rect 589464 169600 589516 169652
rect 671804 169464 671856 169516
rect 675484 169464 675536 169516
rect 670608 169056 670660 169108
rect 675484 169056 675536 169108
rect 673184 168648 673236 168700
rect 675484 168648 675536 168700
rect 578240 168376 578292 168428
rect 580448 168376 580500 168428
rect 580264 168240 580316 168292
rect 589464 168240 589516 168292
rect 672632 167016 672684 167068
rect 675484 167016 675536 167068
rect 669964 166812 670016 166864
rect 675484 166812 675536 166864
rect 579620 166268 579672 166320
rect 590384 166268 590436 166320
rect 579068 165588 579120 165640
rect 584588 165588 584640 165640
rect 584404 165452 584456 165504
rect 589464 165520 589516 165572
rect 579528 164296 579580 164348
rect 583024 164296 583076 164348
rect 578700 162868 578752 162920
rect 581644 162868 581696 162920
rect 583208 162800 583260 162852
rect 589464 162800 589516 162852
rect 671804 162052 671856 162104
rect 673552 162052 673604 162104
rect 581828 161372 581880 161424
rect 589464 161372 589516 161424
rect 578516 160216 578568 160268
rect 580264 160216 580316 160268
rect 579528 158720 579580 158772
rect 588544 158720 588596 158772
rect 580448 158584 580500 158636
rect 589464 158584 589516 158636
rect 579620 156612 579672 156664
rect 589924 156612 589976 156664
rect 673552 155796 673604 155848
rect 675392 155796 675444 155848
rect 670424 154912 670476 154964
rect 675116 154912 675168 154964
rect 579252 154572 579304 154624
rect 587348 154572 587400 154624
rect 584588 154436 584640 154488
rect 589372 154436 589424 154488
rect 579252 153280 579304 153332
rect 585784 153280 585836 153332
rect 583024 153076 583076 153128
rect 589464 153076 589516 153128
rect 578700 152260 578752 152312
rect 584404 152260 584456 152312
rect 673184 151716 673236 151768
rect 675116 151716 675168 151768
rect 581644 151648 581696 151700
rect 589464 151648 589516 151700
rect 579160 150424 579212 150476
rect 583208 150424 583260 150476
rect 670608 150356 670660 150408
rect 674932 150356 674984 150408
rect 578884 150288 578936 150340
rect 589464 150288 589516 150340
rect 578884 149064 578936 149116
rect 581644 149064 581696 149116
rect 674472 148928 674524 148980
rect 675300 148928 675352 148980
rect 668768 148180 668820 148232
rect 674104 148180 674156 148232
rect 579528 147636 579580 147688
rect 588728 147636 588780 147688
rect 579252 147500 579304 147552
rect 591304 147500 591356 147552
rect 580264 147364 580316 147416
rect 589464 147364 589516 147416
rect 668768 146208 668820 146260
rect 671436 146208 671488 146260
rect 579620 144168 579672 144220
rect 590384 144168 590436 144220
rect 668768 144168 668820 144220
rect 674288 144168 674340 144220
rect 578516 143624 578568 143676
rect 580264 143624 580316 143676
rect 587348 143488 587400 143540
rect 590016 143488 590068 143540
rect 579528 142128 579580 142180
rect 587164 142128 587216 142180
rect 585784 141992 585836 142044
rect 589464 141992 589516 142044
rect 584404 140700 584456 140752
rect 589464 140700 589516 140752
rect 668768 140700 668820 140752
rect 671620 140700 671672 140752
rect 579528 139408 579580 139460
rect 584588 139408 584640 139460
rect 668768 139340 668820 139392
rect 671160 139340 671212 139392
rect 668032 137980 668084 138032
rect 672172 137980 672224 138032
rect 579252 137912 579304 137964
rect 583024 137912 583076 137964
rect 583208 137912 583260 137964
rect 589464 137912 589516 137964
rect 668584 137300 668636 137352
rect 669136 137300 669188 137352
rect 581644 136484 581696 136536
rect 589372 136484 589424 136536
rect 579068 135328 579120 135380
rect 581092 135328 581144 135380
rect 578240 134512 578292 134564
rect 585968 134512 586020 134564
rect 669228 133764 669280 133816
rect 672816 133764 672868 133816
rect 669412 133356 669464 133408
rect 675484 133356 675536 133408
rect 581092 133152 581144 133204
rect 589924 133152 589976 133204
rect 578516 132880 578568 132932
rect 581644 132880 581696 132932
rect 667204 132880 667256 132932
rect 675484 132880 675536 132932
rect 667572 132744 667624 132796
rect 675484 132744 675536 132796
rect 580264 132336 580316 132388
rect 589464 132336 589516 132388
rect 673920 132132 673972 132184
rect 675484 132132 675536 132184
rect 668400 131180 668452 131232
rect 668768 131180 668820 131232
rect 675484 131180 675536 131232
rect 668308 131044 668360 131096
rect 670240 131044 670292 131096
rect 671344 130840 671396 130892
rect 675484 130840 675536 130892
rect 673368 130500 673420 130552
rect 675484 130500 675536 130552
rect 578424 130364 578476 130416
rect 588544 130364 588596 130416
rect 578608 129888 578660 129940
rect 580448 129888 580500 129940
rect 668584 129888 668636 129940
rect 675484 129888 675536 129940
rect 584588 129684 584640 129736
rect 589464 129684 589516 129736
rect 673000 129684 673052 129736
rect 675484 129684 675536 129736
rect 669228 129616 669280 129668
rect 672356 129616 672408 129668
rect 668216 129208 668268 129260
rect 669780 129208 669832 129260
rect 578884 128324 578936 128376
rect 668952 128324 669004 128376
rect 675484 128324 675536 128376
rect 589464 128188 589516 128240
rect 578332 126964 578384 127016
rect 580264 126964 580316 127016
rect 587164 126896 587216 126948
rect 589740 126896 589792 126948
rect 579436 126216 579488 126268
rect 587348 126216 587400 126268
rect 675024 126148 675076 126200
rect 675484 126148 675536 126200
rect 675852 126148 675904 126200
rect 676404 126148 676456 126200
rect 673184 125944 673236 125996
rect 675484 125944 675536 125996
rect 578516 125808 578568 125860
rect 584404 125808 584456 125860
rect 673000 125740 673052 125792
rect 675484 125740 675536 125792
rect 585968 124856 586020 124908
rect 590384 124856 590436 124908
rect 578884 124176 578936 124228
rect 585784 124176 585836 124228
rect 583024 124040 583076 124092
rect 589464 124040 589516 124092
rect 673368 123904 673420 123956
rect 675484 123904 675536 123956
rect 674012 123088 674064 123140
rect 675484 123088 675536 123140
rect 670148 122408 670200 122460
rect 675484 122408 675536 122460
rect 579528 121456 579580 121508
rect 583024 121456 583076 121508
rect 671528 121388 671580 121440
rect 675484 121388 675536 121440
rect 580264 120708 580316 120760
rect 589924 120708 589976 120760
rect 581644 120028 581696 120080
rect 589464 120028 589516 120080
rect 669228 120028 669280 120080
rect 671804 120028 671856 120080
rect 579252 118668 579304 118720
rect 587164 118668 587216 118720
rect 579068 117308 579120 117360
rect 581644 117308 581696 117360
rect 675852 117240 675904 117292
rect 679624 117240 679676 117292
rect 580448 117172 580500 117224
rect 589464 117172 589516 117224
rect 578332 116968 578384 117020
rect 580264 116968 580316 117020
rect 587348 115880 587400 115932
rect 589280 115880 589332 115932
rect 669228 115812 669280 115864
rect 672632 115812 672684 115864
rect 675024 115472 675076 115524
rect 675392 115472 675444 115524
rect 585784 114452 585836 114504
rect 589464 114452 589516 114504
rect 669228 114112 669280 114164
rect 674012 114112 674064 114164
rect 668308 112820 668360 112872
rect 670148 112820 670200 112872
rect 584404 111732 584456 111784
rect 589464 111732 589516 111784
rect 669044 111732 669096 111784
rect 671528 111732 671580 111784
rect 673184 111732 673236 111784
rect 675116 111732 675168 111784
rect 673000 111120 673052 111172
rect 675392 111120 675444 111172
rect 578884 108944 578936 108996
rect 589464 108944 589516 108996
rect 669136 108944 669188 108996
rect 671344 108944 671396 108996
rect 583024 107584 583076 107636
rect 589372 107584 589424 107636
rect 674196 106972 674248 107024
rect 675300 106972 675352 107024
rect 673368 106496 673420 106548
rect 675116 106496 675168 106548
rect 587164 106224 587216 106276
rect 589280 106224 589332 106276
rect 581644 104796 581696 104848
rect 589372 104796 589424 104848
rect 580264 102076 580316 102128
rect 589464 102076 589516 102128
rect 623688 99152 623740 99204
rect 632152 99152 632204 99204
rect 625068 99016 625120 99068
rect 634452 99016 634504 99068
rect 629760 98880 629812 98932
rect 640984 98880 641036 98932
rect 621664 98744 621716 98796
rect 628380 98744 628432 98796
rect 629024 98744 629076 98796
rect 639880 98744 639932 98796
rect 622308 98608 622360 98660
rect 629484 98608 629536 98660
rect 630496 98608 630548 98660
rect 642088 98608 642140 98660
rect 577504 97928 577556 97980
rect 594064 97928 594116 97980
rect 596180 97928 596232 97980
rect 624608 97928 624660 97980
rect 632980 97928 633032 97980
rect 634176 97928 634228 97980
rect 643376 97928 643428 97980
rect 595260 97792 595312 97844
rect 595628 97792 595680 97844
rect 626080 97792 626132 97844
rect 635280 97792 635332 97844
rect 592684 97656 592736 97708
rect 597560 97656 597612 97708
rect 620192 97656 620244 97708
rect 626080 97656 626132 97708
rect 633348 97656 633400 97708
rect 643560 97792 643612 97844
rect 639328 97656 639380 97708
rect 595444 97520 595496 97572
rect 600412 97520 600464 97572
rect 623136 97520 623188 97572
rect 630680 97520 630732 97572
rect 632704 97520 632756 97572
rect 618720 97384 618772 97436
rect 626264 97384 626316 97436
rect 627552 97384 627604 97436
rect 637580 97384 637632 97436
rect 578884 97248 578936 97300
rect 598940 97248 598992 97300
rect 605472 97248 605524 97300
rect 611912 97248 611964 97300
rect 628196 97248 628248 97300
rect 639052 97248 639104 97300
rect 647148 97656 647200 97708
rect 659752 97928 659804 97980
rect 659936 97928 659988 97980
rect 665180 97928 665232 97980
rect 655428 97792 655480 97844
rect 662512 97792 662564 97844
rect 651840 97656 651892 97708
rect 659568 97656 659620 97708
rect 659752 97656 659804 97708
rect 661960 97656 662012 97708
rect 644296 97520 644348 97572
rect 646504 97384 646556 97436
rect 658832 97520 658884 97572
rect 658188 97384 658240 97436
rect 663064 97384 663116 97436
rect 644756 97248 644808 97300
rect 656808 97248 656860 97300
rect 661408 97248 661460 97300
rect 651104 97180 651156 97232
rect 654324 97180 654376 97232
rect 626816 97112 626868 97164
rect 636384 97112 636436 97164
rect 650368 96976 650420 97028
rect 658280 96976 658332 97028
rect 601056 96908 601108 96960
rect 601884 96908 601936 96960
rect 606208 96908 606260 96960
rect 606944 96908 606996 96960
rect 612648 96908 612700 96960
rect 613384 96908 613436 96960
rect 614028 96908 614080 96960
rect 614764 96908 614816 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 645216 96908 645268 96960
rect 645768 96908 645820 96960
rect 609152 96840 609204 96892
rect 609704 96840 609756 96892
rect 646688 96840 646740 96892
rect 647148 96840 647200 96892
rect 654784 96840 654836 96892
rect 655244 96840 655296 96892
rect 656716 96840 656768 96892
rect 660120 96908 660172 96960
rect 613568 96772 613620 96824
rect 614028 96772 614080 96824
rect 641536 96772 641588 96824
rect 642824 96772 642876 96824
rect 612096 96704 612148 96756
rect 612556 96704 612608 96756
rect 617248 96704 617300 96756
rect 618076 96704 618128 96756
rect 643008 96704 643060 96756
rect 660120 96704 660172 96756
rect 642272 96568 642324 96620
rect 644112 96568 644164 96620
rect 638592 96432 638644 96484
rect 651288 96568 651340 96620
rect 652576 96568 652628 96620
rect 654968 96568 655020 96620
rect 653312 96432 653364 96484
rect 663984 96432 664036 96484
rect 631232 96296 631284 96348
rect 642640 96296 642692 96348
rect 642824 96296 642876 96348
rect 648804 96296 648856 96348
rect 648988 96296 649040 96348
rect 620928 96228 620980 96280
rect 626448 96228 626500 96280
rect 631876 96160 631928 96212
rect 644480 96160 644532 96212
rect 610624 96024 610676 96076
rect 621664 96024 621716 96076
rect 635648 96024 635700 96076
rect 608416 95888 608468 95940
rect 620284 95888 620336 95940
rect 637764 95888 637816 95940
rect 634728 95548 634780 95600
rect 640064 96024 640116 96076
rect 652024 96160 652076 96212
rect 654968 96296 655020 96348
rect 665548 96296 665600 96348
rect 663800 96160 663852 96212
rect 649264 96024 649316 96076
rect 660672 96024 660724 96076
rect 640800 95888 640852 95940
rect 665364 95888 665416 95940
rect 642824 95752 642876 95804
rect 645584 95616 645636 95668
rect 656164 95616 656216 95668
rect 659200 95616 659252 95668
rect 664168 95616 664220 95668
rect 649264 95480 649316 95532
rect 643100 95344 643152 95396
rect 616512 95140 616564 95192
rect 623044 95140 623096 95192
rect 649632 95140 649684 95192
rect 650644 95140 650696 95192
rect 643744 94596 643796 94648
rect 653404 94596 653456 94648
rect 607680 94460 607732 94512
rect 624976 94460 625028 94512
rect 642916 94460 642968 94512
rect 663248 94460 663300 94512
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 644112 93780 644164 93832
rect 654140 93712 654192 93764
rect 609704 93100 609756 93152
rect 618904 93100 618956 93152
rect 617892 92420 617944 92472
rect 625436 92420 625488 92472
rect 651288 92420 651340 92472
rect 654324 92420 654376 92472
rect 611268 90992 611320 91044
rect 617340 90992 617392 91044
rect 618076 90992 618128 91044
rect 626448 90992 626500 91044
rect 646504 90992 646556 91044
rect 654140 90992 654192 91044
rect 623044 89632 623096 89684
rect 626448 89632 626500 89684
rect 647148 88952 647200 89004
rect 656900 88952 656952 89004
rect 656164 88748 656216 88800
rect 657452 88748 657504 88800
rect 662328 88748 662380 88800
rect 664168 88748 664220 88800
rect 656716 88612 656768 88664
rect 659292 88612 659344 88664
rect 607312 88272 607364 88324
rect 626448 88272 626500 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 617340 88136 617392 88188
rect 625620 88136 625672 88188
rect 648160 87116 648212 87168
rect 662512 87116 662564 87168
rect 645768 86980 645820 87032
rect 660672 86980 660724 87032
rect 652024 86708 652076 86760
rect 660120 86708 660172 86760
rect 653404 86572 653456 86624
rect 661408 86572 661460 86624
rect 650644 86436 650696 86488
rect 658832 86436 658884 86488
rect 621664 86232 621716 86284
rect 626448 86232 626500 86284
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 620284 84124 620336 84176
rect 626264 84124 626316 84176
rect 618904 83988 618956 84040
rect 626448 83920 626500 83972
rect 628564 80928 628616 80980
rect 642456 80928 642508 80980
rect 612556 80792 612608 80844
rect 645860 80792 645912 80844
rect 595628 80656 595680 80708
rect 636108 80656 636160 80708
rect 629208 79432 629260 79484
rect 637488 79432 637540 79484
rect 616788 79296 616840 79348
rect 647424 79296 647476 79348
rect 637488 78208 637540 78260
rect 645308 78208 645360 78260
rect 631048 78072 631100 78124
rect 638960 78072 639012 78124
rect 614028 77936 614080 77988
rect 647608 77936 647660 77988
rect 591304 77392 591356 77444
rect 631048 77664 631100 77716
rect 628288 77528 628340 77580
rect 631508 77528 631560 77580
rect 625804 77392 625856 77444
rect 633900 77392 633952 77444
rect 577504 77256 577556 77308
rect 637120 77256 637172 77308
rect 639604 77256 639656 77308
rect 614764 76644 614816 76696
rect 646320 76644 646372 76696
rect 613384 76508 613436 76560
rect 649172 76508 649224 76560
rect 580264 75896 580316 75948
rect 628288 75896 628340 75948
rect 615408 75284 615460 75336
rect 646136 75284 646188 75336
rect 607128 75148 607180 75200
rect 646872 75148 646924 75200
rect 612004 57196 612056 57248
rect 662420 57196 662472 57248
rect 145380 52912 145432 52964
rect 580264 53048 580316 53100
rect 288164 52368 288216 52420
rect 625804 52368 625856 52420
rect 391940 52232 391992 52284
rect 392584 52232 392636 52284
rect 577504 52232 577556 52284
rect 235816 51008 235868 51060
rect 288164 51008 288216 51060
rect 340512 51008 340564 51060
rect 391940 51008 391992 51060
rect 405096 50464 405148 50516
rect 578884 50464 578936 50516
rect 183468 50328 183520 50380
rect 406384 50328 406436 50380
rect 461032 47200 461084 47252
rect 465908 47200 465960 47252
rect 194048 44820 194100 44872
rect 661592 44820 661644 44872
rect 315948 43392 316000 43444
rect 661132 43392 661184 43444
rect 464896 42328 464948 42380
rect 315948 42173 316000 42225
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366180 1027880 366232 1027886
rect 366180 1027822 366232 1027828
rect 366548 1027880 366600 1027886
rect 366548 1027822 366600 1027828
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366192 1027752 366220 1027822
rect 366560 1027752 366588 1027822
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366192 1024418 366220 1024488
rect 366560 1024418 366588 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366180 1024412 366232 1024418
rect 366180 1024354 366232 1024360
rect 366548 1024412 366600 1024418
rect 366548 1024354 366600 1024360
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 505008 1007208 505060 1007214
rect 357714 1007176 357770 1007185
rect 505006 1007176 505008 1007185
rect 513840 1007208 513892 1007214
rect 505060 1007176 505062 1007185
rect 357714 1007111 357716 1007120
rect 357768 1007111 357770 1007120
rect 368940 1007140 368992 1007146
rect 357716 1007082 357768 1007088
rect 513840 1007150 513892 1007156
rect 505006 1007111 505062 1007120
rect 368940 1007082 368992 1007088
rect 357716 1006936 357768 1006942
rect 357714 1006904 357716 1006913
rect 357768 1006904 357770 1006913
rect 357714 1006839 357770 1006848
rect 358544 1006800 358596 1006806
rect 358542 1006768 358544 1006777
rect 358596 1006768 358598 1006777
rect 358542 1006703 358598 1006712
rect 103150 1006632 103206 1006641
rect 94688 1006596 94740 1006602
rect 153750 1006632 153806 1006641
rect 103150 1006567 103152 1006576
rect 94688 1006538 94740 1006544
rect 103204 1006567 103206 1006576
rect 145564 1006596 145616 1006602
rect 103152 1006538 103204 1006544
rect 306930 1006632 306986 1006641
rect 153750 1006567 153752 1006576
rect 145564 1006538 145616 1006544
rect 153804 1006567 153806 1006576
rect 298836 1006596 298888 1006602
rect 153752 1006538 153804 1006544
rect 306930 1006567 306932 1006576
rect 298836 1006538 298888 1006544
rect 306984 1006567 306986 1006576
rect 306932 1006538 306984 1006544
rect 93124 1006324 93176 1006330
rect 93124 1006266 93176 1006272
rect 92664 999796 92716 999802
rect 92664 999738 92716 999744
rect 92296 998028 92348 998034
rect 92296 997970 92348 997976
rect 85946 995752 86002 995761
rect 85698 995710 85946 995738
rect 85946 995687 86002 995696
rect 84658 995480 84714 995489
rect 77036 995042 77064 995452
rect 77680 995178 77708 995452
rect 77668 995172 77720 995178
rect 77668 995114 77720 995120
rect 77024 995036 77076 995042
rect 77024 994978 77076 994984
rect 78324 994906 78352 995452
rect 78312 994900 78364 994906
rect 78312 994842 78364 994848
rect 80164 994770 80192 995452
rect 80152 994764 80204 994770
rect 80152 994706 80204 994712
rect 80716 994537 80744 995452
rect 81360 994634 81388 995452
rect 81348 994628 81400 994634
rect 81348 994570 81400 994576
rect 80702 994528 80758 994537
rect 82004 994498 82032 995452
rect 84502 995438 84658 995466
rect 86590 995480 86646 995489
rect 84658 995415 84714 995424
rect 85040 995217 85068 995452
rect 86342 995438 86590 995466
rect 90178 995480 90234 995489
rect 86590 995415 86646 995424
rect 85026 995208 85082 995217
rect 85026 995143 85082 995152
rect 80702 994463 80758 994472
rect 81992 994492 82044 994498
rect 81992 994434 82044 994440
rect 87524 994129 87552 995452
rect 88734 995438 89024 995466
rect 88996 995382 89024 995438
rect 88984 995376 89036 995382
rect 88984 995318 89036 995324
rect 89364 994809 89392 995452
rect 90022 995438 90178 995466
rect 91218 995438 91692 995466
rect 90178 995415 90234 995424
rect 91664 995330 91692 995438
rect 92308 995330 92336 997970
rect 92480 996396 92532 996402
rect 92480 996338 92532 996344
rect 92492 995382 92520 996338
rect 91664 995302 92336 995330
rect 92480 995376 92532 995382
rect 92480 995318 92532 995324
rect 89350 994800 89406 994809
rect 89350 994735 89406 994744
rect 92676 994129 92704 999738
rect 93136 994498 93164 1006266
rect 94504 1006188 94556 1006194
rect 94504 1006130 94556 1006136
rect 93308 1006052 93360 1006058
rect 93308 1005994 93360 1006000
rect 93320 996441 93348 1005994
rect 93306 996432 93362 996441
rect 93306 996367 93362 996376
rect 93490 995752 93546 995761
rect 93490 995687 93546 995696
rect 93504 995081 93532 995687
rect 93490 995072 93546 995081
rect 93490 995007 93546 995016
rect 93124 994492 93176 994498
rect 93124 994434 93176 994440
rect 94516 994401 94544 1006130
rect 94700 998034 94728 1006538
rect 103978 1006496 104034 1006505
rect 102784 1006460 102836 1006466
rect 103978 1006431 103980 1006440
rect 102784 1006402 102836 1006408
rect 104032 1006431 104034 1006440
rect 103980 1006402 104032 1006408
rect 100298 1006360 100354 1006369
rect 100298 1006295 100300 1006304
rect 100352 1006295 100354 1006304
rect 100300 1006266 100352 1006272
rect 101954 1006224 102010 1006233
rect 101954 1006159 101956 1006168
rect 102008 1006159 102010 1006168
rect 101956 1006130 102008 1006136
rect 98274 1006088 98330 1006097
rect 98274 1006023 98276 1006032
rect 98328 1006023 98330 1006032
rect 101404 1006052 101456 1006058
rect 98276 1005994 98328 1006000
rect 101404 1005994 101456 1006000
rect 98644 1002788 98696 1002794
rect 98644 1002730 98696 1002736
rect 97264 1002652 97316 1002658
rect 97264 1002594 97316 1002600
rect 96528 1002380 96580 1002386
rect 96528 1002322 96580 1002328
rect 96344 1001972 96396 1001978
rect 96344 1001914 96396 1001920
rect 94688 998028 94740 998034
rect 94688 997970 94740 997976
rect 94502 994392 94558 994401
rect 94502 994327 94558 994336
rect 87510 994120 87566 994129
rect 87510 994055 87566 994064
rect 92662 994120 92718 994129
rect 92662 994055 92718 994064
rect 51724 993064 51776 993070
rect 51724 993006 51776 993012
rect 46204 992928 46256 992934
rect 46204 992870 46256 992876
rect 42524 969468 42576 969474
rect 42524 969410 42576 969416
rect 41800 968833 41828 969272
rect 41786 968824 41842 968833
rect 41786 968759 41842 968768
rect 42182 968034 42288 968062
rect 41984 967201 42012 967405
rect 41970 967192 42026 967201
rect 41970 967127 42026 967136
rect 42260 966890 42288 968034
rect 42248 966884 42300 966890
rect 42248 966826 42300 966832
rect 42536 966770 42564 969410
rect 42708 966884 42760 966890
rect 42708 966826 42760 966832
rect 42182 966742 42564 966770
rect 42182 965551 42472 965579
rect 42444 964714 42472 965551
rect 42432 964708 42484 964714
rect 42432 964650 42484 964656
rect 42182 964362 42472 964390
rect 42444 963898 42472 964362
rect 42432 963892 42484 963898
rect 42432 963834 42484 963840
rect 42182 963711 42472 963739
rect 42444 963490 42472 963711
rect 42432 963484 42484 963490
rect 42432 963426 42484 963432
rect 42182 963070 42472 963098
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 42444 961926 42472 963070
rect 42432 961920 42484 961926
rect 42432 961862 42484 961868
rect 42168 960078 42288 960106
rect 42168 960024 42196 960078
rect 42260 960038 42288 960078
rect 42260 960010 42472 960038
rect 41800 959177 41828 959412
rect 41786 959168 41842 959177
rect 42444 959138 42472 960010
rect 41786 959103 41842 959112
rect 42432 959132 42484 959138
rect 42432 959074 42484 959080
rect 42168 958854 42288 958882
rect 42168 958732 42196 958854
rect 42260 958746 42288 958854
rect 42260 958718 42472 958746
rect 42168 958310 42288 958338
rect 42444 958322 42472 958718
rect 42168 958188 42196 958310
rect 42260 958202 42288 958310
rect 42432 958316 42484 958322
rect 42432 958258 42484 958264
rect 42260 958174 42380 958202
rect 41786 956584 41842 956593
rect 41786 956519 41842 956528
rect 41800 956352 41828 956519
rect 41800 955505 41828 955740
rect 41786 955496 41842 955505
rect 41786 955431 41842 955440
rect 42168 955182 42288 955210
rect 42168 955060 42196 955182
rect 42260 954122 42288 955182
rect 41708 954094 42288 954122
rect 39302 952504 39358 952513
rect 39302 952439 39358 952448
rect 37922 952232 37978 952241
rect 37922 952167 37978 952176
rect 35164 951516 35216 951522
rect 35164 951458 35216 951464
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 35176 938471 35204 951458
rect 35162 938462 35218 938471
rect 35162 938397 35218 938406
rect 37936 937009 37964 952167
rect 39316 937417 39344 952439
rect 40038 951688 40094 951697
rect 40038 951623 40094 951632
rect 41510 951688 41566 951697
rect 41510 951623 41566 951632
rect 39302 937408 39358 937417
rect 39302 937343 39358 937352
rect 37922 937000 37978 937009
rect 37922 936935 37978 936944
rect 40052 935785 40080 951623
rect 41326 941896 41382 941905
rect 41326 941831 41382 941840
rect 41340 941526 41368 941831
rect 41328 941520 41380 941526
rect 41328 941462 41380 941468
rect 40958 941080 41014 941089
rect 40958 941015 41014 941024
rect 40972 940166 41000 941015
rect 40960 940160 41012 940166
rect 40960 940102 41012 940108
rect 41142 939448 41198 939457
rect 41142 939383 41198 939392
rect 40960 938596 41012 938602
rect 40960 938538 41012 938544
rect 40972 938471 41000 938538
rect 40958 938462 41014 938471
rect 41156 938466 41184 939383
rect 41524 938602 41552 951623
rect 41708 951522 41736 954094
rect 42352 953594 42380 958174
rect 42720 953594 42748 966826
rect 42892 964708 42944 964714
rect 42892 964650 42944 964656
rect 42904 953594 42932 964650
rect 44180 963892 44232 963898
rect 44180 963834 44232 963840
rect 43076 963484 43128 963490
rect 43076 963426 43128 963432
rect 42260 953566 42380 953594
rect 42536 953566 42748 953594
rect 42812 953566 42932 953594
rect 41696 951516 41748 951522
rect 41696 951458 41748 951464
rect 41696 941520 41748 941526
rect 41748 941468 41920 941474
rect 41696 941462 41920 941468
rect 41708 941446 41920 941462
rect 41696 940160 41748 940166
rect 41696 940102 41748 940108
rect 41512 938596 41564 938602
rect 41512 938538 41564 938544
rect 40958 938397 41014 938406
rect 41144 938460 41196 938466
rect 41144 938402 41196 938408
rect 41512 938460 41564 938466
rect 41512 938402 41564 938408
rect 40038 935776 40094 935785
rect 40038 935711 40094 935720
rect 40682 881920 40738 881929
rect 40682 881855 40738 881864
rect 39946 819088 40002 819097
rect 39946 819023 40002 819032
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35622 818000 35678 818009
rect 35622 817935 35678 817944
rect 35636 817018 35664 817935
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817154 35848 817255
rect 35808 817148 35860 817154
rect 35808 817090 35860 817096
rect 39960 817018 39988 819023
rect 40314 818000 40370 818009
rect 40314 817935 40370 817944
rect 35624 817012 35676 817018
rect 35624 816954 35676 816960
rect 39948 817012 40000 817018
rect 39948 816954 40000 816960
rect 35254 816912 35310 816921
rect 35254 816847 35310 816856
rect 35268 815658 35296 816847
rect 35438 816504 35494 816513
rect 35438 816439 35494 816448
rect 35452 815930 35480 816439
rect 35806 816096 35862 816105
rect 35624 816060 35676 816066
rect 35806 816031 35862 816040
rect 35624 816002 35676 816008
rect 35440 815924 35492 815930
rect 35440 815866 35492 815872
rect 35636 815697 35664 816002
rect 35820 815794 35848 816031
rect 35808 815788 35860 815794
rect 35808 815730 35860 815736
rect 35622 815688 35678 815697
rect 35256 815652 35308 815658
rect 35622 815623 35678 815632
rect 35256 815594 35308 815600
rect 35438 815280 35494 815289
rect 35438 815215 35494 815224
rect 35452 814298 35480 815215
rect 35622 814872 35678 814881
rect 35622 814807 35678 814816
rect 35636 814434 35664 814807
rect 35808 814700 35860 814706
rect 35808 814642 35860 814648
rect 35820 814473 35848 814642
rect 35806 814464 35862 814473
rect 35624 814428 35676 814434
rect 40328 814434 40356 817935
rect 40696 817154 40724 881855
rect 40684 817148 40736 817154
rect 40684 817090 40736 817096
rect 41328 815788 41380 815794
rect 41328 815730 41380 815736
rect 35806 814399 35862 814408
rect 40316 814428 40368 814434
rect 35624 814370 35676 814376
rect 40316 814370 40368 814376
rect 35440 814292 35492 814298
rect 35440 814234 35492 814240
rect 41142 814056 41198 814065
rect 41142 813991 41198 814000
rect 41156 813006 41184 813991
rect 41144 813000 41196 813006
rect 41144 812942 41196 812948
rect 41142 812832 41198 812841
rect 41340 812818 41368 815730
rect 41524 813006 41552 938402
rect 41708 816066 41736 940102
rect 41696 816060 41748 816066
rect 41696 816002 41748 816008
rect 41892 815946 41920 941446
rect 42062 940264 42118 940273
rect 42062 940199 42118 940208
rect 42076 823874 42104 940199
rect 42260 937825 42288 953566
rect 42246 937816 42302 937825
rect 42246 937751 42302 937760
rect 42536 932929 42564 953566
rect 42812 935377 42840 953566
rect 42798 935368 42854 935377
rect 42798 935303 42854 935312
rect 43088 934969 43116 963426
rect 43260 959132 43312 959138
rect 43260 959074 43312 959080
rect 43074 934960 43130 934969
rect 43074 934895 43130 934904
rect 43272 934561 43300 959074
rect 43536 946008 43588 946014
rect 43536 945950 43588 945956
rect 43548 943537 43576 945950
rect 43534 943528 43590 943537
rect 43534 943463 43590 943472
rect 43442 942304 43498 942313
rect 43442 942239 43498 942248
rect 43456 941254 43484 942239
rect 43628 941384 43680 941390
rect 43626 941352 43628 941361
rect 43680 941352 43682 941361
rect 43626 941287 43682 941296
rect 43444 941248 43496 941254
rect 43444 941190 43496 941196
rect 43442 939856 43498 939865
rect 43442 939791 43444 939800
rect 43496 939791 43498 939800
rect 43444 939762 43496 939768
rect 43258 934552 43314 934561
rect 43258 934487 43314 934496
rect 44192 933745 44220 963834
rect 44456 961920 44508 961926
rect 44456 961862 44508 961868
rect 44468 934153 44496 961862
rect 44640 958316 44692 958322
rect 44640 958258 44692 958264
rect 44652 949454 44680 958258
rect 44652 949426 44864 949454
rect 44638 943120 44694 943129
rect 44638 943055 44694 943064
rect 44652 937038 44680 943055
rect 44640 937032 44692 937038
rect 44640 936974 44692 936980
rect 44836 936193 44864 949426
rect 46216 940681 46244 992870
rect 50344 991500 50396 991506
rect 50344 991442 50396 991448
rect 48964 990140 49016 990146
rect 48964 990082 49016 990088
rect 47584 961920 47636 961926
rect 47584 961862 47636 961868
rect 47596 942721 47624 961862
rect 47582 942712 47638 942721
rect 47582 942647 47638 942656
rect 48976 941390 49004 990082
rect 48964 941384 49016 941390
rect 48964 941326 49016 941332
rect 50356 941254 50384 991442
rect 50344 941248 50396 941254
rect 50344 941190 50396 941196
rect 46202 940672 46258 940681
rect 46202 940607 46258 940616
rect 51736 939826 51764 993006
rect 73436 991636 73488 991642
rect 73436 991578 73488 991584
rect 73448 983620 73476 991578
rect 96356 987426 96384 1001914
rect 96344 987420 96396 987426
rect 96344 987362 96396 987368
rect 89628 985992 89680 985998
rect 89628 985934 89680 985940
rect 89640 983620 89668 985934
rect 96540 984638 96568 1002322
rect 97080 997280 97132 997286
rect 97078 997248 97080 997257
rect 97132 997248 97134 997257
rect 97078 997183 97134 997192
rect 97276 995353 97304 1002594
rect 97448 1002108 97500 1002114
rect 97448 1002050 97500 1002056
rect 97460 995625 97488 1002050
rect 98274 1002008 98330 1002017
rect 98274 1001943 98276 1001952
rect 98328 1001943 98330 1001952
rect 98276 1001914 98328 1001920
rect 97446 995616 97502 995625
rect 97446 995551 97502 995560
rect 97262 995344 97318 995353
rect 97262 995279 97318 995288
rect 98656 994634 98684 1002730
rect 100298 1002688 100354 1002697
rect 100298 1002623 100300 1002632
rect 100352 1002623 100354 1002632
rect 100300 1002594 100352 1002600
rect 101126 1002552 101182 1002561
rect 98828 1002516 98880 1002522
rect 101126 1002487 101128 1002496
rect 98828 1002458 98880 1002464
rect 101180 1002487 101182 1002496
rect 101128 1002458 101180 1002464
rect 98840 997286 98868 1002458
rect 99102 1002416 99158 1002425
rect 99102 1002351 99104 1002360
rect 99156 1002351 99158 1002360
rect 99104 1002322 99156 1002328
rect 101126 1002280 101182 1002289
rect 99012 1002244 99064 1002250
rect 101126 1002215 101128 1002224
rect 99012 1002186 99064 1002192
rect 101180 1002215 101182 1002224
rect 101128 1002186 101180 1002192
rect 99024 999802 99052 1002186
rect 99470 1002144 99526 1002153
rect 99470 1002079 99472 1002088
rect 99524 1002079 99526 1002088
rect 100024 1002108 100076 1002114
rect 99472 1002050 99524 1002056
rect 100024 1002050 100076 1002056
rect 99012 999796 99064 999802
rect 99012 999738 99064 999744
rect 98828 997280 98880 997286
rect 98828 997222 98880 997228
rect 100036 995081 100064 1002050
rect 100208 1001972 100260 1001978
rect 100208 1001914 100260 1001920
rect 100220 995178 100248 1001914
rect 100208 995172 100260 995178
rect 100208 995114 100260 995120
rect 100022 995072 100078 995081
rect 100022 995007 100078 995016
rect 101416 994770 101444 1005994
rect 101954 1002824 102010 1002833
rect 101954 1002759 101956 1002768
rect 102008 1002759 102010 1002768
rect 101956 1002730 102008 1002736
rect 102322 1002008 102378 1002017
rect 102322 1001943 102324 1001952
rect 102376 1001943 102378 1001952
rect 102324 1001914 102376 1001920
rect 102796 995042 102824 1006402
rect 144276 1006324 144328 1006330
rect 144276 1006266 144328 1006272
rect 106830 1006224 106886 1006233
rect 106830 1006159 106832 1006168
rect 106884 1006159 106886 1006168
rect 124864 1006188 124916 1006194
rect 106832 1006130 106884 1006136
rect 124864 1006130 124916 1006136
rect 103978 1006088 104034 1006097
rect 103978 1006023 103980 1006032
rect 104032 1006023 104034 1006032
rect 107658 1006088 107714 1006097
rect 107658 1006023 107660 1006032
rect 103980 1005994 104032 1006000
rect 107712 1006023 107714 1006032
rect 107660 1005994 107712 1006000
rect 108486 1004728 108542 1004737
rect 106188 1004692 106240 1004698
rect 108486 1004663 108488 1004672
rect 106188 1004634 106240 1004640
rect 108540 1004663 108542 1004672
rect 108488 1004634 108540 1004640
rect 106002 1002552 106058 1002561
rect 106002 1002487 106004 1002496
rect 106056 1002487 106058 1002496
rect 106004 1002458 106056 1002464
rect 105634 1002416 105690 1002425
rect 105634 1002351 105636 1002360
rect 105688 1002351 105690 1002360
rect 105636 1002322 105688 1002328
rect 104806 1002280 104862 1002289
rect 104806 1002215 104808 1002224
rect 104860 1002215 104862 1002224
rect 104808 1002186 104860 1002192
rect 103150 1002144 103206 1002153
rect 103150 1002079 103152 1002088
rect 103204 1002079 103206 1002088
rect 103152 1002050 103204 1002056
rect 104806 1002008 104862 1002017
rect 104176 1001966 104806 1001994
rect 102784 995036 102836 995042
rect 102784 994978 102836 994984
rect 104176 994906 104204 1001966
rect 104806 1001943 104862 1001952
rect 106002 1002008 106058 1002017
rect 106002 1001943 106004 1001952
rect 106056 1001943 106058 1001952
rect 106004 1001914 106056 1001920
rect 104164 994900 104216 994906
rect 104164 994842 104216 994848
rect 101404 994764 101456 994770
rect 101404 994706 101456 994712
rect 98644 994628 98696 994634
rect 98644 994570 98696 994576
rect 96528 984632 96580 984638
rect 96528 984574 96580 984580
rect 106200 983634 106228 1004634
rect 109500 1002516 109552 1002522
rect 109500 1002458 109552 1002464
rect 108026 1002416 108082 1002425
rect 107752 1002380 107804 1002386
rect 108026 1002351 108028 1002360
rect 107752 1002322 107804 1002328
rect 108080 1002351 108082 1002360
rect 108028 1002322 108080 1002328
rect 106464 1002244 106516 1002250
rect 106464 1002186 106516 1002192
rect 106476 994809 106504 1002186
rect 106830 1002144 106886 1002153
rect 106830 1002079 106832 1002088
rect 106884 1002079 106886 1002088
rect 106832 1002050 106884 1002056
rect 106924 996940 106976 996946
rect 106924 996882 106976 996888
rect 106462 994800 106518 994809
rect 106462 994735 106518 994744
rect 106936 985998 106964 996882
rect 107764 993070 107792 1002322
rect 108486 1002280 108542 1002289
rect 108486 1002215 108488 1002224
rect 108540 1002215 108542 1002224
rect 108488 1002186 108540 1002192
rect 109040 1002108 109092 1002114
rect 109040 1002050 109092 1002056
rect 108854 1002008 108910 1002017
rect 108120 1001972 108172 1001978
rect 108854 1001943 108856 1001952
rect 108120 1001914 108172 1001920
rect 108908 1001943 108910 1001952
rect 108856 1001914 108908 1001920
rect 107752 993064 107804 993070
rect 107752 993006 107804 993012
rect 108132 992934 108160 1001914
rect 108120 992928 108172 992934
rect 108120 992870 108172 992876
rect 109052 990146 109080 1002050
rect 109512 996130 109540 1002458
rect 110420 1002380 110472 1002386
rect 110420 1002322 110472 1002328
rect 109682 1002144 109738 1002153
rect 109682 1002079 109684 1002088
rect 109736 1002079 109738 1002088
rect 109684 1002050 109736 1002056
rect 109500 996124 109552 996130
rect 109500 996066 109552 996072
rect 110432 991506 110460 1002322
rect 111064 1002244 111116 1002250
rect 111064 1002186 111116 1002192
rect 111076 995994 111104 1002186
rect 111892 1002108 111944 1002114
rect 111892 1002050 111944 1002056
rect 111904 996946 111932 1002050
rect 112076 1001972 112128 1001978
rect 112076 1001914 112128 1001920
rect 111892 996940 111944 996946
rect 111892 996882 111944 996888
rect 111064 995988 111116 995994
rect 111064 995930 111116 995936
rect 112088 991642 112116 1001914
rect 121736 996396 121788 996402
rect 121736 996338 121788 996344
rect 112076 991636 112128 991642
rect 112076 991578 112128 991584
rect 110420 991500 110472 991506
rect 110420 991442 110472 991448
rect 109040 990140 109092 990146
rect 109040 990082 109092 990088
rect 106924 985992 106976 985998
rect 106924 985934 106976 985940
rect 105846 983606 106228 983634
rect 121748 983634 121776 996338
rect 124876 995858 124904 1006130
rect 126244 1006052 126296 1006058
rect 126244 1005994 126296 1006000
rect 124864 995852 124916 995858
rect 124864 995794 124916 995800
rect 126256 995450 126284 1005994
rect 143724 998096 143776 998102
rect 143724 998038 143776 998044
rect 143736 995761 143764 998038
rect 143908 997892 143960 997898
rect 143908 997834 143960 997840
rect 133050 995752 133106 995761
rect 137374 995752 137430 995761
rect 133106 995710 133446 995738
rect 137126 995710 137374 995738
rect 133050 995687 133106 995696
rect 139122 995752 139178 995761
rect 138966 995710 139122 995738
rect 137374 995687 137430 995696
rect 140962 995752 141018 995761
rect 140806 995710 140962 995738
rect 139122 995687 139178 995696
rect 141790 995752 141846 995761
rect 141450 995710 141790 995738
rect 140962 995687 141018 995696
rect 141790 995687 141846 995696
rect 143722 995752 143778 995761
rect 143722 995687 143778 995696
rect 143920 995602 143948 997834
rect 144288 996985 144316 1006266
rect 144460 1006188 144512 1006194
rect 144460 1006130 144512 1006136
rect 144274 996976 144330 996985
rect 144274 996911 144330 996920
rect 144472 995994 144500 1006130
rect 144736 1002380 144788 1002386
rect 144736 1002322 144788 1002328
rect 144748 1001894 144776 1002322
rect 144656 1001866 144776 1001894
rect 144460 995988 144512 995994
rect 144460 995930 144512 995936
rect 143460 995574 143948 995602
rect 136638 995480 136694 995489
rect 126244 995444 126296 995450
rect 126244 995386 126296 995392
rect 128464 994974 128492 995452
rect 128452 994968 128504 994974
rect 128452 994910 128504 994916
rect 129108 994809 129136 995452
rect 129094 994800 129150 994809
rect 129094 994735 129150 994744
rect 129752 994537 129780 995452
rect 131592 994566 131620 995452
rect 132144 994838 132172 995452
rect 132802 995438 133184 995466
rect 132406 995344 132462 995353
rect 132406 995279 132462 995288
rect 132132 994832 132184 994838
rect 132132 994774 132184 994780
rect 132420 994702 132448 995279
rect 132408 994696 132460 994702
rect 132408 994638 132460 994644
rect 131580 994560 131632 994566
rect 129738 994528 129794 994537
rect 131580 994502 131632 994508
rect 129738 994463 129794 994472
rect 133156 993993 133184 995438
rect 135916 995081 135944 995452
rect 136482 995438 136638 995466
rect 137770 995438 137968 995466
rect 136638 995415 136694 995424
rect 137940 995178 137968 995438
rect 137928 995172 137980 995178
rect 137928 995114 137980 995120
rect 135902 995072 135958 995081
rect 135902 995007 135958 995016
rect 140148 994294 140176 995452
rect 142646 995438 143028 995466
rect 143000 995330 143028 995438
rect 143460 995330 143488 995574
rect 142804 995308 142856 995314
rect 143000 995302 143488 995330
rect 142804 995250 142856 995256
rect 140136 994288 140188 994294
rect 140136 994230 140188 994236
rect 142816 993993 142844 995250
rect 144656 995178 144684 1001866
rect 144828 997756 144880 997762
rect 144828 997698 144880 997704
rect 144840 996441 144868 997698
rect 144826 996432 144882 996441
rect 144826 996367 144882 996376
rect 144644 995172 144696 995178
rect 144644 995114 144696 995120
rect 145576 994838 145604 1006538
rect 152922 1006496 152978 1006505
rect 145748 1006460 145800 1006466
rect 152922 1006431 152924 1006440
rect 145748 1006402 145800 1006408
rect 152976 1006431 152978 1006440
rect 152924 1006402 152976 1006408
rect 145760 996713 145788 1006402
rect 210424 1006392 210476 1006398
rect 152094 1006360 152150 1006369
rect 152094 1006295 152096 1006304
rect 152148 1006295 152150 1006304
rect 158258 1006360 158314 1006369
rect 210422 1006360 210424 1006369
rect 228364 1006392 228416 1006398
rect 210476 1006360 210478 1006369
rect 158258 1006295 158260 1006304
rect 152096 1006266 152148 1006272
rect 158312 1006295 158314 1006304
rect 175924 1006324 175976 1006330
rect 158260 1006266 158312 1006272
rect 228364 1006334 228416 1006340
rect 256146 1006360 256202 1006369
rect 210422 1006295 210478 1006304
rect 175924 1006266 175976 1006272
rect 159454 1006224 159510 1006233
rect 159454 1006159 159456 1006168
rect 159508 1006159 159510 1006168
rect 160282 1006224 160338 1006233
rect 160282 1006159 160284 1006168
rect 159456 1006130 159508 1006136
rect 160336 1006159 160338 1006168
rect 164884 1006188 164936 1006194
rect 160284 1006130 160336 1006136
rect 164884 1006130 164936 1006136
rect 146942 1006088 146998 1006097
rect 146942 1006023 146998 1006032
rect 148874 1006088 148930 1006097
rect 148874 1006023 148876 1006032
rect 146956 998102 146984 1006023
rect 148928 1006023 148930 1006032
rect 150070 1006088 150126 1006097
rect 155774 1006088 155830 1006097
rect 150070 1006023 150072 1006032
rect 148876 1005994 148928 1006000
rect 150124 1006023 150126 1006032
rect 152648 1006052 152700 1006058
rect 150072 1005994 150124 1006000
rect 155774 1006023 155776 1006032
rect 152648 1005994 152700 1006000
rect 155828 1006023 155830 1006032
rect 158626 1006088 158682 1006097
rect 158626 1006023 158628 1006032
rect 155776 1005994 155828 1006000
rect 158680 1006023 158682 1006032
rect 158628 1005994 158680 1006000
rect 149888 1005372 149940 1005378
rect 149888 1005314 149940 1005320
rect 149704 1004692 149756 1004698
rect 149704 1004634 149756 1004640
rect 148324 1002244 148376 1002250
rect 148324 1002186 148376 1002192
rect 147588 1001972 147640 1001978
rect 147588 1001914 147640 1001920
rect 146944 998096 146996 998102
rect 146944 998038 146996 998044
rect 145746 996704 145802 996713
rect 145746 996639 145802 996648
rect 145564 994832 145616 994838
rect 145564 994774 145616 994780
rect 133142 993984 133198 993993
rect 133142 993919 133198 993928
rect 142802 993984 142858 993993
rect 142802 993919 142858 993928
rect 147600 993070 147628 1001914
rect 148336 995489 148364 1002186
rect 148968 1002108 149020 1002114
rect 148968 1002050 149020 1002056
rect 148322 995480 148378 995489
rect 148322 995415 148378 995424
rect 147588 993064 147640 993070
rect 147588 993006 147640 993012
rect 148980 992934 149008 1002050
rect 149242 1002008 149298 1002017
rect 149242 1001943 149244 1001952
rect 149296 1001943 149298 1001952
rect 149244 1001914 149296 1001920
rect 149716 994702 149744 1004634
rect 149900 995314 149928 1005314
rect 151084 1004964 151136 1004970
rect 151084 1004906 151136 1004912
rect 150898 1002416 150954 1002425
rect 150898 1002351 150900 1002360
rect 150952 1002351 150954 1002360
rect 150900 1002322 150952 1002328
rect 150898 1002144 150954 1002153
rect 150898 1002079 150900 1002088
rect 150952 1002079 150954 1002088
rect 150900 1002050 150952 1002056
rect 149888 995308 149940 995314
rect 149888 995250 149940 995256
rect 151096 994809 151124 1004906
rect 151268 1004828 151320 1004834
rect 151268 1004770 151320 1004776
rect 151280 997898 151308 1004770
rect 151726 1004728 151782 1004737
rect 151726 1004663 151728 1004672
rect 151780 1004663 151782 1004672
rect 151728 1004634 151780 1004640
rect 151726 1002280 151782 1002289
rect 151726 1002215 151728 1002224
rect 151780 1002215 151782 1002224
rect 151728 1002186 151780 1002192
rect 152464 1002040 152516 1002046
rect 152464 1001982 152516 1001988
rect 151268 997892 151320 997898
rect 151268 997834 151320 997840
rect 152476 995081 152504 1001982
rect 152660 997762 152688 1005994
rect 152922 1005408 152978 1005417
rect 152922 1005343 152924 1005352
rect 152976 1005343 152978 1005352
rect 152924 1005314 152976 1005320
rect 153750 1005000 153806 1005009
rect 160650 1005000 160706 1005009
rect 153750 1004935 153752 1004944
rect 153804 1004935 153806 1004944
rect 154396 1004964 154448 1004970
rect 153752 1004906 153804 1004912
rect 160650 1004935 160652 1004944
rect 154396 1004906 154448 1004912
rect 160704 1004935 160706 1004944
rect 160652 1004906 160704 1004912
rect 154118 1004864 154174 1004873
rect 154118 1004799 154120 1004808
rect 154172 1004799 154174 1004808
rect 154120 1004770 154172 1004776
rect 154408 1001894 154436 1004906
rect 159454 1004864 159510 1004873
rect 159454 1004799 159456 1004808
rect 159508 1004799 159510 1004808
rect 162124 1004828 162176 1004834
rect 159456 1004770 159508 1004776
rect 162124 1004770 162176 1004776
rect 160650 1004728 160706 1004737
rect 160650 1004663 160652 1004672
rect 160704 1004663 160706 1004672
rect 160652 1004634 160704 1004640
rect 157430 1002688 157486 1002697
rect 157430 1002623 157432 1002632
rect 157484 1002623 157486 1002632
rect 159364 1002652 159416 1002658
rect 157432 1002594 157484 1002600
rect 159364 1002594 159416 1002600
rect 158626 1002552 158682 1002561
rect 158626 1002487 158628 1002496
rect 158680 1002487 158682 1002496
rect 158628 1002458 158680 1002464
rect 156602 1002416 156658 1002425
rect 156602 1002351 156604 1002360
rect 156656 1002351 156658 1002360
rect 158720 1002380 158772 1002386
rect 156604 1002322 156656 1002328
rect 158720 1002322 158772 1002328
rect 155774 1002280 155830 1002289
rect 155774 1002215 155776 1002224
rect 155828 1002215 155830 1002224
rect 157340 1002244 157392 1002250
rect 155776 1002186 155828 1002192
rect 157340 1002186 157392 1002192
rect 156602 1002144 156658 1002153
rect 155224 1002108 155276 1002114
rect 156602 1002079 156604 1002088
rect 155224 1002050 155276 1002056
rect 156656 1002079 156658 1002088
rect 156604 1002050 156656 1002056
rect 154580 1002040 154632 1002046
rect 154578 1002008 154580 1002017
rect 154632 1002008 154634 1002017
rect 154578 1001943 154634 1001952
rect 154946 1002008 155002 1002017
rect 154946 1001943 154948 1001952
rect 155000 1001943 155002 1001952
rect 154948 1001914 155000 1001920
rect 154408 1001866 154528 1001894
rect 152648 997756 152700 997762
rect 152648 997698 152700 997704
rect 152462 995072 152518 995081
rect 152462 995007 152518 995016
rect 151082 994800 151138 994809
rect 151082 994735 151138 994744
rect 149704 994696 149756 994702
rect 149704 994638 149756 994644
rect 148968 992928 149020 992934
rect 148968 992870 149020 992876
rect 138296 991500 138348 991506
rect 138296 991442 138348 991448
rect 121748 983606 122130 983634
rect 138308 983620 138336 991442
rect 154500 983620 154528 1001866
rect 155236 994537 155264 1002050
rect 155960 1001972 156012 1001978
rect 155960 1001914 156012 1001920
rect 155972 994838 156000 1001914
rect 157352 994974 157380 1002186
rect 157798 1002008 157854 1002017
rect 157798 1001943 157800 1001952
rect 157852 1001943 157854 1001952
rect 157800 1001914 157852 1001920
rect 158732 996130 158760 1002322
rect 159376 996130 159404 1002594
rect 160192 1002516 160244 1002522
rect 160192 1002458 160244 1002464
rect 158720 996124 158772 996130
rect 158720 996066 158772 996072
rect 159364 996124 159416 996130
rect 159364 996066 159416 996072
rect 160204 995450 160232 1002458
rect 160376 1001972 160428 1001978
rect 160376 1001914 160428 1001920
rect 160388 995858 160416 1001914
rect 162136 995994 162164 1004770
rect 162860 1004692 162912 1004698
rect 162860 1004634 162912 1004640
rect 162124 995988 162176 995994
rect 162124 995930 162176 995936
rect 160376 995852 160428 995858
rect 160376 995794 160428 995800
rect 160192 995444 160244 995450
rect 160192 995386 160244 995392
rect 157340 994968 157392 994974
rect 157340 994910 157392 994916
rect 155960 994832 156012 994838
rect 155960 994774 156012 994780
rect 155222 994528 155278 994537
rect 155222 994463 155278 994472
rect 162872 991506 162900 1004634
rect 164896 997694 164924 1006130
rect 164884 997688 164936 997694
rect 164884 997630 164936 997636
rect 170312 997688 170364 997694
rect 170312 997630 170364 997636
rect 162860 991500 162912 991506
rect 162860 991442 162912 991448
rect 170324 983634 170352 997630
rect 175936 995858 175964 1006266
rect 208400 1006256 208452 1006262
rect 208398 1006224 208400 1006233
rect 208452 1006224 208454 1006233
rect 208398 1006159 208454 1006168
rect 201038 1006088 201094 1006097
rect 177304 1006052 177356 1006058
rect 177304 1005994 177356 1006000
rect 198648 1006052 198700 1006058
rect 201038 1006023 201040 1006032
rect 198648 1005994 198700 1006000
rect 201092 1006023 201094 1006032
rect 201040 1005994 201092 1006000
rect 175924 995852 175976 995858
rect 175924 995794 175976 995800
rect 177316 995518 177344 1005994
rect 195704 1005304 195756 1005310
rect 195704 1005246 195756 1005252
rect 195152 1001972 195204 1001978
rect 195152 1001914 195204 1001920
rect 195164 997754 195192 1001914
rect 195520 999796 195572 999802
rect 195520 999738 195572 999744
rect 195072 997726 195192 997754
rect 195072 995761 195100 997726
rect 195242 996704 195298 996713
rect 195242 996639 195298 996648
rect 188066 995752 188122 995761
rect 187864 995710 188066 995738
rect 189354 995752 189410 995761
rect 189152 995710 189354 995738
rect 188066 995687 188122 995696
rect 192482 995752 192538 995761
rect 192188 995710 192482 995738
rect 189354 995687 189410 995696
rect 193126 995752 193182 995761
rect 192832 995710 193126 995738
rect 192482 995687 192538 995696
rect 193126 995687 193182 995696
rect 195058 995752 195114 995761
rect 195058 995687 195114 995696
rect 195060 995580 195112 995586
rect 195060 995522 195112 995528
rect 177304 995512 177356 995518
rect 183834 995480 183890 995489
rect 177304 995454 177356 995460
rect 179860 995438 180380 995466
rect 180504 995438 180656 995466
rect 180352 994650 180380 995438
rect 180628 994838 180656 995438
rect 180812 995438 181148 995466
rect 182988 995438 183324 995466
rect 183540 995438 183834 995466
rect 180812 995246 180840 995438
rect 180800 995240 180852 995246
rect 180800 995182 180852 995188
rect 183296 994974 183324 995438
rect 184184 995438 184520 995466
rect 184828 995438 184888 995466
rect 187312 995438 187648 995466
rect 188508 995438 188844 995466
rect 190348 995438 190408 995466
rect 191544 995438 191880 995466
rect 194028 995438 194364 995466
rect 183834 995415 183890 995424
rect 183284 994968 183336 994974
rect 183284 994910 183336 994916
rect 180616 994832 180668 994838
rect 180616 994774 180668 994780
rect 180616 994696 180668 994702
rect 180352 994644 180616 994650
rect 180352 994638 180668 994644
rect 180352 994622 180656 994638
rect 184492 994158 184520 995438
rect 184860 994401 184888 995438
rect 187620 994945 187648 995438
rect 187606 994936 187662 994945
rect 187606 994871 187662 994880
rect 188816 994673 188844 995438
rect 188802 994664 188858 994673
rect 188802 994599 188858 994608
rect 184846 994392 184902 994401
rect 184846 994327 184902 994336
rect 186504 994288 186556 994294
rect 186504 994230 186556 994236
rect 184480 994152 184532 994158
rect 184480 994094 184532 994100
rect 186516 983634 186544 994230
rect 190380 994129 190408 995438
rect 191852 994294 191880 995438
rect 194336 995314 194364 995438
rect 194324 995308 194376 995314
rect 194324 995250 194376 995256
rect 194692 995172 194744 995178
rect 194692 995114 194744 995120
rect 192852 994832 192904 994838
rect 192852 994774 192904 994780
rect 192864 994430 192892 994774
rect 194704 994673 194732 995114
rect 194690 994664 194746 994673
rect 194690 994599 194746 994608
rect 192852 994424 192904 994430
rect 195072 994401 195100 995522
rect 195256 995314 195284 996639
rect 195532 996033 195560 999738
rect 195716 997257 195744 1005246
rect 198660 1001978 198688 1005994
rect 202696 1005304 202748 1005310
rect 202694 1005272 202696 1005281
rect 202748 1005272 202750 1005281
rect 202694 1005207 202750 1005216
rect 209226 1005136 209282 1005145
rect 209226 1005071 209228 1005080
rect 209280 1005071 209282 1005080
rect 211804 1005100 211856 1005106
rect 209228 1005042 209280 1005048
rect 211804 1005042 211856 1005048
rect 207570 1005000 207626 1005009
rect 207570 1004935 207572 1004944
rect 207624 1004935 207626 1004944
rect 209872 1004964 209924 1004970
rect 207572 1004906 207624 1004912
rect 209872 1004906 209924 1004912
rect 209226 1004728 209282 1004737
rect 209226 1004663 209228 1004672
rect 209280 1004663 209282 1004672
rect 209228 1004634 209280 1004640
rect 206374 1002280 206430 1002289
rect 203340 1002244 203392 1002250
rect 206374 1002215 206376 1002224
rect 203340 1002186 203392 1002192
rect 206428 1002215 206430 1002224
rect 206376 1002186 206428 1002192
rect 198648 1001972 198700 1001978
rect 198648 1001914 198700 1001920
rect 196624 998708 196676 998714
rect 196624 998650 196676 998656
rect 195702 997248 195758 997257
rect 195702 997183 195758 997192
rect 195518 996024 195574 996033
rect 195518 995959 195574 995968
rect 195244 995308 195296 995314
rect 195244 995250 195296 995256
rect 195244 994832 195296 994838
rect 195244 994774 195296 994780
rect 195256 994566 195284 994774
rect 195244 994560 195296 994566
rect 195244 994502 195296 994508
rect 192852 994366 192904 994372
rect 195058 994392 195114 994401
rect 195058 994327 195114 994336
rect 191840 994288 191892 994294
rect 191840 994230 191892 994236
rect 196636 994158 196664 998650
rect 199384 998572 199436 998578
rect 199384 998514 199436 998520
rect 196808 998300 196860 998306
rect 196808 998242 196860 998248
rect 196820 996441 196848 998242
rect 198648 998164 198700 998170
rect 198648 998106 198700 998112
rect 196806 996432 196862 996441
rect 196806 996367 196862 996376
rect 196624 994152 196676 994158
rect 190366 994120 190422 994129
rect 196624 994094 196676 994100
rect 190366 994055 190422 994064
rect 198660 991506 198688 998106
rect 199396 995178 199424 998514
rect 200856 998436 200908 998442
rect 200856 998378 200908 998384
rect 200670 998200 200726 998209
rect 200670 998135 200672 998144
rect 200724 998135 200726 998144
rect 200672 998106 200724 998112
rect 200028 998028 200080 998034
rect 200028 997970 200080 997976
rect 199384 995172 199436 995178
rect 199384 995114 199436 995120
rect 200040 991642 200068 997970
rect 200868 997914 200896 998378
rect 202694 998336 202750 998345
rect 202694 998271 202696 998280
rect 202748 998271 202750 998280
rect 202696 998242 202748 998248
rect 202144 998164 202196 998170
rect 202144 998106 202196 998112
rect 201866 998064 201922 998073
rect 201866 997999 201868 998008
rect 201920 997999 201922 998008
rect 201868 997970 201920 997976
rect 200776 997886 200896 997914
rect 200212 996464 200264 996470
rect 200210 996432 200212 996441
rect 200264 996432 200266 996441
rect 200210 996367 200266 996376
rect 200776 994129 200804 997886
rect 200948 997824 201000 997830
rect 200948 997766 201000 997772
rect 200960 995586 200988 997766
rect 200948 995580 201000 995586
rect 200948 995522 201000 995528
rect 202156 994430 202184 998106
rect 202328 997960 202380 997966
rect 202328 997902 202380 997908
rect 202340 995489 202368 997902
rect 202326 995480 202382 995489
rect 202326 995415 202382 995424
rect 203352 994945 203380 1002186
rect 205546 1002144 205602 1002153
rect 203708 1002108 203760 1002114
rect 205546 1002079 205548 1002088
rect 203708 1002050 203760 1002056
rect 205600 1002079 205602 1002088
rect 205548 1002050 205600 1002056
rect 203522 998608 203578 998617
rect 203522 998543 203524 998552
rect 203576 998543 203578 998552
rect 203524 998514 203576 998520
rect 203524 997824 203576 997830
rect 203522 997792 203524 997801
rect 203576 997792 203578 997801
rect 203522 997727 203578 997736
rect 203720 996470 203748 1002050
rect 206374 1002008 206430 1002017
rect 204904 1001972 204956 1001978
rect 204904 1001914 204956 1001920
rect 205652 1001966 206374 1001994
rect 204350 998744 204406 998753
rect 204350 998679 204352 998688
rect 204404 998679 204406 998688
rect 204352 998650 204404 998656
rect 203890 998472 203946 998481
rect 203890 998407 203892 998416
rect 203944 998407 203946 998416
rect 203892 998378 203944 998384
rect 204076 998164 204128 998170
rect 204076 998106 204128 998112
rect 203708 996464 203760 996470
rect 203708 996406 203760 996412
rect 204088 995897 204116 998106
rect 204720 997960 204772 997966
rect 204718 997928 204720 997937
rect 204772 997928 204774 997937
rect 204718 997863 204774 997872
rect 204074 995888 204130 995897
rect 204074 995823 204130 995832
rect 203338 994936 203394 994945
rect 203338 994871 203394 994880
rect 204916 994702 204944 1001914
rect 205652 994974 205680 1001966
rect 206374 1001943 206430 1001952
rect 206742 1002008 206798 1002017
rect 207570 1002008 207626 1002017
rect 206742 1001943 206744 1001952
rect 206796 1001943 206798 1001952
rect 207032 1001966 207570 1001994
rect 206744 1001914 206796 1001920
rect 205640 994968 205692 994974
rect 205640 994910 205692 994916
rect 207032 994838 207060 1001966
rect 207570 1001943 207626 1001952
rect 208398 1002008 208454 1002017
rect 208398 1001943 208454 1001952
rect 208412 996130 208440 1001943
rect 209884 999802 209912 1004906
rect 211160 1004692 211212 1004698
rect 211160 1004634 211212 1004640
rect 211172 1002538 211200 1004634
rect 211080 1002510 211200 1002538
rect 210054 1002280 210110 1002289
rect 210054 1002215 210056 1002224
rect 210108 1002215 210110 1002224
rect 210056 1002186 210108 1002192
rect 210422 1002008 210478 1002017
rect 210252 1001966 210422 1001994
rect 209872 999796 209924 999802
rect 209872 999738 209924 999744
rect 208400 996124 208452 996130
rect 208400 996066 208452 996072
rect 210252 995994 210280 1001966
rect 211080 1001994 211108 1002510
rect 211250 1002416 211306 1002425
rect 211250 1002351 211252 1002360
rect 211304 1002351 211306 1002360
rect 211252 1002322 211304 1002328
rect 211250 1002144 211306 1002153
rect 211250 1002079 211252 1002088
rect 211304 1002079 211306 1002088
rect 211252 1002050 211304 1002056
rect 211080 1001966 211200 1001994
rect 210422 1001943 210478 1001952
rect 210240 995988 210292 995994
rect 210240 995930 210292 995936
rect 211172 995858 211200 1001966
rect 211160 995852 211212 995858
rect 211160 995794 211212 995800
rect 211816 995314 211844 1005042
rect 212538 1004728 212594 1004737
rect 212538 1004663 212540 1004672
rect 212592 1004663 212594 1004672
rect 217324 1004692 217376 1004698
rect 212540 1004634 212592 1004640
rect 217324 1004634 217376 1004640
rect 215944 1002380 215996 1002386
rect 215944 1002322 215996 1002328
rect 212540 1002244 212592 1002250
rect 212540 1002186 212592 1002192
rect 212078 1002008 212134 1002017
rect 212078 1001943 212080 1001952
rect 212132 1001943 212134 1001952
rect 212080 1001914 212132 1001920
rect 212552 995450 212580 1002186
rect 213184 1002108 213236 1002114
rect 213184 1002050 213236 1002056
rect 213196 995858 213224 1002050
rect 213920 1001972 213972 1001978
rect 213920 1001914 213972 1001920
rect 213184 995852 213236 995858
rect 213184 995794 213236 995800
rect 212540 995444 212592 995450
rect 212540 995386 212592 995392
rect 211804 995308 211856 995314
rect 211804 995250 211856 995256
rect 207020 994832 207072 994838
rect 207020 994774 207072 994780
rect 204904 994696 204956 994702
rect 204904 994638 204956 994644
rect 213932 994430 213960 1001914
rect 202144 994424 202196 994430
rect 202144 994366 202196 994372
rect 207020 994424 207072 994430
rect 207020 994366 207072 994372
rect 213920 994424 213972 994430
rect 213920 994366 213972 994372
rect 200762 994120 200818 994129
rect 200762 994055 200818 994064
rect 200028 991636 200080 991642
rect 200028 991578 200080 991584
rect 198648 991500 198700 991506
rect 198648 991442 198700 991448
rect 207032 986678 207060 994366
rect 203156 986672 203208 986678
rect 203156 986614 203208 986620
rect 207020 986672 207072 986678
rect 207020 986614 207072 986620
rect 170324 983606 170798 983634
rect 186516 983606 186990 983634
rect 203168 983620 203196 986614
rect 215956 985998 215984 1002322
rect 217336 986678 217364 1004634
rect 228376 995994 228404 1006334
rect 249064 1006324 249116 1006330
rect 256146 1006295 256148 1006304
rect 249064 1006266 249116 1006272
rect 256200 1006295 256202 1006304
rect 256148 1006266 256200 1006272
rect 247040 1006188 247092 1006194
rect 247040 1006130 247092 1006136
rect 229744 1006052 229796 1006058
rect 229744 1005994 229796 1006000
rect 229006 997248 229062 997257
rect 229006 997183 229062 997192
rect 229190 997248 229246 997257
rect 229190 997183 229246 997192
rect 228364 995988 228416 995994
rect 228364 995930 228416 995936
rect 229020 994566 229048 997183
rect 229204 994974 229232 997183
rect 229756 996130 229784 1005994
rect 246764 1002584 246816 1002590
rect 246764 1002526 246816 1002532
rect 246580 1001224 246632 1001230
rect 246580 1001166 246632 1001172
rect 229744 996124 229796 996130
rect 229744 996066 229796 996072
rect 238574 995752 238630 995761
rect 239586 995752 239642 995761
rect 238630 995710 238740 995738
rect 239292 995710 239586 995738
rect 238574 995687 238630 995696
rect 242070 995752 242126 995761
rect 241776 995710 242070 995738
rect 239586 995687 239642 995696
rect 243266 995752 243322 995761
rect 242972 995710 243266 995738
rect 242070 995687 242126 995696
rect 243266 995687 243322 995696
rect 243818 995616 243874 995625
rect 243616 995574 243818 995602
rect 243818 995551 243874 995560
rect 244094 995616 244150 995625
rect 244150 995574 244260 995602
rect 246212 995580 246264 995586
rect 244094 995551 244150 995560
rect 246212 995522 246264 995528
rect 235906 995480 235962 995489
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 234416 995438 234568 995466
rect 229192 994968 229244 994974
rect 229192 994910 229244 994916
rect 231596 994838 231624 995438
rect 231584 994832 231636 994838
rect 231584 994774 231636 994780
rect 229008 994560 229060 994566
rect 229008 994502 229060 994508
rect 232240 994430 232268 995438
rect 232884 994702 232912 995438
rect 234540 994974 234568 995438
rect 234724 995438 234968 995466
rect 235612 995438 235906 995466
rect 234724 995110 234752 995438
rect 236256 995438 236592 995466
rect 239936 995438 240088 995466
rect 240580 995438 240916 995466
rect 245456 995438 245608 995466
rect 235906 995415 235962 995424
rect 234712 995104 234764 995110
rect 234712 995046 234764 995052
rect 234528 994968 234580 994974
rect 236564 994945 236592 995438
rect 234528 994910 234580 994916
rect 236550 994936 236606 994945
rect 236550 994871 236606 994880
rect 232872 994696 232924 994702
rect 232872 994638 232924 994644
rect 239404 994560 239456 994566
rect 239404 994502 239456 994508
rect 232228 994424 232280 994430
rect 232228 994366 232280 994372
rect 239416 994158 239444 994502
rect 239404 994152 239456 994158
rect 239404 994094 239456 994100
rect 240060 994022 240088 995438
rect 240888 994673 240916 995438
rect 245580 995353 245608 995438
rect 245566 995344 245622 995353
rect 244372 995308 244424 995314
rect 245566 995279 245622 995288
rect 244372 995250 244424 995256
rect 244096 995240 244148 995246
rect 244384 995194 244412 995250
rect 244148 995188 244412 995194
rect 244096 995182 244412 995188
rect 244108 995166 244412 995182
rect 240874 994664 240930 994673
rect 240874 994599 240930 994608
rect 246224 994022 246252 995522
rect 246592 995353 246620 1001166
rect 246776 996441 246804 1002526
rect 246762 996432 246818 996441
rect 246762 996367 246818 996376
rect 247052 995625 247080 1006130
rect 247868 998436 247920 998442
rect 247868 998378 247920 998384
rect 247684 998164 247736 998170
rect 247684 998106 247736 998112
rect 247224 997756 247276 997762
rect 247224 997698 247276 997704
rect 247236 997121 247264 997698
rect 247222 997112 247278 997121
rect 247222 997047 247278 997056
rect 247038 995616 247094 995625
rect 247038 995551 247094 995560
rect 246578 995344 246634 995353
rect 246578 995279 246634 995288
rect 247696 994673 247724 998106
rect 247880 996169 247908 998378
rect 247866 996160 247922 996169
rect 247866 996095 247922 996104
rect 247682 994664 247738 994673
rect 247682 994599 247738 994608
rect 249076 994158 249104 1006266
rect 252466 1006224 252522 1006233
rect 252466 1006159 252468 1006168
rect 252520 1006159 252522 1006168
rect 262678 1006224 262734 1006233
rect 262678 1006159 262680 1006168
rect 252468 1006130 252520 1006136
rect 262732 1006159 262734 1006168
rect 278044 1006188 278096 1006194
rect 262680 1006130 262732 1006136
rect 278044 1006130 278096 1006136
rect 254122 1006088 254178 1006097
rect 249800 1006052 249852 1006058
rect 254122 1006023 254124 1006032
rect 249800 1005994 249852 1006000
rect 254176 1006023 254178 1006032
rect 261850 1006088 261906 1006097
rect 261850 1006023 261852 1006032
rect 254124 1005994 254176 1006000
rect 261904 1006023 261906 1006032
rect 261852 1005994 261904 1006000
rect 249812 1004654 249840 1005994
rect 263048 1005304 263100 1005310
rect 263046 1005272 263048 1005281
rect 263100 1005272 263102 1005281
rect 263046 1005207 263102 1005216
rect 256514 1004728 256570 1004737
rect 250444 1004692 250496 1004698
rect 249812 1004626 249932 1004654
rect 256514 1004663 256516 1004672
rect 250444 1004634 250496 1004640
rect 256568 1004663 256570 1004672
rect 256516 1004634 256568 1004640
rect 249708 997892 249760 997898
rect 249708 997834 249760 997840
rect 249064 994152 249116 994158
rect 249064 994094 249116 994100
rect 240048 994016 240100 994022
rect 240048 993958 240100 993964
rect 246212 994016 246264 994022
rect 246212 993958 246264 993964
rect 249720 990146 249748 997834
rect 249904 996849 249932 1004626
rect 249890 996840 249946 996849
rect 249890 996775 249946 996784
rect 250456 994430 250484 1004634
rect 255318 1002824 255374 1002833
rect 252008 1002788 252060 1002794
rect 255318 1002759 255320 1002768
rect 252008 1002730 252060 1002736
rect 255372 1002759 255374 1002768
rect 255320 1002730 255372 1002736
rect 251824 1002244 251876 1002250
rect 251824 1002186 251876 1002192
rect 250996 998028 251048 998034
rect 250996 997970 251048 997976
rect 250444 994424 250496 994430
rect 250444 994366 250496 994372
rect 249708 990140 249760 990146
rect 249708 990082 249760 990088
rect 251008 988786 251036 997970
rect 251836 994945 251864 1002186
rect 252020 995586 252048 1002730
rect 255320 1002584 255372 1002590
rect 255318 1002552 255320 1002561
rect 255372 1002552 255374 1002561
rect 255318 1002487 255374 1002496
rect 261022 1002552 261078 1002561
rect 261022 1002487 261024 1002496
rect 261076 1002487 261078 1002496
rect 264244 1002516 264296 1002522
rect 261024 1002458 261076 1002464
rect 264244 1002458 264296 1002464
rect 254490 1002280 254546 1002289
rect 254490 1002215 254492 1002224
rect 254544 1002215 254546 1002224
rect 254492 1002186 254544 1002192
rect 256146 1002144 256202 1002153
rect 253480 1002108 253532 1002114
rect 256146 1002079 256148 1002088
rect 253480 1002050 253532 1002056
rect 256200 1002079 256202 1002088
rect 263506 1002144 263562 1002153
rect 263506 1002079 263508 1002088
rect 256148 1002050 256200 1002056
rect 263560 1002079 263562 1002088
rect 263508 1002050 263560 1002056
rect 253294 998064 253350 998073
rect 253294 997999 253296 998008
rect 253348 997999 253350 998008
rect 253296 997970 253348 997976
rect 252466 997928 252522 997937
rect 252466 997863 252468 997872
rect 252520 997863 252522 997872
rect 252468 997834 252520 997840
rect 253492 995897 253520 1002050
rect 261022 1002008 261078 1002017
rect 263874 1002008 263930 1002017
rect 261022 1001943 261024 1001952
rect 261076 1001943 261078 1001952
rect 263600 1001972 263652 1001978
rect 261024 1001914 261076 1001920
rect 263874 1001943 263876 1001952
rect 263600 1001914 263652 1001920
rect 263928 1001943 263930 1001952
rect 263876 1001914 263928 1001920
rect 256976 1001224 257028 1001230
rect 256974 1001192 256976 1001201
rect 257028 1001192 257030 1001201
rect 256974 1001127 257030 1001136
rect 258998 998472 259054 998481
rect 258998 998407 259000 998416
rect 259052 998407 259054 998416
rect 259000 998378 259052 998384
rect 254584 998232 254636 998238
rect 253662 998200 253718 998209
rect 257344 998232 257396 998238
rect 254584 998174 254636 998180
rect 257342 998200 257344 998209
rect 257396 998200 257398 998209
rect 253662 998135 253664 998144
rect 253716 998135 253718 998144
rect 253664 998106 253716 998112
rect 254596 997762 254624 998174
rect 257342 998135 257398 998144
rect 255964 998096 256016 998102
rect 258172 998096 258224 998102
rect 255964 998038 256016 998044
rect 258170 998064 258172 998073
rect 260196 998096 260248 998102
rect 258224 998064 258226 998073
rect 254584 997756 254636 997762
rect 254584 997698 254636 997704
rect 253478 995888 253534 995897
rect 253478 995823 253534 995832
rect 252008 995580 252060 995586
rect 252008 995522 252060 995528
rect 251822 994936 251878 994945
rect 251822 994871 251878 994880
rect 255976 994838 256004 998038
rect 258170 997999 258226 998008
rect 260194 998064 260196 998073
rect 262864 998096 262916 998102
rect 260248 998064 260250 998073
rect 262864 998038 262916 998044
rect 260194 997999 260250 998008
rect 257344 997960 257396 997966
rect 259000 997960 259052 997966
rect 257344 997902 257396 997908
rect 258998 997928 259000 997937
rect 259828 997960 259880 997966
rect 259052 997928 259054 997937
rect 255964 994832 256016 994838
rect 255964 994774 256016 994780
rect 257356 994702 257384 997902
rect 258998 997863 259054 997872
rect 259826 997928 259828 997937
rect 262220 997960 262272 997966
rect 259880 997928 259882 997937
rect 262220 997902 262272 997908
rect 259826 997863 259882 997872
rect 258172 997824 258224 997830
rect 258170 997792 258172 997801
rect 259460 997824 259512 997830
rect 258224 997792 258226 997801
rect 260196 997824 260248 997830
rect 259460 997766 259512 997772
rect 260194 997792 260196 997801
rect 260932 997824 260984 997830
rect 260248 997792 260250 997801
rect 258170 997727 258226 997736
rect 259472 994974 259500 997766
rect 260932 997766 260984 997772
rect 261850 997792 261906 997801
rect 260194 997727 260250 997736
rect 260944 995314 260972 997766
rect 261128 997736 261850 997754
rect 261128 997727 261906 997736
rect 261128 997726 261892 997727
rect 261128 995858 261156 997726
rect 262232 996130 262260 997902
rect 262220 996124 262272 996130
rect 262220 996066 262272 996072
rect 261116 995852 261168 995858
rect 261116 995794 261168 995800
rect 262876 995450 262904 998038
rect 263612 995994 263640 1001914
rect 264256 995994 264284 1002458
rect 265624 1002108 265676 1002114
rect 265624 1002050 265676 1002056
rect 263600 995988 263652 995994
rect 263600 995930 263652 995936
rect 264244 995988 264296 995994
rect 264244 995930 264296 995936
rect 262864 995444 262916 995450
rect 262864 995386 262916 995392
rect 260932 995308 260984 995314
rect 260932 995250 260984 995256
rect 259460 994968 259512 994974
rect 259460 994910 259512 994916
rect 257344 994696 257396 994702
rect 257344 994638 257396 994644
rect 251456 994288 251508 994294
rect 251456 994230 251508 994236
rect 250996 988780 251048 988786
rect 250996 988722 251048 988728
rect 217324 986672 217376 986678
rect 217324 986614 217376 986620
rect 219440 986672 219492 986678
rect 219440 986614 219492 986620
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 219452 983620 219480 986614
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 235644 983620 235672 985934
rect 251468 983634 251496 994230
rect 265636 994158 265664 1002050
rect 267004 1001972 267056 1001978
rect 267004 1001914 267056 1001920
rect 265624 994152 265676 994158
rect 265624 994094 265676 994100
rect 267016 991778 267044 1001914
rect 278056 996130 278084 1006130
rect 280804 1006052 280856 1006058
rect 280804 1005994 280856 1006000
rect 279424 1005304 279476 1005310
rect 279424 1005246 279476 1005252
rect 278044 996124 278096 996130
rect 278044 996066 278096 996072
rect 267740 994152 267792 994158
rect 267740 994094 267792 994100
rect 267004 991772 267056 991778
rect 267004 991714 267056 991720
rect 267752 983634 267780 994094
rect 279436 985998 279464 1005246
rect 280816 995858 280844 1005994
rect 298652 1003332 298704 1003338
rect 298652 1003274 298704 1003280
rect 298098 1002280 298154 1002289
rect 298098 1002215 298154 1002224
rect 280804 995852 280856 995858
rect 280804 995794 280856 995800
rect 298112 995761 298140 1002215
rect 298282 997928 298338 997937
rect 298282 997863 298338 997872
rect 292486 995752 292542 995761
rect 292146 995710 292486 995738
rect 292486 995687 292542 995696
rect 295062 995752 295118 995761
rect 296166 995752 296222 995761
rect 295118 995710 295182 995738
rect 295826 995710 296166 995738
rect 295062 995687 295118 995696
rect 296166 995687 296222 995696
rect 298098 995752 298154 995761
rect 298098 995687 298154 995696
rect 280710 995616 280766 995625
rect 298296 995602 298324 997863
rect 280710 995551 280766 995560
rect 297836 995574 298324 995602
rect 298468 995580 298520 995586
rect 280724 993206 280752 995551
rect 294878 995480 294934 995489
rect 282840 994430 282868 995452
rect 283484 994566 283512 995452
rect 283472 994560 283524 994566
rect 283472 994502 283524 994508
rect 282828 994424 282880 994430
rect 282828 994366 282880 994372
rect 284128 994294 284156 995452
rect 285968 994702 285996 995452
rect 286520 994974 286548 995452
rect 287178 995438 287560 995466
rect 286508 994968 286560 994974
rect 286508 994910 286560 994916
rect 285956 994696 286008 994702
rect 285956 994638 286008 994644
rect 284116 994288 284168 994294
rect 284116 994230 284168 994236
rect 287532 993993 287560 995438
rect 287808 994809 287836 995452
rect 290292 995081 290320 995452
rect 290858 995438 291148 995466
rect 291120 995314 291148 995438
rect 291108 995308 291160 995314
rect 291108 995250 291160 995256
rect 290278 995072 290334 995081
rect 290278 995007 290334 995016
rect 287794 994800 287850 994809
rect 287794 994735 287850 994744
rect 289452 994696 289504 994702
rect 289452 994638 289504 994644
rect 289464 994158 289492 994638
rect 291488 994265 291516 995452
rect 293342 995438 293632 995466
rect 294538 995438 294878 995466
rect 293604 995178 293632 995438
rect 297022 995438 297404 995466
rect 294878 995415 294934 995424
rect 297376 995330 297404 995438
rect 297836 995330 297864 995574
rect 298468 995522 298520 995528
rect 298480 995466 298508 995522
rect 298664 995489 298692 1003274
rect 298848 1001894 298876 1006538
rect 307758 1006496 307814 1006505
rect 300308 1006460 300360 1006466
rect 307758 1006431 307760 1006440
rect 300308 1006402 300360 1006408
rect 307812 1006431 307814 1006440
rect 360198 1006496 360254 1006505
rect 360198 1006431 360200 1006440
rect 307760 1006402 307812 1006408
rect 360252 1006431 360254 1006440
rect 360200 1006402 360252 1006408
rect 299296 1006324 299348 1006330
rect 299296 1006266 299348 1006272
rect 298756 1001866 298876 1001894
rect 298756 995602 298784 1001866
rect 298928 999184 298980 999190
rect 298928 999126 298980 999132
rect 298940 996033 298968 999126
rect 299112 997756 299164 997762
rect 299112 997698 299164 997704
rect 299124 996441 299152 997698
rect 299110 996432 299166 996441
rect 299110 996367 299166 996376
rect 298926 996024 298982 996033
rect 299308 995994 299336 1006266
rect 300124 1006188 300176 1006194
rect 300124 1006130 300176 1006136
rect 298926 995959 298982 995968
rect 299296 995988 299348 995994
rect 299296 995930 299348 995936
rect 298756 995574 298876 995602
rect 297376 995302 297864 995330
rect 298020 995438 298508 995466
rect 298650 995480 298706 995489
rect 293592 995172 293644 995178
rect 293592 995114 293644 995120
rect 291474 994256 291530 994265
rect 291474 994191 291530 994200
rect 289452 994152 289504 994158
rect 289452 994094 289504 994100
rect 298020 993993 298048 995438
rect 298650 995415 298706 995424
rect 298848 995178 298876 995574
rect 298836 995172 298888 995178
rect 298836 995114 298888 995120
rect 300136 994809 300164 1006130
rect 300320 994974 300348 1006402
rect 314658 1006360 314714 1006369
rect 311808 1006324 311860 1006330
rect 360566 1006360 360622 1006369
rect 314658 1006295 314660 1006304
rect 311808 1006266 311860 1006272
rect 314712 1006295 314714 1006304
rect 319444 1006324 319496 1006330
rect 314660 1006266 314712 1006272
rect 360566 1006295 360568 1006304
rect 319444 1006266 319496 1006272
rect 360620 1006295 360622 1006304
rect 360568 1006266 360620 1006272
rect 306102 1006224 306158 1006233
rect 306102 1006159 306104 1006168
rect 306156 1006159 306158 1006168
rect 306104 1006130 306156 1006136
rect 311820 1006097 311848 1006266
rect 304078 1006088 304134 1006097
rect 302148 1006052 302200 1006058
rect 304078 1006023 304080 1006032
rect 302148 1005994 302200 1006000
rect 304132 1006023 304134 1006032
rect 311806 1006088 311862 1006097
rect 311806 1006023 311862 1006032
rect 314658 1006088 314714 1006097
rect 314658 1006023 314660 1006032
rect 304080 1005994 304132 1006000
rect 314712 1006023 314714 1006032
rect 314660 1005994 314712 1006000
rect 302160 1002289 302188 1005994
rect 313830 1004864 313886 1004873
rect 313830 1004799 313832 1004808
rect 313884 1004799 313886 1004808
rect 316040 1004828 316092 1004834
rect 313832 1004770 313884 1004776
rect 316040 1004770 316092 1004776
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 302146 1002280 302202 1002289
rect 302146 1002215 302202 1002224
rect 310978 1002144 311034 1002153
rect 310978 1002079 310980 1002088
rect 311032 1002079 311034 1002088
rect 313280 1002108 313332 1002114
rect 310980 1002050 311032 1002056
rect 313280 1002050 313332 1002056
rect 310150 1002008 310206 1002017
rect 312634 1002008 312690 1002017
rect 310150 1001943 310152 1001952
rect 310204 1001943 310206 1001952
rect 311900 1001972 311952 1001978
rect 310152 1001914 310204 1001920
rect 312634 1001943 312636 1001952
rect 311900 1001914 311952 1001920
rect 312688 1001943 312690 1001952
rect 312636 1001914 312688 1001920
rect 305276 999184 305328 999190
rect 305274 999152 305276 999161
rect 305328 999152 305330 999161
rect 305274 999087 305330 999096
rect 308954 998608 309010 998617
rect 303252 998572 303304 998578
rect 308954 998543 308956 998552
rect 303252 998514 303304 998520
rect 309008 998543 309010 998552
rect 308956 998514 309008 998520
rect 302884 998300 302936 998306
rect 302884 998242 302936 998248
rect 302146 995616 302202 995625
rect 302146 995551 302202 995560
rect 300308 994968 300360 994974
rect 300308 994910 300360 994916
rect 300122 994800 300178 994809
rect 300122 994735 300178 994744
rect 301504 994560 301556 994566
rect 301504 994502 301556 994508
rect 301516 994158 301544 994502
rect 301504 994152 301556 994158
rect 301504 994094 301556 994100
rect 287518 993984 287574 993993
rect 287518 993919 287574 993928
rect 298006 993984 298062 993993
rect 298006 993919 298062 993928
rect 280712 993200 280764 993206
rect 280712 993142 280764 993148
rect 284300 991772 284352 991778
rect 284300 991714 284352 991720
rect 279424 985992 279476 985998
rect 279424 985934 279476 985940
rect 251468 983606 251850 983634
rect 267752 983606 268134 983634
rect 284312 983620 284340 991714
rect 300492 985992 300544 985998
rect 300492 985934 300544 985940
rect 300504 983620 300532 985934
rect 302160 984774 302188 995551
rect 302896 995314 302924 998242
rect 303264 997937 303292 998514
rect 307298 998472 307354 998481
rect 304448 998436 304500 998442
rect 307298 998407 307300 998416
rect 304448 998378 304500 998384
rect 307352 998407 307354 998416
rect 307300 998378 307352 998384
rect 304264 998028 304316 998034
rect 304264 997970 304316 997976
rect 303250 997928 303306 997937
rect 303250 997863 303306 997872
rect 303528 997892 303580 997898
rect 303528 997834 303580 997840
rect 302884 995308 302936 995314
rect 302884 995250 302936 995256
rect 303540 990282 303568 997834
rect 304276 994265 304304 997970
rect 304460 995586 304488 998378
rect 306102 998336 306158 998345
rect 306102 998271 306104 998280
rect 306156 998271 306158 998280
rect 310610 998336 310666 998345
rect 310610 998271 310666 998280
rect 306104 998242 306156 998248
rect 308126 998200 308182 998209
rect 305644 998164 305696 998170
rect 310624 998186 310652 998271
rect 308126 998135 308128 998144
rect 305644 998106 305696 998112
rect 308180 998135 308182 998144
rect 310440 998158 310652 998186
rect 308128 998106 308180 998112
rect 304906 997928 304962 997937
rect 304906 997863 304908 997872
rect 304960 997863 304962 997872
rect 304908 997834 304960 997840
rect 304448 995580 304500 995586
rect 304448 995522 304500 995528
rect 305656 994838 305684 998106
rect 306930 998064 306986 998073
rect 306930 997999 306932 998008
rect 306984 997999 306986 998008
rect 308404 998028 308456 998034
rect 306932 997970 306984 997976
rect 308404 997970 308456 997976
rect 307024 997892 307076 997898
rect 307024 997834 307076 997840
rect 307036 995081 307064 997834
rect 307022 995072 307078 995081
rect 307022 995007 307078 995016
rect 305644 994832 305696 994838
rect 305644 994774 305696 994780
rect 308416 994430 308444 997970
rect 308954 997928 309010 997937
rect 308954 997863 308956 997872
rect 309008 997863 309010 997872
rect 308956 997834 309008 997840
rect 309782 997792 309838 997801
rect 310440 997762 310468 998158
rect 310610 998064 310666 998073
rect 310610 997999 310612 998008
rect 310664 997999 310666 998008
rect 310612 997970 310664 997976
rect 309782 997727 309838 997736
rect 310428 997756 310480 997762
rect 309796 994566 309824 997727
rect 310428 997698 310480 997704
rect 311912 994702 311940 1001914
rect 313292 995450 313320 1002050
rect 314660 1001972 314712 1001978
rect 314660 1001914 314712 1001920
rect 314672 995858 314700 1001914
rect 316052 996130 316080 1004770
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 318076 997082 318104 1004634
rect 319456 997354 319484 1006266
rect 365260 1006188 365312 1006194
rect 365260 1006130 365312 1006136
rect 354862 1006088 354918 1006097
rect 323584 1006052 323636 1006058
rect 323584 1005994 323636 1006000
rect 354588 1006052 354640 1006058
rect 354862 1006023 354864 1006032
rect 354588 1005994 354640 1006000
rect 354916 1006023 354918 1006032
rect 355690 1006088 355746 1006097
rect 361394 1006088 361450 1006097
rect 355690 1006023 355692 1006032
rect 354864 1005994 354916 1006000
rect 355744 1006023 355746 1006032
rect 359556 1006052 359608 1006058
rect 355692 1005994 355744 1006000
rect 361394 1006023 361396 1006032
rect 359556 1005994 359608 1006000
rect 361448 1006023 361450 1006032
rect 365074 1006088 365130 1006097
rect 365074 1006023 365076 1006032
rect 361396 1005994 361448 1006000
rect 365128 1006023 365130 1006032
rect 365076 1005994 365128 1006000
rect 319444 997348 319496 997354
rect 319444 997290 319496 997296
rect 318064 997076 318116 997082
rect 318064 997018 318116 997024
rect 316040 996124 316092 996130
rect 316040 996066 316092 996072
rect 314660 995852 314712 995858
rect 314660 995794 314712 995800
rect 323596 995586 323624 1005994
rect 352840 1004828 352892 1004834
rect 352840 1004770 352892 1004776
rect 331128 1003332 331180 1003338
rect 331128 1003274 331180 1003280
rect 331140 997218 331168 1003274
rect 351828 1001972 351880 1001978
rect 351828 1001914 351880 1001920
rect 332600 997348 332652 997354
rect 332600 997290 332652 997296
rect 331128 997212 331180 997218
rect 331128 997154 331180 997160
rect 323584 995580 323636 995586
rect 323584 995522 323636 995528
rect 313280 995444 313332 995450
rect 313280 995386 313332 995392
rect 311900 994696 311952 994702
rect 311900 994638 311952 994644
rect 309784 994560 309836 994566
rect 309784 994502 309836 994508
rect 308404 994424 308456 994430
rect 308404 994366 308456 994372
rect 304262 994256 304318 994265
rect 304262 994191 304318 994200
rect 316408 993200 316460 993206
rect 316408 993142 316460 993148
rect 303528 990276 303580 990282
rect 303528 990218 303580 990224
rect 302148 984768 302200 984774
rect 302148 984710 302200 984716
rect 316420 983634 316448 993142
rect 332612 983634 332640 997290
rect 349160 997076 349212 997082
rect 349160 997018 349212 997024
rect 316420 983606 316802 983634
rect 332612 983606 332994 983634
rect 349172 983620 349200 997018
rect 351840 993206 351868 1001914
rect 351828 993200 351880 993206
rect 351828 993142 351880 993148
rect 352852 987562 352880 1004770
rect 354600 1002862 354628 1005994
rect 355690 1004864 355746 1004873
rect 355690 1004799 355692 1004808
rect 355744 1004799 355746 1004808
rect 355692 1004770 355744 1004776
rect 356520 1003944 356572 1003950
rect 356518 1003912 356520 1003921
rect 356572 1003912 356574 1003921
rect 356518 1003847 356574 1003856
rect 354588 1002856 354640 1002862
rect 354588 1002798 354640 1002804
rect 355140 1002856 355192 1002862
rect 355140 1002798 355192 1002804
rect 354034 1002008 354090 1002017
rect 354034 1001943 354036 1001952
rect 354088 1001943 354090 1001952
rect 354036 1001914 354088 1001920
rect 355152 998578 355180 1002798
rect 358542 1002144 358598 1002153
rect 355784 1002108 355836 1002114
rect 358542 1002079 358544 1002088
rect 355784 1002050 355836 1002056
rect 358596 1002079 358598 1002088
rect 358544 1002050 358596 1002056
rect 355796 1001230 355824 1002050
rect 356518 1002008 356574 1002017
rect 356060 1001972 356112 1001978
rect 356518 1001943 356520 1001952
rect 356060 1001914 356112 1001920
rect 356572 1001943 356574 1001952
rect 357346 1002008 357402 1002017
rect 359370 1002008 359426 1002017
rect 357346 1001943 357348 1001952
rect 356520 1001914 356572 1001920
rect 357400 1001943 357402 1001952
rect 358740 1001966 359370 1001994
rect 357348 1001914 357400 1001920
rect 355784 1001224 355836 1001230
rect 355784 1001166 355836 1001172
rect 355140 998572 355192 998578
rect 355140 998514 355192 998520
rect 356072 998442 356100 1001914
rect 356060 998436 356112 998442
rect 356060 998378 356112 998384
rect 357348 997212 357400 997218
rect 357348 997154 357400 997160
rect 357360 994294 357388 997154
rect 358740 995042 358768 1001966
rect 359370 1001943 359426 1001952
rect 358728 995036 358780 995042
rect 358728 994978 358780 994984
rect 359568 994906 359596 1005994
rect 360568 1005304 360620 1005310
rect 360566 1005272 360568 1005281
rect 360620 1005272 360622 1005281
rect 360566 1005207 360622 1005216
rect 363418 1005136 363474 1005145
rect 363418 1005071 363420 1005080
rect 363472 1005071 363474 1005080
rect 363420 1005042 363472 1005048
rect 365074 1005000 365130 1005009
rect 365074 1004935 365076 1004944
rect 365128 1004935 365130 1004944
rect 365076 1004906 365128 1004912
rect 362590 1004864 362646 1004873
rect 362590 1004799 362592 1004808
rect 362644 1004799 362646 1004808
rect 364984 1004828 365036 1004834
rect 362592 1004770 362644 1004776
rect 364984 1004770 365036 1004776
rect 364246 1004728 364302 1004737
rect 364246 1004663 364248 1004672
rect 364300 1004663 364302 1004672
rect 364248 1004634 364300 1004640
rect 359738 1002144 359794 1002153
rect 359738 1002079 359740 1002088
rect 359792 1002079 359794 1002088
rect 362224 1002108 362276 1002114
rect 359740 1002050 359792 1002056
rect 362224 1002050 362276 1002056
rect 361394 1002008 361450 1002017
rect 360844 1001972 360896 1001978
rect 361394 1001943 361396 1001952
rect 360844 1001914 360896 1001920
rect 361448 1001943 361450 1001952
rect 361396 1001914 361448 1001920
rect 360856 997082 360884 1001914
rect 360844 997076 360896 997082
rect 360844 997018 360896 997024
rect 359556 994900 359608 994906
rect 359556 994842 359608 994848
rect 362236 994634 362264 1002050
rect 363604 1001972 363656 1001978
rect 363604 1001914 363656 1001920
rect 363616 997762 363644 1001914
rect 363604 997756 363656 997762
rect 363604 997698 363656 997704
rect 364996 995858 365024 1004770
rect 365272 995994 365300 1006130
rect 368952 1006058 368980 1007082
rect 505376 1007072 505428 1007078
rect 425518 1007040 425574 1007049
rect 373264 1007004 373316 1007010
rect 505374 1007040 505376 1007049
rect 505428 1007040 505430 1007049
rect 425518 1006975 425520 1006984
rect 373264 1006946 373316 1006952
rect 425572 1006975 425574 1006984
rect 439688 1007004 439740 1007010
rect 425520 1006946 425572 1006952
rect 505374 1006975 505430 1006984
rect 439688 1006946 439740 1006952
rect 369124 1006800 369176 1006806
rect 369124 1006742 369176 1006748
rect 369136 1006330 369164 1006742
rect 369124 1006324 369176 1006330
rect 369124 1006266 369176 1006272
rect 371884 1006188 371936 1006194
rect 371884 1006130 371936 1006136
rect 367744 1006052 367796 1006058
rect 367744 1005994 367796 1006000
rect 368940 1006052 368992 1006058
rect 368940 1005994 368992 1006000
rect 366364 1005100 366416 1005106
rect 366364 1005042 366416 1005048
rect 365902 1002008 365958 1002017
rect 365902 1001943 365904 1001952
rect 365956 1001943 365958 1001952
rect 365904 1001914 365956 1001920
rect 365260 995988 365312 995994
rect 365260 995930 365312 995936
rect 364984 995852 365036 995858
rect 364984 995794 365036 995800
rect 366376 995586 366404 1005042
rect 366548 1004692 366600 1004698
rect 366548 1004634 366600 1004640
rect 366560 996130 366588 1004634
rect 366548 996124 366600 996130
rect 366548 996066 366600 996072
rect 364984 995580 365036 995586
rect 364984 995522 365036 995528
rect 366364 995580 366416 995586
rect 366364 995522 366416 995528
rect 362224 994628 362276 994634
rect 362224 994570 362276 994576
rect 357348 994288 357400 994294
rect 357348 994230 357400 994236
rect 352840 987556 352892 987562
rect 352840 987498 352892 987504
rect 364996 983634 365024 995522
rect 367756 991778 367784 1005994
rect 370504 1004964 370556 1004970
rect 370504 1004906 370556 1004912
rect 369124 1001972 369176 1001978
rect 369124 1001914 369176 1001920
rect 367744 991772 367796 991778
rect 367744 991714 367796 991720
rect 369136 985998 369164 1001914
rect 370516 986134 370544 1004906
rect 371896 994770 371924 1006130
rect 373276 999122 373304 1006946
rect 427542 1006904 427598 1006913
rect 427542 1006839 427544 1006848
rect 427596 1006839 427598 1006848
rect 438124 1006868 438176 1006874
rect 427544 1006810 427596 1006816
rect 438124 1006810 438176 1006816
rect 430854 1006768 430910 1006777
rect 400864 1006732 400916 1006738
rect 430854 1006703 430856 1006712
rect 400864 1006674 400916 1006680
rect 430908 1006703 430910 1006712
rect 430856 1006674 430908 1006680
rect 376024 1006460 376076 1006466
rect 376024 1006402 376076 1006408
rect 374644 1006324 374696 1006330
rect 374644 1006266 374696 1006272
rect 373264 999116 373316 999122
rect 373264 999058 373316 999064
rect 372344 997756 372396 997762
rect 372344 997698 372396 997704
rect 372356 996441 372384 997698
rect 372342 996432 372398 996441
rect 372342 996367 372398 996376
rect 374656 995081 374684 1006266
rect 375564 999116 375616 999122
rect 375564 999058 375616 999064
rect 374642 995072 374698 995081
rect 374642 995007 374698 995016
rect 375576 994809 375604 999058
rect 376036 996985 376064 1006402
rect 378140 1006052 378192 1006058
rect 378140 1005994 378192 1006000
rect 377404 1005304 377456 1005310
rect 377404 1005246 377456 1005252
rect 377416 998646 377444 1005246
rect 378152 999190 378180 1005994
rect 381452 1003944 381504 1003950
rect 381452 1003886 381504 1003892
rect 378784 1001224 378836 1001230
rect 378784 1001166 378836 1001172
rect 378140 999184 378192 999190
rect 378140 999126 378192 999132
rect 378600 998776 378652 998782
rect 378600 998718 378652 998724
rect 377404 998640 377456 998646
rect 377404 998582 377456 998588
rect 376022 996976 376078 996985
rect 376022 996911 376078 996920
rect 375562 994800 375618 994809
rect 371884 994764 371936 994770
rect 375562 994735 375618 994744
rect 371884 994706 371936 994712
rect 378612 994158 378640 998718
rect 378796 997830 378824 1001166
rect 378784 997824 378836 997830
rect 378784 997766 378836 997772
rect 380900 997076 380952 997082
rect 380900 997018 380952 997024
rect 380912 994498 380940 997018
rect 381464 995353 381492 1003886
rect 383292 999184 383344 999190
rect 383292 999126 383344 999132
rect 383108 997824 383160 997830
rect 383108 997766 383160 997772
rect 383120 995761 383148 997766
rect 383304 997665 383332 999126
rect 383568 998640 383620 998646
rect 383620 998588 383700 998594
rect 383568 998582 383700 998588
rect 383580 998566 383700 998582
rect 383476 998436 383528 998442
rect 383476 998378 383528 998384
rect 383290 997656 383346 997665
rect 383290 997591 383346 997600
rect 383488 997257 383516 998378
rect 383474 997248 383530 997257
rect 383474 997183 383530 997192
rect 383106 995752 383162 995761
rect 383106 995687 383162 995696
rect 381450 995344 381506 995353
rect 383672 995330 383700 998566
rect 385038 995752 385094 995761
rect 385774 995752 385830 995761
rect 385094 995710 385342 995738
rect 385038 995687 385094 995696
rect 387890 995752 387946 995761
rect 385830 995710 385986 995738
rect 387826 995710 387890 995738
rect 385774 995687 385830 995696
rect 387890 995687 387946 995696
rect 388718 995752 388774 995761
rect 389362 995752 389418 995761
rect 388774 995710 389022 995738
rect 388718 995687 388774 995696
rect 392398 995752 392454 995761
rect 389418 995710 389666 995738
rect 392150 995710 392398 995738
rect 389362 995687 389418 995696
rect 396538 995752 396594 995761
rect 396382 995710 396538 995738
rect 392398 995687 392454 995696
rect 396538 995687 396594 995696
rect 384316 995438 384698 995466
rect 384316 995330 384344 995438
rect 383672 995302 384344 995330
rect 381450 995279 381506 995288
rect 388364 995081 388392 995452
rect 392320 995438 392702 995466
rect 392320 995353 392348 995438
rect 392306 995344 392362 995353
rect 392306 995279 392362 995288
rect 388350 995072 388406 995081
rect 388350 995007 388406 995016
rect 393332 994770 393360 995452
rect 393502 995344 393558 995353
rect 393502 995279 393558 995288
rect 388076 994764 388128 994770
rect 388076 994706 388128 994712
rect 388260 994764 388312 994770
rect 388260 994706 388312 994712
rect 393320 994764 393372 994770
rect 393320 994706 393372 994712
rect 380900 994492 380952 994498
rect 380900 994434 380952 994440
rect 381176 994288 381228 994294
rect 381176 994230 381228 994236
rect 378600 994152 378652 994158
rect 378600 994094 378652 994100
rect 370504 986128 370556 986134
rect 370504 986070 370556 986076
rect 369124 985992 369176 985998
rect 369124 985934 369176 985940
rect 381188 983634 381216 994230
rect 388088 994226 388116 994706
rect 388272 994498 388300 994706
rect 393516 994634 393544 995279
rect 393976 994906 394004 995452
rect 393964 994900 394016 994906
rect 393964 994842 394016 994848
rect 395172 994809 395200 995452
rect 397012 994974 397040 995452
rect 397000 994968 397052 994974
rect 397000 994910 397052 994916
rect 395158 994800 395214 994809
rect 395158 994735 395214 994744
rect 393504 994628 393556 994634
rect 393504 994570 393556 994576
rect 397656 994498 397684 995452
rect 398852 995110 398880 995452
rect 400876 995382 400904 1006674
rect 429198 1006632 429254 1006641
rect 429198 1006567 429200 1006576
rect 429252 1006567 429254 1006576
rect 429200 1006538 429252 1006544
rect 425150 1006360 425206 1006369
rect 425150 1006295 425152 1006304
rect 425204 1006295 425206 1006304
rect 425152 1006266 425204 1006272
rect 423494 1006224 423550 1006233
rect 422024 1006188 422076 1006194
rect 423494 1006159 423496 1006168
rect 422024 1006130 422076 1006136
rect 423548 1006159 423550 1006168
rect 423496 1006130 423548 1006136
rect 422036 1003950 422064 1006130
rect 422666 1006088 422722 1006097
rect 430026 1006088 430082 1006097
rect 422666 1006023 422668 1006032
rect 422720 1006023 422722 1006032
rect 429844 1006052 429896 1006058
rect 422668 1005994 422720 1006000
rect 430026 1006023 430028 1006032
rect 429844 1005994 429896 1006000
rect 430080 1006023 430082 1006032
rect 430028 1005994 430080 1006000
rect 423496 1005712 423548 1005718
rect 423494 1005680 423496 1005689
rect 423548 1005680 423550 1005689
rect 423494 1005615 423550 1005624
rect 428372 1005576 428424 1005582
rect 428370 1005544 428372 1005553
rect 428424 1005544 428426 1005553
rect 428370 1005479 428426 1005488
rect 427174 1005408 427230 1005417
rect 427174 1005343 427176 1005352
rect 427228 1005343 427230 1005352
rect 427176 1005314 427228 1005320
rect 429198 1005000 429254 1005009
rect 429198 1004935 429200 1004944
rect 429252 1004935 429254 1004944
rect 429200 1004906 429252 1004912
rect 422666 1004728 422722 1004737
rect 422220 1004686 422666 1004714
rect 422024 1003944 422076 1003950
rect 422024 1003886 422076 1003892
rect 421470 1002008 421526 1002017
rect 419448 1001972 419500 1001978
rect 421470 1001943 421472 1001952
rect 419448 1001914 419500 1001920
rect 421524 1001943 421526 1001952
rect 421472 1001914 421524 1001920
rect 400864 995376 400916 995382
rect 400864 995318 400916 995324
rect 402980 995376 403032 995382
rect 402980 995318 403032 995324
rect 398840 995104 398892 995110
rect 398840 995046 398892 995052
rect 402992 994498 403020 995318
rect 388260 994492 388312 994498
rect 388260 994434 388312 994440
rect 397644 994492 397696 994498
rect 397644 994434 397696 994440
rect 402980 994492 403032 994498
rect 402980 994434 403032 994440
rect 388076 994220 388128 994226
rect 388076 994162 388128 994168
rect 419460 991778 419488 1001914
rect 421012 996464 421064 996470
rect 421010 996432 421012 996441
rect 421064 996432 421066 996441
rect 421010 996367 421066 996376
rect 415032 991772 415084 991778
rect 415032 991714 415084 991720
rect 419448 991772 419500 991778
rect 419448 991714 419500 991720
rect 397828 986128 397880 986134
rect 397828 986070 397880 986076
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 986070
rect 415044 985998 415072 991714
rect 422220 988922 422248 1004686
rect 422666 1004663 422722 1004672
rect 424692 1002720 424744 1002726
rect 424690 1002688 424692 1002697
rect 424744 1002688 424746 1002697
rect 424690 1002623 424746 1002632
rect 426348 1002584 426400 1002590
rect 426346 1002552 426348 1002561
rect 426400 1002552 426402 1002561
rect 426346 1002487 426402 1002496
rect 428002 1002280 428058 1002289
rect 428002 1002215 428004 1002224
rect 428056 1002215 428058 1002224
rect 428004 1002186 428056 1002192
rect 425150 1002144 425206 1002153
rect 423588 1002108 423640 1002114
rect 425150 1002079 425152 1002088
rect 423588 1002050 423640 1002056
rect 425204 1002079 425206 1002088
rect 428370 1002144 428426 1002153
rect 428370 1002079 428372 1002088
rect 425152 1002050 425204 1002056
rect 428424 1002079 428426 1002088
rect 428372 1002050 428424 1002056
rect 423600 998442 423628 1002050
rect 424322 1002008 424378 1002017
rect 426346 1002008 426402 1002017
rect 424322 1001943 424324 1001952
rect 424376 1001943 424378 1001952
rect 425060 1001972 425112 1001978
rect 424324 1001914 424376 1001920
rect 426346 1001943 426348 1001952
rect 425060 1001914 425112 1001920
rect 426400 1001943 426402 1001952
rect 428464 1001972 428516 1001978
rect 426348 1001914 426400 1001920
rect 428464 1001914 428516 1001920
rect 425072 998578 425100 1001914
rect 428476 998850 428504 1001914
rect 428464 998844 428516 998850
rect 428464 998786 428516 998792
rect 425060 998572 425112 998578
rect 425060 998514 425112 998520
rect 423588 998436 423640 998442
rect 423588 998378 423640 998384
rect 426440 996464 426492 996470
rect 426440 996406 426492 996412
rect 426452 994294 426480 996406
rect 429856 994974 429884 1005994
rect 432052 1005848 432104 1005854
rect 432050 1005816 432052 1005825
rect 433524 1005848 433576 1005854
rect 432104 1005816 432106 1005825
rect 433524 1005790 433576 1005796
rect 432050 1005751 432106 1005760
rect 430854 1005272 430910 1005281
rect 431926 1005242 432276 1005258
rect 430854 1005207 430856 1005216
rect 430908 1005207 430910 1005216
rect 431914 1005236 432276 1005242
rect 430856 1005178 430908 1005184
rect 431966 1005230 432276 1005236
rect 431914 1005178 431966 1005184
rect 432052 1005168 432104 1005174
rect 432050 1005136 432052 1005145
rect 432104 1005136 432106 1005145
rect 432248 1005122 432276 1005230
rect 432248 1005094 432460 1005122
rect 432050 1005071 432106 1005080
rect 432432 1005038 432460 1005094
rect 432420 1005032 432472 1005038
rect 432420 1004974 432472 1004980
rect 432236 1004964 432288 1004970
rect 432236 1004906 432288 1004912
rect 431682 1004864 431738 1004873
rect 431682 1004799 431684 1004808
rect 431736 1004799 431738 1004808
rect 431684 1004770 431736 1004776
rect 430026 1004728 430082 1004737
rect 430026 1004663 430028 1004672
rect 430080 1004663 430082 1004672
rect 431868 1004692 431920 1004698
rect 430028 1004634 430080 1004640
rect 431920 1004640 432092 1004654
rect 431868 1004634 432092 1004640
rect 431880 1004626 432092 1004634
rect 431132 1002244 431184 1002250
rect 431132 1002186 431184 1002192
rect 431144 997762 431172 1002186
rect 431316 1002108 431368 1002114
rect 431316 1002050 431368 1002056
rect 431328 998714 431356 1002050
rect 431316 998708 431368 998714
rect 431316 998650 431368 998656
rect 431132 997756 431184 997762
rect 431132 997698 431184 997704
rect 432064 995858 432092 1004626
rect 432248 995994 432276 1004906
rect 433338 1002144 433394 1002153
rect 433338 1002079 433340 1002088
rect 433392 1002079 433394 1002088
rect 433340 1002050 433392 1002056
rect 432878 1002008 432934 1002017
rect 432878 1001943 432880 1001952
rect 432932 1001943 432934 1001952
rect 432880 1001914 432932 1001920
rect 433536 996130 433564 1005790
rect 436928 1005440 436980 1005446
rect 436928 1005382 436980 1005388
rect 436940 1005174 436968 1005382
rect 436928 1005168 436980 1005174
rect 436928 1005110 436980 1005116
rect 434168 1005032 434220 1005038
rect 434168 1004974 434220 1004980
rect 433984 1004692 434036 1004698
rect 433984 1004634 434036 1004640
rect 433996 996130 434024 1004634
rect 433524 996124 433576 996130
rect 433524 996066 433576 996072
rect 433984 996124 434036 996130
rect 433984 996066 434036 996072
rect 434180 995994 434208 1004974
rect 435364 1002108 435416 1002114
rect 435364 1002050 435416 1002056
rect 432236 995988 432288 995994
rect 432236 995930 432288 995936
rect 434168 995988 434220 995994
rect 434168 995930 434220 995936
rect 432052 995852 432104 995858
rect 432052 995794 432104 995800
rect 429844 994968 429896 994974
rect 429844 994910 429896 994916
rect 426440 994288 426492 994294
rect 426440 994230 426492 994236
rect 435376 990418 435404 1002050
rect 436744 1001972 436796 1001978
rect 436744 1001914 436796 1001920
rect 435364 990412 435416 990418
rect 435364 990354 435416 990360
rect 422208 988916 422260 988922
rect 422208 988858 422260 988864
rect 436756 985998 436784 1001914
rect 438136 997626 438164 1006810
rect 439700 998345 439728 1006946
rect 503352 1006936 503404 1006942
rect 503350 1006904 503352 1006913
rect 503404 1006904 503406 1006913
rect 503350 1006839 503406 1006848
rect 506204 1006664 506256 1006670
rect 506202 1006632 506204 1006641
rect 506256 1006632 506258 1006641
rect 471244 1006596 471296 1006602
rect 506202 1006567 506258 1006576
rect 471244 1006538 471296 1006544
rect 443644 1006324 443696 1006330
rect 443644 1006266 443696 1006272
rect 439686 998336 439742 998345
rect 443656 998306 443684 1006266
rect 446404 1005712 446456 1005718
rect 446404 1005654 446456 1005660
rect 446416 999122 446444 1005654
rect 460204 1005576 460256 1005582
rect 460204 1005518 460256 1005524
rect 456064 1005304 456116 1005310
rect 456064 1005246 456116 1005252
rect 456076 1002862 456104 1005246
rect 456064 1002856 456116 1002862
rect 456064 1002798 456116 1002804
rect 449164 1002720 449216 1002726
rect 449164 1002662 449216 1002668
rect 446404 999116 446456 999122
rect 446404 999058 446456 999064
rect 439686 998271 439742 998280
rect 443644 998300 443696 998306
rect 443644 998242 443696 998248
rect 446864 998300 446916 998306
rect 446864 998242 446916 998248
rect 439688 997756 439740 997762
rect 439688 997698 439740 997704
rect 438124 997620 438176 997626
rect 438124 997562 438176 997568
rect 439700 996713 439728 997698
rect 439872 997620 439924 997626
rect 439872 997562 439924 997568
rect 439686 996704 439742 996713
rect 439686 996639 439742 996648
rect 439884 996441 439912 997562
rect 439870 996432 439926 996441
rect 439870 996367 439926 996376
rect 446876 994945 446904 998242
rect 449176 996169 449204 1002662
rect 458088 1002584 458140 1002590
rect 458088 1002526 458140 1002532
rect 458100 999190 458128 1002526
rect 458088 999184 458140 999190
rect 458088 999126 458140 999132
rect 452292 999116 452344 999122
rect 452292 999058 452344 999064
rect 449162 996160 449218 996169
rect 449162 996095 449218 996104
rect 446862 994936 446918 994945
rect 446862 994871 446918 994880
rect 452304 994673 452332 999058
rect 460216 994838 460244 1005518
rect 465724 1005440 465776 1005446
rect 465724 1005382 465776 1005388
rect 462320 1002856 462372 1002862
rect 462320 1002798 462372 1002804
rect 462332 995897 462360 1002798
rect 462318 995888 462374 995897
rect 462318 995823 462374 995832
rect 460204 994832 460256 994838
rect 460204 994774 460256 994780
rect 452290 994664 452346 994673
rect 452290 994599 452346 994608
rect 446128 994288 446180 994294
rect 446128 994230 446180 994236
rect 414112 985992 414164 985998
rect 414112 985934 414164 985940
rect 415032 985992 415084 985998
rect 415032 985934 415084 985940
rect 430304 985992 430356 985998
rect 430304 985934 430356 985940
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 414124 983620 414152 985934
rect 430316 983620 430344 985934
rect 446140 983634 446168 994230
rect 463608 990412 463660 990418
rect 463608 990354 463660 990360
rect 463620 986134 463648 990354
rect 463608 986128 463660 986134
rect 463608 986070 463660 986076
rect 465736 985998 465764 1005382
rect 469864 1003944 469916 1003950
rect 469864 1003886 469916 1003892
rect 466460 998844 466512 998850
rect 466460 998786 466512 998792
rect 466472 994401 466500 998786
rect 469876 994702 469904 1003886
rect 471256 995858 471284 1006538
rect 505376 1006528 505428 1006534
rect 505374 1006496 505376 1006505
rect 505428 1006496 505430 1006505
rect 505374 1006431 505430 1006440
rect 502154 1006360 502210 1006369
rect 502154 1006295 502156 1006304
rect 502208 1006295 502210 1006304
rect 502156 1006266 502208 1006272
rect 508226 1006224 508282 1006233
rect 508226 1006159 508228 1006168
rect 508280 1006159 508282 1006168
rect 508228 1006130 508280 1006136
rect 498842 1006088 498898 1006097
rect 471428 1006052 471480 1006058
rect 471428 1005994 471480 1006000
rect 497924 1006052 497976 1006058
rect 498842 1006023 498844 1006032
rect 497924 1005994 497976 1006000
rect 498896 1006023 498898 1006032
rect 501326 1006088 501382 1006097
rect 509054 1006088 509110 1006097
rect 501326 1006023 501328 1006032
rect 498844 1005994 498896 1006000
rect 501380 1006023 501382 1006032
rect 506480 1006052 506532 1006058
rect 501328 1005994 501380 1006000
rect 509054 1006023 509056 1006032
rect 506480 1005994 506532 1006000
rect 509108 1006023 509110 1006032
rect 509056 1005994 509108 1006000
rect 471244 995852 471296 995858
rect 471244 995794 471296 995800
rect 471440 995314 471468 1005994
rect 496728 1001972 496780 1001978
rect 496728 1001914 496780 1001920
rect 472624 998980 472676 998986
rect 472624 998922 472676 998928
rect 472440 998708 472492 998714
rect 472440 998650 472492 998656
rect 472072 998572 472124 998578
rect 472072 998514 472124 998520
rect 471428 995308 471480 995314
rect 471428 995250 471480 995256
rect 472084 995217 472112 998514
rect 472256 998436 472308 998442
rect 472256 998378 472308 998384
rect 472070 995208 472126 995217
rect 472268 995178 472296 998378
rect 472452 995450 472480 998650
rect 472636 995586 472664 998922
rect 488908 997824 488960 997830
rect 488908 997766 488960 997772
rect 493508 997824 493560 997830
rect 493508 997766 493560 997772
rect 488920 995761 488948 997766
rect 473358 995752 473414 995761
rect 475934 995752 475990 995761
rect 473414 995710 473662 995738
rect 473358 995687 473414 995696
rect 475934 995687 475990 995696
rect 476486 995752 476542 995761
rect 477038 995752 477094 995761
rect 476542 995710 476790 995738
rect 476486 995687 476542 995696
rect 485686 995752 485742 995761
rect 477094 995710 477342 995738
rect 485346 995710 485686 995738
rect 477038 995687 477094 995696
rect 485686 995687 485742 995696
rect 488906 995752 488962 995761
rect 488906 995687 488962 995696
rect 474016 995586 474306 995602
rect 472624 995580 472676 995586
rect 472624 995522 472676 995528
rect 474004 995580 474306 995586
rect 474056 995574 474306 995580
rect 474004 995522 474056 995528
rect 475948 995518 475976 995687
rect 493520 995586 493548 997766
rect 493508 995580 493560 995586
rect 493508 995522 493560 995528
rect 475936 995512 475988 995518
rect 474752 995450 474950 995466
rect 478788 995512 478840 995518
rect 475936 995454 475988 995460
rect 472440 995444 472492 995450
rect 472440 995386 472492 995392
rect 474740 995444 474950 995450
rect 474792 995438 474950 995444
rect 477696 995438 477986 995466
rect 478248 995438 478630 995466
rect 478788 995454 478840 995460
rect 480810 995480 480866 995489
rect 474740 995386 474792 995392
rect 477696 995178 477724 995438
rect 478248 995217 478276 995438
rect 478800 995217 478828 995454
rect 480866 995438 481114 995466
rect 481376 995438 481666 995466
rect 481836 995438 482310 995466
rect 480810 995415 480866 995424
rect 478234 995208 478290 995217
rect 472070 995143 472126 995152
rect 472256 995172 472308 995178
rect 472256 995114 472308 995120
rect 477684 995172 477736 995178
rect 478234 995143 478290 995152
rect 478786 995208 478842 995217
rect 478786 995143 478842 995152
rect 477684 995114 477736 995120
rect 475750 994936 475806 994945
rect 475750 994871 475806 994880
rect 469864 994696 469916 994702
rect 469864 994638 469916 994644
rect 466458 994392 466514 994401
rect 466458 994327 466514 994336
rect 475764 994129 475792 994871
rect 481376 994702 481404 995438
rect 481836 995228 481864 995438
rect 481560 995217 481864 995228
rect 481546 995208 481864 995217
rect 481602 995200 481864 995208
rect 481546 995143 481602 995152
rect 481364 994696 481416 994702
rect 481364 994638 481416 994644
rect 482940 994401 482968 995452
rect 484136 994673 484164 995452
rect 485976 994838 486004 995452
rect 486620 994838 486648 995452
rect 487816 994945 487844 995452
rect 489736 995240 489788 995246
rect 489736 995182 489788 995188
rect 487802 994936 487858 994945
rect 487802 994871 487858 994880
rect 489748 994838 489776 995182
rect 485964 994832 486016 994838
rect 485964 994774 486016 994780
rect 486608 994832 486660 994838
rect 486608 994774 486660 994780
rect 489736 994832 489788 994838
rect 489736 994774 489788 994780
rect 484122 994664 484178 994673
rect 484122 994599 484178 994608
rect 482926 994392 482982 994401
rect 482926 994327 482982 994336
rect 475750 994120 475806 994129
rect 475750 994055 475806 994064
rect 496740 993342 496768 1001914
rect 497936 994498 497964 1005994
rect 499670 1004864 499726 1004873
rect 498108 1004828 498160 1004834
rect 499670 1004799 499672 1004808
rect 498108 1004770 498160 1004776
rect 499724 1004799 499726 1004808
rect 499672 1004770 499724 1004776
rect 497924 994492 497976 994498
rect 497924 994434 497976 994440
rect 496728 993336 496780 993342
rect 496728 993278 496780 993284
rect 498120 990418 498148 1004770
rect 500498 1004728 500554 1004737
rect 499488 1004692 499540 1004698
rect 500498 1004663 500500 1004672
rect 499488 1004634 499540 1004640
rect 500552 1004663 500554 1004672
rect 500500 1004634 500552 1004640
rect 498474 1002008 498530 1002017
rect 498474 1001943 498476 1001952
rect 498528 1001943 498530 1001952
rect 498476 1001914 498528 1001920
rect 499500 998714 499528 1004634
rect 504548 1004488 504600 1004494
rect 504546 1004456 504548 1004465
rect 504600 1004456 504602 1004465
rect 504546 1004391 504602 1004400
rect 501694 1002552 501750 1002561
rect 501694 1002487 501696 1002496
rect 501748 1002487 501750 1002496
rect 504364 1002516 504416 1002522
rect 501696 1002458 501748 1002464
rect 504364 1002458 504416 1002464
rect 502154 1002416 502210 1002425
rect 500224 1002380 500276 1002386
rect 502154 1002351 502156 1002360
rect 500224 1002322 500276 1002328
rect 502208 1002351 502210 1002360
rect 502156 1002322 502208 1002328
rect 499488 998708 499540 998714
rect 499488 998650 499540 998656
rect 500236 998442 500264 1002322
rect 500498 1002280 500554 1002289
rect 500498 1002215 500500 1002224
rect 500552 1002215 500554 1002224
rect 502984 1002244 503036 1002250
rect 500500 1002186 500552 1002192
rect 502984 1002186 503036 1002192
rect 502522 1002144 502578 1002153
rect 500684 1002108 500736 1002114
rect 502522 1002079 502524 1002088
rect 500684 1002050 500736 1002056
rect 502576 1002079 502578 1002088
rect 502524 1002050 502576 1002056
rect 500224 998436 500276 998442
rect 500224 998378 500276 998384
rect 500696 995042 500724 1002050
rect 502248 1001972 502300 1001978
rect 502248 1001914 502300 1001920
rect 500684 995036 500736 995042
rect 500684 994978 500736 994984
rect 502260 994634 502288 1001914
rect 502996 994770 503024 1002186
rect 503350 1002008 503406 1002017
rect 503350 1001943 503352 1001952
rect 503404 1001943 503406 1001952
rect 504178 1002008 504234 1002017
rect 504178 1001943 504180 1001952
rect 503352 1001914 503404 1001920
rect 504232 1001943 504234 1001952
rect 504180 1001914 504232 1001920
rect 504376 998850 504404 1002458
rect 506202 1002008 506258 1002017
rect 505744 1001972 505796 1001978
rect 506202 1001943 506204 1001952
rect 505744 1001914 505796 1001920
rect 506256 1001943 506258 1001952
rect 506204 1001914 506256 1001920
rect 504364 998844 504416 998850
rect 504364 998786 504416 998792
rect 505756 995314 505784 1001914
rect 506492 998578 506520 1005994
rect 507030 1005272 507086 1005281
rect 507030 1005207 507032 1005216
rect 507084 1005207 507086 1005216
rect 509976 1005236 510028 1005242
rect 507032 1005178 507084 1005184
rect 509976 1005178 510028 1005184
rect 508226 1005136 508282 1005145
rect 508226 1005071 508228 1005080
rect 508280 1005071 508282 1005080
rect 508228 1005042 508280 1005048
rect 507858 1005000 507914 1005009
rect 507858 1004935 507860 1004944
rect 507912 1004935 507914 1004944
rect 509700 1004964 509752 1004970
rect 507860 1004906 507912 1004912
rect 509700 1004906 509752 1004912
rect 507398 1004864 507454 1004873
rect 507398 1004799 507400 1004808
rect 507452 1004799 507454 1004808
rect 509240 1004828 509292 1004834
rect 507400 1004770 507452 1004776
rect 509240 1004770 509292 1004776
rect 509054 1004728 509110 1004737
rect 509054 1004663 509056 1004672
rect 509108 1004663 509110 1004672
rect 509056 1004634 509108 1004640
rect 507860 1001972 507912 1001978
rect 507860 1001914 507912 1001920
rect 506480 998572 506532 998578
rect 506480 998514 506532 998520
rect 507872 995858 507900 1001914
rect 507860 995852 507912 995858
rect 507860 995794 507912 995800
rect 509252 995450 509280 1004770
rect 509712 995858 509740 1004906
rect 509988 1004306 510016 1005178
rect 510896 1005100 510948 1005106
rect 510896 1005042 510948 1005048
rect 510712 1004692 510764 1004698
rect 510712 1004634 510764 1004640
rect 510160 1004488 510212 1004494
rect 510160 1004430 510212 1004436
rect 509988 1004278 510108 1004306
rect 509882 1002280 509938 1002289
rect 509882 1002215 509884 1002224
rect 509936 1002215 509938 1002224
rect 509884 1002186 509936 1002192
rect 510080 1001894 510108 1004278
rect 509896 1001866 510108 1001894
rect 509700 995852 509752 995858
rect 509700 995794 509752 995800
rect 509896 995450 509924 1001866
rect 510172 1000958 510200 1004430
rect 510342 1002144 510398 1002153
rect 510342 1002079 510344 1002088
rect 510396 1002079 510398 1002088
rect 510344 1002050 510396 1002056
rect 510160 1000952 510212 1000958
rect 510160 1000894 510212 1000900
rect 510068 998708 510120 998714
rect 510068 998650 510120 998656
rect 510080 998306 510108 998650
rect 510068 998300 510120 998306
rect 510068 998242 510120 998248
rect 510724 996130 510752 1004634
rect 510712 996124 510764 996130
rect 510712 996066 510764 996072
rect 510908 995994 510936 1005042
rect 512644 1002244 512696 1002250
rect 512644 1002186 512696 1002192
rect 510896 995988 510948 995994
rect 510896 995930 510948 995936
rect 511080 995580 511132 995586
rect 511080 995522 511132 995528
rect 509240 995444 509292 995450
rect 509240 995386 509292 995392
rect 509884 995444 509936 995450
rect 509884 995386 509936 995392
rect 505744 995308 505796 995314
rect 505744 995250 505796 995256
rect 502984 994764 503036 994770
rect 502984 994706 503036 994712
rect 502248 994628 502300 994634
rect 502248 994570 502300 994576
rect 498108 990412 498160 990418
rect 498108 990354 498160 990360
rect 478972 986128 479024 986134
rect 478972 986070 479024 986076
rect 462780 985992 462832 985998
rect 462780 985934 462832 985940
rect 465724 985992 465776 985998
rect 465724 985934 465776 985940
rect 446140 983606 446522 983634
rect 462792 983620 462820 985934
rect 478984 983620 479012 986070
rect 495164 985992 495216 985998
rect 495164 985934 495216 985940
rect 495176 983620 495204 985934
rect 511092 983634 511120 995522
rect 512656 991914 512684 1002186
rect 512828 1002108 512880 1002114
rect 512828 1002050 512880 1002056
rect 512840 1001434 512868 1002050
rect 512828 1001428 512880 1001434
rect 512828 1001370 512880 1001376
rect 513852 998986 513880 1007150
rect 515588 1007072 515640 1007078
rect 515588 1007014 515640 1007020
rect 551098 1007040 551154 1007049
rect 514024 1006664 514076 1006670
rect 514024 1006606 514076 1006612
rect 514036 1006058 514064 1006606
rect 514024 1006052 514076 1006058
rect 514024 1005994 514076 1006000
rect 515404 1005916 515456 1005922
rect 515404 1005858 515456 1005864
rect 513840 998980 513892 998986
rect 513840 998922 513892 998928
rect 512644 991908 512696 991914
rect 512644 991850 512696 991856
rect 515416 985998 515444 1005858
rect 515600 997762 515628 1007014
rect 520924 1007004 520976 1007010
rect 551098 1006975 551100 1006984
rect 520924 1006946 520976 1006952
rect 551152 1006975 551154 1006984
rect 569224 1007004 569276 1007010
rect 551100 1006946 551152 1006952
rect 569224 1006946 569276 1006952
rect 516784 1006528 516836 1006534
rect 516784 1006470 516836 1006476
rect 516796 999122 516824 1006470
rect 518164 1006324 518216 1006330
rect 518164 1006266 518216 1006272
rect 517244 1000952 517296 1000958
rect 517244 1000894 517296 1000900
rect 516784 999116 516836 999122
rect 516784 999058 516836 999064
rect 516692 998844 516744 998850
rect 516692 998786 516744 998792
rect 515588 997756 515640 997762
rect 515588 997698 515640 997704
rect 516704 996169 516732 998786
rect 517256 998617 517284 1000894
rect 517242 998608 517298 998617
rect 517242 998543 517298 998552
rect 516876 997756 516928 997762
rect 516876 997698 516928 997704
rect 516888 996441 516916 997698
rect 516874 996432 516930 996441
rect 516874 996367 516930 996376
rect 516690 996160 516746 996169
rect 516690 996095 516746 996104
rect 518176 994809 518204 1006266
rect 519544 1001428 519596 1001434
rect 519544 1001370 519596 1001376
rect 518162 994800 518218 994809
rect 518162 994735 518218 994744
rect 519556 986134 519584 1001370
rect 520556 998300 520608 998306
rect 520556 998242 520608 998248
rect 520568 994906 520596 998242
rect 520936 997830 520964 1006946
rect 559654 1006904 559710 1006913
rect 554136 1006868 554188 1006874
rect 559654 1006839 559656 1006848
rect 554136 1006810 554188 1006816
rect 559708 1006839 559710 1006848
rect 559656 1006810 559708 1006816
rect 553122 1006496 553178 1006505
rect 553122 1006431 553124 1006440
rect 553176 1006431 553178 1006440
rect 553124 1006402 553176 1006408
rect 522304 1006188 522356 1006194
rect 522304 1006130 522356 1006136
rect 520924 997824 520976 997830
rect 520924 997766 520976 997772
rect 522316 995994 522344 1006130
rect 522488 1006052 522540 1006058
rect 522488 1005994 522540 1006000
rect 522500 996130 522528 1005994
rect 553952 1005440 554004 1005446
rect 553950 1005408 553952 1005417
rect 554004 1005408 554006 1005417
rect 553950 1005343 554006 1005352
rect 552296 1005304 552348 1005310
rect 552294 1005272 552296 1005281
rect 552348 1005272 552350 1005281
rect 552294 1005207 552350 1005216
rect 553124 1002244 553176 1002250
rect 553124 1002186 553176 1002192
rect 523316 999116 523368 999122
rect 523316 999058 523368 999064
rect 523132 998436 523184 998442
rect 523132 998378 523184 998384
rect 522488 996124 522540 996130
rect 522488 996066 522540 996072
rect 522304 995988 522356 995994
rect 522304 995930 522356 995936
rect 523144 995217 523172 998378
rect 523130 995208 523186 995217
rect 523328 995178 523356 999058
rect 523684 998980 523736 998986
rect 523684 998922 523736 998928
rect 523498 998608 523554 998617
rect 523498 998543 523554 998552
rect 523512 995489 523540 998543
rect 523696 995761 523724 998922
rect 524052 998572 524104 998578
rect 524052 998514 524104 998520
rect 523868 997824 523920 997830
rect 523868 997766 523920 997772
rect 523682 995752 523738 995761
rect 523682 995687 523738 995696
rect 523880 995586 523908 997766
rect 524064 996713 524092 998514
rect 551098 998064 551154 998073
rect 549168 998028 549220 998034
rect 551098 997999 551100 998008
rect 549168 997970 549220 997976
rect 551152 997999 551154 998008
rect 551100 997970 551152 997976
rect 547788 997892 547840 997898
rect 547788 997834 547840 997840
rect 524050 996704 524106 996713
rect 524050 996639 524106 996648
rect 524786 995752 524842 995761
rect 529846 995752 529902 995761
rect 524842 995710 525090 995738
rect 524786 995687 524842 995696
rect 536562 995752 536618 995761
rect 529902 995710 530058 995738
rect 529846 995687 529902 995696
rect 537206 995752 537262 995761
rect 536618 995710 536774 995738
rect 536562 995687 536618 995696
rect 537262 995710 537418 995738
rect 537206 995687 537262 995696
rect 525352 995586 525734 995602
rect 523868 995580 523920 995586
rect 523868 995522 523920 995528
rect 525340 995580 525734 995586
rect 525392 995574 525734 995580
rect 525340 995522 525392 995528
rect 523498 995480 523554 995489
rect 527914 995480 527970 995489
rect 523498 995415 523554 995424
rect 526088 995438 526378 995466
rect 526088 995178 526116 995438
rect 533434 995480 533490 995489
rect 527970 995438 528218 995466
rect 527914 995415 527970 995424
rect 526258 995208 526314 995217
rect 523130 995143 523186 995152
rect 523316 995172 523368 995178
rect 523316 995114 523368 995120
rect 526076 995172 526128 995178
rect 526258 995143 526260 995152
rect 526076 995114 526128 995120
rect 526312 995143 526314 995152
rect 526260 995114 526312 995120
rect 528756 995042 528784 995452
rect 529032 995438 529414 995466
rect 532160 995438 532542 995466
rect 529032 995178 529060 995438
rect 532160 995314 532188 995438
rect 532148 995308 532200 995314
rect 532148 995250 532200 995256
rect 529020 995172 529072 995178
rect 529020 995114 529072 995120
rect 528744 995036 528796 995042
rect 528744 994978 528796 994984
rect 533080 994974 533108 995452
rect 537850 995480 537906 995489
rect 533490 995438 533738 995466
rect 534092 995438 534382 995466
rect 533434 995415 533490 995424
rect 534092 995110 534120 995438
rect 534080 995104 534132 995110
rect 534080 995046 534132 995052
rect 533068 994968 533120 994974
rect 533068 994910 533120 994916
rect 520556 994900 520608 994906
rect 520556 994842 520608 994848
rect 535564 994809 535592 995452
rect 538218 995480 538274 995489
rect 537850 995415 537906 995424
rect 537864 994974 537892 995415
rect 537852 994968 537904 994974
rect 537852 994910 537904 994916
rect 535550 994800 535606 994809
rect 535550 994735 535606 994744
rect 538048 994498 538076 995452
rect 538218 995415 538274 995424
rect 538232 994770 538260 995415
rect 538220 994764 538272 994770
rect 538220 994706 538272 994712
rect 539244 994634 539272 995452
rect 539232 994628 539284 994634
rect 539232 994570 539284 994576
rect 538036 994492 538088 994498
rect 538036 994434 538088 994440
rect 547800 994294 547828 997834
rect 549180 994430 549208 997970
rect 550270 997928 550326 997937
rect 550270 997863 550272 997872
rect 550324 997863 550326 997872
rect 550548 997892 550600 997898
rect 550272 997834 550324 997840
rect 550548 997834 550600 997840
rect 550560 997754 550588 997834
rect 551466 997792 551522 997801
rect 550376 997726 550588 997754
rect 550652 997736 551466 997754
rect 552294 997792 552350 997801
rect 550652 997727 551522 997736
rect 551940 997750 552294 997778
rect 550652 997726 551508 997727
rect 550376 994906 550404 997726
rect 550652 995042 550680 997726
rect 551940 996266 551968 997750
rect 552294 997727 552350 997736
rect 553136 997422 553164 1002186
rect 553306 997928 553362 997937
rect 553306 997863 553308 997872
rect 553360 997863 553362 997872
rect 553308 997834 553360 997840
rect 553124 997416 553176 997422
rect 553124 997358 553176 997364
rect 551928 996260 551980 996266
rect 551928 996202 551980 996208
rect 554148 995858 554176 1006810
rect 555974 1006768 556030 1006777
rect 555974 1006703 555976 1006712
rect 556028 1006703 556030 1006712
rect 566464 1006732 566516 1006738
rect 555976 1006674 556028 1006680
rect 566464 1006674 566516 1006680
rect 556802 1006360 556858 1006369
rect 556802 1006295 556804 1006304
rect 556856 1006295 556858 1006304
rect 560208 1006324 560260 1006330
rect 556804 1006266 556856 1006272
rect 560208 1006266 560260 1006272
rect 557170 1006224 557226 1006233
rect 557170 1006159 557172 1006168
rect 557224 1006159 557226 1006168
rect 557172 1006130 557224 1006136
rect 555148 1005576 555200 1005582
rect 555146 1005544 555148 1005553
rect 555200 1005544 555202 1005553
rect 555146 1005479 555202 1005488
rect 555974 1004864 556030 1004873
rect 555974 1004799 555976 1004808
rect 556028 1004799 556030 1004808
rect 558184 1004828 558236 1004834
rect 555976 1004770 556028 1004776
rect 558184 1004770 558236 1004776
rect 557630 1004728 557686 1004737
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 557632 1004634 557684 1004640
rect 557998 1002416 558054 1002425
rect 557998 1002351 558000 1002360
rect 558052 1002351 558054 1002360
rect 558000 1002322 558052 1002328
rect 554318 1002280 554374 1002289
rect 554318 1002215 554320 1002224
rect 554372 1002215 554374 1002224
rect 554320 1002186 554372 1002192
rect 555146 1002144 555202 1002153
rect 557998 1002144 558054 1002153
rect 555146 1002079 555148 1002088
rect 555200 1002079 555202 1002088
rect 556804 1002108 556856 1002114
rect 555148 1002050 555200 1002056
rect 557998 1002079 558000 1002088
rect 556804 1002050 556856 1002056
rect 558052 1002079 558054 1002088
rect 558000 1002050 558052 1002056
rect 554318 1002008 554374 1002017
rect 554318 1001943 554320 1001952
rect 554372 1001943 554374 1001952
rect 555424 1001972 555476 1001978
rect 554320 1001914 554372 1001920
rect 555424 1001914 555476 1001920
rect 555436 996334 555464 1001914
rect 555424 996328 555476 996334
rect 555424 996270 555476 996276
rect 554320 996260 554372 996266
rect 554320 996202 554372 996208
rect 554332 995858 554360 996202
rect 554136 995852 554188 995858
rect 554136 995794 554188 995800
rect 554320 995852 554372 995858
rect 554320 995794 554372 995800
rect 556816 995178 556844 1002050
rect 558196 997082 558224 1004770
rect 559564 1004692 559616 1004698
rect 559564 1004634 559616 1004640
rect 558826 1002552 558882 1002561
rect 558826 1002487 558828 1002496
rect 558880 1002487 558882 1002496
rect 558828 1002458 558880 1002464
rect 558826 1002008 558882 1002017
rect 558826 1001943 558828 1001952
rect 558880 1001943 558882 1001952
rect 558828 1001914 558880 1001920
rect 558184 997076 558236 997082
rect 558184 997018 558236 997024
rect 556804 995172 556856 995178
rect 556804 995114 556856 995120
rect 550640 995036 550692 995042
rect 550640 994978 550692 994984
rect 550364 994900 550416 994906
rect 550364 994842 550416 994848
rect 549168 994424 549220 994430
rect 549168 994366 549220 994372
rect 547788 994288 547840 994294
rect 547788 994230 547840 994236
rect 527640 991908 527692 991914
rect 527640 991850 527692 991856
rect 519544 986128 519596 986134
rect 519544 986070 519596 986076
rect 515404 985992 515456 985998
rect 515404 985934 515456 985940
rect 511092 983606 511474 983634
rect 527652 983620 527680 991850
rect 559576 987698 559604 1004634
rect 560220 1002658 560248 1006266
rect 560852 1005712 560904 1005718
rect 560850 1005680 560852 1005689
rect 560904 1005680 560906 1005689
rect 560850 1005615 560906 1005624
rect 560208 1002652 560260 1002658
rect 560208 1002594 560260 1002600
rect 562324 1002516 562376 1002522
rect 562324 1002458 562376 1002464
rect 560482 1002416 560538 1002425
rect 560300 1002380 560352 1002386
rect 560482 1002351 560484 1002360
rect 560300 1002322 560352 1002328
rect 560536 1002351 560538 1002360
rect 560484 1002322 560536 1002328
rect 560022 1002280 560078 1002289
rect 560022 1002215 560024 1002224
rect 560076 1002215 560078 1002224
rect 560024 1002186 560076 1002192
rect 560312 1002130 560340 1002322
rect 560850 1002144 560906 1002153
rect 560312 1002102 560524 1002130
rect 560496 1001994 560524 1002102
rect 560668 1002108 560720 1002114
rect 560850 1002079 560852 1002088
rect 560668 1002050 560720 1002056
rect 560904 1002079 560906 1002088
rect 560852 1002050 560904 1002056
rect 560208 1001972 560260 1001978
rect 560496 1001966 560616 1001994
rect 560208 1001914 560260 1001920
rect 560220 1001858 560248 1001914
rect 560220 1001830 560340 1001858
rect 560312 995450 560340 1001830
rect 560588 996130 560616 1001966
rect 560680 1001894 560708 1002050
rect 561678 1002008 561734 1002017
rect 561678 1001943 561680 1001952
rect 561732 1001943 561734 1001952
rect 561680 1001914 561732 1001920
rect 560680 1001866 560984 1001894
rect 560576 996124 560628 996130
rect 560576 996066 560628 996072
rect 560300 995444 560352 995450
rect 560300 995386 560352 995392
rect 559564 987692 559616 987698
rect 559564 987634 559616 987640
rect 543832 986128 543884 986134
rect 543832 986070 543884 986076
rect 543844 983620 543872 986070
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 560128 983620 560156 985934
rect 560956 984910 560984 1001866
rect 562336 985998 562364 1002458
rect 563060 1002380 563112 1002386
rect 563060 1002322 563112 1002328
rect 562508 1002244 562560 1002250
rect 562508 1002186 562560 1002192
rect 562520 990554 562548 1002186
rect 563072 995994 563100 1002322
rect 563704 1002108 563756 1002114
rect 563704 1002050 563756 1002056
rect 563060 995988 563112 995994
rect 563060 995930 563112 995936
rect 563716 994566 563744 1002050
rect 565084 1001972 565136 1001978
rect 565084 1001914 565136 1001920
rect 563704 994560 563756 994566
rect 563704 994502 563756 994508
rect 562508 990548 562560 990554
rect 562508 990490 562560 990496
rect 565096 986134 565124 1001914
rect 566476 997694 566504 1006674
rect 567844 1005576 567896 1005582
rect 567844 1005518 567896 1005524
rect 567200 1002652 567252 1002658
rect 567200 1002594 567252 1002600
rect 566464 997688 566516 997694
rect 566464 997630 566516 997636
rect 567212 995314 567240 1002594
rect 567200 995308 567252 995314
rect 567200 995250 567252 995256
rect 567856 993721 567884 1005518
rect 569236 997218 569264 1006946
rect 571984 1006324 572036 1006330
rect 571984 1006266 572036 1006272
rect 570604 1005712 570656 1005718
rect 570604 1005654 570656 1005660
rect 569224 997212 569276 997218
rect 569224 997154 569276 997160
rect 567842 993712 567898 993721
rect 567842 993647 567898 993656
rect 570616 986270 570644 1005654
rect 570788 1005304 570840 1005310
rect 570788 1005246 570840 1005252
rect 570800 996946 570828 1005246
rect 570788 996940 570840 996946
rect 570788 996882 570840 996888
rect 571996 994770 572024 1006266
rect 574744 1006052 574796 1006058
rect 574744 1005994 574796 1006000
rect 573364 1005440 573416 1005446
rect 573364 1005382 573416 1005388
rect 573376 997558 573404 1005382
rect 573364 997552 573416 997558
rect 573364 997494 573416 997500
rect 574756 996810 574784 1005994
rect 591304 999320 591356 999326
rect 591304 999262 591356 999268
rect 616788 999320 616840 999326
rect 616788 999262 616840 999268
rect 591120 999184 591172 999190
rect 591120 999126 591172 999132
rect 581828 997552 581880 997558
rect 581472 997500 581828 997506
rect 581472 997494 581880 997500
rect 581472 997478 581868 997494
rect 581276 997416 581328 997422
rect 581276 997358 581328 997364
rect 574744 996804 574796 996810
rect 574744 996746 574796 996752
rect 581288 996674 581316 997358
rect 581472 996946 581500 997478
rect 590384 997416 590436 997422
rect 590384 997358 590436 997364
rect 581460 996940 581512 996946
rect 581460 996882 581512 996888
rect 581276 996668 581328 996674
rect 581276 996610 581328 996616
rect 590396 996418 590424 997358
rect 590566 996704 590622 996713
rect 590566 996639 590568 996648
rect 590620 996639 590622 996648
rect 590568 996610 590620 996616
rect 590566 996432 590622 996441
rect 590396 996390 590566 996418
rect 590566 996367 590622 996376
rect 591132 996334 591160 999126
rect 591316 997558 591344 999262
rect 616800 998442 616828 999262
rect 625620 999184 625672 999190
rect 625620 999126 625672 999132
rect 616788 998436 616840 998442
rect 616788 998378 616840 998384
rect 625436 998436 625488 998442
rect 625436 998378 625488 998384
rect 592040 997824 592092 997830
rect 592040 997766 592092 997772
rect 591304 997552 591356 997558
rect 591304 997494 591356 997500
rect 592052 996946 592080 997766
rect 623688 997688 623740 997694
rect 623688 997630 623740 997636
rect 620284 997212 620336 997218
rect 620284 997154 620336 997160
rect 617340 997076 617392 997082
rect 617340 997018 617392 997024
rect 592040 996940 592092 996946
rect 592040 996882 592092 996888
rect 591120 996328 591172 996334
rect 591120 996270 591172 996276
rect 617352 995081 617380 997018
rect 620296 995450 620324 997154
rect 623700 995761 623728 997630
rect 625448 996033 625476 998378
rect 625434 996024 625490 996033
rect 625434 995959 625490 995968
rect 625436 995852 625488 995858
rect 625436 995794 625488 995800
rect 623686 995752 623742 995761
rect 623686 995687 623742 995696
rect 620284 995444 620336 995450
rect 620284 995386 620336 995392
rect 617338 995072 617394 995081
rect 617338 995007 617394 995016
rect 625448 994809 625476 995794
rect 625632 995489 625660 999126
rect 625804 997824 625856 997830
rect 625804 997766 625856 997772
rect 625816 995586 625844 997766
rect 626538 995752 626594 995761
rect 627182 995752 627238 995761
rect 626594 995710 626888 995738
rect 626538 995687 626594 995696
rect 631506 995752 631562 995761
rect 627238 995710 627532 995738
rect 627182 995687 627238 995696
rect 631562 995710 631856 995738
rect 631506 995687 631562 995696
rect 627932 995586 628176 995602
rect 625804 995580 625856 995586
rect 625804 995522 625856 995528
rect 627920 995580 628176 995586
rect 627972 995574 628176 995580
rect 627920 995522 627972 995528
rect 625618 995480 625674 995489
rect 630218 995480 630274 995489
rect 625618 995415 625674 995424
rect 629680 995438 630016 995466
rect 629680 995081 629708 995438
rect 630862 995480 630918 995489
rect 630274 995438 630568 995466
rect 630218 995415 630274 995424
rect 630918 995438 631212 995466
rect 634004 995438 634340 995466
rect 634740 995438 634892 995466
rect 635200 995438 635536 995466
rect 635844 995438 636180 995466
rect 637040 995438 637376 995466
rect 638512 995438 638572 995466
rect 638972 995438 639216 995466
rect 639524 995438 639860 995466
rect 640720 995438 641056 995466
rect 630862 995415 630918 995424
rect 630600 995314 630812 995330
rect 630588 995308 630812 995314
rect 630640 995302 630812 995308
rect 630588 995250 630640 995256
rect 629666 995072 629722 995081
rect 629666 995007 629722 995016
rect 630784 994906 630812 995302
rect 625804 994900 625856 994906
rect 625804 994842 625856 994848
rect 630772 994900 630824 994906
rect 630772 994842 630824 994848
rect 625434 994800 625490 994809
rect 571984 994764 572036 994770
rect 625434 994735 625490 994744
rect 571984 994706 572036 994712
rect 625816 994634 625844 994842
rect 625804 994628 625856 994634
rect 625804 994570 625856 994576
rect 624608 994560 624660 994566
rect 624608 994502 624660 994508
rect 576306 989496 576362 989505
rect 576306 989431 576362 989440
rect 570604 986264 570656 986270
rect 570604 986206 570656 986212
rect 565084 986128 565136 986134
rect 565084 986070 565136 986076
rect 562324 985992 562376 985998
rect 562324 985934 562376 985940
rect 560944 984904 560996 984910
rect 560944 984846 560996 984852
rect 576320 983620 576348 989431
rect 592500 986264 592552 986270
rect 592500 986206 592552 986212
rect 592512 983620 592540 986206
rect 608784 986128 608836 986134
rect 608784 986070 608836 986076
rect 608796 983620 608824 986070
rect 624620 983634 624648 994502
rect 634004 993721 634032 995438
rect 634740 994809 634768 995438
rect 634726 994800 634782 994809
rect 635200 994770 635228 995438
rect 635844 995042 635872 995438
rect 635832 995036 635884 995042
rect 635832 994978 635884 994984
rect 634726 994735 634782 994744
rect 635188 994764 635240 994770
rect 635188 994706 635240 994712
rect 637040 994634 637068 995438
rect 638512 994906 638540 995438
rect 638972 995058 639000 995438
rect 639524 995382 639552 995438
rect 639512 995376 639564 995382
rect 639512 995318 639564 995324
rect 640720 995178 640748 995438
rect 640708 995172 640760 995178
rect 640708 995114 640760 995120
rect 638696 995042 639000 995058
rect 638684 995036 639000 995042
rect 638736 995030 639000 995036
rect 638684 994978 638736 994984
rect 640800 994968 640852 994974
rect 640800 994910 640852 994916
rect 638500 994900 638552 994906
rect 638500 994842 638552 994848
rect 637028 994628 637080 994634
rect 637028 994570 637080 994576
rect 633990 993712 634046 993721
rect 633990 993647 634046 993656
rect 640812 983634 640840 994910
rect 667112 994424 667164 994430
rect 667112 994366 667164 994372
rect 666560 994288 666612 994294
rect 666560 994230 666612 994236
rect 665180 993200 665232 993206
rect 665180 993142 665232 993148
rect 650000 993064 650052 993070
rect 650000 993006 650052 993012
rect 648896 990140 648948 990146
rect 648896 990082 648948 990088
rect 624620 983606 625002 983634
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 55864 975724 55916 975730
rect 55864 975666 55916 975672
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 55876 969474 55904 975666
rect 55864 969468 55916 969474
rect 55864 969410 55916 969416
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 51724 939820 51776 939826
rect 51724 939762 51776 939768
rect 62120 937032 62172 937038
rect 62118 937000 62120 937009
rect 62172 937000 62174 937009
rect 62118 936935 62174 936944
rect 44822 936184 44878 936193
rect 44822 936119 44878 936128
rect 44454 934144 44510 934153
rect 44454 934079 44510 934088
rect 44178 933736 44234 933745
rect 44178 933671 44234 933680
rect 43442 933328 43498 933337
rect 43442 933263 43498 933272
rect 43456 932958 43484 933263
rect 43444 932952 43496 932958
rect 42522 932920 42578 932929
rect 43444 932894 43496 932900
rect 54484 932952 54536 932958
rect 54484 932894 54536 932900
rect 42522 932855 42578 932864
rect 42798 932104 42854 932113
rect 42798 932039 42854 932048
rect 42812 931598 42840 932039
rect 42800 931592 42852 931598
rect 42800 931534 42852 931540
rect 53104 931592 53156 931598
rect 53104 931534 53156 931540
rect 47584 923296 47636 923302
rect 47584 923238 47636 923244
rect 46204 897048 46256 897054
rect 46204 896990 46256 896996
rect 42432 884740 42484 884746
rect 42432 884682 42484 884688
rect 42444 881929 42472 884682
rect 42430 881920 42486 881929
rect 42430 881855 42486 881864
rect 43444 870868 43496 870874
rect 43444 870810 43496 870816
rect 41984 823846 42104 823874
rect 41984 821114 42012 823846
rect 41984 821086 42104 821114
rect 42076 818009 42104 821086
rect 42062 818000 42118 818009
rect 42062 817935 42118 817944
rect 41708 815930 41920 815946
rect 41696 815924 41920 815930
rect 41748 815918 41920 815924
rect 41696 815866 41748 815872
rect 41708 815658 42196 815674
rect 41696 815652 42208 815658
rect 41748 815646 42156 815652
rect 41696 815594 41748 815600
rect 42156 815594 42208 815600
rect 41696 814768 41748 814774
rect 41748 814745 41920 814756
rect 41748 814736 41934 814745
rect 41748 814728 41878 814736
rect 41696 814710 41748 814716
rect 41878 814671 41934 814680
rect 42890 814736 42946 814745
rect 42890 814671 42946 814680
rect 41708 814298 42104 814314
rect 41696 814292 42116 814298
rect 41748 814286 42064 814292
rect 41696 814234 41748 814240
rect 42064 814234 42116 814240
rect 41512 813000 41564 813006
rect 41512 812942 41564 812948
rect 41786 812832 41842 812841
rect 41340 812790 41786 812818
rect 41142 812767 41198 812776
rect 41786 812767 41842 812776
rect 35162 812424 35218 812433
rect 35162 812359 35218 812368
rect 32402 811200 32458 811209
rect 32402 811135 32458 811144
rect 31666 809976 31722 809985
rect 31666 809911 31722 809920
rect 31680 802330 31708 809911
rect 32416 802602 32444 811135
rect 33782 809568 33838 809577
rect 33782 809503 33838 809512
rect 32404 802596 32456 802602
rect 32404 802538 32456 802544
rect 31668 802324 31720 802330
rect 31668 802266 31720 802272
rect 33796 800970 33824 809503
rect 35176 803865 35204 812359
rect 40958 812016 41014 812025
rect 40958 811951 41014 811960
rect 36542 809160 36598 809169
rect 36542 809095 36598 809104
rect 35162 803856 35218 803865
rect 35162 803791 35218 803800
rect 36556 801786 36584 809095
rect 40972 804817 41000 811951
rect 41156 811454 41184 812767
rect 41328 811640 41380 811646
rect 41326 811608 41328 811617
rect 41696 811640 41748 811646
rect 41380 811608 41382 811617
rect 41748 811588 42288 811594
rect 41696 811582 42288 811588
rect 41708 811566 42288 811582
rect 41326 811543 41382 811552
rect 42260 811454 42288 811566
rect 41156 811426 41276 811454
rect 42260 811426 42380 811454
rect 40958 804808 41014 804817
rect 40958 804743 41014 804752
rect 39764 802324 39816 802330
rect 39764 802266 39816 802272
rect 39776 801961 39804 802266
rect 39762 801952 39818 801961
rect 39762 801887 39818 801896
rect 36544 801780 36596 801786
rect 36544 801722 36596 801728
rect 39856 801780 39908 801786
rect 39856 801722 39908 801728
rect 39868 801009 39896 801722
rect 39854 801000 39910 801009
rect 33784 800964 33836 800970
rect 39854 800935 39910 800944
rect 40040 800964 40092 800970
rect 33784 800906 33836 800912
rect 40040 800906 40092 800912
rect 40052 800737 40080 800906
rect 41248 800873 41276 811426
rect 41970 810384 42026 810393
rect 41970 810319 42026 810328
rect 41984 806834 42012 810319
rect 41800 806806 42012 806834
rect 41800 805361 41828 806806
rect 42062 806712 42118 806721
rect 42062 806647 42118 806656
rect 41786 805352 41842 805361
rect 41786 805287 41842 805296
rect 41696 802596 41748 802602
rect 41696 802538 41748 802544
rect 41708 802482 41736 802538
rect 41708 802454 41828 802482
rect 41234 800864 41290 800873
rect 41234 800799 41290 800808
rect 40038 800728 40094 800737
rect 40038 800663 40094 800672
rect 41800 800329 41828 802454
rect 42076 800578 42104 806647
rect 42352 801145 42380 811426
rect 42614 801952 42670 801961
rect 42670 801910 42840 801938
rect 42614 801887 42670 801896
rect 42338 801136 42394 801145
rect 42338 801071 42394 801080
rect 42338 800864 42394 800873
rect 42338 800799 42394 800808
rect 42076 800550 42288 800578
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 798266 42288 800550
rect 42352 800442 42380 800799
rect 42812 800442 42840 801910
rect 42352 800414 42656 800442
rect 42182 798238 42288 798266
rect 42628 797619 42656 800414
rect 42182 797591 42656 797619
rect 42720 800414 42840 800442
rect 42154 797328 42210 797337
rect 42154 797263 42210 797272
rect 42168 796960 42196 797263
rect 41786 796240 41842 796249
rect 41786 796175 41842 796184
rect 41800 795765 41828 796175
rect 42062 795016 42118 795025
rect 42062 794951 42118 794960
rect 42076 794894 42104 794951
rect 42076 794866 42196 794894
rect 42168 794580 42196 794866
rect 41786 794472 41842 794481
rect 41786 794407 41842 794416
rect 41800 793900 41828 794407
rect 41786 793520 41842 793529
rect 41786 793455 41842 793464
rect 41800 793288 41828 793455
rect 42154 792976 42210 792985
rect 42154 792911 42210 792920
rect 42168 792744 42196 792911
rect 42248 792600 42300 792606
rect 42248 792542 42300 792548
rect 42260 791738 42288 792542
rect 42430 792024 42486 792033
rect 42430 791959 42486 791968
rect 42260 791710 42380 791738
rect 42352 790650 42380 791710
rect 42168 790622 42380 790650
rect 42168 790228 42196 790622
rect 42156 790016 42208 790022
rect 42156 789958 42208 789964
rect 42168 789616 42196 789958
rect 42444 789426 42472 791959
rect 42720 790294 42748 800414
rect 42708 790288 42760 790294
rect 42708 790230 42760 790236
rect 42614 790120 42670 790129
rect 42614 790055 42670 790064
rect 42168 789398 42472 789426
rect 42168 788936 42196 789398
rect 42338 789168 42394 789177
rect 42338 789103 42394 789112
rect 42352 788950 42380 789103
rect 42260 788922 42380 788950
rect 42260 788406 42288 788922
rect 42182 788378 42288 788406
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 42260 786570 42288 788151
rect 42628 788066 42656 790055
rect 42182 786542 42288 786570
rect 42352 788038 42656 788066
rect 42352 785958 42380 788038
rect 42522 787944 42578 787953
rect 42522 787879 42578 787888
rect 42168 785890 42196 785944
rect 42260 785930 42380 785958
rect 42260 785890 42288 785930
rect 42168 785862 42288 785890
rect 42536 785278 42564 787879
rect 42182 785250 42564 785278
rect 39762 775296 39818 775305
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 39762 775231 39818 775240
rect 39776 774382 39804 775231
rect 35808 774376 35860 774382
rect 35806 774344 35808 774353
rect 39764 774376 39816 774382
rect 35860 774344 35862 774353
rect 39764 774318 39816 774324
rect 35806 774279 35862 774288
rect 35806 773936 35862 773945
rect 35806 773871 35862 773880
rect 35346 773528 35402 773537
rect 35346 773463 35402 773472
rect 35360 772886 35388 773463
rect 35532 773424 35584 773430
rect 35532 773366 35584 773372
rect 35544 773129 35572 773366
rect 35820 773294 35848 773871
rect 40868 773424 40920 773430
rect 40868 773366 40920 773372
rect 35808 773288 35860 773294
rect 35808 773230 35860 773236
rect 35808 773152 35860 773158
rect 35530 773120 35586 773129
rect 35530 773055 35586 773064
rect 35806 773120 35808 773129
rect 40880 773129 40908 773366
rect 41696 773152 41748 773158
rect 35860 773120 35862 773129
rect 35806 773055 35862 773064
rect 40866 773120 40922 773129
rect 42064 773152 42116 773158
rect 41748 773100 42064 773106
rect 41696 773094 42116 773100
rect 41708 773078 42104 773094
rect 40866 773055 40922 773064
rect 41696 773016 41748 773022
rect 42064 773016 42116 773022
rect 41748 772964 42064 772970
rect 41696 772958 42116 772964
rect 41708 772942 42104 772958
rect 35348 772880 35400 772886
rect 35348 772822 35400 772828
rect 41696 772744 41748 772750
rect 42064 772744 42116 772750
rect 41748 772692 42064 772698
rect 41696 772686 42116 772692
rect 41708 772670 42104 772686
rect 35346 772304 35402 772313
rect 35346 772239 35402 772248
rect 35360 771458 35388 772239
rect 35530 771896 35586 771905
rect 35530 771831 35586 771840
rect 35806 771896 35862 771905
rect 35806 771831 35862 771840
rect 35544 771730 35572 771831
rect 35532 771724 35584 771730
rect 35532 771666 35584 771672
rect 35820 771594 35848 771831
rect 39856 771724 39908 771730
rect 39856 771666 39908 771672
rect 35808 771588 35860 771594
rect 35808 771530 35860 771536
rect 35348 771452 35400 771458
rect 35348 771394 35400 771400
rect 35806 771080 35862 771089
rect 35806 771015 35862 771024
rect 35622 770672 35678 770681
rect 35622 770607 35678 770616
rect 35636 770234 35664 770607
rect 35820 770506 35848 771015
rect 39868 770681 39896 771666
rect 41708 771594 42104 771610
rect 42904 771594 42932 814671
rect 43258 813648 43314 813657
rect 43258 813583 43314 813592
rect 43074 808752 43130 808761
rect 43074 808687 43130 808696
rect 43088 792606 43116 808687
rect 43076 792600 43128 792606
rect 43076 792542 43128 792548
rect 43074 773120 43130 773129
rect 43074 773055 43130 773064
rect 41696 771588 42116 771594
rect 41748 771582 42064 771588
rect 41696 771530 41748 771536
rect 42064 771530 42116 771536
rect 42892 771588 42944 771594
rect 42892 771530 42944 771536
rect 41708 771458 42104 771474
rect 41696 771452 42116 771458
rect 41748 771446 42064 771452
rect 41696 771394 41748 771400
rect 42064 771394 42116 771400
rect 39854 770672 39910 770681
rect 39854 770607 39910 770616
rect 42890 770672 42946 770681
rect 42890 770607 42946 770616
rect 35808 770500 35860 770506
rect 35808 770442 35860 770448
rect 39856 770500 39908 770506
rect 39856 770442 39908 770448
rect 39868 770273 39896 770442
rect 41696 770296 41748 770302
rect 35806 770264 35862 770273
rect 35624 770228 35676 770234
rect 35806 770199 35862 770208
rect 39854 770264 39910 770273
rect 42064 770296 42116 770302
rect 41748 770244 42064 770250
rect 41696 770238 42116 770244
rect 41708 770222 42104 770238
rect 39854 770199 39910 770208
rect 35624 770170 35676 770176
rect 35820 770098 35848 770199
rect 41708 770098 42104 770114
rect 35808 770092 35860 770098
rect 35808 770034 35860 770040
rect 41696 770092 42116 770098
rect 41748 770086 42064 770092
rect 41696 770034 41748 770040
rect 42064 770034 42116 770040
rect 35622 769448 35678 769457
rect 35622 769383 35678 769392
rect 35636 768738 35664 769383
rect 35806 769040 35862 769049
rect 35806 768975 35862 768984
rect 35820 768874 35848 768975
rect 35808 768868 35860 768874
rect 35808 768810 35860 768816
rect 39304 768868 39356 768874
rect 39304 768810 39356 768816
rect 35624 768732 35676 768738
rect 35624 768674 35676 768680
rect 35806 768224 35862 768233
rect 35806 768159 35862 768168
rect 35622 767816 35678 767825
rect 35622 767751 35678 767760
rect 35636 767514 35664 767751
rect 35820 767650 35848 768159
rect 35808 767644 35860 767650
rect 35808 767586 35860 767592
rect 35624 767508 35676 767514
rect 35624 767450 35676 767456
rect 36544 767508 36596 767514
rect 36544 767450 36596 767456
rect 32402 767408 32458 767417
rect 32402 767343 32458 767352
rect 32416 759665 32444 767343
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 32402 759656 32458 759665
rect 32402 759591 32458 759600
rect 35176 758198 35204 766935
rect 35806 766592 35862 766601
rect 35806 766527 35862 766536
rect 35820 766358 35848 766527
rect 35808 766352 35860 766358
rect 35808 766294 35860 766300
rect 35806 766184 35862 766193
rect 35806 766119 35862 766128
rect 35820 765950 35848 766119
rect 35808 765944 35860 765950
rect 35808 765886 35860 765892
rect 35808 764720 35860 764726
rect 35808 764662 35860 764668
rect 35820 764561 35848 764662
rect 35806 764552 35862 764561
rect 35806 764487 35862 764496
rect 35622 764144 35678 764153
rect 35622 764079 35678 764088
rect 35636 763230 35664 764079
rect 35808 763360 35860 763366
rect 35806 763328 35808 763337
rect 35860 763328 35862 763337
rect 35806 763263 35862 763272
rect 35624 763224 35676 763230
rect 35624 763166 35676 763172
rect 35806 762920 35862 762929
rect 35806 762855 35862 762864
rect 35820 761938 35848 762855
rect 35808 761932 35860 761938
rect 35808 761874 35860 761880
rect 36556 759082 36584 767450
rect 39120 764720 39172 764726
rect 39120 764662 39172 764668
rect 39132 763745 39160 764662
rect 39118 763736 39174 763745
rect 39118 763671 39174 763680
rect 37924 763360 37976 763366
rect 37924 763302 37976 763308
rect 36544 759076 36596 759082
rect 36544 759018 36596 759024
rect 35164 758192 35216 758198
rect 35164 758134 35216 758140
rect 37936 757790 37964 763302
rect 37924 757784 37976 757790
rect 39316 757761 39344 768810
rect 42522 768768 42578 768777
rect 41328 768732 41380 768738
rect 42522 768703 42578 768712
rect 41328 768674 41380 768680
rect 40040 767644 40092 767650
rect 40040 767586 40092 767592
rect 39764 766216 39816 766222
rect 39764 766158 39816 766164
rect 39776 764561 39804 766158
rect 40052 765202 40080 767586
rect 41340 765898 41368 768674
rect 41696 766012 41748 766018
rect 41696 765954 41748 765960
rect 41708 765898 41736 765954
rect 42076 765950 42104 765981
rect 42064 765944 42116 765950
rect 41800 765898 42064 765914
rect 41340 765870 41552 765898
rect 41708 765892 42064 765898
rect 41708 765886 42116 765892
rect 42536 765914 42564 768703
rect 42536 765886 42748 765914
rect 41708 765870 41828 765886
rect 40040 765196 40092 765202
rect 40040 765138 40092 765144
rect 41524 764946 41552 765870
rect 41696 765196 41748 765202
rect 41696 765138 41748 765144
rect 41708 765082 41736 765138
rect 41708 765066 42104 765082
rect 41708 765060 42116 765066
rect 41708 765054 42064 765060
rect 42064 765002 42116 765008
rect 42524 765060 42576 765066
rect 42524 765002 42576 765008
rect 42536 764946 42564 765002
rect 41524 764918 42288 764946
rect 39762 764552 39818 764561
rect 39762 764487 39818 764496
rect 41694 763328 41750 763337
rect 41694 763263 41696 763272
rect 41748 763263 41750 763272
rect 41696 763234 41748 763240
rect 40224 761932 40276 761938
rect 40224 761874 40276 761880
rect 39948 759076 40000 759082
rect 39948 759018 40000 759024
rect 37924 757726 37976 757732
rect 39302 757752 39358 757761
rect 39302 757687 39358 757696
rect 39960 757489 39988 759018
rect 40236 758169 40264 761874
rect 42260 758441 42288 764918
rect 42444 764918 42564 764946
rect 42246 758432 42302 758441
rect 42246 758367 42302 758376
rect 42444 758198 42472 764918
rect 41696 758192 41748 758198
rect 40222 758160 40278 758169
rect 41696 758134 41748 758140
rect 42432 758192 42484 758198
rect 42432 758134 42484 758140
rect 40222 758095 40278 758104
rect 41708 757874 41736 758134
rect 41970 757888 42026 757897
rect 41708 757846 41970 757874
rect 41970 757823 42026 757832
rect 42430 757888 42486 757897
rect 42486 757846 42656 757874
rect 42430 757823 42486 757832
rect 41604 757784 41656 757790
rect 41656 757732 41828 757738
rect 41604 757726 41828 757732
rect 41616 757710 41828 757726
rect 39946 757480 40002 757489
rect 39946 757415 40002 757424
rect 41800 757081 41828 757710
rect 42432 757648 42484 757654
rect 42432 757590 42484 757596
rect 42246 757480 42302 757489
rect 42246 757415 42302 757424
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 42260 756786 42288 757415
rect 42168 756758 42288 756786
rect 42168 756228 42196 756758
rect 41970 755440 42026 755449
rect 41970 755375 42026 755384
rect 41984 755072 42012 755375
rect 42154 754896 42210 754905
rect 42154 754831 42210 754840
rect 42168 754392 42196 754831
rect 42248 754316 42300 754322
rect 42248 754258 42300 754264
rect 42062 754080 42118 754089
rect 42062 754015 42118 754024
rect 42076 753780 42104 754015
rect 42260 753250 42288 754258
rect 42444 753494 42472 757590
rect 42444 753466 42564 753494
rect 42260 753222 42380 753250
rect 42352 752978 42380 753222
rect 42168 752950 42380 752978
rect 42168 752556 42196 752950
rect 42246 752176 42302 752185
rect 42246 752111 42302 752120
rect 42062 751768 42118 751777
rect 42062 751703 42118 751712
rect 42076 751369 42104 751703
rect 41786 751088 41842 751097
rect 41786 751023 41842 751032
rect 41800 750720 41828 751023
rect 42168 749986 42196 750108
rect 42260 749986 42288 752111
rect 42168 749958 42288 749986
rect 42168 749550 42380 749578
rect 42168 749529 42196 749550
rect 42352 749543 42380 749550
rect 42536 749543 42564 753466
rect 42352 749515 42564 749543
rect 42246 749456 42302 749465
rect 42246 749391 42302 749400
rect 42260 747062 42288 749391
rect 42432 749352 42484 749358
rect 42432 749294 42484 749300
rect 42182 747034 42288 747062
rect 42444 746722 42472 749294
rect 42076 746694 42472 746722
rect 42076 746401 42104 746694
rect 42246 746600 42302 746609
rect 42246 746535 42302 746544
rect 42062 746056 42118 746065
rect 42062 745991 42118 746000
rect 42076 745756 42104 745991
rect 42062 745512 42118 745521
rect 42062 745447 42118 745456
rect 42076 745212 42104 745447
rect 42260 743390 42288 746535
rect 42430 746328 42486 746337
rect 42430 746263 42486 746272
rect 42182 743362 42288 743390
rect 42168 742750 42288 742778
rect 42168 742696 42196 742750
rect 42260 742710 42288 742750
rect 42444 742710 42472 746263
rect 42628 746065 42656 757846
rect 42720 746178 42748 765886
rect 42720 746150 42840 746178
rect 42614 746056 42670 746065
rect 42614 745991 42670 746000
rect 42812 745906 42840 746150
rect 42720 745878 42840 745906
rect 42720 745521 42748 745878
rect 42706 745512 42762 745521
rect 42706 745447 42762 745456
rect 42614 745104 42670 745113
rect 42614 745039 42670 745048
rect 42260 742682 42472 742710
rect 42628 742098 42656 745039
rect 42182 742070 42656 742098
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42904 729337 42932 770607
rect 43088 730153 43116 773055
rect 43272 770302 43300 813583
rect 43260 770296 43312 770302
rect 43260 770238 43312 770244
rect 43258 764552 43314 764561
rect 43258 764487 43314 764496
rect 43272 749358 43300 764487
rect 43456 754089 43484 870810
rect 44824 844620 44876 844626
rect 44824 844562 44876 844568
rect 44180 814292 44232 814298
rect 44180 814234 44232 814240
rect 43628 807492 43680 807498
rect 43628 807434 43680 807440
rect 43640 807265 43668 807434
rect 43626 807256 43682 807265
rect 43626 807191 43682 807200
rect 43628 799060 43680 799066
rect 43628 799002 43680 799008
rect 43640 797337 43668 799002
rect 43626 797328 43682 797337
rect 43626 797263 43682 797272
rect 44192 771458 44220 814234
rect 44454 812832 44510 812841
rect 44454 812767 44510 812776
rect 44468 773158 44496 812767
rect 44638 807936 44694 807945
rect 44638 807871 44694 807880
rect 44652 795025 44680 807871
rect 44638 795016 44694 795025
rect 44638 794951 44694 794960
rect 44836 775305 44864 844562
rect 46216 819097 46244 896990
rect 46202 819088 46258 819097
rect 46202 819023 46258 819032
rect 46202 806304 46258 806313
rect 46202 806239 46258 806248
rect 44822 775296 44878 775305
rect 44822 775231 44878 775240
rect 44456 773152 44508 773158
rect 44456 773094 44508 773100
rect 44180 771452 44232 771458
rect 44180 771394 44232 771400
rect 44270 770264 44326 770273
rect 44270 770199 44326 770208
rect 43628 767372 43680 767378
rect 43628 767314 43680 767320
rect 43442 754080 43498 754089
rect 43442 754015 43498 754024
rect 43444 753568 43496 753574
rect 43444 753510 43496 753516
rect 43456 751777 43484 753510
rect 43442 751768 43498 751777
rect 43442 751703 43498 751712
rect 43260 749352 43312 749358
rect 43260 749294 43312 749300
rect 43444 731196 43496 731202
rect 43444 731138 43496 731144
rect 43258 730960 43314 730969
rect 43258 730895 43314 730904
rect 43272 730182 43300 730895
rect 43456 730561 43484 731138
rect 43442 730552 43498 730561
rect 43442 730487 43498 730496
rect 43260 730176 43312 730182
rect 43074 730144 43130 730153
rect 43260 730118 43312 730124
rect 43074 730079 43130 730088
rect 42890 729328 42946 729337
rect 42890 729263 42946 729272
rect 40866 728682 40922 728691
rect 40866 728617 40922 728626
rect 41326 728682 41382 728691
rect 41326 728617 41382 728626
rect 41696 728680 41748 728686
rect 42064 728680 42116 728686
rect 41748 728640 42064 728668
rect 41696 728622 41748 728628
rect 42064 728622 42116 728628
rect 40880 727326 40908 728617
rect 42890 728104 42946 728113
rect 42890 728039 42946 728048
rect 41050 727458 41106 727467
rect 41050 727393 41106 727402
rect 41696 727456 41748 727462
rect 42064 727456 42116 727462
rect 41748 727416 42064 727444
rect 41696 727398 41748 727404
rect 42064 727398 42116 727404
rect 40868 727320 40920 727326
rect 40868 727262 40920 727268
rect 41696 727320 41748 727326
rect 42064 727320 42116 727326
rect 41748 727268 42064 727274
rect 41696 727262 42116 727268
rect 41708 727246 42104 727262
rect 41326 726880 41382 726889
rect 41326 726815 41382 726824
rect 41340 726374 41368 726815
rect 42522 726472 42578 726481
rect 42522 726407 42578 726416
rect 41328 726368 41380 726374
rect 41328 726310 41380 726316
rect 41604 726368 41656 726374
rect 41604 726310 41656 726316
rect 40958 726234 41014 726243
rect 40958 726169 41014 726178
rect 37922 725248 37978 725257
rect 37922 725183 37978 725192
rect 35162 724840 35218 724849
rect 35162 724775 35218 724784
rect 33046 724432 33102 724441
rect 33046 724367 33102 724376
rect 31758 720352 31814 720361
rect 31758 720287 31760 720296
rect 31812 720287 31814 720296
rect 31760 720258 31812 720264
rect 33060 716825 33088 724367
rect 33782 723786 33838 723795
rect 33782 723721 33838 723730
rect 33046 716816 33102 716825
rect 33046 716751 33102 716760
rect 33796 715426 33824 723721
rect 35176 715698 35204 724775
rect 37936 716106 37964 725183
rect 40682 723208 40738 723217
rect 40682 723143 40738 723152
rect 40040 720316 40092 720322
rect 40040 720258 40092 720264
rect 37924 716100 37976 716106
rect 37924 716042 37976 716048
rect 35164 715692 35216 715698
rect 35164 715634 35216 715640
rect 33784 715420 33836 715426
rect 33784 715362 33836 715368
rect 40052 714542 40080 720258
rect 40316 716100 40368 716106
rect 40316 716042 40368 716048
rect 40328 714921 40356 716042
rect 40314 714912 40370 714921
rect 40314 714847 40370 714856
rect 40040 714536 40092 714542
rect 40040 714478 40092 714484
rect 40696 714241 40724 723143
rect 40972 721754 41000 726169
rect 41616 725778 41644 726310
rect 41786 725792 41842 725801
rect 41616 725750 41786 725778
rect 41786 725727 41842 725736
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41142 721768 41198 721777
rect 40972 721726 41142 721754
rect 41142 721703 41198 721712
rect 41340 718321 41368 725591
rect 41786 722392 41842 722401
rect 41786 722327 41842 722336
rect 41800 718593 41828 722327
rect 42338 719944 42394 719953
rect 42338 719879 42394 719888
rect 42352 719166 42380 719879
rect 42340 719160 42392 719166
rect 42340 719102 42392 719108
rect 41786 718584 41842 718593
rect 41786 718519 41842 718528
rect 41326 718312 41382 718321
rect 41326 718247 41382 718256
rect 42338 718312 42394 718321
rect 42338 718247 42394 718256
rect 41328 715692 41380 715698
rect 41328 715634 41380 715640
rect 41340 714854 41368 715634
rect 41696 715420 41748 715426
rect 41696 715362 41748 715368
rect 41708 715306 41736 715362
rect 41708 715290 42104 715306
rect 41708 715284 42116 715290
rect 41708 715278 42064 715284
rect 42064 715226 42116 715232
rect 42352 715034 42380 718247
rect 42536 715193 42564 726407
rect 42708 715284 42760 715290
rect 42708 715226 42760 715232
rect 42522 715184 42578 715193
rect 42720 715170 42748 715226
rect 42720 715142 42840 715170
rect 42522 715119 42578 715128
rect 42352 715006 42656 715034
rect 42338 714912 42394 714921
rect 41340 714826 41460 714854
rect 42338 714847 42394 714856
rect 40682 714232 40738 714241
rect 41432 714218 41460 714826
rect 41696 714536 41748 714542
rect 41748 714484 42288 714490
rect 41696 714478 42288 714484
rect 41708 714462 42288 714478
rect 41432 714190 41828 714218
rect 40682 714167 40738 714176
rect 41800 713969 41828 714190
rect 41786 713960 41842 713969
rect 41786 713895 41842 713904
rect 41786 713552 41842 713561
rect 41786 713487 41842 713496
rect 41800 713048 41828 713487
rect 42260 712314 42288 714462
rect 42168 712286 42288 712314
rect 42168 711824 42196 712286
rect 42154 711648 42210 711657
rect 42154 711583 42210 711592
rect 42168 711212 42196 711583
rect 42352 711090 42380 714847
rect 42352 711062 42564 711090
rect 42248 711000 42300 711006
rect 42076 710948 42248 710954
rect 42076 710942 42300 710948
rect 42076 710926 42288 710942
rect 42076 710561 42104 710926
rect 41786 709880 41842 709889
rect 41786 709815 41842 709824
rect 41800 709376 41828 709815
rect 41786 708520 41842 708529
rect 41786 708455 41842 708464
rect 41800 708152 41828 708455
rect 42340 708416 42392 708422
rect 42340 708358 42392 708364
rect 42352 707554 42380 708358
rect 42182 707526 42380 707554
rect 41878 707160 41934 707169
rect 41878 707095 41934 707104
rect 41892 706860 41920 707095
rect 42536 706330 42564 711062
rect 42182 706302 42564 706330
rect 42246 706208 42302 706217
rect 42246 706143 42302 706152
rect 42260 704290 42288 706143
rect 42628 705194 42656 715006
rect 42812 713474 42840 715142
rect 42076 704262 42288 704290
rect 42444 705166 42656 705194
rect 42720 713446 42840 713474
rect 42076 703868 42104 704262
rect 42246 703760 42302 703769
rect 42246 703695 42302 703704
rect 42062 703488 42118 703497
rect 42062 703423 42118 703432
rect 42076 703188 42104 703423
rect 42062 703080 42118 703089
rect 42062 703015 42118 703024
rect 42076 702576 42104 703015
rect 42260 702166 42288 703695
rect 42248 702160 42300 702166
rect 42248 702102 42300 702108
rect 42444 702046 42472 705166
rect 42720 703089 42748 713446
rect 42904 712722 42932 728039
rect 43076 727456 43128 727462
rect 43076 727398 43128 727404
rect 43088 712858 43116 727398
rect 43258 723616 43314 723625
rect 43258 723551 43314 723560
rect 43272 714854 43300 723551
rect 43272 714826 43484 714854
rect 43088 712830 43208 712858
rect 42904 712694 43116 712722
rect 42892 712292 42944 712298
rect 42892 712234 42944 712240
rect 42904 711006 42932 712234
rect 42892 711000 42944 711006
rect 42892 710942 42944 710948
rect 43088 707954 43116 712694
rect 43180 709866 43208 712830
rect 43180 709838 43300 709866
rect 42904 707926 43116 707954
rect 42706 703080 42762 703089
rect 42706 703015 42762 703024
rect 42614 702400 42670 702409
rect 42614 702335 42670 702344
rect 42168 701978 42196 702032
rect 42260 702018 42472 702046
rect 42260 701978 42288 702018
rect 42168 701950 42288 701978
rect 42248 701888 42300 701894
rect 42248 701830 42300 701836
rect 42430 701856 42486 701865
rect 42260 700179 42288 701830
rect 42430 701791 42486 701800
rect 42182 700151 42288 700179
rect 42444 699530 42472 701791
rect 42182 699502 42472 699530
rect 42628 698918 42656 702335
rect 42168 698850 42196 698904
rect 42260 698890 42656 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 40958 688392 41014 688401
rect 40958 688327 41014 688336
rect 40972 687274 41000 688327
rect 40960 687268 41012 687274
rect 40960 687210 41012 687216
rect 41696 687268 41748 687274
rect 42064 687268 42116 687274
rect 41748 687228 42064 687256
rect 41696 687210 41748 687216
rect 42064 687210 42116 687216
rect 41142 686896 41198 686905
rect 41142 686831 41198 686840
rect 41156 686050 41184 686831
rect 41696 686112 41748 686118
rect 42064 686112 42116 686118
rect 41748 686060 42064 686066
rect 41696 686054 42116 686060
rect 41144 686044 41196 686050
rect 41708 686038 42104 686054
rect 41144 685986 41196 685992
rect 40866 685910 40922 685919
rect 40866 685845 40922 685854
rect 41326 685910 41382 685919
rect 41326 685845 41382 685854
rect 41696 685908 41748 685914
rect 42064 685908 42116 685914
rect 41748 685868 42064 685896
rect 41696 685850 41748 685856
rect 42064 685850 42116 685856
rect 40880 684826 40908 685845
rect 41142 685264 41198 685273
rect 41142 685199 41198 685208
rect 40868 684820 40920 684826
rect 40868 684762 40920 684768
rect 41156 684690 41184 685199
rect 42706 684856 42762 684865
rect 42706 684791 42762 684800
rect 41696 684752 41748 684758
rect 42064 684752 42116 684758
rect 41748 684700 42064 684706
rect 41696 684694 42116 684700
rect 41144 684684 41196 684690
rect 41708 684678 42104 684694
rect 41144 684626 41196 684632
rect 41708 684554 42104 684570
rect 41696 684548 42116 684554
rect 41748 684542 42064 684548
rect 41696 684490 41748 684496
rect 42064 684490 42116 684496
rect 40958 683632 41014 683641
rect 40958 683567 41014 683576
rect 40774 682816 40830 682825
rect 40774 682751 40830 682760
rect 40590 682408 40646 682417
rect 40590 682343 40646 682352
rect 37922 682000 37978 682009
rect 37922 681935 37978 681944
rect 36542 681592 36598 681601
rect 36542 681527 36598 681536
rect 32402 681184 32458 681193
rect 32402 681119 32458 681128
rect 32416 672761 32444 681119
rect 33782 680776 33838 680785
rect 33782 680711 33838 680720
rect 33796 672790 33824 680711
rect 33784 672784 33836 672790
rect 32402 672752 32458 672761
rect 33784 672726 33836 672732
rect 32402 672687 32458 672696
rect 36556 672110 36584 681527
rect 36544 672104 36596 672110
rect 36544 672046 36596 672052
rect 37936 671294 37964 681935
rect 40604 679250 40632 682343
rect 40788 679386 40816 682751
rect 40972 682394 41000 683567
rect 41328 683528 41380 683534
rect 41328 683470 41380 683476
rect 41696 683528 41748 683534
rect 41748 683476 42012 683482
rect 41696 683470 42012 683476
rect 41340 683233 41368 683470
rect 41708 683454 42012 683470
rect 41326 683224 41382 683233
rect 41326 683159 41382 683168
rect 41786 682408 41842 682417
rect 40972 682366 41786 682394
rect 41786 682343 41842 682352
rect 41984 681578 42012 683454
rect 41984 681550 42472 681578
rect 40776 679380 40828 679386
rect 40776 679322 40828 679328
rect 41328 679380 41380 679386
rect 41328 679322 41380 679328
rect 40592 679244 40644 679250
rect 40592 679186 40644 679192
rect 41340 678858 41368 679322
rect 41696 679244 41748 679250
rect 41696 679186 41748 679192
rect 41708 678974 41736 679186
rect 41708 678946 42380 678974
rect 41786 678872 41842 678881
rect 41340 678830 41786 678858
rect 41786 678807 41842 678816
rect 41142 677104 41198 677113
rect 41142 677039 41198 677048
rect 39488 672784 39540 672790
rect 39488 672726 39540 672732
rect 39500 671537 39528 672726
rect 41156 672489 41184 677039
rect 42352 676214 42380 678946
rect 42260 676186 42380 676214
rect 41142 672480 41198 672489
rect 41142 672415 41198 672424
rect 42260 672217 42288 676186
rect 42246 672208 42302 672217
rect 42246 672143 42302 672152
rect 41696 672104 41748 672110
rect 41748 672052 42288 672058
rect 41696 672046 42288 672052
rect 41708 672030 42288 672046
rect 39486 671528 39542 671537
rect 39486 671463 39542 671472
rect 37924 671288 37976 671294
rect 40040 671288 40092 671294
rect 37924 671230 37976 671236
rect 40038 671256 40040 671265
rect 40092 671256 40094 671265
rect 40038 671191 40094 671200
rect 42168 669746 42196 669868
rect 42260 669746 42288 672030
rect 42444 670970 42472 681550
rect 42720 676214 42748 684791
rect 42904 684758 42932 707926
rect 43076 707804 43128 707810
rect 43076 707746 43128 707752
rect 43088 705194 43116 707746
rect 43272 705194 43300 709838
rect 43456 707810 43484 714826
rect 43444 707804 43496 707810
rect 43444 707746 43496 707752
rect 43088 705166 43208 705194
rect 43272 705166 43392 705194
rect 43180 703497 43208 705166
rect 43166 703488 43222 703497
rect 43166 703423 43222 703432
rect 43364 698294 43392 705166
rect 43088 698266 43392 698294
rect 42892 684752 42944 684758
rect 42892 684694 42944 684700
rect 43088 684457 43116 698266
rect 43444 687744 43496 687750
rect 43258 687712 43314 687721
rect 43444 687686 43496 687692
rect 43258 687647 43314 687656
rect 43272 687410 43300 687647
rect 43260 687404 43312 687410
rect 43260 687346 43312 687352
rect 43456 687313 43484 687686
rect 43442 687304 43498 687313
rect 43442 687239 43498 687248
rect 43074 684448 43130 684457
rect 43074 684383 43130 684392
rect 43258 684040 43314 684049
rect 43258 683975 43314 683984
rect 43272 683210 43300 683975
rect 43088 683182 43300 683210
rect 42720 676186 42932 676214
rect 42706 671528 42762 671537
rect 42536 671486 42706 671514
rect 42536 671106 42564 671486
rect 42706 671463 42762 671472
rect 42706 671256 42762 671265
rect 42706 671191 42762 671200
rect 42536 671078 42656 671106
rect 42444 670942 42564 670970
rect 42168 669718 42288 669746
rect 41786 669080 41842 669089
rect 41786 669015 41842 669024
rect 41800 668644 41828 669015
rect 42536 668046 42564 670942
rect 42168 667978 42196 668032
rect 42260 668018 42564 668046
rect 42260 667978 42288 668018
rect 42168 667950 42288 667978
rect 42248 667820 42300 667826
rect 42248 667762 42300 667768
rect 42062 667720 42118 667729
rect 42062 667655 42118 667664
rect 42076 667352 42104 667655
rect 42260 666179 42288 667762
rect 42430 667448 42486 667457
rect 42430 667383 42486 667392
rect 42182 666151 42288 666179
rect 42248 666052 42300 666058
rect 42248 665994 42300 666000
rect 42062 665136 42118 665145
rect 42062 665071 42118 665080
rect 42076 664972 42104 665071
rect 42260 664850 42288 665994
rect 42168 664822 42288 664850
rect 42168 664325 42196 664822
rect 42444 664442 42472 667383
rect 42444 664414 42564 664442
rect 41786 664184 41842 664193
rect 42536 664170 42564 664414
rect 41786 664119 41842 664128
rect 42352 664142 42564 664170
rect 41800 663680 41828 664119
rect 42352 663270 42380 664142
rect 42628 663354 42656 671078
rect 42536 663338 42656 663354
rect 42524 663332 42656 663338
rect 42576 663326 42656 663332
rect 42524 663274 42576 663280
rect 42340 663264 42392 663270
rect 42340 663206 42392 663212
rect 42720 663150 42748 671191
rect 42182 663122 42748 663150
rect 42708 663060 42760 663066
rect 42708 663002 42760 663008
rect 42524 662992 42576 662998
rect 42352 662940 42524 662946
rect 42352 662934 42576 662940
rect 42352 662918 42564 662934
rect 42154 662824 42210 662833
rect 42154 662759 42210 662768
rect 42168 662674 42196 662759
rect 42168 662646 42288 662674
rect 42260 661042 42288 662646
rect 42168 661014 42288 661042
rect 42168 660620 42196 661014
rect 42156 660544 42208 660550
rect 42156 660486 42208 660492
rect 42168 660008 42196 660486
rect 42352 659371 42380 662918
rect 42524 662720 42576 662726
rect 42524 662662 42576 662668
rect 42536 662402 42564 662662
rect 42182 659343 42380 659371
rect 42444 662374 42564 662402
rect 42444 659002 42472 662374
rect 42720 660550 42748 663002
rect 42708 660544 42760 660550
rect 42708 660486 42760 660492
rect 42614 660376 42670 660385
rect 42614 660311 42670 660320
rect 42168 658974 42472 659002
rect 42168 658784 42196 658974
rect 42430 658880 42486 658889
rect 42430 658815 42486 658824
rect 42246 658608 42302 658617
rect 42246 658543 42302 658552
rect 42064 657416 42116 657422
rect 42064 657358 42116 657364
rect 42076 656948 42104 657358
rect 42260 656350 42288 658543
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42444 655670 42472 658815
rect 42628 657422 42656 660311
rect 42616 657416 42668 657422
rect 42616 657358 42668 657364
rect 42260 655642 42472 655670
rect 39394 646096 39450 646105
rect 39394 646031 39450 646040
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 39408 644774 39436 646031
rect 35808 644768 35860 644774
rect 35530 644736 35586 644745
rect 35530 644671 35586 644680
rect 35806 644736 35808 644745
rect 39396 644768 39448 644774
rect 35860 644736 35862 644745
rect 39396 644710 39448 644716
rect 39762 644736 39818 644745
rect 35806 644671 35862 644680
rect 39762 644671 39818 644680
rect 35544 644502 35572 644671
rect 39776 644502 39804 644671
rect 35532 644496 35584 644502
rect 35532 644438 35584 644444
rect 39764 644496 39816 644502
rect 39764 644438 39816 644444
rect 35346 643920 35402 643929
rect 35346 643855 35402 643864
rect 39854 643920 39910 643929
rect 39854 643855 39910 643864
rect 35360 643142 35388 643855
rect 35808 643544 35860 643550
rect 35530 643512 35586 643521
rect 35530 643447 35586 643456
rect 35806 643512 35808 643521
rect 39672 643544 39724 643550
rect 35860 643512 35862 643521
rect 35806 643447 35862 643456
rect 39670 643512 39672 643521
rect 39724 643512 39726 643521
rect 39670 643447 39726 643456
rect 35544 643278 35572 643447
rect 35532 643272 35584 643278
rect 35532 643214 35584 643220
rect 35348 643136 35400 643142
rect 35348 643078 35400 643084
rect 39578 643104 39634 643113
rect 39578 643039 39634 643048
rect 35438 642696 35494 642705
rect 35438 642631 35494 642640
rect 35452 641918 35480 642631
rect 35622 642288 35678 642297
rect 35622 642223 35678 642232
rect 38934 642288 38990 642297
rect 38934 642223 38936 642232
rect 35440 641912 35492 641918
rect 35440 641854 35492 641860
rect 35636 641782 35664 642223
rect 38988 642223 38990 642232
rect 38936 642194 38988 642200
rect 35808 642184 35860 642190
rect 35808 642126 35860 642132
rect 35820 641889 35848 642126
rect 39592 642054 39620 643039
rect 39580 642048 39632 642054
rect 39580 641990 39632 641996
rect 35806 641880 35862 641889
rect 35806 641815 35862 641824
rect 35624 641776 35676 641782
rect 35624 641718 35676 641724
rect 35806 641472 35862 641481
rect 35806 641407 35862 641416
rect 35622 641064 35678 641073
rect 35622 640999 35678 641008
rect 35636 640490 35664 640999
rect 35820 640830 35848 641407
rect 35808 640824 35860 640830
rect 35808 640766 35860 640772
rect 39672 640756 39724 640762
rect 39672 640698 39724 640704
rect 35806 640656 35862 640665
rect 35806 640591 35862 640600
rect 35624 640484 35676 640490
rect 35624 640426 35676 640432
rect 35820 640354 35848 640591
rect 35808 640348 35860 640354
rect 35808 640290 35860 640296
rect 39684 640257 39712 640698
rect 39868 640490 39896 643855
rect 41708 643346 42104 643362
rect 41696 643340 42116 643346
rect 41748 643334 42064 643340
rect 41696 643282 41748 643288
rect 42064 643282 42116 643288
rect 41696 643136 41748 643142
rect 42064 643136 42116 643142
rect 41748 643084 42064 643090
rect 41696 643078 42116 643084
rect 41708 643062 42104 643078
rect 42904 642297 42932 676186
rect 43088 643929 43116 683182
rect 43442 680368 43498 680377
rect 43442 680303 43498 680312
rect 43258 678328 43314 678337
rect 43258 678263 43314 678272
rect 43272 665145 43300 678263
rect 43258 665136 43314 665145
rect 43258 665071 43314 665080
rect 43456 663066 43484 680303
rect 43640 667729 43668 767314
rect 44284 727326 44312 770199
rect 44640 770092 44692 770098
rect 44640 770034 44692 770040
rect 44456 765944 44508 765950
rect 44456 765886 44508 765892
rect 44468 754934 44496 765886
rect 44456 754928 44508 754934
rect 44456 754870 44508 754876
rect 44454 729736 44510 729745
rect 44454 729671 44510 729680
rect 44272 727320 44324 727326
rect 44272 727262 44324 727268
rect 44178 722800 44234 722809
rect 44178 722735 44234 722744
rect 44192 709374 44220 722735
rect 44180 709368 44232 709374
rect 44180 709310 44232 709316
rect 43812 688696 43864 688702
rect 43812 688638 43864 688644
rect 43626 667720 43682 667729
rect 43626 667655 43682 667664
rect 43444 663060 43496 663066
rect 43444 663002 43496 663008
rect 43444 662448 43496 662454
rect 43444 662390 43496 662396
rect 43074 643920 43130 643929
rect 43074 643855 43130 643864
rect 42890 642288 42946 642297
rect 42890 642223 42946 642232
rect 41696 641776 41748 641782
rect 42064 641776 42116 641782
rect 41748 641724 42064 641730
rect 41696 641718 42116 641724
rect 41708 641702 42104 641718
rect 39856 640484 39908 640490
rect 39856 640426 39908 640432
rect 41696 640348 41748 640354
rect 42064 640348 42116 640354
rect 41748 640306 42064 640334
rect 41696 640290 41748 640296
rect 42064 640290 42116 640296
rect 43076 640348 43128 640354
rect 43076 640290 43128 640296
rect 39670 640248 39726 640257
rect 39670 640183 39726 640192
rect 35346 639840 35402 639849
rect 35346 639775 35402 639784
rect 33782 638616 33838 638625
rect 33782 638551 33838 638560
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 33796 630086 33824 638551
rect 35360 638246 35388 639775
rect 35530 639432 35586 639441
rect 35530 639367 35586 639376
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 35544 638994 35572 639367
rect 35820 639130 35848 639367
rect 35808 639124 35860 639130
rect 35808 639066 35860 639072
rect 40224 639124 40276 639130
rect 40224 639066 40276 639072
rect 35532 638988 35584 638994
rect 35532 638930 35584 638936
rect 40040 638988 40092 638994
rect 40040 638930 40092 638936
rect 35348 638240 35400 638246
rect 35348 638182 35400 638188
rect 35532 637968 35584 637974
rect 35532 637910 35584 637916
rect 35544 637809 35572 637910
rect 35530 637800 35586 637809
rect 35530 637735 35586 637744
rect 35806 637800 35862 637809
rect 35806 637735 35808 637744
rect 35860 637735 35862 637744
rect 35808 637706 35860 637712
rect 40052 637401 40080 638930
rect 40038 637392 40094 637401
rect 40038 637327 40094 637336
rect 35806 636576 35862 636585
rect 35806 636511 35862 636520
rect 35820 636410 35848 636511
rect 35808 636404 35860 636410
rect 35808 636346 35860 636352
rect 40236 635361 40264 639066
rect 41696 638240 41748 638246
rect 41510 638208 41566 638217
rect 41696 638182 41748 638188
rect 41510 638143 41566 638152
rect 40960 637968 41012 637974
rect 40960 637910 41012 637916
rect 40972 637809 41000 637910
rect 40958 637800 41014 637809
rect 41524 637770 41552 638143
rect 40958 637735 41014 637744
rect 41512 637764 41564 637770
rect 41512 637706 41564 637712
rect 40684 636404 40736 636410
rect 40684 636346 40736 636352
rect 35622 635352 35678 635361
rect 35622 635287 35678 635296
rect 40222 635352 40278 635361
rect 40222 635287 40278 635296
rect 35636 634846 35664 635287
rect 35808 635112 35860 635118
rect 35808 635054 35860 635060
rect 39580 635112 39632 635118
rect 39580 635054 39632 635060
rect 35820 634953 35848 635054
rect 39592 634953 39620 635054
rect 35806 634944 35862 634953
rect 35806 634879 35862 634888
rect 39578 634944 39634 634953
rect 39578 634879 39634 634888
rect 35624 634840 35676 634846
rect 35624 634782 35676 634788
rect 40500 634840 40552 634846
rect 40500 634782 40552 634788
rect 35806 634536 35862 634545
rect 35806 634471 35862 634480
rect 35820 633894 35848 634471
rect 35808 633888 35860 633894
rect 35808 633830 35860 633836
rect 35806 633720 35862 633729
rect 35806 633655 35862 633664
rect 35820 633554 35848 633655
rect 35808 633548 35860 633554
rect 35808 633490 35860 633496
rect 40512 632097 40540 634782
rect 40696 634545 40724 636346
rect 41708 635202 41736 638182
rect 41708 635174 42564 635202
rect 40682 634536 40738 634545
rect 40682 634471 40738 634480
rect 42338 633856 42394 633865
rect 42338 633791 42394 633800
rect 41696 633752 41748 633758
rect 42064 633752 42116 633758
rect 41748 633700 42064 633706
rect 41696 633694 42116 633700
rect 41708 633678 42104 633694
rect 41708 633554 42104 633570
rect 41696 633548 42116 633554
rect 41748 633542 42064 633548
rect 41696 633490 41748 633496
rect 42064 633490 42116 633496
rect 40498 632088 40554 632097
rect 40498 632023 40554 632032
rect 33784 630080 33836 630086
rect 33784 630022 33836 630028
rect 41696 630080 41748 630086
rect 41748 630028 42104 630034
rect 41696 630022 42104 630028
rect 41708 630018 42104 630022
rect 41708 630012 42116 630018
rect 41708 630006 42064 630012
rect 42064 629954 42116 629960
rect 32404 629944 32456 629950
rect 32404 629886 32456 629892
rect 41696 629944 41748 629950
rect 41748 629892 42288 629898
rect 41696 629886 42288 629892
rect 41708 629870 42288 629886
rect 42260 627178 42288 629870
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42352 625818 42380 633791
rect 42168 625790 42380 625818
rect 42168 625464 42196 625790
rect 42338 625424 42394 625433
rect 42536 625394 42564 635174
rect 42708 630012 42760 630018
rect 42708 629954 42760 629960
rect 42338 625359 42394 625368
rect 42524 625388 42576 625394
rect 42352 625274 42380 625359
rect 42524 625330 42576 625336
rect 42352 625246 42656 625274
rect 42248 625184 42300 625190
rect 42248 625126 42300 625132
rect 42260 624866 42288 625126
rect 42168 624838 42288 624866
rect 42168 624784 42196 624838
rect 42340 624708 42392 624714
rect 42340 624650 42392 624656
rect 42154 624608 42210 624617
rect 42154 624543 42210 624552
rect 42168 624172 42196 624543
rect 42154 623384 42210 623393
rect 42154 623319 42210 623328
rect 42168 622948 42196 623319
rect 42352 622146 42380 624650
rect 42628 623234 42656 625246
rect 42076 622118 42380 622146
rect 42536 623206 42656 623234
rect 42076 621792 42104 622118
rect 42536 621126 42564 623206
rect 42182 621098 42564 621126
rect 42062 620936 42118 620945
rect 42062 620871 42118 620880
rect 42076 620500 42104 620871
rect 42720 620265 42748 629954
rect 42892 626680 42944 626686
rect 42892 626622 42944 626628
rect 42904 624617 42932 626622
rect 42890 624608 42946 624617
rect 42890 624543 42946 624552
rect 43088 621014 43116 640290
rect 43258 640248 43314 640257
rect 43258 640183 43314 640192
rect 43272 621014 43300 640183
rect 42904 620986 43116 621014
rect 43180 620986 43300 621014
rect 42062 620256 42118 620265
rect 42062 620191 42118 620200
rect 42706 620256 42762 620265
rect 42706 620191 42762 620200
rect 42076 619956 42104 620191
rect 42246 619848 42302 619857
rect 42246 619783 42302 619792
rect 42260 617454 42288 619783
rect 42430 619032 42486 619041
rect 42430 618967 42486 618976
rect 42182 617426 42288 617454
rect 42444 616842 42472 618967
rect 42616 618928 42668 618934
rect 42168 616706 42196 616828
rect 42260 616814 42472 616842
rect 42536 618876 42616 618882
rect 42536 618870 42668 618876
rect 42536 618854 42656 618870
rect 42260 616706 42288 616814
rect 42168 616678 42288 616706
rect 42536 616434 42564 618854
rect 42706 618760 42762 618769
rect 42706 618695 42762 618704
rect 42168 616406 42564 616434
rect 42168 616148 42196 616406
rect 42246 616040 42302 616049
rect 42246 615975 42302 615984
rect 42260 615738 42288 615975
rect 42248 615732 42300 615738
rect 42248 615674 42300 615680
rect 42720 615618 42748 618695
rect 42182 615590 42748 615618
rect 42248 615528 42300 615534
rect 42248 615470 42300 615476
rect 42260 613782 42288 615470
rect 42182 613754 42288 613782
rect 42156 613624 42208 613630
rect 42156 613566 42208 613572
rect 42168 613121 42196 613566
rect 41786 612776 41842 612785
rect 41786 612711 41842 612720
rect 41800 612476 41828 612711
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 35806 601760 35862 601769
rect 41708 601730 42104 601746
rect 35806 601695 35808 601704
rect 35860 601695 35862 601704
rect 41696 601724 42116 601730
rect 35808 601666 35860 601672
rect 41748 601718 42064 601724
rect 41696 601666 41748 601672
rect 42064 601666 42116 601672
rect 41326 599312 41382 599321
rect 41326 599247 41382 599256
rect 41340 599010 41368 599247
rect 41328 599004 41380 599010
rect 41328 598946 41380 598952
rect 41696 599004 41748 599010
rect 42064 599004 42116 599010
rect 41748 598964 42064 598992
rect 41696 598946 41748 598952
rect 42064 598946 42116 598952
rect 40866 598904 40922 598913
rect 40866 598839 40922 598848
rect 40880 597718 40908 598839
rect 42706 598496 42762 598505
rect 42706 598431 42762 598440
rect 41708 597922 42104 597938
rect 41696 597916 42116 597922
rect 41748 597910 42064 597916
rect 41050 597850 41106 597859
rect 41050 597785 41106 597794
rect 41326 597850 41382 597859
rect 41696 597858 41748 597864
rect 42064 597858 42116 597864
rect 41326 597785 41382 597794
rect 41708 597786 42104 597802
rect 40868 597712 40920 597718
rect 40868 597654 40920 597660
rect 41340 597582 41368 597785
rect 41696 597780 42116 597786
rect 41748 597774 42064 597780
rect 41696 597722 41748 597728
rect 42064 597722 42116 597728
rect 41328 597576 41380 597582
rect 41328 597518 41380 597524
rect 41696 597576 41748 597582
rect 42064 597576 42116 597582
rect 41748 597536 42064 597564
rect 41696 597518 41748 597524
rect 42064 597518 42116 597524
rect 41142 597272 41198 597281
rect 41142 597207 41198 597216
rect 41156 595950 41184 597207
rect 42246 596864 42302 596873
rect 42246 596799 42302 596808
rect 42062 596048 42118 596057
rect 42062 595983 42118 595992
rect 41144 595944 41196 595950
rect 41144 595886 41196 595892
rect 41696 595944 41748 595950
rect 41696 595886 41748 595892
rect 41708 595785 41736 595886
rect 41694 595776 41750 595785
rect 41694 595711 41750 595720
rect 33046 595640 33102 595649
rect 33046 595575 33102 595584
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585614 31064 594351
rect 33060 587178 33088 595575
rect 35162 595232 35218 595241
rect 35162 595167 35218 595176
rect 34426 594824 34482 594833
rect 34426 594759 34482 594768
rect 34440 587217 34468 594759
rect 34426 587208 34482 587217
rect 33048 587172 33100 587178
rect 34426 587143 34482 587152
rect 33048 587114 33100 587120
rect 35176 585954 35204 595167
rect 36542 593600 36598 593609
rect 36542 593535 36598 593544
rect 36556 586430 36584 593535
rect 41694 592920 41750 592929
rect 40776 592884 40828 592890
rect 41694 592855 41696 592864
rect 40776 592826 40828 592832
rect 41748 592855 41750 592864
rect 41696 592826 41748 592832
rect 39946 590744 40002 590753
rect 39946 590679 40002 590688
rect 39580 587172 39632 587178
rect 39580 587114 39632 587120
rect 39592 586673 39620 587114
rect 39578 586664 39634 586673
rect 39578 586599 39634 586608
rect 36544 586424 36596 586430
rect 36544 586366 36596 586372
rect 39580 586424 39632 586430
rect 39580 586366 39632 586372
rect 35164 585948 35216 585954
rect 35164 585890 35216 585896
rect 39592 585857 39620 586366
rect 39578 585848 39634 585857
rect 39578 585783 39634 585792
rect 31024 585608 31076 585614
rect 31024 585550 31076 585556
rect 39672 585608 39724 585614
rect 39960 585585 39988 590679
rect 40788 589665 40816 592826
rect 41786 592376 41842 592385
rect 41786 592311 41842 592320
rect 40774 589656 40830 589665
rect 40774 589591 40830 589600
rect 41800 589529 41828 592311
rect 42076 591938 42104 595983
rect 42064 591932 42116 591938
rect 42064 591874 42116 591880
rect 41786 589520 41842 589529
rect 41786 589455 41842 589464
rect 40500 585948 40552 585954
rect 40500 585890 40552 585896
rect 39672 585550 39724 585556
rect 39946 585576 40002 585585
rect 39684 584633 39712 585550
rect 39946 585511 40002 585520
rect 40512 584769 40540 585890
rect 42260 585188 42288 596799
rect 42432 591932 42484 591938
rect 42432 591874 42484 591880
rect 42444 585449 42472 591874
rect 42720 589274 42748 598431
rect 42904 597922 42932 620986
rect 42892 597916 42944 597922
rect 42892 597858 42944 597864
rect 43180 597786 43208 620986
rect 43168 597780 43220 597786
rect 43168 597722 43220 597728
rect 42982 593192 43038 593201
rect 42982 593127 43038 593136
rect 42720 589246 42932 589274
rect 42430 585440 42486 585449
rect 42430 585375 42486 585384
rect 42260 585160 42380 585188
rect 40498 584760 40554 584769
rect 40498 584695 40554 584704
rect 42062 584760 42118 584769
rect 42118 584718 42288 584746
rect 42062 584695 42118 584704
rect 39670 584624 39726 584633
rect 39670 584559 39726 584568
rect 42260 583454 42288 584718
rect 42182 583426 42288 583454
rect 41786 582584 41842 582593
rect 41786 582519 41842 582528
rect 41800 582249 41828 582519
rect 42352 581754 42380 585160
rect 42260 581726 42380 581754
rect 42260 581618 42288 581726
rect 42182 581590 42288 581618
rect 42430 581632 42486 581641
rect 42430 581567 42486 581576
rect 42246 581496 42302 581505
rect 42246 581431 42302 581440
rect 42062 581224 42118 581233
rect 42062 581159 42118 581168
rect 42076 580961 42104 581159
rect 42260 580258 42288 581431
rect 42076 580230 42288 580258
rect 42076 579768 42104 580230
rect 42246 580136 42302 580145
rect 42246 580071 42302 580080
rect 42062 578912 42118 578921
rect 42062 578847 42118 578856
rect 42076 578544 42104 578847
rect 42260 578474 42288 580071
rect 42248 578468 42300 578474
rect 42248 578410 42300 578416
rect 42154 578232 42210 578241
rect 42154 578167 42210 578176
rect 42168 577932 42196 578167
rect 42248 577856 42300 577862
rect 42248 577798 42300 577804
rect 42260 577295 42288 577798
rect 42182 577267 42288 577295
rect 42154 577008 42210 577017
rect 42154 576943 42210 576952
rect 42168 576708 42196 576943
rect 42246 575648 42302 575657
rect 42246 575583 42302 575592
rect 42062 574696 42118 574705
rect 42062 574631 42118 574640
rect 42076 574260 42104 574631
rect 42260 573866 42288 575583
rect 42168 573838 42288 573866
rect 42168 573580 42196 573838
rect 42156 573504 42208 573510
rect 42156 573446 42208 573452
rect 42168 572968 42196 573446
rect 42444 573322 42472 581567
rect 42614 579864 42670 579873
rect 42614 579799 42670 579808
rect 42628 573510 42656 579799
rect 42904 579614 42932 589246
rect 42812 579586 42932 579614
rect 42616 573504 42668 573510
rect 42616 573446 42668 573452
rect 42352 573294 42472 573322
rect 42352 572438 42380 573294
rect 42614 572792 42670 572801
rect 42614 572727 42670 572736
rect 42168 572370 42196 572424
rect 42260 572410 42380 572438
rect 42260 572370 42288 572410
rect 42168 572342 42288 572370
rect 42628 572234 42656 572727
rect 42352 572206 42656 572234
rect 42352 571010 42380 572206
rect 42522 572112 42578 572121
rect 42522 572047 42578 572056
rect 42076 570982 42380 571010
rect 42076 570588 42104 570982
rect 41786 570208 41842 570217
rect 41786 570143 41842 570152
rect 41800 569908 41828 570143
rect 42536 569310 42564 572047
rect 42168 569242 42196 569296
rect 42260 569282 42564 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 40590 556064 40646 556073
rect 40590 555999 40646 556008
rect 40604 554810 40632 555999
rect 40866 555656 40922 555665
rect 40866 555591 40922 555600
rect 40880 554946 40908 555591
rect 41708 554946 42104 554962
rect 42812 554946 42840 579586
rect 42996 578241 43024 593127
rect 43258 591560 43314 591569
rect 43258 591495 43314 591504
rect 43272 590850 43300 591495
rect 43260 590844 43312 590850
rect 43260 590786 43312 590792
rect 43456 581233 43484 662390
rect 43824 644745 43852 688638
rect 44270 686488 44326 686497
rect 44270 686423 44326 686432
rect 44284 685874 44312 686423
rect 44468 686118 44496 729671
rect 44652 727705 44680 770034
rect 45006 763736 45062 763745
rect 45006 763671 45062 763680
rect 44822 758160 44878 758169
rect 44822 758095 44878 758104
rect 44638 727696 44694 727705
rect 44638 727631 44694 727640
rect 44456 686112 44508 686118
rect 44456 686054 44508 686060
rect 44284 685846 44496 685874
rect 44272 684548 44324 684554
rect 44272 684490 44324 684496
rect 43994 676696 44050 676705
rect 43994 676631 44050 676640
rect 44008 676462 44036 676631
rect 43996 676456 44048 676462
rect 43996 676398 44048 676404
rect 43810 644736 43866 644745
rect 43810 644671 43866 644680
rect 44284 643113 44312 684490
rect 44468 643346 44496 685846
rect 44638 679552 44694 679561
rect 44638 679487 44694 679496
rect 44652 666602 44680 679487
rect 44640 666596 44692 666602
rect 44640 666538 44692 666544
rect 44638 643512 44694 643521
rect 44638 643447 44694 643456
rect 44456 643340 44508 643346
rect 44456 643282 44508 643288
rect 44270 643104 44326 643113
rect 44270 643039 44326 643048
rect 44180 641776 44232 641782
rect 44180 641718 44232 641724
rect 43626 637800 43682 637809
rect 43626 637735 43682 637744
rect 43640 618934 43668 637735
rect 43810 634944 43866 634953
rect 43810 634879 43866 634888
rect 43824 624714 43852 634879
rect 43994 634536 44050 634545
rect 43994 634471 44050 634480
rect 43812 624708 43864 624714
rect 43812 624650 43864 624656
rect 44008 623393 44036 634471
rect 43994 623384 44050 623393
rect 43994 623319 44050 623328
rect 43628 618928 43680 618934
rect 43628 618870 43680 618876
rect 43628 609272 43680 609278
rect 43628 609214 43680 609220
rect 43442 581224 43498 581233
rect 43442 581159 43498 581168
rect 43168 581052 43220 581058
rect 43168 580994 43220 581000
rect 43180 578921 43208 580994
rect 43166 578912 43222 578921
rect 43166 578847 43222 578856
rect 42982 578232 43038 578241
rect 42982 578167 43038 578176
rect 43444 571396 43496 571402
rect 43444 571338 43496 571344
rect 43258 558512 43314 558521
rect 43258 558447 43314 558456
rect 43272 557598 43300 558447
rect 43456 558113 43484 571338
rect 43442 558104 43498 558113
rect 43442 558039 43498 558048
rect 43444 557864 43496 557870
rect 43444 557806 43496 557812
rect 43456 557705 43484 557806
rect 43442 557696 43498 557705
rect 43442 557631 43498 557640
rect 43260 557592 43312 557598
rect 43260 557534 43312 557540
rect 42982 555248 43038 555257
rect 42982 555183 43038 555192
rect 40868 554940 40920 554946
rect 40868 554882 40920 554888
rect 41696 554940 42116 554946
rect 41748 554934 42064 554940
rect 41696 554882 41748 554888
rect 42064 554882 42116 554888
rect 42800 554940 42852 554946
rect 42800 554882 42852 554888
rect 41708 554810 42104 554826
rect 40592 554804 40644 554810
rect 40592 554746 40644 554752
rect 41696 554804 42116 554810
rect 41748 554798 42064 554804
rect 41696 554746 41748 554752
rect 42064 554746 42116 554752
rect 40038 553408 40094 553417
rect 40038 553343 40094 553352
rect 40866 553408 40922 553417
rect 40866 553343 40922 553352
rect 34426 551984 34482 551993
rect 34426 551919 34482 551928
rect 31758 547496 31814 547505
rect 31758 547431 31760 547440
rect 31812 547431 31814 547440
rect 31760 547402 31812 547408
rect 34440 544406 34468 551919
rect 40052 550458 40080 553343
rect 40040 550452 40092 550458
rect 40040 550394 40092 550400
rect 38476 547460 38528 547466
rect 38476 547402 38528 547408
rect 34428 544400 34480 544406
rect 34428 544342 34480 544348
rect 38488 542230 38516 547402
rect 40880 545873 40908 553343
rect 42064 550724 42116 550730
rect 42064 550666 42116 550672
rect 41878 550624 41934 550633
rect 42076 550610 42104 550666
rect 41934 550582 42104 550610
rect 41878 550559 41934 550568
rect 41708 550458 42104 550474
rect 41696 550452 42104 550458
rect 41748 550446 42104 550452
rect 41696 550394 41748 550400
rect 42076 550390 42104 550446
rect 42064 550384 42116 550390
rect 42064 550326 42116 550332
rect 42524 550384 42576 550390
rect 42524 550326 42576 550332
rect 42154 549944 42210 549953
rect 42154 549879 42210 549888
rect 41970 549536 42026 549545
rect 41970 549471 42026 549480
rect 41142 548142 41198 548151
rect 41142 548077 41198 548086
rect 41696 548140 41748 548146
rect 41696 548082 41748 548088
rect 41708 547777 41736 548082
rect 41694 547768 41750 547777
rect 41694 547703 41750 547712
rect 40866 545864 40922 545873
rect 40866 545799 40922 545808
rect 41984 545329 42012 549471
rect 42168 545601 42196 549879
rect 42154 545592 42210 545601
rect 42154 545527 42210 545536
rect 41970 545320 42026 545329
rect 41970 545255 42026 545264
rect 39488 544400 39540 544406
rect 39488 544342 39540 544348
rect 38476 542224 38528 542230
rect 38476 542166 38528 542172
rect 39500 541929 39528 544342
rect 39764 542224 39816 542230
rect 39762 542192 39764 542201
rect 39816 542192 39818 542201
rect 39762 542127 39818 542136
rect 42338 542192 42394 542201
rect 42338 542127 42394 542136
rect 39486 541920 39542 541929
rect 39486 541855 39542 541864
rect 42062 541920 42118 541929
rect 42118 541878 42288 541906
rect 42062 541855 42118 541864
rect 42260 540682 42288 541878
rect 42168 540654 42288 540682
rect 42168 540260 42196 540654
rect 42352 539050 42380 542127
rect 42182 539022 42380 539050
rect 42536 538438 42564 550326
rect 42996 543734 43024 555183
rect 43350 551576 43406 551585
rect 43350 551511 43406 551520
rect 43168 550724 43220 550730
rect 43168 550666 43220 550672
rect 42904 543706 43024 543734
rect 42708 540728 42760 540734
rect 42708 540670 42760 540676
rect 42168 538370 42196 538424
rect 42260 538410 42564 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42338 538248 42394 538257
rect 42338 538183 42394 538192
rect 42154 537976 42210 537985
rect 42154 537911 42210 537920
rect 42168 537744 42196 537911
rect 42352 537758 42380 538183
rect 42720 537985 42748 540670
rect 42706 537976 42762 537985
rect 42706 537911 42762 537920
rect 42260 537730 42380 537758
rect 42168 536466 42196 536588
rect 42260 536466 42288 537730
rect 42432 537668 42484 537674
rect 42432 537610 42484 537616
rect 42168 536438 42288 536466
rect 42444 535378 42472 537610
rect 42708 536648 42760 536654
rect 42708 536590 42760 536596
rect 42182 535350 42472 535378
rect 42340 535288 42392 535294
rect 41786 535256 41842 535265
rect 42340 535230 42392 535236
rect 41786 535191 41842 535200
rect 41800 534752 41828 535191
rect 42352 534086 42380 535230
rect 42182 534058 42380 534086
rect 42720 534074 42748 536590
rect 42444 534046 42748 534074
rect 42444 533542 42472 534046
rect 42182 533514 42472 533542
rect 42432 533452 42484 533458
rect 42432 533394 42484 533400
rect 42246 533352 42302 533361
rect 42246 533287 42302 533296
rect 42260 531434 42288 533287
rect 42168 531406 42288 531434
rect 42168 531045 42196 531406
rect 42444 530482 42472 533394
rect 42708 532704 42760 532710
rect 42708 532646 42760 532652
rect 42260 530454 42472 530482
rect 42260 530414 42288 530454
rect 42182 530386 42288 530414
rect 42720 530346 42748 532646
rect 42904 531434 42932 543706
rect 43180 540974 43208 550666
rect 43364 549254 43392 551511
rect 43088 540946 43208 540974
rect 43272 549226 43392 549254
rect 43088 533458 43116 540946
rect 43076 533452 43128 533458
rect 43076 533394 43128 533400
rect 42812 531406 42932 531434
rect 42812 531162 42840 531406
rect 42812 531134 42932 531162
rect 42352 530318 42748 530346
rect 42352 529771 42380 530318
rect 42614 530224 42670 530233
rect 42182 529743 42380 529771
rect 42444 530182 42614 530210
rect 42444 529666 42472 530182
rect 42614 530159 42670 530168
rect 42706 529816 42762 529825
rect 42706 529751 42762 529760
rect 42352 529638 42472 529666
rect 41786 529408 41842 529417
rect 41786 529343 41842 529352
rect 41800 529205 41828 529343
rect 42352 528554 42380 529638
rect 42524 529100 42576 529106
rect 42524 529042 42576 529048
rect 42352 528526 42472 528554
rect 42168 527462 42288 527490
rect 42168 527340 42196 527462
rect 42260 527354 42288 527462
rect 42444 527354 42472 528526
rect 42260 527326 42472 527354
rect 42536 526742 42564 529042
rect 42182 526714 42564 526742
rect 42720 526091 42748 529751
rect 42182 526063 42748 526091
rect 40682 522744 40738 522753
rect 40682 522679 40738 522688
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 40696 431225 40724 522679
rect 42064 518968 42116 518974
rect 42064 518910 42116 518916
rect 42076 437474 42104 518910
rect 41708 437446 42104 437474
rect 40682 431216 40738 431225
rect 40682 431151 40738 431160
rect 41326 430536 41382 430545
rect 41326 430471 41382 430480
rect 41142 430128 41198 430137
rect 41142 430063 41198 430072
rect 40958 429482 41014 429491
rect 40958 429417 41014 429426
rect 40972 429214 41000 429417
rect 41156 429350 41184 430063
rect 41340 429622 41368 430471
rect 41708 429622 41736 437446
rect 41328 429616 41380 429622
rect 41328 429558 41380 429564
rect 41696 429616 41748 429622
rect 41696 429558 41748 429564
rect 41326 429482 41382 429491
rect 41326 429417 41382 429426
rect 41696 429480 41748 429486
rect 42064 429480 42116 429486
rect 41748 429440 42064 429468
rect 41696 429422 41748 429428
rect 42064 429422 42116 429428
rect 41144 429344 41196 429350
rect 41144 429286 41196 429292
rect 41696 429344 41748 429350
rect 42064 429344 42116 429350
rect 41748 429304 42064 429332
rect 41696 429286 41748 429292
rect 42064 429286 42116 429292
rect 40960 429208 41012 429214
rect 40960 429150 41012 429156
rect 41696 429208 41748 429214
rect 42064 429208 42116 429214
rect 41748 429168 42064 429196
rect 41696 429150 41748 429156
rect 42064 429150 42116 429156
rect 41142 428904 41198 428913
rect 41142 428839 41198 428848
rect 41156 427854 41184 428839
rect 42706 428496 42762 428505
rect 42064 428460 42116 428466
rect 42904 428466 42932 531134
rect 43272 529106 43300 549226
rect 43444 547936 43496 547942
rect 43444 547878 43496 547884
rect 43456 547777 43484 547878
rect 43442 547768 43498 547777
rect 43442 547703 43498 547712
rect 43442 547088 43498 547097
rect 43442 547023 43498 547032
rect 43456 546582 43484 547023
rect 43444 546576 43496 546582
rect 43444 546518 43496 546524
rect 43444 545148 43496 545154
rect 43444 545090 43496 545096
rect 43260 529100 43312 529106
rect 43260 529042 43312 529048
rect 43260 523728 43312 523734
rect 43260 523670 43312 523676
rect 43272 522753 43300 523670
rect 43258 522744 43314 522753
rect 43258 522679 43314 522688
rect 43260 429480 43312 429486
rect 43260 429422 43312 429428
rect 42706 428431 42762 428440
rect 42892 428460 42944 428466
rect 42064 428402 42116 428408
rect 42076 428074 42104 428402
rect 41708 428058 42104 428074
rect 41696 428052 42104 428058
rect 41748 428046 42104 428052
rect 41696 427994 41748 428000
rect 41328 427984 41380 427990
rect 41328 427926 41380 427932
rect 41340 427859 41368 427926
rect 41144 427848 41196 427854
rect 41144 427790 41196 427796
rect 41326 427850 41382 427859
rect 41326 427785 41382 427794
rect 41696 427848 41748 427854
rect 42064 427848 42116 427854
rect 41748 427808 42064 427836
rect 41696 427790 41748 427796
rect 42064 427790 42116 427796
rect 40958 427680 41014 427689
rect 40958 427615 41014 427624
rect 40972 426494 41000 427615
rect 41142 427272 41198 427281
rect 41142 427207 41198 427216
rect 41156 426630 41184 427207
rect 41708 426698 42104 426714
rect 41696 426692 42116 426698
rect 41748 426686 42064 426692
rect 41696 426634 41748 426640
rect 42064 426634 42116 426640
rect 41144 426624 41196 426630
rect 41144 426566 41196 426572
rect 40960 426488 41012 426494
rect 40960 426430 41012 426436
rect 41696 426488 41748 426494
rect 42064 426488 42116 426494
rect 41748 426448 42064 426476
rect 41696 426430 41748 426436
rect 42064 426430 42116 426436
rect 41326 426048 41382 426057
rect 41326 425983 41382 425992
rect 40774 425232 40830 425241
rect 40774 425167 40830 425176
rect 40788 421138 40816 425167
rect 41340 424386 41368 425983
rect 42720 425054 42748 428431
rect 42892 428402 42944 428408
rect 42720 425026 42932 425054
rect 42614 424416 42670 424425
rect 41328 424380 41380 424386
rect 41328 424322 41380 424328
rect 41696 424380 41748 424386
rect 41748 424340 42104 424368
rect 42614 424351 42670 424360
rect 41696 424322 41748 424328
rect 41786 421152 41842 421161
rect 40788 421110 41786 421138
rect 41786 421087 41842 421096
rect 41878 419928 41934 419937
rect 41878 419863 41934 419872
rect 41892 414882 41920 419863
rect 42076 418154 42104 424340
rect 42430 420744 42486 420753
rect 42430 420679 42486 420688
rect 42444 419558 42472 420679
rect 42432 419552 42484 419558
rect 42432 419494 42484 419500
rect 42076 418126 42472 418154
rect 41892 414854 42288 414882
rect 42062 412992 42118 413001
rect 42062 412927 42118 412936
rect 42076 412624 42104 412927
rect 42168 411346 42196 411468
rect 42260 411346 42288 414854
rect 42168 411318 42288 411346
rect 42168 410910 42288 410938
rect 42168 410788 42196 410910
rect 42260 410802 42288 410910
rect 42444 410802 42472 418126
rect 42628 413001 42656 424351
rect 42614 412992 42670 413001
rect 42614 412927 42670 412936
rect 42260 410774 42472 410802
rect 42182 410162 42472 410190
rect 42248 409828 42300 409834
rect 42248 409770 42300 409776
rect 42260 408966 42288 409770
rect 42182 408938 42288 408966
rect 42444 408474 42472 410162
rect 42432 408468 42484 408474
rect 42432 408410 42484 408416
rect 42432 408332 42484 408338
rect 42432 408274 42484 408280
rect 42444 407810 42472 408274
rect 42168 407674 42196 407796
rect 42260 407782 42472 407810
rect 42260 407674 42288 407782
rect 42168 407646 42288 407674
rect 41786 407552 41842 407561
rect 41786 407487 41842 407496
rect 41800 407116 41828 407487
rect 42432 407108 42484 407114
rect 42432 407050 42484 407056
rect 42444 406518 42472 407050
rect 42168 406450 42196 406504
rect 42260 406490 42472 406518
rect 42260 406450 42288 406490
rect 42168 406422 42288 406450
rect 42340 406020 42392 406026
rect 42168 405980 42340 406008
rect 42168 405929 42196 405980
rect 42340 405962 42392 405968
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42248 402960 42300 402966
rect 42248 402902 42300 402908
rect 42260 402815 42288 402902
rect 42182 402787 42288 402815
rect 42432 402552 42484 402558
rect 42432 402494 42484 402500
rect 42444 402166 42472 402494
rect 42182 402138 42472 402166
rect 41786 401976 41842 401985
rect 41786 401911 41842 401920
rect 41800 401608 41828 401911
rect 42432 400172 42484 400178
rect 42432 400114 42484 400120
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 42444 399135 42472 400114
rect 42182 399107 42472 399135
rect 41878 398848 41934 398857
rect 41878 398783 41934 398792
rect 41892 398480 41920 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 35808 387592 35860 387598
rect 35438 387560 35494 387569
rect 35438 387495 35494 387504
rect 35806 387560 35808 387569
rect 41696 387592 41748 387598
rect 35860 387560 35862 387569
rect 41748 387540 42104 387546
rect 41696 387534 42104 387540
rect 41708 387530 42104 387534
rect 41708 387524 42116 387530
rect 41708 387518 42064 387524
rect 35806 387495 35862 387504
rect 35452 386442 35480 387495
rect 42064 387466 42116 387472
rect 39946 387152 40002 387161
rect 39946 387087 40002 387096
rect 39960 386850 39988 387087
rect 35624 386844 35676 386850
rect 35624 386786 35676 386792
rect 39948 386844 40000 386850
rect 39948 386786 40000 386792
rect 35440 386436 35492 386442
rect 35440 386378 35492 386384
rect 35636 386345 35664 386786
rect 35806 386744 35862 386753
rect 35806 386679 35862 386688
rect 40130 386744 40186 386753
rect 40130 386679 40132 386688
rect 35820 386578 35848 386679
rect 40184 386679 40186 386688
rect 40132 386650 40184 386656
rect 35808 386572 35860 386578
rect 35808 386514 35860 386520
rect 41696 386504 41748 386510
rect 42064 386504 42116 386510
rect 41748 386452 42064 386458
rect 41696 386446 42116 386452
rect 41708 386430 42104 386446
rect 35622 386336 35678 386345
rect 35622 386271 35678 386280
rect 35346 385928 35402 385937
rect 35346 385863 35402 385872
rect 35360 385082 35388 385863
rect 35530 385520 35586 385529
rect 35530 385455 35586 385464
rect 35806 385520 35862 385529
rect 35806 385455 35808 385464
rect 35544 385218 35572 385455
rect 35860 385455 35862 385464
rect 40132 385484 40184 385490
rect 35808 385426 35860 385432
rect 40132 385426 40184 385432
rect 35532 385212 35584 385218
rect 35532 385154 35584 385160
rect 39946 385112 40002 385121
rect 35348 385076 35400 385082
rect 39946 385047 40002 385056
rect 35348 385018 35400 385024
rect 35622 384704 35678 384713
rect 35622 384639 35678 384648
rect 35636 383858 35664 384639
rect 35806 384296 35862 384305
rect 35806 384231 35862 384240
rect 35820 384130 35848 384231
rect 35808 384124 35860 384130
rect 35808 384066 35860 384072
rect 39764 384124 39816 384130
rect 39764 384066 39816 384072
rect 39776 383897 39804 384066
rect 39960 383926 39988 385047
rect 39948 383920 40000 383926
rect 35806 383888 35862 383897
rect 35624 383852 35676 383858
rect 35806 383823 35862 383832
rect 39762 383888 39818 383897
rect 39948 383862 40000 383868
rect 39762 383823 39818 383832
rect 35624 383794 35676 383800
rect 35820 383722 35848 383823
rect 35808 383716 35860 383722
rect 35808 383658 35860 383664
rect 40144 383489 40172 385426
rect 42904 385286 42932 425026
rect 43074 421560 43130 421569
rect 43074 421495 43130 421504
rect 43088 407114 43116 421495
rect 43076 407108 43128 407114
rect 43076 407050 43128 407056
rect 43272 387161 43300 429422
rect 43456 429350 43484 545090
rect 43640 540734 43668 609214
rect 43810 600944 43866 600953
rect 43810 600879 43866 600888
rect 43824 600438 43852 600879
rect 43812 600432 43864 600438
rect 43812 600374 43864 600380
rect 44192 599729 44220 641718
rect 44362 638208 44418 638217
rect 44362 638143 44418 638152
rect 44376 613630 44404 638143
rect 44652 621014 44680 643447
rect 44560 620986 44680 621014
rect 44364 613624 44416 613630
rect 44364 613566 44416 613572
rect 44560 600545 44588 620986
rect 44546 600536 44602 600545
rect 44546 600471 44602 600480
rect 44362 600128 44418 600137
rect 44362 600063 44418 600072
rect 44178 599720 44234 599729
rect 44178 599655 44234 599664
rect 44376 599536 44404 600063
rect 44284 599508 44404 599536
rect 43812 597576 43864 597582
rect 43812 597518 43864 597524
rect 43824 554849 43852 597518
rect 44284 557297 44312 599508
rect 44456 599004 44508 599010
rect 44456 598946 44508 598952
rect 44270 557288 44326 557297
rect 44270 557223 44326 557232
rect 44468 556481 44496 598946
rect 44638 591968 44694 591977
rect 44638 591903 44694 591912
rect 44652 581058 44680 591903
rect 44640 581052 44692 581058
rect 44640 580994 44692 581000
rect 44638 556880 44694 556889
rect 44638 556815 44694 556824
rect 44454 556472 44510 556481
rect 44454 556407 44510 556416
rect 43810 554840 43866 554849
rect 43810 554775 43866 554784
rect 44364 554804 44416 554810
rect 44364 554746 44416 554752
rect 43810 554432 43866 554441
rect 43810 554367 43866 554376
rect 43628 540728 43680 540734
rect 43628 540670 43680 540676
rect 43824 537010 43852 554367
rect 43994 549128 44050 549137
rect 43994 549063 44050 549072
rect 44008 540974 44036 549063
rect 44178 548720 44234 548729
rect 44178 548655 44234 548664
rect 44192 540974 44220 548655
rect 44376 543734 44404 554746
rect 44652 550634 44680 556815
rect 43548 536982 43852 537010
rect 43916 540946 44036 540974
rect 44100 540946 44220 540974
rect 44284 543706 44404 543734
rect 44560 550606 44680 550634
rect 43548 531314 43576 536982
rect 43916 535294 43944 540946
rect 44100 537674 44128 540946
rect 44088 537668 44140 537674
rect 44088 537610 44140 537616
rect 43904 535288 43956 535294
rect 43904 535230 43956 535236
rect 43548 531286 43852 531314
rect 43628 491972 43680 491978
rect 43628 491914 43680 491920
rect 43444 429344 43496 429350
rect 43444 429286 43496 429292
rect 43442 422784 43498 422793
rect 43442 422719 43498 422728
rect 43456 409834 43484 422719
rect 43444 409828 43496 409834
rect 43444 409770 43496 409776
rect 43444 401668 43496 401674
rect 43444 401610 43496 401616
rect 43258 387152 43314 387161
rect 43258 387087 43314 387096
rect 41696 385280 41748 385286
rect 42064 385280 42116 385286
rect 41748 385228 42064 385234
rect 41696 385222 42116 385228
rect 42892 385280 42944 385286
rect 42892 385222 42944 385228
rect 41708 385206 42104 385222
rect 41708 385082 42104 385098
rect 41696 385076 42116 385082
rect 41748 385070 42064 385076
rect 41696 385018 41748 385024
rect 42064 385018 42116 385024
rect 42798 383888 42854 383897
rect 42798 383823 42854 383832
rect 42064 383784 42116 383790
rect 41708 383732 42064 383738
rect 41708 383726 42116 383732
rect 41708 383722 42104 383726
rect 41696 383716 42104 383722
rect 41748 383710 42104 383716
rect 41696 383658 41748 383664
rect 35254 383480 35310 383489
rect 35254 383415 35310 383424
rect 40130 383480 40186 383489
rect 40130 383415 40186 383424
rect 35268 382294 35296 383415
rect 35438 383072 35494 383081
rect 35438 383007 35494 383016
rect 35452 382430 35480 383007
rect 35808 382696 35860 382702
rect 35806 382664 35808 382673
rect 41696 382696 41748 382702
rect 35860 382664 35862 382673
rect 41696 382638 41748 382644
rect 35806 382599 35862 382608
rect 35624 382560 35676 382566
rect 35624 382502 35676 382508
rect 40224 382560 40276 382566
rect 40224 382502 40276 382508
rect 35440 382424 35492 382430
rect 35440 382366 35492 382372
rect 35256 382288 35308 382294
rect 35636 382265 35664 382502
rect 40040 382424 40092 382430
rect 40040 382366 40092 382372
rect 39028 382288 39080 382294
rect 35256 382230 35308 382236
rect 35622 382256 35678 382265
rect 40052 382265 40080 382366
rect 39028 382230 39080 382236
rect 40038 382256 40094 382265
rect 35622 382191 35678 382200
rect 39040 381857 39068 382230
rect 40038 382191 40094 382200
rect 35622 381848 35678 381857
rect 35622 381783 35678 381792
rect 39026 381848 39082 381857
rect 39026 381783 39082 381792
rect 32402 381440 32458 381449
rect 32402 381375 32458 381384
rect 28814 376544 28870 376553
rect 28814 376479 28870 376488
rect 28828 375902 28856 376479
rect 28816 375896 28868 375902
rect 28816 375838 28868 375844
rect 32416 371890 32444 381375
rect 35636 381070 35664 381783
rect 35808 381200 35860 381206
rect 35808 381142 35860 381148
rect 35624 381064 35676 381070
rect 35820 381041 35848 381142
rect 40040 381064 40092 381070
rect 35624 381006 35676 381012
rect 35806 381032 35862 381041
rect 40040 381006 40092 381012
rect 35806 380967 35862 380976
rect 35622 380624 35678 380633
rect 35622 380559 35678 380568
rect 35636 379710 35664 380559
rect 40052 380225 40080 381006
rect 35806 380216 35862 380225
rect 35806 380151 35862 380160
rect 40038 380216 40094 380225
rect 40038 380151 40094 380160
rect 35820 379982 35848 380151
rect 35808 379976 35860 379982
rect 35808 379918 35860 379924
rect 35806 379808 35862 379817
rect 35806 379743 35862 379752
rect 35624 379704 35676 379710
rect 35624 379646 35676 379652
rect 35820 379574 35848 379743
rect 39948 379704 40000 379710
rect 39948 379646 40000 379652
rect 35808 379568 35860 379574
rect 35808 379510 35860 379516
rect 39580 379568 39632 379574
rect 39580 379510 39632 379516
rect 35806 378992 35862 379001
rect 35806 378927 35862 378936
rect 35820 378350 35848 378927
rect 35808 378344 35860 378350
rect 35808 378286 35860 378292
rect 35622 377768 35678 377777
rect 35622 377703 35678 377712
rect 35636 377058 35664 377703
rect 39592 377369 39620 379510
rect 39960 377777 39988 379646
rect 40236 379001 40264 382502
rect 41420 381200 41472 381206
rect 41420 381142 41472 381148
rect 41432 381041 41460 381142
rect 41418 381032 41474 381041
rect 41418 380967 41474 380976
rect 41512 379976 41564 379982
rect 41512 379918 41564 379924
rect 40222 378992 40278 379001
rect 40222 378927 40278 378936
rect 41524 378593 41552 379918
rect 41708 379514 41736 382638
rect 41708 379486 42472 379514
rect 41510 378584 41566 378593
rect 41510 378519 41566 378528
rect 41236 378344 41288 378350
rect 41236 378286 41288 378292
rect 41248 378185 41276 378286
rect 41234 378176 41290 378185
rect 41234 378111 41290 378120
rect 39946 377768 40002 377777
rect 39946 377703 40002 377712
rect 35806 377360 35862 377369
rect 35806 377295 35862 377304
rect 39578 377360 39634 377369
rect 39578 377295 39634 377304
rect 35624 377052 35676 377058
rect 35624 376994 35676 377000
rect 35820 376786 35848 377295
rect 41696 376984 41748 376990
rect 41694 376952 41696 376961
rect 41748 376952 41750 376961
rect 41694 376887 41750 376896
rect 42064 376848 42116 376854
rect 41708 376796 42064 376802
rect 41708 376790 42116 376796
rect 41708 376786 42104 376790
rect 35808 376780 35860 376786
rect 35808 376722 35860 376728
rect 41696 376780 42104 376786
rect 41748 376774 42104 376780
rect 41696 376722 41748 376728
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 33784 375896 33836 375902
rect 33784 375838 33836 375844
rect 33796 373318 33824 375838
rect 35820 375630 35848 376071
rect 35808 375624 35860 375630
rect 35808 375566 35860 375572
rect 41696 375624 41748 375630
rect 41748 375572 42104 375578
rect 41696 375566 42104 375572
rect 41708 375562 42104 375566
rect 41708 375556 42116 375562
rect 41708 375550 42064 375556
rect 42064 375498 42116 375504
rect 33784 373312 33836 373318
rect 33784 373254 33836 373260
rect 41696 373312 41748 373318
rect 41696 373254 41748 373260
rect 41708 372858 41736 373254
rect 41708 372830 42288 372858
rect 32404 371884 32456 371890
rect 32404 371826 32456 371832
rect 41696 371884 41748 371890
rect 41696 371826 41748 371832
rect 41708 371770 41736 371826
rect 41708 371754 42104 371770
rect 41708 371748 42116 371754
rect 41708 371742 42064 371748
rect 42064 371690 42116 371696
rect 42062 369744 42118 369753
rect 42062 369679 42118 369688
rect 42076 369444 42104 369679
rect 42260 368263 42288 372830
rect 42182 368235 42288 368263
rect 42444 367622 42472 379486
rect 42616 371748 42668 371754
rect 42616 371690 42668 371696
rect 42182 367594 42472 367622
rect 42182 366947 42472 366975
rect 41800 365673 41828 365772
rect 42248 365696 42300 365702
rect 41786 365664 41842 365673
rect 42248 365638 42300 365644
rect 41786 365599 41842 365608
rect 42260 364698 42288 365638
rect 42168 364670 42288 364698
rect 42168 364548 42196 364670
rect 42444 364290 42472 366947
rect 42628 364334 42656 371690
rect 42352 364274 42472 364290
rect 42340 364268 42472 364274
rect 42392 364262 42472 364268
rect 42536 364306 42656 364334
rect 42340 364210 42392 364216
rect 42340 364132 42392 364138
rect 42340 364074 42392 364080
rect 42352 363950 42380 364074
rect 42182 363922 42380 363950
rect 41786 363760 41842 363769
rect 41786 363695 41842 363704
rect 41800 363256 41828 363695
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42536 362726 42564 364306
rect 42260 362698 42564 362726
rect 41786 360632 41842 360641
rect 41786 360567 41842 360576
rect 41800 360264 41828 360567
rect 42432 360188 42484 360194
rect 42432 360130 42484 360136
rect 42156 359984 42208 359990
rect 42156 359926 42208 359932
rect 42168 359584 42196 359926
rect 42444 358986 42472 360130
rect 42182 358958 42472 358986
rect 41878 358728 41934 358737
rect 41878 358663 41934 358672
rect 41892 358428 41920 358663
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42432 356040 42484 356046
rect 42432 355982 42484 355988
rect 42444 355926 42472 355982
rect 42182 355898 42472 355926
rect 41970 355736 42026 355745
rect 41970 355671 42026 355680
rect 41984 355300 42012 355671
rect 39210 345944 39266 345953
rect 39210 345879 39266 345888
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 35806 344312 35862 344321
rect 35806 344247 35862 344256
rect 35820 344078 35848 344247
rect 39224 344078 39252 345879
rect 35808 344072 35860 344078
rect 35808 344014 35860 344020
rect 39212 344072 39264 344078
rect 39212 344014 39264 344020
rect 35622 343904 35678 343913
rect 41708 343874 42104 343890
rect 35622 343839 35678 343848
rect 41696 343868 42116 343874
rect 35636 343670 35664 343839
rect 41748 343862 42064 343868
rect 41696 343810 41748 343816
rect 42064 343810 42116 343816
rect 35808 343800 35860 343806
rect 35808 343742 35860 343748
rect 35624 343664 35676 343670
rect 35624 343606 35676 343612
rect 35820 343505 35848 343742
rect 41696 343664 41748 343670
rect 42064 343664 42116 343670
rect 41748 343612 42064 343618
rect 41696 343606 42116 343612
rect 41708 343590 42104 343606
rect 35806 343496 35862 343505
rect 35806 343431 35862 343440
rect 35622 343088 35678 343097
rect 35622 343023 35678 343032
rect 40038 343088 40094 343097
rect 40038 343023 40094 343032
rect 35636 342446 35664 343023
rect 35808 342712 35860 342718
rect 35806 342680 35808 342689
rect 35860 342680 35862 342689
rect 35806 342615 35862 342624
rect 40052 342446 40080 343023
rect 40316 342712 40368 342718
rect 40314 342680 40316 342689
rect 40368 342680 40370 342689
rect 40314 342615 40370 342624
rect 35624 342440 35676 342446
rect 35624 342382 35676 342388
rect 40040 342440 40092 342446
rect 40040 342382 40092 342388
rect 35624 342304 35676 342310
rect 35622 342272 35624 342281
rect 41696 342304 41748 342310
rect 35676 342272 35678 342281
rect 42064 342304 42116 342310
rect 41748 342252 42064 342258
rect 41696 342246 42116 342252
rect 41708 342230 42104 342246
rect 35622 342207 35678 342216
rect 35806 341864 35862 341873
rect 35806 341799 35862 341808
rect 35820 341494 35848 341799
rect 42812 341578 42840 383823
rect 42982 377768 43038 377777
rect 42982 377703 43038 377712
rect 42996 356046 43024 377703
rect 43258 377360 43314 377369
rect 43258 377295 43314 377304
rect 43272 359990 43300 377295
rect 43260 359984 43312 359990
rect 43260 359926 43312 359932
rect 42984 356040 43036 356046
rect 42984 355982 43036 355988
rect 43258 342680 43314 342689
rect 43258 342615 43314 342624
rect 42720 341550 42840 341578
rect 35808 341488 35860 341494
rect 35346 341456 35402 341465
rect 35346 341391 35402 341400
rect 35622 341456 35678 341465
rect 35808 341430 35860 341436
rect 41696 341488 41748 341494
rect 41748 341436 42104 341442
rect 41696 341430 42104 341436
rect 41708 341426 42104 341430
rect 41708 341420 42116 341426
rect 41708 341414 42064 341420
rect 35622 341391 35678 341400
rect 35360 341222 35388 341391
rect 35348 341216 35400 341222
rect 35348 341158 35400 341164
rect 35636 340950 35664 341391
rect 42064 341362 42116 341368
rect 41708 341290 42104 341306
rect 42720 341290 42748 341550
rect 42892 341420 42944 341426
rect 42892 341362 42944 341368
rect 41696 341284 42116 341290
rect 41748 341278 42064 341284
rect 41696 341226 41748 341232
rect 42064 341226 42116 341232
rect 42708 341284 42760 341290
rect 42708 341226 42760 341232
rect 35808 341080 35860 341086
rect 35806 341048 35808 341057
rect 41696 341080 41748 341086
rect 35860 341048 35862 341057
rect 42064 341080 42116 341086
rect 41748 341028 42064 341034
rect 41696 341022 42116 341028
rect 41708 341006 42104 341022
rect 35806 340983 35862 340992
rect 35624 340944 35676 340950
rect 35624 340886 35676 340892
rect 41696 340944 41748 340950
rect 42064 340944 42116 340950
rect 41748 340892 42064 340898
rect 41696 340886 42116 340892
rect 41708 340870 42104 340886
rect 35806 340232 35862 340241
rect 35806 340167 35862 340176
rect 35820 339658 35848 340167
rect 35808 339652 35860 339658
rect 35808 339594 35860 339600
rect 41420 339652 41472 339658
rect 41420 339594 41472 339600
rect 41432 339017 41460 339594
rect 35622 339008 35678 339017
rect 35622 338943 35678 338952
rect 41418 339008 41474 339017
rect 41418 338943 41474 338952
rect 35636 338162 35664 338943
rect 41786 338736 41842 338745
rect 41524 338694 41786 338722
rect 35806 338600 35862 338609
rect 35806 338535 35862 338544
rect 35820 338434 35848 338535
rect 35808 338428 35860 338434
rect 35808 338370 35860 338376
rect 41524 338162 41552 338694
rect 41786 338671 41842 338680
rect 41696 338428 41748 338434
rect 41696 338370 41748 338376
rect 41708 338201 41736 338370
rect 41694 338192 41750 338201
rect 35624 338156 35676 338162
rect 35624 338098 35676 338104
rect 41512 338156 41564 338162
rect 41694 338127 41750 338136
rect 41512 338098 41564 338104
rect 35806 337784 35862 337793
rect 35806 337719 35862 337728
rect 35820 337142 35848 337719
rect 35808 337136 35860 337142
rect 35808 337078 35860 337084
rect 39856 337136 39908 337142
rect 39856 337078 39908 337084
rect 35530 336968 35586 336977
rect 35530 336903 35586 336912
rect 35806 336968 35862 336977
rect 35806 336903 35808 336912
rect 35544 336802 35572 336903
rect 35860 336903 35862 336912
rect 35808 336874 35860 336880
rect 35532 336796 35584 336802
rect 35532 336738 35584 336744
rect 35622 335744 35678 335753
rect 35622 335679 35678 335688
rect 35636 335374 35664 335679
rect 35808 335640 35860 335646
rect 35806 335608 35808 335617
rect 35860 335608 35862 335617
rect 35806 335543 35862 335552
rect 35624 335368 35676 335374
rect 35624 335310 35676 335316
rect 35622 334928 35678 334937
rect 35622 334863 35678 334872
rect 35438 334520 35494 334529
rect 35438 334455 35494 334464
rect 35452 334150 35480 334455
rect 35636 334422 35664 334863
rect 35806 334520 35862 334529
rect 35806 334455 35862 334464
rect 35624 334416 35676 334422
rect 35624 334358 35676 334364
rect 35440 334144 35492 334150
rect 35440 334086 35492 334092
rect 35820 334014 35848 334455
rect 35808 334008 35860 334014
rect 35808 333950 35860 333956
rect 35806 333296 35862 333305
rect 35806 333231 35862 333240
rect 35820 333062 35848 333231
rect 35808 333056 35860 333062
rect 35808 332998 35860 333004
rect 39304 332920 39356 332926
rect 35806 332888 35862 332897
rect 39868 332897 39896 337078
rect 40316 336932 40368 336938
rect 40316 336874 40368 336880
rect 40328 335753 40356 336874
rect 41708 336802 42104 336818
rect 41696 336796 42116 336802
rect 41748 336790 42064 336796
rect 41696 336738 41748 336744
rect 42064 336738 42116 336744
rect 40314 335744 40370 335753
rect 40314 335679 40370 335688
rect 40868 335640 40920 335646
rect 40868 335582 40920 335588
rect 40224 335368 40276 335374
rect 40224 335310 40276 335316
rect 40236 334937 40264 335310
rect 40222 334928 40278 334937
rect 40222 334863 40278 334872
rect 40316 334416 40368 334422
rect 40316 334358 40368 334364
rect 40132 334144 40184 334150
rect 40132 334086 40184 334092
rect 39304 332862 39356 332868
rect 39854 332888 39910 332897
rect 35806 332823 35862 332832
rect 35820 332654 35848 332823
rect 35808 332648 35860 332654
rect 35808 332590 35860 332596
rect 39316 330721 39344 332862
rect 39854 332823 39910 332832
rect 40144 331265 40172 334086
rect 40328 333713 40356 334358
rect 40314 333704 40370 333713
rect 40314 333639 40370 333648
rect 40880 332489 40908 335582
rect 41696 334008 41748 334014
rect 42064 334008 42116 334014
rect 41748 333956 42064 333962
rect 41696 333950 42116 333956
rect 41708 333934 42104 333950
rect 41696 332648 41748 332654
rect 42064 332648 42116 332654
rect 41748 332596 42064 332602
rect 41696 332590 42116 332596
rect 41708 332574 42104 332590
rect 40866 332480 40922 332489
rect 40866 332415 40922 332424
rect 40130 331256 40186 331265
rect 40130 331191 40186 331200
rect 39302 330712 39358 330721
rect 39302 330647 39358 330656
rect 42432 327072 42484 327078
rect 42432 327014 42484 327020
rect 42444 326278 42472 327014
rect 42168 326210 42196 326264
rect 42260 326250 42472 326278
rect 42260 326210 42288 326250
rect 42168 326182 42288 326210
rect 42432 325372 42484 325378
rect 42432 325314 42484 325320
rect 42444 325054 42472 325314
rect 42182 325026 42472 325054
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42182 323734 42472 323762
rect 41786 322824 41842 322833
rect 41786 322759 41842 322768
rect 41800 322592 41828 322759
rect 42444 321570 42472 323734
rect 42432 321564 42484 321570
rect 42432 321506 42484 321512
rect 42182 321354 42656 321382
rect 42432 321292 42484 321298
rect 42432 321234 42484 321240
rect 42444 320739 42472 321234
rect 42182 320711 42472 320739
rect 42182 320062 42472 320090
rect 42248 320000 42300 320006
rect 42248 319942 42300 319948
rect 42260 319546 42288 319942
rect 42182 319518 42288 319546
rect 42444 319190 42472 320062
rect 42432 319184 42484 319190
rect 42432 319126 42484 319132
rect 42628 318782 42656 321354
rect 42616 318776 42668 318782
rect 42616 318718 42668 318724
rect 42432 317416 42484 317422
rect 42432 317358 42484 317364
rect 42444 317059 42472 317358
rect 42182 317031 42472 317059
rect 42432 316940 42484 316946
rect 42432 316882 42484 316888
rect 42444 316418 42472 316882
rect 42182 316390 42472 316418
rect 42432 315920 42484 315926
rect 42432 315862 42484 315868
rect 42444 315771 42472 315862
rect 42182 315743 42472 315771
rect 41786 315616 41842 315625
rect 41786 315551 41842 315560
rect 41800 315180 41828 315551
rect 41786 313712 41842 313721
rect 41786 313647 41842 313656
rect 41800 313344 41828 313647
rect 41786 313032 41842 313041
rect 41786 312967 41842 312976
rect 41800 312732 41828 312967
rect 42168 312174 42288 312202
rect 42168 312052 42196 312174
rect 42260 312066 42288 312174
rect 42260 312038 42472 312066
rect 42444 310486 42472 312038
rect 42432 310480 42484 310486
rect 42432 310422 42484 310428
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 40958 300520 41014 300529
rect 40958 300455 41014 300464
rect 40972 299538 41000 300455
rect 41142 300112 41198 300121
rect 41142 300047 41198 300056
rect 41156 299674 41184 300047
rect 41696 299736 41748 299742
rect 42064 299736 42116 299742
rect 41748 299684 42064 299690
rect 41696 299678 42116 299684
rect 41144 299668 41196 299674
rect 41708 299662 42104 299678
rect 41144 299610 41196 299616
rect 40960 299532 41012 299538
rect 40960 299474 41012 299480
rect 41696 299532 41748 299538
rect 42064 299532 42116 299538
rect 41748 299492 42064 299520
rect 41696 299474 41748 299480
rect 42064 299474 42116 299480
rect 41142 299296 41198 299305
rect 41142 299231 41198 299240
rect 40958 298480 41014 298489
rect 40958 298415 41014 298424
rect 40972 298314 41000 298415
rect 41156 298314 41184 299231
rect 42706 298888 42762 298897
rect 42706 298823 42762 298832
rect 41696 298376 41748 298382
rect 42064 298376 42116 298382
rect 41748 298324 42064 298330
rect 41696 298318 42116 298324
rect 40960 298308 41012 298314
rect 40960 298250 41012 298256
rect 41144 298308 41196 298314
rect 41708 298302 42104 298318
rect 41144 298250 41196 298256
rect 42064 298240 42116 298246
rect 41708 298188 42064 298194
rect 41708 298182 42116 298188
rect 41708 298178 42104 298182
rect 41696 298172 42104 298178
rect 41748 298166 42104 298172
rect 41696 298114 41748 298120
rect 40958 298072 41014 298081
rect 40958 298007 41014 298016
rect 40972 296750 41000 298007
rect 41142 297664 41198 297673
rect 41142 297599 41198 297608
rect 41156 296886 41184 297599
rect 41708 296954 42104 296970
rect 41696 296948 42116 296954
rect 41748 296942 42064 296948
rect 41696 296890 41748 296896
rect 42064 296890 42116 296896
rect 41144 296880 41196 296886
rect 41144 296822 41196 296828
rect 40960 296744 41012 296750
rect 40960 296686 41012 296692
rect 41696 296744 41748 296750
rect 42064 296744 42116 296750
rect 41748 296704 42064 296732
rect 41696 296686 41748 296692
rect 42064 296686 42116 296692
rect 40774 295624 40830 295633
rect 40774 295559 40830 295568
rect 37922 294808 37978 294817
rect 37922 294743 37978 294752
rect 37936 285054 37964 294743
rect 40500 292597 40552 292602
rect 40498 292596 40554 292597
rect 40498 292588 40500 292596
rect 40552 292588 40554 292596
rect 40788 292574 40816 295559
rect 41786 295216 41842 295225
rect 41786 295151 41842 295160
rect 41800 294545 41828 295151
rect 41786 294536 41842 294545
rect 41786 294471 41842 294480
rect 41326 294400 41382 294409
rect 41326 294335 41382 294344
rect 41340 294030 41368 294335
rect 41328 294024 41380 294030
rect 41328 293966 41380 293972
rect 41696 294024 41748 294030
rect 42064 294024 42116 294030
rect 41748 293984 42064 294012
rect 41696 293966 41748 293972
rect 42064 293966 42116 293972
rect 41786 293584 41842 293593
rect 41616 293542 41786 293570
rect 41616 292602 41644 293542
rect 41786 293519 41842 293528
rect 41604 292596 41656 292602
rect 40788 292546 41368 292574
rect 40498 292523 40554 292532
rect 41340 292074 41368 292546
rect 41604 292538 41656 292544
rect 41786 292088 41842 292097
rect 41340 292046 41786 292074
rect 41786 292023 41842 292032
rect 41142 291952 41198 291961
rect 41142 291887 41198 291896
rect 41156 291242 41184 291887
rect 41144 291236 41196 291242
rect 41144 291178 41196 291184
rect 41696 291236 41748 291242
rect 42064 291236 42116 291242
rect 41748 291196 42064 291224
rect 41696 291178 41748 291184
rect 42064 291178 42116 291184
rect 40958 291136 41014 291145
rect 40958 291071 41014 291080
rect 40972 289882 41000 291071
rect 41142 290320 41198 290329
rect 41142 290255 41198 290264
rect 40960 289876 41012 289882
rect 40960 289818 41012 289824
rect 41156 289134 41184 290255
rect 42064 290080 42116 290086
rect 41340 290028 42064 290034
rect 41340 290022 42116 290028
rect 41340 290006 42104 290022
rect 41340 289814 41368 290006
rect 41696 289876 41748 289882
rect 42064 289876 42116 289882
rect 41748 289836 42064 289864
rect 41696 289818 41748 289824
rect 42064 289818 42116 289824
rect 42720 289814 42748 298823
rect 42904 298382 42932 341362
rect 43074 332480 43130 332489
rect 43074 332415 43130 332424
rect 43088 317422 43116 332415
rect 43076 317416 43128 317422
rect 43076 317358 43128 317364
rect 43074 301336 43130 301345
rect 43074 301271 43130 301280
rect 43088 301034 43116 301271
rect 43076 301028 43128 301034
rect 43076 300970 43128 300976
rect 43272 299742 43300 342615
rect 43260 299736 43312 299742
rect 43074 299704 43130 299713
rect 43260 299678 43312 299684
rect 43074 299639 43130 299648
rect 43088 299474 43116 299639
rect 43088 299446 43208 299474
rect 42892 298376 42944 298382
rect 42892 298318 42944 298324
rect 42982 293176 43038 293185
rect 42982 293111 43038 293120
rect 41340 289786 41552 289814
rect 42720 289786 42840 289814
rect 41524 289762 41552 289786
rect 41524 289734 42012 289762
rect 41984 289649 42012 289734
rect 41970 289640 42026 289649
rect 41970 289575 42026 289584
rect 41144 289128 41196 289134
rect 41144 289070 41196 289076
rect 41696 289128 41748 289134
rect 41696 289070 41748 289076
rect 41708 288946 41736 289070
rect 41708 288918 42380 288946
rect 37924 285048 37976 285054
rect 37924 284990 37976 284996
rect 41696 285048 41748 285054
rect 41748 284996 42288 285002
rect 41696 284990 42288 284996
rect 41708 284974 42288 284990
rect 42260 283059 42288 284974
rect 42182 283031 42288 283059
rect 42352 281874 42380 288918
rect 42182 281846 42380 281874
rect 42432 281512 42484 281518
rect 41970 281480 42026 281489
rect 42432 281454 42484 281460
rect 41970 281415 42026 281424
rect 41984 281180 42012 281415
rect 42444 280582 42472 281454
rect 42182 280554 42472 280582
rect 42432 280152 42484 280158
rect 42432 280094 42484 280100
rect 42168 279398 42288 279426
rect 42168 279344 42196 279398
rect 42260 279358 42288 279398
rect 42444 279358 42472 280094
rect 42260 279330 42472 279358
rect 42522 278760 42578 278769
rect 42522 278695 42578 278704
rect 42168 277930 42196 278188
rect 42168 277902 42288 277930
rect 41800 277409 41828 277508
rect 41786 277400 41842 277409
rect 42260 277394 42288 277902
rect 42260 277366 42380 277394
rect 41786 277335 41842 277344
rect 42352 277234 42380 277366
rect 42340 277228 42392 277234
rect 42340 277170 42392 277176
rect 42340 277092 42392 277098
rect 42340 277034 42392 277040
rect 42352 276910 42380 277034
rect 42182 276882 42380 276910
rect 42168 276298 42196 276352
rect 42168 276270 42288 276298
rect 42260 274650 42288 276270
rect 42248 274644 42300 274650
rect 42248 274586 42300 274592
rect 42536 273850 42564 278695
rect 42182 273822 42564 273850
rect 41800 273057 41828 273224
rect 42432 273216 42484 273222
rect 42432 273158 42484 273164
rect 41786 273048 41842 273057
rect 41786 272983 41842 272992
rect 42444 272558 42472 273158
rect 42182 272530 42472 272558
rect 41786 272368 41842 272377
rect 41786 272303 41842 272312
rect 41800 272000 41828 272303
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 42182 269507 42656 269535
rect 42432 269068 42484 269074
rect 42432 269010 42484 269016
rect 42444 268886 42472 269010
rect 42182 268858 42472 268886
rect 42628 267714 42656 269507
rect 42616 267708 42668 267714
rect 42616 267650 42668 267656
rect 39946 259584 40002 259593
rect 39946 259519 40002 259528
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 39960 258262 39988 259519
rect 35808 258256 35860 258262
rect 35808 258198 35860 258204
rect 39948 258256 40000 258262
rect 39948 258198 40000 258204
rect 35820 258097 35848 258198
rect 35806 258088 35862 258097
rect 35806 258023 35862 258032
rect 35622 257544 35678 257553
rect 35622 257479 35678 257488
rect 39578 257544 39634 257553
rect 39578 257479 39634 257488
rect 35438 257136 35494 257145
rect 35438 257071 35494 257080
rect 35452 256766 35480 257071
rect 35636 256902 35664 257479
rect 39592 257174 39620 257479
rect 35808 257168 35860 257174
rect 35806 257136 35808 257145
rect 39580 257168 39632 257174
rect 35860 257136 35862 257145
rect 39580 257110 39632 257116
rect 35806 257071 35862 257080
rect 42064 257032 42116 257038
rect 41708 256980 42064 256986
rect 41708 256974 42116 256980
rect 41708 256970 42104 256974
rect 41696 256964 42104 256970
rect 41748 256958 42104 256964
rect 41696 256906 41748 256912
rect 35624 256896 35676 256902
rect 35624 256838 35676 256844
rect 35440 256760 35492 256766
rect 35440 256702 35492 256708
rect 41696 256760 41748 256766
rect 42064 256760 42116 256766
rect 41748 256708 42064 256714
rect 41696 256702 42116 256708
rect 41708 256686 42104 256702
rect 35438 256320 35494 256329
rect 35438 256255 35494 256264
rect 35452 255338 35480 256255
rect 35622 255912 35678 255921
rect 35622 255847 35678 255856
rect 35636 255474 35664 255847
rect 35808 255740 35860 255746
rect 35808 255682 35860 255688
rect 40408 255740 40460 255746
rect 40408 255682 40460 255688
rect 35820 255513 35848 255682
rect 35806 255504 35862 255513
rect 35624 255468 35676 255474
rect 35806 255439 35862 255448
rect 35624 255410 35676 255416
rect 35440 255332 35492 255338
rect 35440 255274 35492 255280
rect 35438 255096 35494 255105
rect 35438 255031 35494 255040
rect 35806 255096 35862 255105
rect 35806 255031 35862 255040
rect 35452 253978 35480 255031
rect 35622 254688 35678 254697
rect 35622 254623 35678 254632
rect 35636 254182 35664 254623
rect 35820 254590 35848 255031
rect 35808 254584 35860 254590
rect 35808 254526 35860 254532
rect 39764 254584 39816 254590
rect 39764 254526 39816 254532
rect 35808 254312 35860 254318
rect 35806 254280 35808 254289
rect 35860 254280 35862 254289
rect 35806 254215 35862 254224
rect 35624 254176 35676 254182
rect 35624 254118 35676 254124
rect 35440 253972 35492 253978
rect 35440 253914 35492 253920
rect 35530 253056 35586 253065
rect 35530 252991 35586 253000
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 35544 252618 35572 252991
rect 35820 252754 35848 252991
rect 35808 252748 35860 252754
rect 35808 252690 35860 252696
rect 39776 252657 39804 254526
rect 40040 254312 40092 254318
rect 40040 254254 40092 254260
rect 40052 253881 40080 254254
rect 40038 253872 40094 253881
rect 40038 253807 40094 253816
rect 40420 253065 40448 255682
rect 42812 255542 42840 289786
rect 42996 280158 43024 293111
rect 42984 280152 43036 280158
rect 42984 280094 43036 280100
rect 43180 257553 43208 299446
rect 43456 281518 43484 401610
rect 43640 386753 43668 491914
rect 43824 426698 43852 531286
rect 44284 427854 44312 543706
rect 44560 429214 44588 550606
rect 44548 429208 44600 429214
rect 44548 429150 44600 429156
rect 44272 427848 44324 427854
rect 44272 427790 44324 427796
rect 44546 426864 44602 426873
rect 44546 426799 44602 426808
rect 43812 426692 43864 426698
rect 43812 426634 43864 426640
rect 44272 426488 44324 426494
rect 44272 426430 44324 426436
rect 43994 424008 44050 424017
rect 43994 423943 44050 423952
rect 43810 423192 43866 423201
rect 43810 423127 43866 423136
rect 43824 402966 43852 423127
rect 43812 402960 43864 402966
rect 43812 402902 43864 402908
rect 44008 400178 44036 423943
rect 44284 402974 44312 426430
rect 44284 402946 44404 402974
rect 43996 400172 44048 400178
rect 43996 400114 44048 400120
rect 43626 386744 43682 386753
rect 43626 386679 43682 386688
rect 44376 385121 44404 402946
rect 44362 385112 44418 385121
rect 44362 385047 44418 385056
rect 44560 383790 44588 426799
rect 44548 383784 44600 383790
rect 44548 383726 44600 383732
rect 44638 383480 44694 383489
rect 44638 383415 44694 383424
rect 43626 381848 43682 381857
rect 43626 381783 43682 381792
rect 43640 341086 43668 381783
rect 44178 381032 44234 381041
rect 44178 380967 44234 380976
rect 43810 378176 43866 378185
rect 43810 378111 43866 378120
rect 43824 364138 43852 378111
rect 44192 369753 44220 380967
rect 44362 378584 44418 378593
rect 44362 378519 44418 378528
rect 44178 369744 44234 369753
rect 44178 369679 44234 369688
rect 43812 364132 43864 364138
rect 43812 364074 43864 364080
rect 44376 360194 44404 378519
rect 44364 360188 44416 360194
rect 44364 360130 44416 360136
rect 44652 342310 44680 383415
rect 44640 342304 44692 342310
rect 44640 342246 44692 342252
rect 43628 341080 43680 341086
rect 43628 341022 43680 341028
rect 44456 340944 44508 340950
rect 44456 340886 44508 340892
rect 44270 339008 44326 339017
rect 44270 338943 44326 338952
rect 43628 336796 43680 336802
rect 43628 336738 43680 336744
rect 43640 315926 43668 336738
rect 43810 335744 43866 335753
rect 43810 335679 43866 335688
rect 43824 316946 43852 335679
rect 43994 334928 44050 334937
rect 43994 334863 44050 334872
rect 44008 321298 44036 334863
rect 43996 321292 44048 321298
rect 43996 321234 44048 321240
rect 43812 316940 43864 316946
rect 43812 316882 43864 316888
rect 43628 315920 43680 315926
rect 43628 315862 43680 315868
rect 43812 313948 43864 313954
rect 43812 313890 43864 313896
rect 43628 301300 43680 301306
rect 43628 301242 43680 301248
rect 43640 300937 43668 301242
rect 43626 300928 43682 300937
rect 43626 300863 43682 300872
rect 43626 290728 43682 290737
rect 43626 290663 43682 290672
rect 43640 290358 43668 290663
rect 43628 290352 43680 290358
rect 43628 290294 43680 290300
rect 43628 284368 43680 284374
rect 43628 284310 43680 284316
rect 43444 281512 43496 281518
rect 43444 281454 43496 281460
rect 43166 257544 43222 257553
rect 43166 257479 43222 257488
rect 41696 255536 41748 255542
rect 42064 255536 42116 255542
rect 41748 255484 42064 255490
rect 41696 255478 42116 255484
rect 42800 255536 42852 255542
rect 42800 255478 42852 255484
rect 41708 255462 42104 255478
rect 41708 255338 42104 255354
rect 41696 255332 42116 255338
rect 41748 255326 42064 255332
rect 41696 255274 41748 255280
rect 42064 255274 42116 255280
rect 41234 254280 41290 254289
rect 41234 254215 41290 254224
rect 41248 254114 41276 254215
rect 41236 254108 41288 254114
rect 41236 254050 41288 254056
rect 41696 253972 41748 253978
rect 42064 253972 42116 253978
rect 41748 253920 42064 253934
rect 41696 253914 42116 253920
rect 41708 253906 42104 253914
rect 42890 253872 42946 253881
rect 42890 253807 42946 253816
rect 42430 253600 42486 253609
rect 42430 253535 42486 253544
rect 40406 253056 40462 253065
rect 40406 252991 40462 253000
rect 41696 252748 41748 252754
rect 41696 252690 41748 252696
rect 39762 252648 39818 252657
rect 35532 252612 35584 252618
rect 39762 252583 39818 252592
rect 40040 252612 40092 252618
rect 35532 252554 35584 252560
rect 40040 252554 40092 252560
rect 31022 252240 31078 252249
rect 31022 252175 31078 252184
rect 31036 242214 31064 252175
rect 35530 251832 35586 251841
rect 35530 251767 35586 251776
rect 35806 251832 35862 251841
rect 35806 251767 35862 251776
rect 35544 251258 35572 251767
rect 35820 251530 35848 251767
rect 35808 251524 35860 251530
rect 35808 251466 35860 251472
rect 35532 251252 35584 251258
rect 35532 251194 35584 251200
rect 35438 251016 35494 251025
rect 35438 250951 35494 250960
rect 35452 249966 35480 250951
rect 35622 250608 35678 250617
rect 35622 250543 35678 250552
rect 35440 249960 35492 249966
rect 35440 249902 35492 249908
rect 35636 249830 35664 250543
rect 35808 250232 35860 250238
rect 35806 250200 35808 250209
rect 39396 250232 39448 250238
rect 35860 250200 35862 250209
rect 35806 250135 35862 250144
rect 39394 250200 39396 250209
rect 39448 250200 39450 250209
rect 39394 250135 39450 250144
rect 39856 249960 39908 249966
rect 39856 249902 39908 249908
rect 35624 249824 35676 249830
rect 35624 249766 35676 249772
rect 35438 249384 35494 249393
rect 35438 249319 35494 249328
rect 35452 248606 35480 249319
rect 35622 248976 35678 248985
rect 35622 248911 35678 248920
rect 35440 248600 35492 248606
rect 35440 248542 35492 248548
rect 35636 248470 35664 248911
rect 35808 248872 35860 248878
rect 35808 248814 35860 248820
rect 35820 248577 35848 248814
rect 39120 248600 39172 248606
rect 35806 248568 35862 248577
rect 35806 248503 35862 248512
rect 39118 248568 39120 248577
rect 39172 248568 39174 248577
rect 39118 248503 39174 248512
rect 35624 248464 35676 248470
rect 35624 248406 35676 248412
rect 35806 248160 35862 248169
rect 35806 248095 35862 248104
rect 35622 247752 35678 247761
rect 35622 247687 35678 247696
rect 35636 247246 35664 247687
rect 35820 247518 35848 248095
rect 35808 247512 35860 247518
rect 35808 247454 35860 247460
rect 35806 247344 35862 247353
rect 35806 247279 35862 247288
rect 35624 247240 35676 247246
rect 35624 247182 35676 247188
rect 35820 247110 35848 247279
rect 35808 247104 35860 247110
rect 35808 247046 35860 247052
rect 39868 245721 39896 249902
rect 40052 249558 40080 252554
rect 41708 252249 41736 252690
rect 41694 252240 41750 252249
rect 41694 252175 41750 252184
rect 41510 251832 41566 251841
rect 41510 251767 41566 251776
rect 41524 251530 41552 251767
rect 41512 251524 41564 251530
rect 41512 251466 41564 251472
rect 41694 251424 41750 251433
rect 41694 251359 41750 251368
rect 41708 251258 41736 251359
rect 41696 251252 41748 251258
rect 41696 251194 41748 251200
rect 41696 249824 41748 249830
rect 42064 249824 42116 249830
rect 41748 249772 42064 249778
rect 41696 249766 42116 249772
rect 41708 249750 42104 249766
rect 40040 249552 40092 249558
rect 40040 249494 40092 249500
rect 41696 249552 41748 249558
rect 41748 249500 42104 249506
rect 41696 249494 42104 249500
rect 41708 249490 42104 249494
rect 41708 249484 42116 249490
rect 41708 249478 42064 249484
rect 42064 249426 42116 249432
rect 40132 248872 40184 248878
rect 40132 248814 40184 248820
rect 39854 245712 39910 245721
rect 39854 245647 39910 245656
rect 40144 245177 40172 248814
rect 41696 248464 41748 248470
rect 42064 248464 42116 248470
rect 41748 248412 42064 248418
rect 41696 248406 42116 248412
rect 41708 248390 42104 248406
rect 40408 247512 40460 247518
rect 40408 247454 40460 247460
rect 40420 247353 40448 247454
rect 40406 247344 40462 247353
rect 40406 247279 40462 247288
rect 41696 247240 41748 247246
rect 42064 247240 42116 247246
rect 41748 247188 42064 247194
rect 41696 247182 42116 247188
rect 41708 247166 42104 247182
rect 41696 247104 41748 247110
rect 42064 247104 42116 247110
rect 41748 247052 42064 247058
rect 41696 247046 42116 247052
rect 41708 247030 42104 247046
rect 40130 245168 40186 245177
rect 40130 245103 40186 245112
rect 31024 242208 31076 242214
rect 31024 242150 31076 242156
rect 41696 242208 41748 242214
rect 41748 242156 42288 242162
rect 41696 242150 42288 242156
rect 41708 242134 42288 242150
rect 42062 240136 42118 240145
rect 42062 240071 42118 240080
rect 42076 239836 42104 240071
rect 41800 238513 41828 238649
rect 41786 238504 41842 238513
rect 41786 238439 41842 238448
rect 42062 238368 42118 238377
rect 42062 238303 42118 238312
rect 42076 238000 42104 238303
rect 42260 237697 42288 242134
rect 42246 237688 42302 237697
rect 42246 237623 42302 237632
rect 42444 237425 42472 253535
rect 42616 249484 42668 249490
rect 42616 249426 42668 249432
rect 42628 238377 42656 249426
rect 42904 238754 42932 253807
rect 43442 252648 43498 252657
rect 43442 252583 43498 252592
rect 43258 250200 43314 250209
rect 43258 250135 43314 250144
rect 43074 245168 43130 245177
rect 43074 245103 43130 245112
rect 43088 238754 43116 245103
rect 43272 238754 43300 250135
rect 43456 238754 43484 252583
rect 42812 238726 42932 238754
rect 42996 238726 43116 238754
rect 43180 238726 43300 238754
rect 43364 238726 43484 238754
rect 42614 238368 42670 238377
rect 42614 238303 42670 238312
rect 42430 237416 42486 237425
rect 42430 237351 42486 237360
rect 41786 236600 41842 236609
rect 41786 236535 41842 236544
rect 41800 236164 41828 236535
rect 42432 235952 42484 235958
rect 42432 235894 42484 235900
rect 42444 234983 42472 235894
rect 42182 234955 42472 234983
rect 42432 234592 42484 234598
rect 42432 234534 42484 234540
rect 42444 234342 42472 234534
rect 42182 234314 42472 234342
rect 42432 234252 42484 234258
rect 42432 234194 42484 234200
rect 42444 233695 42472 234194
rect 42182 233667 42472 233695
rect 42168 233158 42288 233186
rect 42168 233104 42196 233158
rect 42260 233118 42288 233158
rect 42260 233090 42472 233118
rect 42444 231878 42472 233090
rect 42432 231872 42484 231878
rect 42432 231814 42484 231820
rect 42432 231736 42484 231742
rect 42432 231678 42484 231684
rect 42444 230670 42472 231678
rect 42182 230642 42472 230670
rect 42156 230444 42208 230450
rect 42156 230386 42208 230392
rect 42168 229976 42196 230386
rect 42182 229350 42564 229378
rect 41970 228984 42026 228993
rect 41970 228919 42026 228928
rect 41984 228820 42012 228919
rect 42536 227730 42564 229350
rect 42812 229094 42840 238726
rect 42996 234258 43024 238726
rect 42984 234252 43036 234258
rect 42984 234194 43036 234200
rect 43180 230450 43208 238726
rect 43168 230444 43220 230450
rect 43168 230386 43220 230392
rect 42812 229066 42932 229094
rect 42524 227724 42576 227730
rect 42524 227666 42576 227672
rect 42062 227352 42118 227361
rect 42062 227287 42118 227296
rect 42076 226984 42104 227287
rect 42168 226358 42288 226386
rect 42168 226304 42196 226358
rect 42260 226318 42288 226358
rect 42260 226290 42656 226318
rect 42432 226228 42484 226234
rect 42432 226170 42484 226176
rect 42444 225706 42472 226170
rect 42182 225678 42472 225706
rect 42628 224942 42656 226290
rect 42616 224936 42668 224942
rect 42616 224878 42668 224884
rect 28538 223952 28594 223961
rect 28538 223887 28594 223896
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 28552 212673 28580 223887
rect 41694 223680 41750 223689
rect 41694 223615 41750 223624
rect 40682 222320 40738 222329
rect 40682 222255 40738 222264
rect 33048 217252 33100 217258
rect 33048 217194 33100 217200
rect 33060 214305 33088 217194
rect 40314 216744 40370 216753
rect 40314 216679 40370 216688
rect 35806 215112 35862 215121
rect 35806 215047 35862 215056
rect 35820 214878 35848 215047
rect 35808 214872 35860 214878
rect 35808 214814 35860 214820
rect 33046 214296 33102 214305
rect 33046 214231 33102 214240
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 39946 214296 40002 214305
rect 39946 214231 40002 214240
rect 35820 214130 35848 214231
rect 39960 214130 39988 214231
rect 35808 214124 35860 214130
rect 35808 214066 35860 214072
rect 39948 214124 40000 214130
rect 39948 214066 40000 214072
rect 39946 213888 40002 213897
rect 39946 213823 40002 213832
rect 35438 213480 35494 213489
rect 35438 213415 35494 213424
rect 28538 212664 28594 212673
rect 28538 212599 28594 212608
rect 35452 212566 35480 213415
rect 35622 213072 35678 213081
rect 35622 213007 35678 213016
rect 35636 212702 35664 213007
rect 35808 212968 35860 212974
rect 35808 212910 35860 212916
rect 35624 212696 35676 212702
rect 35820 212673 35848 212910
rect 35624 212638 35676 212644
rect 35806 212664 35862 212673
rect 35806 212599 35862 212608
rect 39960 212566 39988 213823
rect 40328 212974 40356 216679
rect 40316 212968 40368 212974
rect 40316 212910 40368 212916
rect 40696 212702 40724 222255
rect 41510 217288 41566 217297
rect 41510 217223 41512 217232
rect 41564 217223 41566 217232
rect 41512 217194 41564 217200
rect 41510 215112 41566 215121
rect 41510 215047 41566 215056
rect 41524 214878 41552 215047
rect 41512 214872 41564 214878
rect 41512 214814 41564 214820
rect 40684 212696 40736 212702
rect 40684 212638 40736 212644
rect 35440 212560 35492 212566
rect 35440 212502 35492 212508
rect 39948 212560 40000 212566
rect 39948 212502 40000 212508
rect 40958 212256 41014 212265
rect 40958 212191 41014 212200
rect 35806 211848 35862 211857
rect 35806 211783 35862 211792
rect 35820 211614 35848 211783
rect 40972 211614 41000 212191
rect 35808 211608 35860 211614
rect 35808 211550 35860 211556
rect 40960 211608 41012 211614
rect 40960 211550 41012 211556
rect 35622 211440 35678 211449
rect 35622 211375 35678 211384
rect 39670 211440 39726 211449
rect 39670 211375 39672 211384
rect 35636 211206 35664 211375
rect 39724 211375 39726 211384
rect 39672 211346 39724 211352
rect 35808 211336 35860 211342
rect 35808 211278 35860 211284
rect 35624 211200 35676 211206
rect 35624 211142 35676 211148
rect 35820 211041 35848 211278
rect 41512 211200 41564 211206
rect 41512 211142 41564 211148
rect 41524 211041 41552 211142
rect 35806 211032 35862 211041
rect 35806 210967 35862 210976
rect 41510 211032 41566 211041
rect 41510 210967 41566 210976
rect 35622 210624 35678 210633
rect 35622 210559 35678 210568
rect 35636 209846 35664 210559
rect 35806 210216 35862 210225
rect 35806 210151 35862 210160
rect 35820 209982 35848 210151
rect 35808 209976 35860 209982
rect 35808 209918 35860 209924
rect 40040 209976 40092 209982
rect 40040 209918 40092 209924
rect 35624 209840 35676 209846
rect 35624 209782 35676 209788
rect 35806 209400 35862 209409
rect 35806 209335 35862 209344
rect 30286 208992 30342 209001
rect 30286 208927 30342 208936
rect 30300 202201 30328 208927
rect 35820 208758 35848 209335
rect 40052 209001 40080 209918
rect 41708 209846 41736 223615
rect 42064 217320 42116 217326
rect 42062 217288 42064 217297
rect 42116 217288 42118 217297
rect 42062 217223 42118 217232
rect 42904 211449 42932 229066
rect 43166 215112 43222 215121
rect 43166 215047 43222 215056
rect 43180 214810 43208 215047
rect 43168 214804 43220 214810
rect 43168 214746 43220 214752
rect 43364 212265 43392 238726
rect 43640 214305 43668 284310
rect 43824 257038 43852 313890
rect 44284 306374 44312 338943
rect 44192 306346 44312 306374
rect 44192 296954 44220 306346
rect 44468 298246 44496 340886
rect 44638 330712 44694 330721
rect 44638 330647 44694 330656
rect 44652 325378 44680 330647
rect 44640 325372 44692 325378
rect 44640 325314 44692 325320
rect 44456 298240 44508 298246
rect 44456 298182 44508 298188
rect 44362 297256 44418 297265
rect 44362 297191 44418 297200
rect 44180 296948 44232 296954
rect 44180 296890 44232 296896
rect 44178 291544 44234 291553
rect 44178 291479 44234 291488
rect 43996 291236 44048 291242
rect 43996 291178 44048 291184
rect 44008 277394 44036 291178
rect 43916 277366 44036 277394
rect 44192 277386 44220 291479
rect 44376 277394 44404 297191
rect 44548 296744 44600 296750
rect 44548 296686 44600 296692
rect 43916 277114 43944 277366
rect 44100 277358 44220 277386
rect 44284 277366 44404 277394
rect 44100 277234 44128 277358
rect 44088 277228 44140 277234
rect 44088 277170 44140 277176
rect 43916 277098 44036 277114
rect 43916 277092 44048 277098
rect 43916 277086 43996 277092
rect 43996 277034 44048 277040
rect 43812 257032 43864 257038
rect 43812 256974 43864 256980
rect 44284 254289 44312 277366
rect 44270 254280 44326 254289
rect 44270 254215 44326 254224
rect 44560 253978 44588 296686
rect 44548 253972 44600 253978
rect 44548 253914 44600 253920
rect 44546 251832 44602 251841
rect 44546 251767 44602 251776
rect 43810 248568 43866 248577
rect 43810 248503 43866 248512
rect 43824 234598 43852 248503
rect 44364 248464 44416 248470
rect 44364 248406 44416 248412
rect 44178 247344 44234 247353
rect 44178 247279 44234 247288
rect 44192 239970 44220 247279
rect 44180 239964 44232 239970
rect 44180 239906 44232 239912
rect 43812 234592 43864 234598
rect 43812 234534 43864 234540
rect 44376 231742 44404 248406
rect 44560 240145 44588 251767
rect 44546 240136 44602 240145
rect 44546 240071 44602 240080
rect 44640 239964 44692 239970
rect 44640 239906 44692 239912
rect 44652 235958 44680 239906
rect 44640 235952 44692 235958
rect 44640 235894 44692 235900
rect 44364 231736 44416 231742
rect 44364 231678 44416 231684
rect 44836 231266 44864 758095
rect 45020 753574 45048 763671
rect 45008 753568 45060 753574
rect 45008 753510 45060 753516
rect 45008 728680 45060 728686
rect 45008 728622 45060 728628
rect 45020 685914 45048 728622
rect 45008 685908 45060 685914
rect 45008 685850 45060 685856
rect 45190 679960 45246 679969
rect 45190 679895 45246 679904
rect 45006 677920 45062 677929
rect 45006 677855 45062 677864
rect 45020 276729 45048 677855
rect 45204 667962 45232 679895
rect 45192 667956 45244 667962
rect 45192 667898 45244 667904
rect 45190 632088 45246 632097
rect 45190 632023 45246 632032
rect 45204 620945 45232 632023
rect 45190 620936 45246 620945
rect 45190 620871 45246 620880
rect 45374 552392 45430 552401
rect 45374 552327 45430 552336
rect 45190 551168 45246 551177
rect 45190 551103 45246 551112
rect 45204 532710 45232 551103
rect 45388 536654 45416 552327
rect 45376 536648 45428 536654
rect 45376 536590 45428 536596
rect 45192 532704 45244 532710
rect 45192 532646 45244 532652
rect 45558 424824 45614 424833
rect 45558 424759 45614 424768
rect 45190 423600 45246 423609
rect 45190 423535 45246 423544
rect 45204 402558 45232 423535
rect 45374 421288 45430 421297
rect 45374 421223 45430 421232
rect 45388 408338 45416 421223
rect 45376 408332 45428 408338
rect 45376 408274 45428 408280
rect 45572 406026 45600 424759
rect 45742 419520 45798 419529
rect 45742 419455 45798 419464
rect 45756 418198 45784 419455
rect 45744 418192 45796 418198
rect 45744 418134 45796 418140
rect 45560 406020 45612 406026
rect 45560 405962 45612 405968
rect 45192 402552 45244 402558
rect 45192 402494 45244 402500
rect 45376 385076 45428 385082
rect 45376 385018 45428 385024
rect 45190 376952 45246 376961
rect 45190 376887 45246 376896
rect 45204 365702 45232 376887
rect 45192 365696 45244 365702
rect 45192 365638 45244 365644
rect 45192 347064 45244 347070
rect 45192 347006 45244 347012
rect 45006 276720 45062 276729
rect 45006 276655 45062 276664
rect 45204 256766 45232 347006
rect 45388 343097 45416 385018
rect 45374 343088 45430 343097
rect 45374 343023 45430 343032
rect 45558 338736 45614 338745
rect 45558 338671 45614 338680
rect 45374 338192 45430 338201
rect 45374 338127 45430 338136
rect 45388 320006 45416 338127
rect 45376 320000 45428 320006
rect 45376 319942 45428 319948
rect 45572 310486 45600 338671
rect 46018 333704 46074 333713
rect 46018 333639 46074 333648
rect 45834 332888 45890 332897
rect 45834 332823 45890 332832
rect 45848 327078 45876 332823
rect 45836 327072 45888 327078
rect 45836 327014 45888 327020
rect 46032 319190 46060 333639
rect 46020 319184 46072 319190
rect 46020 319126 46072 319132
rect 45560 310480 45612 310486
rect 45560 310422 45612 310428
rect 45558 296032 45614 296041
rect 45558 295967 45614 295976
rect 45374 293992 45430 294001
rect 45374 293927 45430 293936
rect 45388 273222 45416 293927
rect 45376 273216 45428 273222
rect 45376 273158 45428 273164
rect 45572 269074 45600 295967
rect 45560 269068 45612 269074
rect 45560 269010 45612 269016
rect 45192 256760 45244 256766
rect 45192 256702 45244 256708
rect 45008 255332 45060 255338
rect 45008 255274 45060 255280
rect 44824 231260 44876 231266
rect 44824 231202 44876 231208
rect 43626 214296 43682 214305
rect 43626 214231 43682 214240
rect 45020 213897 45048 255274
rect 45374 253056 45430 253065
rect 45374 252991 45430 253000
rect 45388 238754 45416 252991
rect 45558 252240 45614 252249
rect 45558 252175 45614 252184
rect 45296 238726 45416 238754
rect 45296 216753 45324 238726
rect 45572 226234 45600 252175
rect 45742 245712 45798 245721
rect 45742 245647 45798 245656
rect 45560 226228 45612 226234
rect 45560 226170 45612 226176
rect 45756 224942 45784 245647
rect 46216 231674 46244 806239
rect 47596 799066 47624 923238
rect 50344 909492 50396 909498
rect 50344 909434 50396 909440
rect 50356 815658 50384 909434
rect 51908 858424 51960 858430
rect 51908 858366 51960 858372
rect 51724 818372 51776 818378
rect 51724 818314 51776 818320
rect 50344 815652 50396 815658
rect 50344 815594 50396 815600
rect 48964 807492 49016 807498
rect 48964 807434 49016 807440
rect 47584 799060 47636 799066
rect 47584 799002 47636 799008
rect 47768 793620 47820 793626
rect 47768 793562 47820 793568
rect 47582 763328 47638 763337
rect 47582 763263 47638 763272
rect 46386 721168 46442 721177
rect 46386 721103 46442 721112
rect 46204 231668 46256 231674
rect 46204 231610 46256 231616
rect 46400 228857 46428 721103
rect 46572 427848 46624 427854
rect 46572 427790 46624 427796
rect 46584 345953 46612 427790
rect 46570 345944 46626 345953
rect 46570 345879 46626 345888
rect 46572 336796 46624 336802
rect 46572 336738 46624 336744
rect 46584 259593 46612 336738
rect 46754 331256 46810 331265
rect 46754 331191 46810 331200
rect 46768 318782 46796 331191
rect 46756 318776 46808 318782
rect 46756 318718 46808 318724
rect 47030 294536 47086 294545
rect 47030 294471 47086 294480
rect 47044 274650 47072 294471
rect 47216 294024 47268 294030
rect 47216 293966 47268 293972
rect 47032 274644 47084 274650
rect 47032 274586 47084 274592
rect 47228 267714 47256 293966
rect 47216 267708 47268 267714
rect 47216 267650 47268 267656
rect 46570 259584 46626 259593
rect 46570 259519 46626 259528
rect 47030 251424 47086 251433
rect 47030 251359 47086 251368
rect 47044 231878 47072 251359
rect 47216 249824 47268 249830
rect 47216 249766 47268 249772
rect 47032 231872 47084 231878
rect 47032 231814 47084 231820
rect 46386 228848 46442 228857
rect 46386 228783 46442 228792
rect 47228 227730 47256 249766
rect 47596 231402 47624 763263
rect 47780 731377 47808 793562
rect 47766 731368 47822 731377
rect 47766 731303 47822 731312
rect 47768 674892 47820 674898
rect 47768 674834 47820 674840
rect 47780 646105 47808 674834
rect 47766 646096 47822 646105
rect 47766 646031 47822 646040
rect 47768 623824 47820 623830
rect 47768 623766 47820 623772
rect 47780 601361 47808 623766
rect 47766 601352 47822 601361
rect 47766 601287 47822 601296
rect 47766 590336 47822 590345
rect 47766 590271 47822 590280
rect 47584 231396 47636 231402
rect 47584 231338 47636 231344
rect 47780 228313 47808 590271
rect 47952 480276 48004 480282
rect 47952 480218 48004 480224
rect 47964 386510 47992 480218
rect 48136 389292 48188 389298
rect 48136 389234 48188 389240
rect 47952 386504 48004 386510
rect 47952 386446 48004 386452
rect 48148 299538 48176 389234
rect 48136 299532 48188 299538
rect 48136 299474 48188 299480
rect 48976 278458 49004 807434
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 50356 731202 50384 805938
rect 50712 753568 50764 753574
rect 50712 753510 50764 753516
rect 50344 731196 50396 731202
rect 50344 731138 50396 731144
rect 50528 714876 50580 714882
rect 50528 714818 50580 714824
rect 50344 676456 50396 676462
rect 50344 676398 50396 676404
rect 49148 636268 49200 636274
rect 49148 636210 49200 636216
rect 49160 601730 49188 636210
rect 49148 601724 49200 601730
rect 49148 601666 49200 601672
rect 49148 597576 49200 597582
rect 49148 597518 49200 597524
rect 49160 557870 49188 597518
rect 49148 557864 49200 557870
rect 49148 557806 49200 557812
rect 49148 546576 49200 546582
rect 49148 546518 49200 546524
rect 48964 278452 49016 278458
rect 48964 278394 49016 278400
rect 49160 228585 49188 546518
rect 49332 466472 49384 466478
rect 49332 466414 49384 466420
rect 49344 387530 49372 466414
rect 49332 387524 49384 387530
rect 49332 387466 49384 387472
rect 49332 375420 49384 375426
rect 49332 375362 49384 375368
rect 49344 301034 49372 375362
rect 49332 301028 49384 301034
rect 49332 300970 49384 300976
rect 49332 298172 49384 298178
rect 49332 298114 49384 298120
rect 49146 228576 49202 228585
rect 49146 228511 49202 228520
rect 47766 228304 47822 228313
rect 47766 228239 47822 228248
rect 47216 227724 47268 227730
rect 47216 227666 47268 227672
rect 45744 224936 45796 224942
rect 45744 224878 45796 224884
rect 47582 222592 47638 222601
rect 47582 222527 47638 222536
rect 45282 216744 45338 216753
rect 45282 216679 45338 216688
rect 45006 213888 45062 213897
rect 45006 213823 45062 213832
rect 43350 212256 43406 212265
rect 43350 212191 43406 212200
rect 42890 211440 42946 211449
rect 42890 211375 42946 211384
rect 42340 211200 42392 211206
rect 42340 211142 42392 211148
rect 42352 211041 42380 211142
rect 42338 211032 42394 211041
rect 42338 210967 42394 210976
rect 41696 209840 41748 209846
rect 41696 209782 41748 209788
rect 40038 208992 40094 209001
rect 40038 208927 40094 208936
rect 35808 208752 35860 208758
rect 35808 208694 35860 208700
rect 39948 208684 40000 208690
rect 39948 208626 40000 208632
rect 35806 208584 35862 208593
rect 35806 208519 35862 208528
rect 35820 208418 35848 208519
rect 35808 208412 35860 208418
rect 35808 208354 35860 208360
rect 35530 207360 35586 207369
rect 35530 207295 35586 207304
rect 35806 207360 35862 207369
rect 35806 207295 35808 207304
rect 35544 207058 35572 207295
rect 35860 207295 35862 207304
rect 35808 207266 35860 207272
rect 35532 207052 35584 207058
rect 35532 206994 35584 207000
rect 35806 206544 35862 206553
rect 35806 206479 35862 206488
rect 35820 205970 35848 206479
rect 35808 205964 35860 205970
rect 35808 205906 35860 205912
rect 39764 205964 39816 205970
rect 39764 205906 39816 205912
rect 35806 205728 35862 205737
rect 35806 205663 35808 205672
rect 35860 205663 35862 205672
rect 35808 205634 35860 205640
rect 35622 205320 35678 205329
rect 35622 205255 35678 205264
rect 35636 204678 35664 205255
rect 35808 204944 35860 204950
rect 35806 204912 35808 204921
rect 35860 204912 35862 204921
rect 35806 204847 35862 204856
rect 35624 204672 35676 204678
rect 35624 204614 35676 204620
rect 35808 204536 35860 204542
rect 35530 204504 35586 204513
rect 35530 204439 35586 204448
rect 35806 204504 35808 204513
rect 35860 204504 35862 204513
rect 35806 204439 35862 204448
rect 35544 204338 35572 204439
rect 35532 204332 35584 204338
rect 35532 204274 35584 204280
rect 39776 204105 39804 205906
rect 39960 205737 39988 208626
rect 41708 208418 42104 208434
rect 41696 208412 42116 208418
rect 41748 208406 42064 208412
rect 41696 208354 41748 208360
rect 42064 208354 42116 208360
rect 43076 208412 43128 208418
rect 43076 208354 43128 208360
rect 40132 207324 40184 207330
rect 40132 207266 40184 207272
rect 40144 206961 40172 207266
rect 40960 207052 41012 207058
rect 40960 206994 41012 207000
rect 40130 206952 40186 206961
rect 40130 206887 40186 206896
rect 39946 205728 40002 205737
rect 39946 205663 40002 205672
rect 40972 205329 41000 206994
rect 42890 206952 42946 206961
rect 42890 206887 42946 206896
rect 41708 205698 42104 205714
rect 41696 205692 42116 205698
rect 41748 205686 42064 205692
rect 41696 205634 41748 205640
rect 42064 205634 42116 205640
rect 40958 205320 41014 205329
rect 40958 205255 41014 205264
rect 40776 204944 40828 204950
rect 40776 204886 40828 204892
rect 40788 204513 40816 204886
rect 41708 204746 42104 204762
rect 41696 204740 42116 204746
rect 41748 204734 42064 204740
rect 41696 204682 41748 204688
rect 42064 204682 42116 204688
rect 42064 204604 42116 204610
rect 42064 204546 42116 204552
rect 41696 204536 41748 204542
rect 40774 204504 40830 204513
rect 42076 204490 42104 204546
rect 41748 204484 42104 204490
rect 41696 204478 42104 204484
rect 41708 204462 42104 204478
rect 40774 204439 40830 204448
rect 41708 204338 42104 204354
rect 41696 204332 42116 204338
rect 41748 204326 42064 204332
rect 41696 204274 41748 204280
rect 42064 204274 42116 204280
rect 39762 204096 39818 204105
rect 39762 204031 39818 204040
rect 35622 203688 35678 203697
rect 35622 203623 35678 203632
rect 35636 203182 35664 203623
rect 35806 203280 35862 203289
rect 35806 203215 35862 203224
rect 40038 203280 40094 203289
rect 40038 203215 40094 203224
rect 35624 203176 35676 203182
rect 35624 203118 35676 203124
rect 35820 202910 35848 203215
rect 40052 202910 40080 203215
rect 41604 203176 41656 203182
rect 41604 203118 41656 203124
rect 41616 202994 41644 203118
rect 41786 203008 41842 203017
rect 41616 202966 41786 202994
rect 41786 202943 41842 202952
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 40040 202904 40092 202910
rect 40040 202846 40092 202852
rect 30286 202192 30342 202201
rect 30286 202127 30342 202136
rect 41786 197160 41842 197169
rect 41786 197095 41842 197104
rect 41800 196656 41828 197095
rect 42904 195974 42932 206887
rect 43088 195974 43116 208354
rect 44178 205728 44234 205737
rect 43444 205692 43496 205698
rect 44178 205663 44234 205672
rect 43444 205634 43496 205640
rect 43258 205320 43314 205329
rect 43258 205255 43314 205264
rect 42812 195946 42932 195974
rect 42996 195946 43116 195974
rect 42432 195696 42484 195702
rect 42432 195638 42484 195644
rect 42168 195486 42288 195514
rect 42168 195432 42196 195486
rect 42260 195446 42288 195486
rect 42444 195446 42472 195638
rect 42260 195418 42472 195446
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42432 193180 42484 193186
rect 42432 193122 42484 193128
rect 42444 192998 42472 193122
rect 42168 192930 42196 192984
rect 42260 192970 42472 192998
rect 42260 192930 42288 192970
rect 42168 192902 42288 192930
rect 42432 191820 42484 191826
rect 42182 191768 42432 191774
rect 42182 191762 42484 191768
rect 42182 191746 42472 191762
rect 42432 191684 42484 191690
rect 42432 191626 42484 191632
rect 41786 191584 41842 191593
rect 41786 191519 41842 191528
rect 41800 191148 41828 191519
rect 42444 190482 42472 191626
rect 42182 190454 42472 190482
rect 42432 190392 42484 190398
rect 42432 190334 42484 190340
rect 42444 189938 42472 190334
rect 42182 189910 42472 189938
rect 42432 187672 42484 187678
rect 42432 187614 42484 187620
rect 42444 187459 42472 187614
rect 42182 187431 42472 187459
rect 42812 186810 42840 195946
rect 42996 190398 43024 195946
rect 42984 190392 43036 190398
rect 42984 190334 43036 190340
rect 42182 186782 42840 186810
rect 43272 186314 43300 205255
rect 43456 187678 43484 205634
rect 43810 204096 43866 204105
rect 43810 204031 43866 204040
rect 43626 203008 43682 203017
rect 43626 202943 43682 202952
rect 43640 195702 43668 202943
rect 43628 195696 43680 195702
rect 43628 195638 43680 195644
rect 43824 193186 43852 204031
rect 43812 193180 43864 193186
rect 43812 193122 43864 193128
rect 43444 187672 43496 187678
rect 43444 187614 43496 187620
rect 43088 186286 43300 186314
rect 43088 186266 43116 186286
rect 42536 186238 43116 186266
rect 42536 186198 42564 186238
rect 42168 186130 42196 186184
rect 42260 186170 42564 186198
rect 42260 186130 42288 186170
rect 42168 186102 42288 186130
rect 41786 185872 41842 185881
rect 41786 185807 41842 185816
rect 41800 185605 41828 185807
rect 41786 184104 41842 184113
rect 41786 184039 41842 184048
rect 41800 183765 41828 184039
rect 44192 183530 44220 205663
rect 44364 204740 44416 204746
rect 44364 204682 44416 204688
rect 44376 191690 44404 204682
rect 44546 204504 44602 204513
rect 44546 204439 44602 204448
rect 44560 191826 44588 204439
rect 47596 203289 47624 222527
rect 48964 215348 49016 215354
rect 48964 215290 49016 215296
rect 48976 204338 49004 215290
rect 49344 214810 49372 298114
rect 49516 290352 49568 290358
rect 49516 290294 49568 290300
rect 49528 278050 49556 290294
rect 49516 278044 49568 278050
rect 49516 277986 49568 277992
rect 50356 227225 50384 676398
rect 50540 626686 50568 714818
rect 50724 687750 50752 753510
rect 51736 712298 51764 818314
rect 51920 772886 51948 858366
rect 51908 772880 51960 772886
rect 51908 772822 51960 772828
rect 51908 727320 51960 727326
rect 51908 727262 51960 727268
rect 51724 712292 51776 712298
rect 51724 712234 51776 712240
rect 51724 701072 51776 701078
rect 51724 701014 51776 701020
rect 50712 687744 50764 687750
rect 50712 687686 50764 687692
rect 51736 643142 51764 701014
rect 51920 687410 51948 727262
rect 51908 687404 51960 687410
rect 51908 687346 51960 687352
rect 51908 647896 51960 647902
rect 51908 647838 51960 647844
rect 51724 643136 51776 643142
rect 51724 643078 51776 643084
rect 51724 633616 51776 633622
rect 51724 633558 51776 633564
rect 50528 626680 50580 626686
rect 50528 626622 50580 626628
rect 50528 590844 50580 590850
rect 50528 590786 50580 590792
rect 50540 231130 50568 590786
rect 50712 440292 50764 440298
rect 50712 440234 50764 440240
rect 50724 343874 50752 440234
rect 50896 356720 50948 356726
rect 50896 356662 50948 356668
rect 50712 343868 50764 343874
rect 50712 343810 50764 343816
rect 50712 334008 50764 334014
rect 50712 333950 50764 333956
rect 50724 265577 50752 333950
rect 50908 301306 50936 356662
rect 50896 301300 50948 301306
rect 50896 301242 50948 301248
rect 50710 265568 50766 265577
rect 50710 265503 50766 265512
rect 51736 231538 51764 633558
rect 51920 600370 51948 647838
rect 51908 600364 51960 600370
rect 51908 600306 51960 600312
rect 51908 583772 51960 583778
rect 51908 583714 51960 583720
rect 51920 557598 51948 583714
rect 51908 557592 51960 557598
rect 51908 557534 51960 557540
rect 52092 506524 52144 506530
rect 52092 506466 52144 506472
rect 51908 419552 51960 419558
rect 51908 419494 51960 419500
rect 51920 264246 51948 419494
rect 52104 364274 52132 506466
rect 52276 375556 52328 375562
rect 52276 375498 52328 375504
rect 52092 364268 52144 364274
rect 52092 364210 52144 364216
rect 52288 276690 52316 375498
rect 52276 276684 52328 276690
rect 52276 276626 52328 276632
rect 51908 264240 51960 264246
rect 51908 264182 51960 264188
rect 51724 231532 51776 231538
rect 51724 231474 51776 231480
rect 50528 231124 50580 231130
rect 50528 231066 50580 231072
rect 53116 230994 53144 931534
rect 53288 633752 53340 633758
rect 53288 633694 53340 633700
rect 53104 230988 53156 230994
rect 53104 230930 53156 230936
rect 53300 227497 53328 633694
rect 53472 376780 53524 376786
rect 53472 376722 53524 376728
rect 53484 277001 53512 376722
rect 54496 278089 54524 932894
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 62120 909492 62172 909498
rect 62120 909434 62172 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 62118 884776 62174 884785
rect 62118 884711 62120 884720
rect 62172 884711 62174 884720
rect 62120 884682 62172 884688
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 62118 858664 62174 858673
rect 62118 858599 62174 858608
rect 62132 858430 62160 858599
rect 62120 858424 62172 858430
rect 62120 858366 62172 858372
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 55864 832176 55916 832182
rect 55864 832118 55916 832124
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 55876 773022 55904 832118
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62118 793656 62174 793665
rect 62118 793591 62120 793600
rect 62172 793591 62174 793600
rect 62120 793562 62172 793568
rect 62118 780464 62174 780473
rect 62118 780399 62174 780408
rect 62132 780094 62160 780399
rect 56232 780088 56284 780094
rect 56232 780030 56284 780036
rect 62120 780088 62172 780094
rect 62120 780030 62172 780036
rect 55864 773016 55916 773022
rect 55864 772958 55916 772964
rect 56048 741124 56100 741130
rect 56048 741066 56100 741072
rect 55864 719160 55916 719166
rect 55864 719102 55916 719108
rect 54852 557592 54904 557598
rect 54852 557534 54904 557540
rect 54668 418192 54720 418198
rect 54668 418134 54720 418140
rect 54482 278080 54538 278089
rect 54482 278015 54538 278024
rect 53470 276992 53526 277001
rect 53470 276927 53526 276936
rect 54680 229809 54708 418134
rect 54864 408474 54892 557534
rect 55036 454096 55088 454102
rect 55036 454038 55088 454044
rect 54852 408468 54904 408474
rect 54852 408410 54904 408416
rect 55048 321570 55076 454038
rect 55036 321564 55088 321570
rect 55036 321506 55088 321512
rect 55876 231810 55904 719102
rect 56060 687274 56088 741066
rect 56244 730114 56272 780030
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 56232 730108 56284 730114
rect 56232 730050 56284 730056
rect 62118 728240 62174 728249
rect 62118 728175 62174 728184
rect 62132 727326 62160 728175
rect 62120 727320 62172 727326
rect 62120 727262 62172 727268
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62118 702264 62174 702273
rect 62118 702199 62174 702208
rect 62132 701078 62160 702199
rect 62120 701072 62172 701078
rect 62120 701014 62172 701020
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 56048 687268 56100 687274
rect 56048 687210 56100 687216
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 609278 62160 610943
rect 62120 609272 62172 609278
rect 62120 609214 62172 609220
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 571402 62160 571775
rect 62120 571396 62172 571402
rect 62120 571338 62172 571344
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 557598 62160 558719
rect 62120 557592 62172 557598
rect 62120 557534 62172 557540
rect 56048 547936 56100 547942
rect 56048 547878 56100 547884
rect 55864 231804 55916 231810
rect 55864 231746 55916 231752
rect 56060 230081 56088 547878
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 62762 532808 62818 532817
rect 62762 532743 62818 532752
rect 62776 523734 62804 532743
rect 62764 523728 62816 523734
rect 62764 523670 62816 523676
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 62120 491972 62172 491978
rect 62120 491914 62172 491920
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 56232 415472 56284 415478
rect 62120 415472 62172 415478
rect 56232 415414 56284 415420
rect 62118 415440 62120 415449
rect 62172 415440 62174 415449
rect 56244 343670 56272 415414
rect 62118 415375 62174 415384
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 62118 389328 62174 389337
rect 62118 389263 62120 389272
rect 62172 389263 62174 389272
rect 62120 389234 62172 389240
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 356726 62160 363287
rect 62120 356720 62172 356726
rect 62120 356662 62172 356668
rect 62118 350296 62174 350305
rect 62118 350231 62174 350240
rect 62132 347070 62160 350231
rect 62120 347064 62172 347070
rect 62120 347006 62172 347012
rect 56232 343664 56284 343670
rect 56232 343606 56284 343612
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 56232 332648 56284 332654
rect 56232 332590 56284 332596
rect 56244 278186 56272 332590
rect 62762 324184 62818 324193
rect 62762 324119 62818 324128
rect 62776 313954 62804 324119
rect 62764 313948 62816 313954
rect 62764 313890 62816 313896
rect 62762 311128 62818 311137
rect 62762 311063 62818 311072
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 60004 290012 60056 290018
rect 60004 289954 60056 289960
rect 56232 278180 56284 278186
rect 56232 278122 56284 278128
rect 56046 230072 56102 230081
rect 56046 230007 56102 230016
rect 54666 229800 54722 229809
rect 54666 229735 54722 229744
rect 53286 227488 53342 227497
rect 53286 227423 53342 227432
rect 50342 227216 50398 227225
rect 50342 227151 50398 227160
rect 60016 226953 60044 289954
rect 62118 285152 62174 285161
rect 62118 285087 62174 285096
rect 62132 284374 62160 285087
rect 62120 284368 62172 284374
rect 62120 284310 62172 284316
rect 61382 230344 61438 230353
rect 61382 230279 61438 230288
rect 60002 226944 60058 226953
rect 60002 226879 60058 226888
rect 59266 226672 59322 226681
rect 59266 226607 59322 226616
rect 56874 226128 56930 226137
rect 56874 226063 56930 226072
rect 50342 222048 50398 222057
rect 50342 221983 50398 221992
rect 49332 214804 49384 214810
rect 49332 214746 49384 214752
rect 50356 204610 50384 221983
rect 51722 221776 51778 221785
rect 51722 221711 51778 221720
rect 51736 211206 51764 221711
rect 56888 220522 56916 226063
rect 57612 220788 57664 220794
rect 57612 220730 57664 220736
rect 55956 220516 56008 220522
rect 55956 220458 56008 220464
rect 56876 220516 56928 220522
rect 56876 220458 56928 220464
rect 55968 217410 55996 220458
rect 56506 220008 56562 220017
rect 56506 219943 56562 219952
rect 56520 217410 56548 219943
rect 57624 217410 57652 220730
rect 58440 220108 58492 220114
rect 58440 220050 58492 220056
rect 58452 217410 58480 220050
rect 59280 217410 59308 226607
rect 60372 222896 60424 222902
rect 60372 222838 60424 222844
rect 60002 222048 60058 222057
rect 60002 221983 60058 221992
rect 59820 221604 59872 221610
rect 59820 221546 59872 221552
rect 59832 217410 59860 221546
rect 60016 221513 60044 221983
rect 60002 221504 60058 221513
rect 60002 221439 60058 221448
rect 60384 220114 60412 222838
rect 61396 220454 61424 230279
rect 62120 225616 62172 225622
rect 62120 225558 62172 225564
rect 61844 224392 61896 224398
rect 61844 224334 61896 224340
rect 60648 220448 60700 220454
rect 60648 220390 60700 220396
rect 61384 220448 61436 220454
rect 61384 220390 61436 220396
rect 60372 220108 60424 220114
rect 60372 220050 60424 220056
rect 60660 217410 60688 220390
rect 61856 217410 61884 224334
rect 62132 220794 62160 225558
rect 62120 220788 62172 220794
rect 62120 220730 62172 220736
rect 62580 220244 62632 220250
rect 62580 220186 62632 220192
rect 62592 217410 62620 220186
rect 55660 217382 55996 217410
rect 56488 217382 56548 217410
rect 57316 217382 57652 217410
rect 58144 217382 58480 217410
rect 58972 217382 59308 217410
rect 59800 217382 59860 217410
rect 60628 217382 60688 217410
rect 61456 217382 61884 217410
rect 62284 217382 62620 217410
rect 62776 217326 62804 311063
rect 64144 289876 64196 289882
rect 64144 289818 64196 289824
rect 64156 278322 64184 289818
rect 499592 278730 499790 278746
rect 406936 278724 406988 278730
rect 406936 278666 406988 278672
rect 499580 278724 499790 278730
rect 499632 278718 499790 278724
rect 499580 278666 499632 278672
rect 64144 278316 64196 278322
rect 64144 278258 64196 278264
rect 65904 271182 65932 277780
rect 67022 277766 67588 277794
rect 65892 271176 65944 271182
rect 65892 271118 65944 271124
rect 67560 270094 67588 277766
rect 68204 275466 68232 277780
rect 68192 275460 68244 275466
rect 68192 275402 68244 275408
rect 67548 270088 67600 270094
rect 67548 270030 67600 270036
rect 69400 269822 69428 277780
rect 70596 275330 70624 277780
rect 70584 275324 70636 275330
rect 70584 275266 70636 275272
rect 71792 274990 71820 277780
rect 71780 274984 71832 274990
rect 71780 274926 71832 274932
rect 72988 273970 73016 277780
rect 74092 275602 74120 277780
rect 75302 277766 75868 277794
rect 76498 277766 77248 277794
rect 74080 275596 74132 275602
rect 74080 275538 74132 275544
rect 73804 274984 73856 274990
rect 73804 274926 73856 274932
rect 72976 273964 73028 273970
rect 72976 273906 73028 273912
rect 69388 269816 69440 269822
rect 69388 269758 69440 269764
rect 73816 267034 73844 274926
rect 75840 269958 75868 277766
rect 75828 269952 75880 269958
rect 75828 269894 75880 269900
rect 77220 268802 77248 277766
rect 77680 277394 77708 277780
rect 77588 277366 77708 277394
rect 77588 274106 77616 277366
rect 77760 275596 77812 275602
rect 77760 275538 77812 275544
rect 77576 274100 77628 274106
rect 77576 274042 77628 274048
rect 77772 272542 77800 275538
rect 77760 272536 77812 272542
rect 77760 272478 77812 272484
rect 78876 270366 78904 277780
rect 78864 270360 78916 270366
rect 78864 270302 78916 270308
rect 80072 270094 80100 277780
rect 81268 274990 81296 277780
rect 82386 277766 82768 277794
rect 83582 277766 84148 277794
rect 81256 274984 81308 274990
rect 81256 274926 81308 274932
rect 78588 270088 78640 270094
rect 78588 270030 78640 270036
rect 80060 270088 80112 270094
rect 80060 270030 80112 270036
rect 77208 268796 77260 268802
rect 77208 268738 77260 268744
rect 73804 267028 73856 267034
rect 73804 266970 73856 266976
rect 78600 266490 78628 270030
rect 82740 268394 82768 277766
rect 84120 269550 84148 277766
rect 84764 271318 84792 277780
rect 85960 275602 85988 277780
rect 85948 275596 86000 275602
rect 85948 275538 86000 275544
rect 86224 274984 86276 274990
rect 86224 274926 86276 274932
rect 84752 271312 84804 271318
rect 84752 271254 84804 271260
rect 84108 269544 84160 269550
rect 84108 269486 84160 269492
rect 82728 268388 82780 268394
rect 82728 268330 82780 268336
rect 86236 267306 86264 274926
rect 87156 268530 87184 277780
rect 88366 277766 88656 277794
rect 88628 271726 88656 277766
rect 89548 274718 89576 277780
rect 90666 277766 91048 277794
rect 89536 274712 89588 274718
rect 89536 274654 89588 274660
rect 88616 271720 88668 271726
rect 88616 271662 88668 271668
rect 87144 268524 87196 268530
rect 87144 268466 87196 268472
rect 86224 267300 86276 267306
rect 86224 267242 86276 267248
rect 91020 267170 91048 277766
rect 91848 272678 91876 277780
rect 92480 274712 92532 274718
rect 92480 274654 92532 274660
rect 91836 272672 91888 272678
rect 91836 272614 91888 272620
rect 92492 271454 92520 274654
rect 93044 272406 93072 277780
rect 93032 272400 93084 272406
rect 93032 272342 93084 272348
rect 92480 271448 92532 271454
rect 92480 271390 92532 271396
rect 94240 270230 94268 277780
rect 94228 270224 94280 270230
rect 94228 270166 94280 270172
rect 95436 268666 95464 277780
rect 96632 274514 96660 277780
rect 96620 274508 96672 274514
rect 96620 274450 96672 274456
rect 97736 272814 97764 277780
rect 97724 272808 97776 272814
rect 97724 272750 97776 272756
rect 98932 271590 98960 277780
rect 100142 277766 100708 277794
rect 98920 271584 98972 271590
rect 98920 271526 98972 271532
rect 95424 268660 95476 268666
rect 95424 268602 95476 268608
rect 100680 267578 100708 277766
rect 101324 271862 101352 277780
rect 102520 274242 102548 277780
rect 103716 275738 103744 277780
rect 103704 275732 103756 275738
rect 103704 275674 103756 275680
rect 102508 274236 102560 274242
rect 102508 274178 102560 274184
rect 101312 271856 101364 271862
rect 101312 271798 101364 271804
rect 104912 268938 104940 277780
rect 106016 274666 106044 277780
rect 107212 275874 107240 277780
rect 108422 277766 108988 277794
rect 107200 275868 107252 275874
rect 107200 275810 107252 275816
rect 106016 274638 106320 274666
rect 104900 268932 104952 268938
rect 104900 268874 104952 268880
rect 106292 268802 106320 274638
rect 108960 270502 108988 277766
rect 109604 272950 109632 277780
rect 110800 276010 110828 277780
rect 110788 276004 110840 276010
rect 110788 275946 110840 275952
rect 111996 274378 112024 277780
rect 113192 275194 113220 277780
rect 113180 275188 113232 275194
rect 113180 275130 113232 275136
rect 111984 274372 112036 274378
rect 111984 274314 112036 274320
rect 109592 272944 109644 272950
rect 109592 272886 109644 272892
rect 114296 271046 114324 277780
rect 115506 277766 115888 277794
rect 114284 271040 114336 271046
rect 114284 270982 114336 270988
rect 108948 270496 109000 270502
rect 108948 270438 109000 270444
rect 104900 268796 104952 268802
rect 104900 268738 104952 268744
rect 106280 268796 106332 268802
rect 106280 268738 106332 268744
rect 100668 267572 100720 267578
rect 100668 267514 100720 267520
rect 91008 267164 91060 267170
rect 91008 267106 91060 267112
rect 104912 266898 104940 268738
rect 115860 268258 115888 277766
rect 116688 272270 116716 277780
rect 117898 277766 118648 277794
rect 116676 272264 116728 272270
rect 116676 272206 116728 272212
rect 118620 269074 118648 277766
rect 119080 274514 119108 277780
rect 120276 274650 120304 277780
rect 119344 274644 119396 274650
rect 119344 274586 119396 274592
rect 120264 274644 120316 274650
rect 120264 274586 120316 274592
rect 119068 274508 119120 274514
rect 119068 274450 119120 274456
rect 118608 269068 118660 269074
rect 118608 269010 118660 269016
rect 115848 268252 115900 268258
rect 115848 268194 115900 268200
rect 104900 266892 104952 266898
rect 104900 266834 104952 266840
rect 119356 266762 119384 274586
rect 121380 273086 121408 277780
rect 122590 277766 122788 277794
rect 121368 273080 121420 273086
rect 121368 273022 121420 273028
rect 122760 269686 122788 277766
rect 123772 270910 123800 277780
rect 124968 273698 124996 277780
rect 126178 277766 126928 277794
rect 124956 273692 125008 273698
rect 124956 273634 125008 273640
rect 123760 270904 123812 270910
rect 123760 270846 123812 270852
rect 122748 269680 122800 269686
rect 122748 269622 122800 269628
rect 126900 269550 126928 277766
rect 127360 273222 127388 277780
rect 127348 273216 127400 273222
rect 127348 273158 127400 273164
rect 126704 269544 126756 269550
rect 126704 269486 126756 269492
rect 126888 269544 126940 269550
rect 126888 269486 126940 269492
rect 119344 266756 119396 266762
rect 119344 266698 119396 266704
rect 126716 266626 126744 269486
rect 128556 269278 128584 277780
rect 129384 277766 129674 277794
rect 129384 269414 129412 277766
rect 130856 273834 130884 277780
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 130844 273828 130896 273834
rect 130844 273770 130896 273776
rect 129372 269408 129424 269414
rect 129372 269350 129424 269356
rect 128544 269272 128596 269278
rect 128544 269214 128596 269220
rect 132420 267714 132448 277766
rect 133800 270366 133828 277766
rect 134444 270774 134472 277780
rect 135260 275460 135312 275466
rect 135260 275402 135312 275408
rect 134432 270768 134484 270774
rect 134432 270710 134484 270716
rect 132592 270360 132644 270366
rect 132592 270302 132644 270308
rect 133788 270360 133840 270366
rect 133788 270302 133840 270308
rect 132408 267708 132460 267714
rect 132408 267650 132460 267656
rect 132604 267442 132632 270302
rect 135272 268122 135300 275402
rect 135640 274922 135668 277780
rect 136836 275466 136864 277780
rect 136824 275460 136876 275466
rect 136824 275402 136876 275408
rect 135628 274916 135680 274922
rect 135628 274858 135680 274864
rect 137940 272406 137968 277780
rect 137560 272400 137612 272406
rect 137560 272342 137612 272348
rect 137928 272400 137980 272406
rect 137928 272342 137980 272348
rect 136640 271176 136692 271182
rect 136640 271118 136692 271124
rect 135260 268116 135312 268122
rect 135260 268058 135312 268064
rect 132592 267436 132644 267442
rect 132592 267378 132644 267384
rect 126704 266620 126756 266626
rect 126704 266562 126756 266568
rect 78588 266484 78640 266490
rect 78588 266426 78640 266432
rect 136652 264316 136680 271118
rect 137572 266490 137600 272342
rect 139136 271182 139164 277780
rect 140346 277766 140728 277794
rect 139308 275324 139360 275330
rect 139308 275266 139360 275272
rect 139124 271176 139176 271182
rect 139124 271118 139176 271124
rect 138848 269816 138900 269822
rect 138848 269758 138900 269764
rect 138112 268116 138164 268122
rect 138112 268058 138164 268064
rect 137376 266484 137428 266490
rect 137376 266426 137428 266432
rect 137560 266484 137612 266490
rect 137560 266426 137612 266432
rect 137388 264316 137416 266426
rect 138124 264316 138152 268058
rect 138860 264316 138888 269758
rect 139320 267734 139348 275266
rect 140504 271176 140556 271182
rect 140504 271118 140556 271124
rect 139320 267706 139440 267734
rect 139412 264330 139440 267706
rect 140516 267034 140544 271118
rect 140700 269822 140728 277766
rect 141528 273970 141556 277780
rect 142724 275058 142752 277780
rect 142988 275188 143040 275194
rect 142988 275130 143040 275136
rect 142712 275052 142764 275058
rect 142712 274994 142764 275000
rect 140964 273964 141016 273970
rect 140964 273906 141016 273912
rect 141516 273964 141568 273970
rect 141516 273906 141568 273912
rect 140688 269816 140740 269822
rect 140688 269758 140740 269764
rect 140320 267028 140372 267034
rect 140320 266970 140372 266976
rect 140504 267028 140556 267034
rect 140504 266970 140556 266976
rect 139412 264302 139610 264330
rect 140332 264316 140360 266970
rect 140976 264330 141004 273906
rect 142160 272536 142212 272542
rect 142160 272478 142212 272484
rect 141792 269952 141844 269958
rect 141792 269894 141844 269900
rect 140976 264302 141082 264330
rect 141804 264316 141832 269894
rect 142172 264330 142200 272478
rect 143000 270638 143028 275130
rect 143632 274100 143684 274106
rect 143632 274042 143684 274048
rect 142988 270632 143040 270638
rect 142988 270574 143040 270580
rect 143264 266892 143316 266898
rect 143264 266834 143316 266840
rect 142172 264302 142554 264330
rect 143276 264316 143304 266834
rect 143644 264330 143672 274042
rect 143920 269958 143948 277780
rect 145024 271182 145052 277780
rect 145656 271720 145708 271726
rect 145656 271662 145708 271668
rect 145012 271176 145064 271182
rect 145012 271118 145064 271124
rect 144460 270088 144512 270094
rect 144460 270030 144512 270036
rect 143908 269952 143960 269958
rect 143908 269894 143960 269900
rect 144472 264330 144500 270030
rect 145668 267442 145696 271662
rect 145472 267436 145524 267442
rect 145472 267378 145524 267384
rect 145656 267436 145708 267442
rect 145656 267378 145708 267384
rect 143644 264302 144026 264330
rect 144472 264302 144762 264330
rect 145484 264316 145512 267378
rect 146220 267306 146248 277780
rect 147416 277394 147444 277780
rect 148626 277766 148916 277794
rect 147416 277366 147536 277394
rect 146944 268388 146996 268394
rect 146944 268330 146996 268336
rect 145932 267300 145984 267306
rect 145932 267242 145984 267248
rect 146208 267300 146260 267306
rect 146208 267242 146260 267248
rect 145944 264330 145972 267242
rect 146760 267164 146812 267170
rect 146760 267106 146812 267112
rect 146772 266898 146800 267106
rect 146760 266892 146812 266898
rect 146760 266834 146812 266840
rect 145944 264302 146234 264330
rect 146956 264316 146984 268330
rect 147508 268122 147536 277366
rect 147680 271312 147732 271318
rect 147680 271254 147732 271260
rect 147496 268116 147548 268122
rect 147496 268058 147548 268064
rect 147692 264316 147720 271254
rect 148888 268394 148916 277766
rect 149808 275602 149836 277780
rect 149060 275596 149112 275602
rect 149060 275538 149112 275544
rect 149796 275596 149848 275602
rect 149796 275538 149848 275544
rect 148876 268388 148928 268394
rect 148876 268330 148928 268336
rect 148416 266620 148468 266626
rect 148416 266562 148468 266568
rect 148428 264316 148456 266562
rect 149072 264330 149100 275538
rect 149704 273692 149756 273698
rect 149704 273634 149756 273640
rect 149716 267442 149744 273634
rect 151004 271454 151032 277780
rect 152200 275330 152228 277780
rect 153304 275466 153332 277780
rect 153844 275868 153896 275874
rect 153844 275810 153896 275816
rect 152740 275460 152792 275466
rect 152740 275402 152792 275408
rect 153292 275460 153344 275466
rect 153292 275402 153344 275408
rect 152188 275324 152240 275330
rect 152188 275266 152240 275272
rect 152372 272672 152424 272678
rect 152372 272614 152424 272620
rect 150440 271448 150492 271454
rect 150440 271390 150492 271396
rect 150992 271448 151044 271454
rect 150992 271390 151044 271396
rect 149888 268524 149940 268530
rect 149888 268466 149940 268472
rect 149520 267436 149572 267442
rect 149520 267378 149572 267384
rect 149704 267436 149756 267442
rect 149704 267378 149756 267384
rect 149532 267170 149560 267378
rect 149520 267164 149572 267170
rect 149520 267106 149572 267112
rect 149072 264302 149178 264330
rect 149900 264316 149928 268466
rect 150452 264330 150480 271390
rect 152384 267734 152412 272614
rect 152752 270094 152780 275402
rect 153568 270224 153620 270230
rect 153568 270166 153620 270172
rect 152740 270088 152792 270094
rect 152740 270030 152792 270036
rect 152384 267706 152504 267734
rect 151360 267164 151412 267170
rect 151360 267106 151412 267112
rect 150452 264302 150650 264330
rect 151372 264316 151400 267106
rect 152096 266892 152148 266898
rect 152096 266834 152148 266840
rect 152108 264316 152136 266834
rect 152476 264330 152504 267706
rect 152476 264302 152858 264330
rect 153580 264316 153608 270166
rect 153856 266898 153884 275810
rect 154500 272542 154528 277780
rect 155408 272808 155460 272814
rect 155408 272750 155460 272756
rect 154488 272536 154540 272542
rect 154488 272478 154540 272484
rect 155040 268660 155092 268666
rect 155040 268602 155092 268608
rect 153844 266892 153896 266898
rect 153844 266834 153896 266840
rect 154304 266484 154356 266490
rect 154304 266426 154356 266432
rect 154316 264316 154344 266426
rect 155052 264316 155080 268602
rect 155420 264330 155448 272750
rect 155696 271318 155724 277780
rect 156696 276004 156748 276010
rect 156696 275946 156748 275952
rect 156512 271584 156564 271590
rect 156512 271526 156564 271532
rect 155684 271312 155736 271318
rect 155684 271254 155736 271260
rect 156524 267734 156552 271526
rect 156708 267734 156736 275946
rect 156892 275194 156920 277780
rect 156880 275188 156932 275194
rect 156880 275130 156932 275136
rect 157892 274236 157944 274242
rect 157892 274178 157944 274184
rect 157616 271856 157668 271862
rect 157616 271798 157668 271804
rect 156524 267706 156644 267734
rect 156708 267706 156828 267734
rect 156236 266756 156288 266762
rect 156236 266698 156288 266704
rect 156248 264330 156276 266698
rect 156616 264602 156644 267706
rect 156800 266762 156828 267706
rect 156788 266756 156840 266762
rect 156788 266698 156840 266704
rect 156616 264574 156920 264602
rect 156892 264330 156920 264574
rect 157628 264330 157656 271798
rect 157904 266422 157932 274178
rect 158088 274106 158116 277780
rect 158720 274916 158772 274922
rect 158720 274858 158772 274864
rect 158076 274100 158128 274106
rect 158076 274042 158128 274048
rect 158732 267986 158760 274858
rect 159284 272678 159312 277780
rect 160480 275874 160508 277780
rect 160468 275868 160520 275874
rect 160468 275810 160520 275816
rect 160560 275732 160612 275738
rect 160560 275674 160612 275680
rect 159272 272672 159324 272678
rect 159272 272614 159324 272620
rect 159640 272264 159692 272270
rect 159640 272206 159692 272212
rect 158720 267980 158772 267986
rect 158720 267922 158772 267928
rect 158720 267572 158772 267578
rect 158720 267514 158772 267520
rect 157892 266416 157944 266422
rect 157892 266358 157944 266364
rect 155420 264302 155802 264330
rect 156248 264302 156538 264330
rect 156892 264302 157274 264330
rect 157628 264302 158010 264330
rect 158732 264316 158760 267514
rect 159652 266626 159680 272206
rect 160192 268932 160244 268938
rect 160192 268874 160244 268880
rect 159640 266620 159692 266626
rect 159640 266562 159692 266568
rect 159456 266416 159508 266422
rect 159456 266358 159508 266364
rect 159468 264316 159496 266358
rect 160204 264316 160232 268874
rect 160572 264330 160600 275674
rect 161584 274718 161612 277780
rect 162584 275324 162636 275330
rect 162584 275266 162636 275272
rect 161572 274712 161624 274718
rect 161572 274654 161624 274660
rect 161434 274644 161486 274650
rect 161434 274586 161486 274592
rect 161446 274530 161474 274586
rect 161446 274502 161520 274530
rect 161492 273698 161520 274502
rect 161480 273692 161532 273698
rect 161480 273634 161532 273640
rect 162400 270496 162452 270502
rect 162400 270438 162452 270444
rect 161664 268796 161716 268802
rect 161664 268738 161716 268744
rect 160572 264302 160954 264330
rect 161676 264316 161704 268738
rect 162412 264316 162440 270438
rect 162596 268666 162624 275266
rect 162584 268660 162636 268666
rect 162584 268602 162636 268608
rect 162780 268530 162808 277780
rect 163976 274718 164004 277780
rect 163688 274712 163740 274718
rect 163688 274654 163740 274660
rect 163964 274712 164016 274718
rect 163964 274654 164016 274660
rect 163412 272944 163464 272950
rect 163412 272886 163464 272892
rect 162768 268524 162820 268530
rect 162768 268466 162820 268472
rect 163424 267734 163452 272886
rect 163700 270230 163728 274654
rect 164240 274372 164292 274378
rect 164240 274314 164292 274320
rect 163688 270224 163740 270230
rect 163688 270166 163740 270172
rect 163596 269272 163648 269278
rect 163596 269214 163648 269220
rect 163608 267734 163636 269214
rect 163424 267706 163544 267734
rect 163608 267706 163728 267734
rect 163136 266892 163188 266898
rect 163136 266834 163188 266840
rect 163148 264316 163176 266834
rect 163516 264330 163544 267706
rect 163700 266898 163728 267706
rect 163688 266892 163740 266898
rect 163688 266834 163740 266840
rect 164252 264330 164280 274314
rect 165172 271590 165200 277780
rect 166172 275188 166224 275194
rect 166172 275130 166224 275136
rect 166184 274122 166212 275130
rect 166368 274242 166396 277780
rect 167564 275330 167592 277780
rect 167552 275324 167604 275330
rect 167552 275266 167604 275272
rect 167644 274712 167696 274718
rect 167644 274654 167696 274660
rect 166356 274236 166408 274242
rect 166356 274178 166408 274184
rect 166184 274094 166304 274122
rect 165160 271584 165212 271590
rect 165160 271526 165212 271532
rect 165712 270632 165764 270638
rect 165712 270574 165764 270580
rect 165344 266756 165396 266762
rect 165344 266698 165396 266704
rect 163516 264302 163898 264330
rect 164252 264302 164634 264330
rect 165356 264316 165384 266698
rect 165724 264330 165752 270574
rect 166080 269544 166132 269550
rect 166080 269486 166132 269492
rect 166092 269278 166120 269486
rect 166080 269272 166132 269278
rect 166080 269214 166132 269220
rect 166276 267578 166304 274094
rect 167184 271040 167236 271046
rect 167184 270982 167236 270988
rect 166448 270224 166500 270230
rect 166448 270166 166500 270172
rect 166460 269686 166488 270166
rect 166448 269680 166500 269686
rect 166448 269622 166500 269628
rect 166816 268252 166868 268258
rect 166816 268194 166868 268200
rect 166264 267572 166316 267578
rect 166264 267514 166316 267520
rect 165724 264302 166106 264330
rect 166828 264316 166856 268194
rect 167196 264330 167224 270982
rect 167656 267170 167684 274654
rect 168472 274508 168524 274514
rect 168472 274450 168524 274456
rect 168484 267734 168512 274450
rect 168668 272814 168696 277780
rect 169878 277766 170168 277794
rect 169760 275052 169812 275058
rect 169760 274994 169812 275000
rect 169772 274514 169800 274994
rect 169760 274508 169812 274514
rect 169760 274450 169812 274456
rect 169944 273692 169996 273698
rect 169944 273634 169996 273640
rect 168656 272808 168708 272814
rect 168656 272750 168708 272756
rect 169760 269068 169812 269074
rect 169760 269010 169812 269016
rect 168484 267706 168696 267734
rect 167644 267164 167696 267170
rect 167644 267106 167696 267112
rect 168288 266620 168340 266626
rect 168288 266562 168340 266568
rect 167196 264302 167578 264330
rect 168300 264316 168328 266562
rect 168668 264330 168696 267706
rect 168668 264302 169050 264330
rect 169772 264316 169800 269010
rect 169956 267734 169984 273634
rect 170140 271726 170168 277766
rect 171060 276010 171088 277780
rect 172270 277766 172468 277794
rect 173466 277766 173848 277794
rect 171048 276004 171100 276010
rect 171048 275946 171100 275952
rect 171600 273080 171652 273086
rect 171600 273022 171652 273028
rect 170128 271720 170180 271726
rect 170128 271662 170180 271668
rect 171232 269544 171284 269550
rect 171232 269486 171284 269492
rect 169956 267706 170168 267734
rect 170140 264330 170168 267706
rect 170140 264302 170522 264330
rect 171244 264316 171272 269486
rect 171612 264330 171640 273022
rect 172440 270230 172468 277766
rect 172704 270904 172756 270910
rect 172704 270846 172756 270852
rect 172428 270224 172480 270230
rect 172428 270166 172480 270172
rect 171612 264302 171994 264330
rect 172716 264316 172744 270846
rect 173532 269816 173584 269822
rect 173532 269758 173584 269764
rect 173820 269770 173848 277766
rect 174452 275868 174504 275874
rect 174452 275810 174504 275816
rect 174464 273086 174492 275810
rect 174648 275738 174676 277780
rect 175844 276010 175872 277780
rect 175832 276004 175884 276010
rect 175832 275946 175884 275952
rect 175924 275868 175976 275874
rect 175924 275810 175976 275816
rect 174636 275732 174688 275738
rect 174636 275674 174688 275680
rect 174636 273216 174688 273222
rect 174636 273158 174688 273164
rect 174452 273080 174504 273086
rect 174452 273022 174504 273028
rect 173544 269550 173572 269758
rect 173820 269742 173940 269770
rect 173912 269686 173940 269742
rect 173900 269680 173952 269686
rect 173900 269622 173952 269628
rect 173532 269544 173584 269550
rect 173532 269486 173584 269492
rect 173440 269272 173492 269278
rect 173440 269214 173492 269220
rect 173452 264316 173480 269214
rect 174176 267436 174228 267442
rect 174176 267378 174228 267384
rect 174188 264316 174216 267378
rect 174648 264330 174676 273158
rect 175648 269408 175700 269414
rect 175648 269350 175700 269356
rect 174648 264302 174938 264330
rect 175660 264316 175688 269350
rect 175936 266762 175964 275810
rect 176752 273828 176804 273834
rect 176752 273770 176804 273776
rect 176384 266892 176436 266898
rect 176384 266834 176436 266840
rect 175924 266756 175976 266762
rect 175924 266698 175976 266704
rect 176396 264316 176424 266834
rect 176764 264330 176792 273770
rect 176948 270502 176976 277780
rect 177856 276004 177908 276010
rect 177856 275946 177908 275952
rect 177868 274378 177896 275946
rect 178144 274718 178172 277780
rect 179156 277766 179354 277794
rect 180550 277766 180748 277794
rect 178132 274712 178184 274718
rect 178132 274654 178184 274660
rect 177856 274372 177908 274378
rect 177856 274314 177908 274320
rect 179156 271862 179184 277766
rect 179972 275596 180024 275602
rect 179972 275538 180024 275544
rect 179328 274712 179380 274718
rect 179328 274654 179380 274660
rect 179144 271856 179196 271862
rect 179144 271798 179196 271804
rect 178960 270768 179012 270774
rect 178960 270710 179012 270716
rect 176936 270496 176988 270502
rect 176936 270438 176988 270444
rect 177580 270360 177632 270366
rect 177580 270302 177632 270308
rect 177592 264330 177620 270302
rect 178592 267708 178644 267714
rect 178592 267650 178644 267656
rect 176764 264302 177146 264330
rect 177592 264302 177882 264330
rect 178604 264316 178632 267650
rect 178972 264330 179000 270710
rect 179144 270496 179196 270502
rect 179144 270438 179196 270444
rect 179156 270230 179184 270438
rect 179144 270224 179196 270230
rect 179144 270166 179196 270172
rect 179340 267442 179368 274654
rect 179512 270224 179564 270230
rect 179512 270166 179564 270172
rect 179524 269686 179552 270166
rect 179788 270088 179840 270094
rect 179788 270030 179840 270036
rect 179512 269680 179564 269686
rect 179512 269622 179564 269628
rect 179328 267436 179380 267442
rect 179328 267378 179380 267384
rect 179800 264330 179828 270030
rect 179984 269686 180012 275538
rect 180720 274666 180748 277766
rect 181732 275602 181760 277780
rect 182942 277766 183508 277794
rect 181720 275596 181772 275602
rect 181720 275538 181772 275544
rect 180720 274638 180840 274666
rect 180812 272950 180840 274638
rect 180800 272944 180852 272950
rect 180800 272886 180852 272892
rect 181168 272400 181220 272406
rect 181168 272342 181220 272348
rect 179972 269680 180024 269686
rect 179972 269622 180024 269628
rect 180800 267980 180852 267986
rect 180800 267922 180852 267928
rect 178972 264302 179354 264330
rect 179800 264302 180090 264330
rect 180812 264316 180840 267922
rect 181180 264330 181208 272342
rect 183480 270094 183508 277766
rect 184124 273970 184152 277780
rect 185228 274718 185256 277780
rect 185584 275460 185636 275466
rect 185584 275402 185636 275408
rect 185216 274712 185268 274718
rect 185216 274654 185268 274660
rect 185124 274508 185176 274514
rect 185124 274450 185176 274456
rect 183744 273964 183796 273970
rect 183744 273906 183796 273912
rect 184112 273964 184164 273970
rect 184112 273906 184164 273912
rect 183468 270088 183520 270094
rect 183468 270030 183520 270036
rect 182272 269544 182324 269550
rect 182272 269486 182324 269492
rect 181180 264302 181562 264330
rect 182284 264316 182312 269486
rect 183008 267028 183060 267034
rect 183008 266970 183060 266976
rect 183020 264316 183048 266970
rect 183756 264316 183784 273906
rect 184940 271176 184992 271182
rect 184940 271118 184992 271124
rect 184480 269952 184532 269958
rect 184480 269894 184532 269900
rect 184492 264316 184520 269894
rect 184952 265946 184980 271118
rect 184940 265940 184992 265946
rect 184940 265882 184992 265888
rect 185136 264330 185164 274450
rect 185596 271182 185624 275402
rect 186424 274990 186452 277780
rect 186412 274984 186464 274990
rect 186412 274926 186464 274932
rect 186964 274712 187016 274718
rect 186964 274654 187016 274660
rect 185584 271176 185636 271182
rect 185584 271118 185636 271124
rect 186688 268116 186740 268122
rect 186688 268058 186740 268064
rect 185676 265940 185728 265946
rect 185676 265882 185728 265888
rect 185688 264330 185716 265882
rect 185136 264302 185242 264330
rect 185688 264302 185978 264330
rect 186700 264316 186728 268058
rect 186976 267034 187004 274654
rect 187620 268802 187648 277780
rect 188816 275466 188844 277780
rect 190026 277766 190408 277794
rect 191222 277766 191696 277794
rect 188804 275460 188856 275466
rect 188804 275402 188856 275408
rect 188068 274984 188120 274990
rect 188068 274926 188120 274932
rect 187608 268796 187660 268802
rect 187608 268738 187660 268744
rect 188080 268394 188108 274926
rect 188252 271448 188304 271454
rect 188252 271390 188304 271396
rect 187884 268388 187936 268394
rect 187884 268330 187936 268336
rect 188068 268388 188120 268394
rect 188068 268330 188120 268336
rect 187424 267300 187476 267306
rect 187424 267242 187476 267248
rect 186964 267028 187016 267034
rect 186964 266970 187016 266976
rect 187436 264316 187464 267242
rect 187896 264330 187924 268330
rect 188264 267734 188292 271390
rect 189632 269680 189684 269686
rect 189632 269622 189684 269628
rect 188264 267706 188568 267734
rect 188540 264330 188568 267706
rect 187896 264302 188186 264330
rect 188540 264302 188922 264330
rect 189644 264316 189672 269622
rect 190380 268666 190408 277766
rect 190736 272536 190788 272542
rect 190736 272478 190788 272484
rect 190092 268660 190144 268666
rect 190092 268602 190144 268608
rect 190368 268660 190420 268666
rect 190368 268602 190420 268608
rect 190104 264330 190132 268602
rect 190748 264330 190776 272478
rect 191668 269958 191696 277766
rect 192312 277394 192340 277780
rect 192312 277366 192432 277394
rect 192208 271312 192260 271318
rect 192208 271254 192260 271260
rect 191840 271176 191892 271182
rect 191840 271118 191892 271124
rect 191656 269952 191708 269958
rect 191656 269894 191708 269900
rect 190104 264302 190394 264330
rect 190748 264302 191130 264330
rect 191852 264316 191880 271118
rect 192220 264330 192248 271254
rect 192404 271182 192432 277366
rect 193312 274100 193364 274106
rect 193312 274042 193364 274048
rect 192392 271176 192444 271182
rect 192392 271118 192444 271124
rect 192220 264302 192602 264330
rect 193324 264316 193352 274042
rect 193508 271318 193536 277780
rect 194704 275126 194732 277780
rect 195716 277766 195914 277794
rect 194692 275120 194744 275126
rect 194692 275062 194744 275068
rect 195716 272678 195744 277766
rect 195888 275120 195940 275126
rect 195888 275062 195940 275068
rect 194784 272672 194836 272678
rect 194784 272614 194836 272620
rect 195704 272672 195756 272678
rect 195704 272614 195756 272620
rect 193496 271312 193548 271318
rect 193496 271254 193548 271260
rect 194508 270088 194560 270094
rect 194508 270030 194560 270036
rect 194048 267572 194100 267578
rect 194048 267514 194100 267520
rect 194060 264316 194088 267514
rect 194520 267306 194548 270030
rect 194508 267300 194560 267306
rect 194508 267242 194560 267248
rect 194796 264316 194824 272614
rect 195900 269822 195928 275062
rect 196164 273080 196216 273086
rect 196164 273022 196216 273028
rect 195520 269816 195572 269822
rect 195520 269758 195572 269764
rect 195888 269816 195940 269822
rect 195888 269758 195940 269764
rect 195532 264316 195560 269758
rect 196176 264330 196204 273022
rect 197096 272542 197124 277780
rect 197544 275732 197596 275738
rect 197544 275674 197596 275680
rect 197084 272536 197136 272542
rect 197084 272478 197136 272484
rect 197360 271584 197412 271590
rect 197360 271526 197412 271532
rect 196992 268524 197044 268530
rect 196992 268466 197044 268472
rect 196176 264302 196282 264330
rect 197004 264316 197032 268466
rect 197372 264330 197400 271526
rect 197556 269686 197584 275674
rect 198292 274106 198320 277780
rect 199488 275738 199516 277780
rect 199476 275732 199528 275738
rect 199476 275674 199528 275680
rect 200028 275324 200080 275330
rect 200028 275266 200080 275272
rect 200040 274530 200068 275266
rect 200040 274502 200252 274530
rect 198924 274236 198976 274242
rect 198924 274178 198976 274184
rect 198280 274100 198332 274106
rect 198280 274042 198332 274048
rect 198740 272808 198792 272814
rect 198740 272750 198792 272756
rect 197544 269680 197596 269686
rect 197544 269622 197596 269628
rect 198464 267164 198516 267170
rect 198464 267106 198516 267112
rect 197372 264302 197754 264330
rect 198476 264316 198504 267106
rect 198752 265946 198780 272750
rect 198740 265940 198792 265946
rect 198740 265882 198792 265888
rect 198936 264330 198964 274178
rect 200224 267734 200252 274502
rect 200592 274242 200620 277780
rect 200580 274236 200632 274242
rect 200580 274178 200632 274184
rect 201040 271720 201092 271726
rect 201040 271662 201092 271668
rect 200224 267706 200344 267734
rect 199660 265940 199712 265946
rect 199660 265882 199712 265888
rect 199672 264330 199700 265882
rect 200316 264330 200344 267706
rect 201052 264330 201080 271662
rect 201788 271454 201816 277780
rect 201776 271448 201828 271454
rect 201776 271390 201828 271396
rect 202144 270496 202196 270502
rect 202144 270438 202196 270444
rect 198936 264302 199226 264330
rect 199672 264302 199962 264330
rect 200316 264302 200698 264330
rect 201052 264302 201434 264330
rect 202156 264316 202184 270438
rect 202984 270094 203012 277780
rect 203904 277766 204194 277794
rect 205390 277766 205588 277794
rect 203616 270224 203668 270230
rect 203616 270166 203668 270172
rect 202972 270088 203024 270094
rect 202972 270030 203024 270036
rect 203340 268660 203392 268666
rect 203340 268602 203392 268608
rect 203352 267578 203380 268602
rect 203340 267572 203392 267578
rect 203340 267514 203392 267520
rect 202880 266892 202932 266898
rect 202880 266834 202932 266840
rect 202892 264316 202920 266834
rect 203628 264316 203656 270166
rect 203904 268938 203932 277766
rect 204260 274372 204312 274378
rect 204260 274314 204312 274320
rect 203892 268932 203944 268938
rect 203892 268874 203944 268880
rect 204272 264330 204300 274314
rect 204904 271856 204956 271862
rect 204904 271798 204956 271804
rect 204916 266422 204944 271798
rect 205560 270230 205588 277766
rect 206572 273970 206600 277780
rect 207020 275596 207072 275602
rect 207020 275538 207072 275544
rect 206284 273964 206336 273970
rect 206284 273906 206336 273912
rect 206560 273964 206612 273970
rect 206560 273906 206612 273912
rect 205824 270360 205876 270366
rect 205824 270302 205876 270308
rect 205548 270224 205600 270230
rect 205548 270166 205600 270172
rect 205088 269680 205140 269686
rect 205088 269622 205140 269628
rect 204904 266416 204956 266422
rect 204904 266358 204956 266364
rect 204272 264302 204378 264330
rect 205100 264316 205128 269622
rect 205836 264316 205864 270302
rect 206296 266694 206324 273906
rect 207032 270502 207060 275538
rect 207768 274990 207796 277780
rect 207756 274984 207808 274990
rect 207756 274926 207808 274932
rect 208400 274984 208452 274990
rect 208400 274926 208452 274932
rect 207480 272944 207532 272950
rect 207480 272886 207532 272892
rect 207020 270496 207072 270502
rect 207020 270438 207072 270444
rect 207492 267734 207520 272886
rect 208412 270366 208440 274926
rect 208400 270360 208452 270366
rect 208400 270302 208452 270308
rect 208492 268796 208544 268802
rect 208492 268738 208544 268744
rect 207492 267706 207704 267734
rect 207296 267436 207348 267442
rect 207296 267378 207348 267384
rect 206284 266688 206336 266694
rect 206284 266630 206336 266636
rect 206560 266416 206612 266422
rect 206560 266358 206612 266364
rect 206572 264316 206600 266358
rect 207308 264316 207336 267378
rect 207676 264330 207704 267706
rect 208504 266422 208532 268738
rect 208872 268530 208900 277780
rect 210068 275398 210096 277780
rect 210884 275732 210936 275738
rect 210884 275674 210936 275680
rect 210056 275392 210108 275398
rect 210056 275334 210108 275340
rect 209504 270496 209556 270502
rect 209504 270438 209556 270444
rect 208860 268524 208912 268530
rect 208860 268466 208912 268472
rect 208768 267300 208820 267306
rect 208768 267242 208820 267248
rect 208492 266416 208544 266422
rect 208492 266358 208544 266364
rect 207676 264302 208058 264330
rect 208780 264316 208808 267242
rect 209516 264316 209544 270438
rect 209872 268864 209924 268870
rect 209872 268806 209924 268812
rect 209884 267170 209912 268806
rect 210896 268394 210924 275674
rect 211264 275262 211292 277780
rect 212276 277766 212474 277794
rect 211252 275256 211304 275262
rect 211252 275198 211304 275204
rect 212276 269958 212304 277766
rect 212448 275256 212500 275262
rect 212448 275198 212500 275204
rect 211160 269952 211212 269958
rect 211160 269894 211212 269900
rect 212264 269952 212316 269958
rect 212264 269894 212316 269900
rect 210884 268388 210936 268394
rect 210884 268330 210936 268336
rect 210976 268252 211028 268258
rect 210976 268194 211028 268200
rect 209872 267164 209924 267170
rect 209872 267106 209924 267112
rect 210240 266688 210292 266694
rect 210240 266630 210292 266636
rect 210252 264316 210280 266630
rect 210988 264316 211016 268194
rect 211172 266558 211200 269894
rect 212460 267034 212488 275198
rect 213184 274236 213236 274242
rect 213184 274178 213236 274184
rect 213196 267714 213224 274178
rect 213656 271590 213684 277780
rect 213920 275528 213972 275534
rect 213920 275470 213972 275476
rect 213644 271584 213696 271590
rect 213644 271526 213696 271532
rect 213184 267708 213236 267714
rect 213184 267650 213236 267656
rect 213184 267572 213236 267578
rect 213184 267514 213236 267520
rect 211712 267028 211764 267034
rect 211712 266970 211764 266976
rect 212448 267028 212500 267034
rect 212448 266970 212500 266976
rect 211160 266552 211212 266558
rect 211160 266494 211212 266500
rect 211724 264316 211752 266970
rect 212448 266416 212500 266422
rect 212448 266358 212500 266364
rect 212460 264316 212488 266358
rect 213196 264316 213224 267514
rect 213932 264316 213960 275470
rect 214852 274854 214880 277780
rect 214840 274848 214892 274854
rect 214840 274790 214892 274796
rect 215760 271312 215812 271318
rect 215760 271254 215812 271260
rect 215300 271176 215352 271182
rect 215300 271118 215352 271124
rect 214656 266552 214708 266558
rect 214656 266494 214708 266500
rect 214668 264316 214696 266494
rect 215312 264330 215340 271118
rect 215772 264330 215800 271254
rect 215956 271182 215984 277780
rect 217166 277766 217456 277794
rect 217428 272678 217456 277766
rect 217232 272672 217284 272678
rect 217232 272614 217284 272620
rect 217416 272672 217468 272678
rect 217416 272614 217468 272620
rect 215944 271176 215996 271182
rect 215944 271118 215996 271124
rect 216864 269816 216916 269822
rect 216864 269758 216916 269764
rect 215312 264302 215418 264330
rect 215772 264302 216154 264330
rect 216876 264316 216904 269758
rect 217244 264330 217272 272614
rect 218348 272542 218376 277780
rect 219544 277394 219572 277780
rect 219544 277366 219664 277394
rect 218704 274100 218756 274106
rect 218704 274042 218756 274048
rect 218060 272536 218112 272542
rect 218060 272478 218112 272484
rect 218336 272536 218388 272542
rect 218336 272478 218388 272484
rect 218072 264330 218100 272478
rect 218716 264330 218744 274042
rect 219636 269958 219664 277366
rect 219440 269952 219492 269958
rect 219440 269894 219492 269900
rect 219624 269952 219676 269958
rect 219624 269894 219676 269900
rect 219452 266422 219480 269894
rect 220740 268394 220768 277780
rect 221740 274848 221792 274854
rect 221740 274790 221792 274796
rect 221004 271448 221056 271454
rect 221004 271390 221056 271396
rect 219808 268388 219860 268394
rect 219808 268330 219860 268336
rect 220728 268388 220780 268394
rect 220728 268330 220780 268336
rect 219440 266416 219492 266422
rect 219440 266358 219492 266364
rect 217244 264302 217626 264330
rect 218072 264302 218362 264330
rect 218716 264302 219098 264330
rect 219820 264316 219848 268330
rect 220544 267708 220596 267714
rect 220544 267650 220596 267656
rect 220556 264316 220584 267650
rect 221016 264330 221044 271390
rect 221752 270502 221780 274790
rect 221936 271318 221964 277780
rect 223146 277766 223344 277794
rect 221924 271312 221976 271318
rect 221924 271254 221976 271260
rect 221740 270496 221792 270502
rect 221740 270438 221792 270444
rect 222016 270088 222068 270094
rect 222016 270030 222068 270036
rect 221016 264302 221306 264330
rect 222028 264316 222056 270030
rect 223316 269822 223344 277766
rect 224236 273970 224264 277780
rect 223856 273964 223908 273970
rect 223856 273906 223908 273912
rect 224224 273964 224276 273970
rect 224224 273906 224276 273912
rect 223488 270224 223540 270230
rect 223488 270166 223540 270172
rect 223304 269816 223356 269822
rect 223304 269758 223356 269764
rect 222752 267164 222804 267170
rect 222752 267106 222804 267112
rect 222764 264316 222792 267106
rect 223500 264316 223528 270166
rect 223868 264330 223896 273906
rect 224960 270360 225012 270366
rect 224960 270302 225012 270308
rect 223868 264302 224250 264330
rect 224972 264316 225000 270302
rect 225432 269074 225460 277780
rect 226432 275392 226484 275398
rect 226432 275334 226484 275340
rect 226444 269906 226472 275334
rect 226628 270094 226656 277780
rect 227824 275330 227852 277780
rect 227812 275324 227864 275330
rect 227812 275266 227864 275272
rect 228272 271584 228324 271590
rect 228272 271526 228324 271532
rect 226616 270088 226668 270094
rect 226616 270030 226668 270036
rect 227720 269952 227772 269958
rect 226444 269878 226564 269906
rect 227720 269894 227772 269900
rect 225420 269068 225472 269074
rect 225420 269010 225472 269016
rect 226340 269068 226392 269074
rect 226340 269010 226392 269016
rect 225696 268524 225748 268530
rect 225696 268466 225748 268472
rect 225708 264316 225736 268466
rect 226352 267034 226380 269010
rect 226340 267028 226392 267034
rect 226340 266970 226392 266976
rect 226536 265962 226564 269878
rect 227732 267170 227760 269894
rect 227720 267164 227772 267170
rect 227720 267106 227772 267112
rect 227168 266892 227220 266898
rect 227168 266834 227220 266840
rect 226444 265934 226564 265962
rect 226444 264316 226472 265934
rect 227180 264316 227208 266834
rect 227904 266416 227956 266422
rect 227904 266358 227956 266364
rect 227916 264316 227944 266358
rect 228284 264330 228312 271526
rect 229020 271454 229048 277780
rect 230230 277766 230428 277794
rect 229008 271448 229060 271454
rect 229008 271390 229060 271396
rect 229744 271176 229796 271182
rect 229744 271118 229796 271124
rect 229376 270496 229428 270502
rect 229376 270438 229428 270444
rect 228284 264302 228666 264330
rect 229388 264316 229416 270438
rect 229756 264330 229784 271118
rect 230400 269958 230428 277766
rect 230664 272672 230716 272678
rect 230664 272614 230716 272620
rect 230388 269952 230440 269958
rect 230388 269894 230440 269900
rect 230676 264330 230704 272614
rect 231412 272542 231440 277780
rect 231216 272536 231268 272542
rect 231216 272478 231268 272484
rect 231400 272536 231452 272542
rect 231400 272478 231452 272484
rect 231228 264330 231256 272478
rect 232516 271862 232544 277780
rect 232504 271856 232556 271862
rect 232504 271798 232556 271804
rect 232504 271312 232556 271318
rect 232504 271254 232556 271260
rect 232320 267164 232372 267170
rect 232320 267106 232372 267112
rect 229756 264302 230138 264330
rect 230676 264302 230874 264330
rect 231228 264302 231610 264330
rect 232332 264316 232360 267106
rect 232516 266422 232544 271254
rect 233712 271182 233740 277780
rect 234908 274174 234936 277780
rect 236104 275466 236132 277780
rect 237300 277394 237328 277780
rect 237208 277366 237328 277394
rect 236092 275460 236144 275466
rect 236092 275402 236144 275408
rect 234896 274168 234948 274174
rect 234896 274110 234948 274116
rect 234896 273964 234948 273970
rect 234896 273906 234948 273912
rect 233884 271856 233936 271862
rect 233884 271798 233936 271804
rect 233700 271176 233752 271182
rect 233700 271118 233752 271124
rect 233056 268388 233108 268394
rect 233056 268330 233108 268336
rect 232504 266416 232556 266422
rect 232504 266358 232556 266364
rect 233068 264316 233096 268330
rect 233896 267442 233924 271798
rect 234528 269816 234580 269822
rect 234528 269758 234580 269764
rect 233884 267436 233936 267442
rect 233884 267378 233936 267384
rect 233792 266416 233844 266422
rect 233792 266358 233844 266364
rect 233804 264316 233832 266358
rect 234540 264316 234568 269758
rect 234908 264330 234936 273906
rect 236736 270088 236788 270094
rect 236736 270030 236788 270036
rect 236000 267028 236052 267034
rect 236000 266970 236052 266976
rect 234908 264302 235290 264330
rect 236012 264316 236040 266970
rect 236748 264316 236776 270030
rect 237208 269822 237236 277366
rect 238496 275330 238524 277780
rect 239600 277394 239628 277780
rect 240810 277766 241376 277794
rect 239600 277366 239720 277394
rect 237380 275324 237432 275330
rect 237380 275266 237432 275272
rect 238484 275324 238536 275330
rect 238484 275266 238536 275272
rect 237196 269816 237248 269822
rect 237196 269758 237248 269764
rect 237392 264330 237420 275266
rect 239496 274168 239548 274174
rect 239496 274110 239548 274116
rect 239312 272536 239364 272542
rect 239312 272478 239364 272484
rect 237840 271448 237892 271454
rect 237840 271390 237892 271396
rect 237852 264330 237880 271390
rect 238944 269952 238996 269958
rect 238944 269894 238996 269900
rect 237392 264302 237498 264330
rect 237852 264302 238234 264330
rect 238956 264316 238984 269894
rect 239324 264330 239352 272478
rect 239508 266422 239536 274110
rect 239692 272610 239720 277366
rect 239680 272604 239732 272610
rect 239680 272546 239732 272552
rect 240784 271176 240836 271182
rect 240784 271118 240836 271124
rect 240416 267436 240468 267442
rect 240416 267378 240468 267384
rect 239496 266416 239548 266422
rect 239496 266358 239548 266364
rect 239324 264302 239706 264330
rect 240428 264316 240456 267378
rect 240796 264330 240824 271118
rect 241348 266558 241376 277766
rect 241992 274718 242020 277780
rect 242256 275460 242308 275466
rect 242256 275402 242308 275408
rect 241980 274712 242032 274718
rect 241980 274654 242032 274660
rect 241336 266552 241388 266558
rect 241336 266494 241388 266500
rect 241888 266416 241940 266422
rect 241888 266358 241940 266364
rect 240796 264302 241178 264330
rect 241900 264316 241928 266358
rect 242268 264330 242296 275402
rect 243188 270366 243216 277780
rect 243728 275324 243780 275330
rect 243728 275266 243780 275272
rect 243176 270360 243228 270366
rect 243176 270302 243228 270308
rect 243360 269816 243412 269822
rect 243360 269758 243412 269764
rect 242268 264302 242650 264330
rect 243372 264316 243400 269758
rect 243740 264330 243768 275266
rect 244384 270502 244412 277780
rect 245580 275194 245608 277780
rect 245568 275188 245620 275194
rect 245568 275130 245620 275136
rect 246304 275188 246356 275194
rect 246304 275130 246356 275136
rect 246028 274712 246080 274718
rect 246028 274654 246080 274660
rect 244556 272604 244608 272610
rect 244556 272546 244608 272552
rect 244372 270496 244424 270502
rect 244372 270438 244424 270444
rect 244568 264330 244596 272546
rect 245568 266552 245620 266558
rect 245568 266494 245620 266500
rect 243740 264302 244122 264330
rect 244568 264302 244858 264330
rect 245580 264316 245608 266494
rect 246040 264330 246068 274654
rect 246316 266626 246344 275130
rect 246776 274718 246804 277780
rect 247894 277766 248368 277794
rect 246764 274712 246816 274718
rect 246764 274654 246816 274660
rect 247776 270496 247828 270502
rect 247776 270438 247828 270444
rect 247040 270360 247092 270366
rect 247040 270302 247092 270308
rect 246304 266620 246356 266626
rect 246304 266562 246356 266568
rect 246040 264302 246330 264330
rect 247052 264316 247080 270302
rect 247788 264316 247816 270438
rect 248340 269142 248368 277766
rect 249076 275058 249104 277780
rect 250272 277394 250300 277780
rect 250180 277366 250300 277394
rect 251192 277766 251482 277794
rect 249064 275052 249116 275058
rect 249064 274994 249116 275000
rect 248880 274712 248932 274718
rect 248880 274654 248932 274660
rect 248328 269136 248380 269142
rect 248328 269078 248380 269084
rect 248512 266620 248564 266626
rect 248512 266562 248564 266568
rect 248524 264316 248552 266562
rect 248892 264330 248920 274654
rect 250180 270502 250208 277366
rect 250352 275052 250404 275058
rect 250352 274994 250404 275000
rect 250168 270496 250220 270502
rect 250168 270438 250220 270444
rect 249984 269136 250036 269142
rect 249984 269078 250036 269084
rect 248892 264302 249274 264330
rect 249996 264316 250024 269078
rect 250364 264330 250392 274994
rect 251192 266422 251220 277766
rect 251456 270496 251508 270502
rect 251456 270438 251508 270444
rect 251180 266416 251232 266422
rect 251180 266358 251232 266364
rect 250364 264302 250746 264330
rect 251468 264316 251496 270438
rect 252192 266416 252244 266422
rect 252192 266358 252244 266364
rect 252204 264316 252232 266358
rect 252664 264330 252692 277780
rect 253032 277766 253874 277794
rect 254412 277766 255070 277794
rect 255332 277766 256174 277794
rect 256712 277766 257370 277794
rect 258092 277766 258566 277794
rect 259472 277766 259762 277794
rect 253032 267734 253060 277766
rect 253032 267706 253336 267734
rect 253308 264330 253336 267706
rect 252664 264302 252954 264330
rect 253308 264302 253690 264330
rect 254412 264316 254440 277766
rect 255332 267734 255360 277766
rect 255148 267706 255360 267734
rect 255148 264316 255176 267706
rect 256516 266892 256568 266898
rect 256516 266834 256568 266840
rect 255872 266416 255924 266422
rect 255872 266358 255924 266364
rect 255884 264316 255912 266358
rect 256528 264330 256556 266834
rect 256712 266422 256740 277766
rect 257344 267300 257396 267306
rect 257344 267242 257396 267248
rect 256700 266416 256752 266422
rect 256700 266358 256752 266364
rect 256528 264302 256634 264330
rect 257356 264316 257384 267242
rect 258092 266898 258120 277766
rect 258816 270496 258868 270502
rect 258816 270438 258868 270444
rect 258080 266892 258132 266898
rect 258080 266834 258132 266840
rect 258080 266416 258132 266422
rect 258080 266358 258132 266364
rect 258092 264316 258120 266358
rect 258828 264316 258856 270438
rect 259472 267306 259500 277766
rect 260944 277394 260972 277780
rect 260852 277366 260972 277394
rect 261312 277766 262154 277794
rect 262600 277766 263258 277794
rect 263612 277766 264454 277794
rect 264992 277766 265650 277794
rect 266372 277766 266846 277794
rect 260852 269482 260880 277366
rect 261312 270502 261340 277766
rect 261300 270496 261352 270502
rect 261300 270438 261352 270444
rect 261024 270360 261076 270366
rect 261024 270302 261076 270308
rect 259736 269476 259788 269482
rect 259736 269418 259788 269424
rect 260840 269476 260892 269482
rect 260840 269418 260892 269424
rect 259460 267300 259512 267306
rect 259460 267242 259512 267248
rect 259552 266552 259604 266558
rect 259552 266494 259604 266500
rect 259564 264316 259592 266494
rect 259748 266422 259776 269418
rect 259736 266416 259788 266422
rect 259736 266358 259788 266364
rect 260288 266416 260340 266422
rect 260288 266358 260340 266364
rect 260300 264316 260328 266358
rect 261036 264316 261064 270302
rect 261760 269816 261812 269822
rect 261760 269758 261812 269764
rect 261772 266422 261800 269758
rect 262600 266558 262628 277766
rect 263416 271788 263468 271794
rect 263416 271730 263468 271736
rect 262864 266892 262916 266898
rect 262864 266834 262916 266840
rect 262588 266552 262640 266558
rect 262588 266494 262640 266500
rect 261760 266416 261812 266422
rect 261760 266358 261812 266364
rect 262128 266416 262180 266422
rect 262128 266358 262180 266364
rect 262140 264330 262168 266358
rect 262876 264330 262904 266834
rect 263428 264330 263456 271730
rect 263612 269822 263640 277766
rect 264992 270366 265020 277766
rect 265900 275324 265952 275330
rect 265900 275266 265952 275272
rect 264980 270360 265032 270366
rect 264980 270302 265032 270308
rect 263600 269816 263652 269822
rect 263600 269758 263652 269764
rect 265440 269816 265492 269822
rect 265440 269758 265492 269764
rect 264704 269340 264756 269346
rect 264704 269282 264756 269288
rect 263968 267776 264020 267782
rect 263968 267718 264020 267724
rect 261786 264302 262168 264330
rect 262522 264302 262904 264330
rect 263258 264302 263456 264330
rect 263980 264316 264008 267718
rect 264716 264316 264744 269282
rect 265452 264316 265480 269758
rect 265912 269346 265940 275266
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 265900 269340 265952 269346
rect 265900 269282 265952 269288
rect 266188 264316 266216 270030
rect 266372 266422 266400 277766
rect 268028 277394 268056 277780
rect 267936 277366 268056 277394
rect 266912 269952 266964 269958
rect 266912 269894 266964 269900
rect 266360 266416 266412 266422
rect 266360 266358 266412 266364
rect 266924 264316 266952 269894
rect 267648 267164 267700 267170
rect 267648 267106 267700 267112
rect 267660 264316 267688 267106
rect 267936 266898 267964 277366
rect 269224 271794 269252 277780
rect 269592 277766 270434 277794
rect 269212 271788 269264 271794
rect 269212 271730 269264 271736
rect 268844 271448 268896 271454
rect 268844 271390 268896 271396
rect 267924 266892 267976 266898
rect 267924 266834 267976 266840
rect 268856 264330 268884 271390
rect 269120 268932 269172 268938
rect 269120 268874 269172 268880
rect 268410 264302 268884 264330
rect 269132 264316 269160 268874
rect 269592 267782 269620 277766
rect 271524 275330 271552 277780
rect 271892 277766 272734 277794
rect 273272 277766 273930 277794
rect 274652 277766 275126 277794
rect 271512 275324 271564 275330
rect 271512 275266 271564 275272
rect 271144 274712 271196 274718
rect 271144 274654 271196 274660
rect 269580 267776 269632 267782
rect 269580 267718 269632 267724
rect 271156 267170 271184 274654
rect 271696 272536 271748 272542
rect 271696 272478 271748 272484
rect 271708 267734 271736 272478
rect 271892 269822 271920 277766
rect 273076 271312 273128 271318
rect 273076 271254 273128 271260
rect 271880 269816 271932 269822
rect 271880 269758 271932 269764
rect 271880 269680 271932 269686
rect 271880 269622 271932 269628
rect 271892 267734 271920 269622
rect 271616 267706 271736 267734
rect 271800 267706 271920 267734
rect 271144 267164 271196 267170
rect 271144 267106 271196 267112
rect 269856 266552 269908 266558
rect 269856 266494 269908 266500
rect 269868 264316 269896 266494
rect 271616 266422 271644 267706
rect 270592 266416 270644 266422
rect 270592 266358 270644 266364
rect 271604 266416 271656 266422
rect 271604 266358 271656 266364
rect 270604 264316 270632 266358
rect 271800 264330 271828 267706
rect 272064 267164 272116 267170
rect 272064 267106 272116 267112
rect 271354 264302 271828 264330
rect 272076 264316 272104 267106
rect 273088 264330 273116 271254
rect 273272 270094 273300 277766
rect 274364 273964 274416 273970
rect 274364 273906 274416 273912
rect 273260 270088 273312 270094
rect 273260 270030 273312 270036
rect 273536 268660 273588 268666
rect 273536 268602 273588 268608
rect 272826 264302 273116 264330
rect 273548 264316 273576 268602
rect 274376 267734 274404 273906
rect 274652 269958 274680 277766
rect 276308 274718 276336 277780
rect 276296 274712 276348 274718
rect 276296 274654 276348 274660
rect 276664 274712 276716 274718
rect 276664 274654 276716 274660
rect 274824 270360 274876 270366
rect 274824 270302 274876 270308
rect 274640 269952 274692 269958
rect 274640 269894 274692 269900
rect 274284 267706 274404 267734
rect 274284 264316 274312 267706
rect 274836 266558 274864 270302
rect 276480 270088 276532 270094
rect 276480 270030 276532 270036
rect 275008 269952 275060 269958
rect 275008 269894 275060 269900
rect 274824 266552 274876 266558
rect 274824 266494 274876 266500
rect 275020 264316 275048 269894
rect 275744 266892 275796 266898
rect 275744 266834 275796 266840
rect 275756 264316 275784 266834
rect 276492 264316 276520 270030
rect 276676 268938 276704 274654
rect 277504 271454 277532 277780
rect 278412 275324 278464 275330
rect 278412 275266 278464 275272
rect 277492 271448 277544 271454
rect 277492 271390 277544 271396
rect 277308 271176 277360 271182
rect 277308 271118 277360 271124
rect 276664 268932 276716 268938
rect 276664 268874 276716 268880
rect 277320 267734 277348 271118
rect 277228 267706 277348 267734
rect 277228 264316 277256 267706
rect 278424 264330 278452 275266
rect 278700 274718 278728 277780
rect 278976 277766 279818 277794
rect 278688 274712 278740 274718
rect 278688 274654 278740 274660
rect 278976 270366 279004 277766
rect 280712 274712 280764 274718
rect 280712 274654 280764 274660
rect 279884 274100 279936 274106
rect 279884 274042 279936 274048
rect 278964 270360 279016 270366
rect 278964 270302 279016 270308
rect 278872 270224 278924 270230
rect 278872 270166 278924 270172
rect 278688 267028 278740 267034
rect 278688 266970 278740 266976
rect 277978 264302 278452 264330
rect 278700 264316 278728 266970
rect 278884 266898 278912 270166
rect 278872 266892 278924 266898
rect 278872 266834 278924 266840
rect 279896 264330 279924 274042
rect 280724 267170 280752 274654
rect 281000 272542 281028 277780
rect 281552 277766 282210 277794
rect 280988 272536 281040 272542
rect 280988 272478 281040 272484
rect 281552 269686 281580 277766
rect 282920 275596 282972 275602
rect 282920 275538 282972 275544
rect 282184 272536 282236 272542
rect 282184 272478 282236 272484
rect 281540 269680 281592 269686
rect 281540 269622 281592 269628
rect 281632 268388 281684 268394
rect 281632 268330 281684 268336
rect 280712 267164 280764 267170
rect 280712 267106 280764 267112
rect 280160 266552 280212 266558
rect 280160 266494 280212 266500
rect 279450 264302 279924 264330
rect 280172 264316 280200 266494
rect 280896 266416 280948 266422
rect 280896 266358 280948 266364
rect 280908 264316 280936 266358
rect 281644 264316 281672 268330
rect 282196 266422 282224 272478
rect 282932 268666 282960 275538
rect 283392 274718 283420 277780
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283932 274236 283984 274242
rect 283932 274178 283984 274184
rect 283104 269816 283156 269822
rect 283104 269758 283156 269764
rect 282920 268660 282972 268666
rect 282920 268602 282972 268608
rect 282368 268524 282420 268530
rect 282368 268466 282420 268472
rect 282184 266416 282236 266422
rect 282184 266358 282236 266364
rect 282380 264316 282408 268466
rect 283116 264316 283144 269758
rect 283944 267734 283972 274178
rect 284588 271318 284616 277780
rect 285784 275602 285812 277780
rect 285772 275596 285824 275602
rect 285772 275538 285824 275544
rect 285680 275460 285732 275466
rect 285680 275402 285732 275408
rect 285692 271538 285720 275402
rect 286888 273970 286916 277780
rect 287072 277766 288098 277794
rect 288452 277766 289294 277794
rect 289832 277766 290490 277794
rect 286876 273964 286928 273970
rect 286876 273906 286928 273912
rect 286876 272672 286928 272678
rect 286876 272614 286928 272620
rect 285508 271510 285720 271538
rect 284576 271312 284628 271318
rect 284576 271254 284628 271260
rect 285312 271312 285364 271318
rect 285312 271254 285364 271260
rect 283852 267706 283972 267734
rect 283852 264316 283880 267706
rect 284576 266416 284628 266422
rect 284576 266358 284628 266364
rect 284588 264316 284616 266358
rect 285324 264316 285352 271254
rect 285508 266422 285536 271510
rect 286324 271448 286376 271454
rect 286324 271390 286376 271396
rect 286336 266558 286364 271390
rect 286692 267572 286744 267578
rect 286692 267514 286744 267520
rect 286324 266552 286376 266558
rect 286324 266494 286376 266500
rect 285496 266416 285548 266422
rect 285496 266358 285548 266364
rect 286048 266416 286100 266422
rect 286048 266358 286100 266364
rect 286060 264316 286088 266358
rect 286704 264330 286732 267514
rect 286888 266422 286916 272614
rect 287072 269958 287100 277766
rect 288072 273964 288124 273970
rect 288072 273906 288124 273912
rect 287060 269952 287112 269958
rect 287060 269894 287112 269900
rect 287520 269952 287572 269958
rect 287520 269894 287572 269900
rect 286876 266416 286928 266422
rect 286876 266358 286928 266364
rect 286704 264302 286810 264330
rect 287532 264316 287560 269894
rect 288084 264330 288112 273906
rect 288452 270230 288480 277766
rect 289636 271584 289688 271590
rect 289636 271526 289688 271532
rect 288440 270224 288492 270230
rect 288440 270166 288492 270172
rect 288992 266892 289044 266898
rect 288992 266834 289044 266840
rect 288084 264302 288282 264330
rect 289004 264316 289032 266834
rect 289648 264330 289676 271526
rect 289832 270094 289860 277766
rect 291672 271182 291700 277780
rect 292868 275330 292896 277780
rect 292856 275324 292908 275330
rect 292856 275266 292908 275272
rect 294064 274718 294092 277780
rect 293224 274712 293276 274718
rect 293224 274654 293276 274660
rect 294052 274712 294104 274718
rect 294052 274654 294104 274660
rect 291660 271176 291712 271182
rect 291660 271118 291712 271124
rect 292396 271176 292448 271182
rect 292396 271118 292448 271124
rect 290464 270224 290516 270230
rect 290464 270166 290516 270172
rect 289820 270088 289872 270094
rect 289820 270030 289872 270036
rect 289648 264302 289754 264330
rect 290476 264316 290504 270166
rect 291200 267164 291252 267170
rect 291200 267106 291252 267112
rect 291212 264316 291240 267106
rect 292408 264330 292436 271118
rect 292672 270496 292724 270502
rect 292672 270438 292724 270444
rect 291962 264302 292436 264330
rect 292684 264316 292712 270438
rect 293236 267034 293264 274654
rect 294604 274508 294656 274514
rect 294604 274450 294656 274456
rect 294616 267578 294644 274450
rect 295168 274106 295196 277780
rect 295340 275324 295392 275330
rect 295340 275266 295392 275272
rect 295156 274100 295208 274106
rect 295156 274042 295208 274048
rect 295064 272944 295116 272950
rect 295064 272886 295116 272892
rect 294880 268660 294932 268666
rect 294880 268602 294932 268608
rect 294604 267572 294656 267578
rect 294604 267514 294656 267520
rect 293408 267436 293460 267442
rect 293408 267378 293460 267384
rect 293224 267028 293276 267034
rect 293224 266970 293276 266976
rect 293420 264316 293448 267378
rect 294144 266416 294196 266422
rect 294144 266358 294196 266364
rect 294156 264316 294184 266358
rect 294892 264316 294920 268602
rect 295076 266422 295104 272886
rect 295352 268530 295380 275266
rect 296364 271454 296392 277780
rect 297272 275732 297324 275738
rect 297272 275674 297324 275680
rect 296628 271720 296680 271726
rect 296628 271662 296680 271668
rect 296352 271448 296404 271454
rect 296352 271390 296404 271396
rect 295340 268524 295392 268530
rect 295340 268466 295392 268472
rect 295616 267572 295668 267578
rect 295616 267514 295668 267520
rect 295064 266416 295116 266422
rect 295064 266358 295116 266364
rect 295628 264316 295656 267514
rect 296640 264330 296668 271662
rect 297284 271590 297312 275674
rect 297560 272542 297588 277780
rect 298112 277766 298770 277794
rect 297548 272536 297600 272542
rect 297548 272478 297600 272484
rect 297272 271584 297324 271590
rect 297272 271526 297324 271532
rect 297824 270088 297876 270094
rect 297824 270030 297876 270036
rect 297088 268524 297140 268530
rect 297088 268466 297140 268472
rect 296378 264302 296668 264330
rect 297100 264316 297128 268466
rect 297836 264316 297864 270030
rect 298112 268394 298140 277766
rect 299952 275330 299980 277780
rect 300872 277766 301162 277794
rect 299940 275324 299992 275330
rect 299940 275266 299992 275272
rect 300124 274100 300176 274106
rect 300124 274042 300176 274048
rect 298744 272808 298796 272814
rect 298744 272750 298796 272756
rect 298100 268388 298152 268394
rect 298100 268330 298152 268336
rect 298756 266898 298784 272750
rect 299296 268932 299348 268938
rect 299296 268874 299348 268880
rect 298744 266892 298796 266898
rect 298744 266834 298796 266840
rect 298560 266416 298612 266422
rect 298560 266358 298612 266364
rect 298572 264316 298600 266358
rect 299308 264316 299336 268874
rect 300136 266422 300164 274042
rect 300676 271448 300728 271454
rect 300676 271390 300728 271396
rect 300400 267028 300452 267034
rect 300400 266970 300452 266976
rect 300124 266416 300176 266422
rect 300124 266358 300176 266364
rect 300412 264330 300440 266970
rect 300058 264302 300440 264330
rect 300688 264330 300716 271390
rect 300872 269822 300900 277766
rect 301136 275324 301188 275330
rect 301136 275266 301188 275272
rect 301148 271726 301176 275266
rect 302344 274242 302372 277780
rect 302516 275596 302568 275602
rect 302516 275538 302568 275544
rect 302332 274236 302384 274242
rect 302332 274178 302384 274184
rect 302528 272950 302556 275538
rect 303448 275466 303476 277780
rect 303436 275460 303488 275466
rect 303436 275402 303488 275408
rect 302884 274372 302936 274378
rect 302884 274314 302936 274320
rect 302516 272944 302568 272950
rect 302516 272886 302568 272892
rect 301136 271720 301188 271726
rect 301136 271662 301188 271668
rect 301504 271584 301556 271590
rect 301504 271526 301556 271532
rect 300860 269816 300912 269822
rect 300860 269758 300912 269764
rect 301516 267170 301544 271526
rect 301964 270360 302016 270366
rect 301964 270302 302016 270308
rect 301976 267578 302004 270302
rect 301964 267572 302016 267578
rect 301964 267514 302016 267520
rect 302896 267442 302924 274314
rect 303436 272536 303488 272542
rect 303436 272478 303488 272484
rect 302884 267436 302936 267442
rect 302884 267378 302936 267384
rect 301504 267164 301556 267170
rect 301504 267106 301556 267112
rect 302240 267164 302292 267170
rect 302240 267106 302292 267112
rect 301504 266552 301556 266558
rect 301504 266494 301556 266500
rect 300688 264302 300794 264330
rect 301516 264316 301544 266494
rect 302252 264316 302280 267106
rect 303448 264330 303476 272478
rect 304644 271318 304672 277780
rect 305092 275868 305144 275874
rect 305092 275810 305144 275816
rect 304908 271856 304960 271862
rect 304908 271798 304960 271804
rect 304632 271312 304684 271318
rect 304632 271254 304684 271260
rect 304172 268388 304224 268394
rect 304172 268330 304224 268336
rect 304184 266558 304212 268330
rect 304172 266552 304224 266558
rect 304172 266494 304224 266500
rect 304448 266552 304500 266558
rect 304448 266494 304500 266500
rect 303712 266416 303764 266422
rect 303712 266358 303764 266364
rect 303002 264302 303476 264330
rect 303724 264316 303752 266358
rect 304460 264316 304488 266494
rect 304920 266422 304948 271798
rect 305104 270502 305132 275810
rect 305840 272678 305868 277780
rect 307036 274514 307064 277780
rect 307772 277766 308246 277794
rect 307024 274508 307076 274514
rect 307024 274450 307076 274456
rect 307576 274236 307628 274242
rect 307576 274178 307628 274184
rect 305828 272672 305880 272678
rect 305828 272614 305880 272620
rect 306288 272672 306340 272678
rect 306288 272614 306340 272620
rect 305092 270496 305144 270502
rect 305092 270438 305144 270444
rect 306104 269816 306156 269822
rect 306104 269758 306156 269764
rect 305920 267708 305972 267714
rect 305920 267650 305972 267656
rect 304908 266416 304960 266422
rect 304908 266358 304960 266364
rect 305184 266416 305236 266422
rect 305184 266358 305236 266364
rect 305196 264316 305224 266358
rect 305932 264316 305960 267650
rect 306116 266558 306144 269758
rect 306104 266552 306156 266558
rect 306104 266494 306156 266500
rect 306300 266422 306328 272614
rect 306288 266416 306340 266422
rect 306288 266358 306340 266364
rect 306656 266416 306708 266422
rect 306656 266358 306708 266364
rect 306668 264316 306696 266358
rect 307588 264330 307616 274178
rect 307772 269958 307800 277766
rect 309428 273970 309456 277780
rect 309416 273964 309468 273970
rect 309416 273906 309468 273912
rect 310060 272944 310112 272950
rect 310060 272886 310112 272892
rect 309048 271720 309100 271726
rect 309048 271662 309100 271668
rect 307760 269952 307812 269958
rect 307760 269894 307812 269900
rect 308128 267572 308180 267578
rect 308128 267514 308180 267520
rect 307418 264302 307616 264330
rect 308140 264316 308168 267514
rect 309060 264330 309088 271662
rect 310072 264330 310100 272886
rect 310532 272814 310560 277780
rect 311728 275738 311756 277780
rect 311912 277766 312938 277794
rect 311716 275732 311768 275738
rect 311716 275674 311768 275680
rect 311072 275460 311124 275466
rect 311072 275402 311124 275408
rect 310520 272808 310572 272814
rect 310520 272750 310572 272756
rect 311084 271454 311112 275402
rect 311072 271448 311124 271454
rect 311072 271390 311124 271396
rect 311716 271448 311768 271454
rect 311716 271390 311768 271396
rect 310336 269952 310388 269958
rect 310336 269894 310388 269900
rect 308890 264302 309088 264330
rect 309626 264302 310100 264330
rect 310348 264316 310376 269894
rect 310796 269544 310848 269550
rect 310796 269486 310848 269492
rect 310808 267034 310836 269486
rect 310796 267028 310848 267034
rect 310796 266970 310848 266976
rect 311072 266892 311124 266898
rect 311072 266834 311124 266840
rect 311084 264316 311112 266834
rect 311728 264330 311756 271390
rect 311912 270230 311940 277766
rect 314120 271590 314148 277780
rect 314476 273964 314528 273970
rect 314476 273906 314528 273912
rect 314108 271584 314160 271590
rect 314108 271526 314160 271532
rect 311900 270224 311952 270230
rect 311900 270166 311952 270172
rect 312820 270224 312872 270230
rect 312820 270166 312872 270172
rect 312832 267170 312860 270166
rect 313924 269680 313976 269686
rect 313924 269622 313976 269628
rect 313280 267436 313332 267442
rect 313280 267378 313332 267384
rect 312820 267164 312872 267170
rect 312820 267106 312872 267112
rect 313004 267164 313056 267170
rect 313004 267106 313056 267112
rect 313016 264330 313044 267106
rect 311728 264302 311834 264330
rect 312570 264302 313044 264330
rect 313292 264316 313320 267378
rect 313936 266422 313964 269622
rect 313924 266416 313976 266422
rect 313924 266358 313976 266364
rect 314488 264330 314516 273906
rect 315316 271182 315344 277780
rect 316512 275874 316540 277780
rect 317144 276004 317196 276010
rect 317144 275946 317196 275952
rect 316500 275868 316552 275874
rect 316500 275810 316552 275816
rect 315948 271584 316000 271590
rect 315948 271526 316000 271532
rect 315304 271176 315356 271182
rect 315304 271118 315356 271124
rect 314752 267028 314804 267034
rect 314752 266970 314804 266976
rect 314042 264302 314516 264330
rect 314764 264316 314792 266970
rect 315960 264330 315988 271526
rect 316960 268796 317012 268802
rect 316960 268738 317012 268744
rect 316224 266416 316276 266422
rect 316224 266358 316276 266364
rect 315514 264302 315988 264330
rect 316236 264316 316264 266358
rect 316972 264316 317000 268738
rect 317156 268666 317184 275946
rect 317328 275868 317380 275874
rect 317328 275810 317380 275816
rect 317340 272678 317368 275810
rect 317708 274378 317736 277780
rect 318812 275602 318840 277780
rect 320008 276010 320036 277780
rect 320192 277766 321218 277794
rect 319996 276004 320048 276010
rect 319996 275946 320048 275952
rect 319996 275732 320048 275738
rect 319996 275674 320048 275680
rect 318800 275596 318852 275602
rect 318800 275538 318852 275544
rect 319628 274712 319680 274718
rect 319628 274654 319680 274660
rect 318708 274508 318760 274514
rect 318708 274450 318760 274456
rect 317696 274372 317748 274378
rect 317696 274314 317748 274320
rect 317512 273080 317564 273086
rect 317512 273022 317564 273028
rect 317328 272672 317380 272678
rect 317328 272614 317380 272620
rect 317524 272490 317552 273022
rect 317340 272462 317552 272490
rect 317144 268660 317196 268666
rect 317144 268602 317196 268608
rect 317340 266422 317368 272462
rect 317696 268252 317748 268258
rect 317696 268194 317748 268200
rect 317328 266416 317380 266422
rect 317328 266358 317380 266364
rect 317708 264316 317736 268194
rect 318720 264330 318748 274450
rect 319640 268938 319668 274654
rect 320008 272950 320036 275674
rect 319996 272944 320048 272950
rect 319996 272886 320048 272892
rect 319996 271312 320048 271318
rect 319996 271254 320048 271260
rect 319628 268932 319680 268938
rect 319628 268874 319680 268880
rect 319812 268932 319864 268938
rect 319812 268874 319864 268880
rect 319824 266898 319852 268874
rect 319812 266892 319864 266898
rect 319812 266834 319864 266840
rect 319168 266756 319220 266762
rect 319168 266698 319220 266704
rect 318458 264302 318748 264330
rect 319180 264316 319208 266698
rect 320008 265962 320036 271254
rect 320192 270366 320220 277766
rect 322400 275330 322428 277780
rect 322952 277766 323610 277794
rect 324332 277766 324806 277794
rect 322388 275324 322440 275330
rect 322388 275266 322440 275272
rect 322572 275324 322624 275330
rect 322572 275266 322624 275272
rect 321468 272944 321520 272950
rect 321468 272886 321520 272892
rect 321284 271176 321336 271182
rect 321284 271118 321336 271124
rect 320180 270360 320232 270366
rect 320180 270302 320232 270308
rect 320640 266416 320692 266422
rect 320640 266358 320692 266364
rect 319916 265934 320036 265962
rect 319916 264316 319944 265934
rect 320652 264316 320680 266358
rect 321296 264330 321324 271118
rect 321480 266422 321508 272886
rect 322584 272542 322612 275266
rect 322756 273828 322808 273834
rect 322756 273770 322808 273776
rect 322572 272536 322624 272542
rect 322572 272478 322624 272484
rect 322112 267300 322164 267306
rect 322112 267242 322164 267248
rect 321468 266416 321520 266422
rect 321468 266358 321520 266364
rect 321296 264302 321402 264330
rect 322124 264316 322152 267242
rect 322768 264330 322796 273770
rect 322952 268530 322980 277766
rect 324044 272808 324096 272814
rect 324044 272750 324096 272756
rect 322940 268524 322992 268530
rect 322940 268466 322992 268472
rect 324056 264330 324084 272750
rect 324332 270094 324360 277766
rect 325988 274106 326016 277780
rect 327092 274718 327120 277780
rect 327552 277766 328302 277794
rect 327080 274712 327132 274718
rect 327080 274654 327132 274660
rect 325976 274100 326028 274106
rect 325976 274042 326028 274048
rect 326988 273216 327040 273222
rect 326988 273158 327040 273164
rect 325516 272672 325568 272678
rect 325516 272614 325568 272620
rect 324320 270088 324372 270094
rect 324320 270030 324372 270036
rect 324320 269068 324372 269074
rect 324320 269010 324372 269016
rect 324332 267714 324360 269010
rect 324688 268524 324740 268530
rect 324688 268466 324740 268472
rect 324320 267708 324372 267714
rect 324320 267650 324372 267656
rect 324700 264330 324728 268466
rect 325528 264330 325556 272614
rect 325792 270496 325844 270502
rect 325792 270438 325844 270444
rect 322768 264302 322874 264330
rect 323610 264302 324084 264330
rect 324346 264302 324728 264330
rect 325082 264302 325556 264330
rect 325804 264316 325832 270438
rect 327000 264330 327028 273158
rect 327552 269550 327580 277766
rect 329196 275596 329248 275602
rect 329196 275538 329248 275544
rect 327540 269544 327592 269550
rect 327540 269486 327592 269492
rect 328000 269272 328052 269278
rect 328000 269214 328052 269220
rect 327264 266892 327316 266898
rect 327264 266834 327316 266840
rect 326554 264302 327028 264330
rect 327276 264316 327304 266834
rect 328012 264316 328040 269214
rect 329208 264330 329236 275538
rect 329484 275466 329512 277780
rect 329852 277766 330694 277794
rect 331416 277766 331890 277794
rect 329472 275460 329524 275466
rect 329472 275402 329524 275408
rect 329656 274644 329708 274650
rect 329656 274586 329708 274592
rect 329472 268660 329524 268666
rect 329472 268602 329524 268608
rect 329484 267578 329512 268602
rect 329472 267572 329524 267578
rect 329472 267514 329524 267520
rect 329668 264330 329696 274586
rect 329852 268394 329880 277766
rect 331220 276004 331272 276010
rect 331220 275946 331272 275952
rect 331232 274242 331260 275946
rect 331220 274236 331272 274242
rect 331220 274178 331272 274184
rect 331416 270230 331444 277766
rect 333072 275330 333100 277780
rect 333612 275460 333664 275466
rect 333612 275402 333664 275408
rect 333060 275324 333112 275330
rect 333060 275266 333112 275272
rect 332508 273420 332560 273426
rect 332508 273362 332560 273368
rect 332324 270360 332376 270366
rect 332324 270302 332376 270308
rect 331404 270224 331456 270230
rect 331404 270166 331456 270172
rect 330208 269544 330260 269550
rect 330208 269486 330260 269492
rect 329840 268388 329892 268394
rect 329840 268330 329892 268336
rect 328762 264302 329236 264330
rect 329498 264302 329696 264330
rect 330220 264316 330248 269486
rect 330944 266552 330996 266558
rect 330944 266494 330996 266500
rect 330956 264316 330984 266494
rect 331680 266416 331732 266422
rect 331680 266358 331732 266364
rect 331692 264316 331720 266358
rect 332336 264330 332364 270302
rect 332520 266422 332548 273362
rect 333244 272536 333296 272542
rect 333244 272478 333296 272484
rect 333256 266558 333284 272478
rect 333428 266892 333480 266898
rect 333428 266834 333480 266840
rect 333440 266626 333468 266834
rect 333428 266620 333480 266626
rect 333428 266562 333480 266568
rect 333244 266552 333296 266558
rect 333244 266494 333296 266500
rect 332508 266416 332560 266422
rect 332508 266358 332560 266364
rect 333624 264330 333652 275402
rect 334176 271862 334204 277780
rect 334164 271856 334216 271862
rect 334164 271798 334216 271804
rect 334624 271856 334676 271862
rect 334624 271798 334676 271804
rect 333888 267708 333940 267714
rect 333888 267650 333940 267656
rect 332336 264302 332442 264330
rect 333178 264302 333652 264330
rect 333900 264316 333928 267650
rect 334636 267442 334664 271798
rect 334992 270088 335044 270094
rect 334992 270030 335044 270036
rect 334624 267436 334676 267442
rect 334624 267378 334676 267384
rect 335004 264330 335032 270030
rect 335372 269822 335400 277780
rect 336568 275874 336596 277780
rect 336752 277766 337778 277794
rect 338132 277766 338974 277794
rect 336556 275868 336608 275874
rect 336556 275810 336608 275816
rect 336556 274372 336608 274378
rect 336556 274314 336608 274320
rect 335360 269816 335412 269822
rect 335360 269758 335412 269764
rect 335360 267436 335412 267442
rect 335360 267378 335412 267384
rect 334650 264302 335032 264330
rect 335372 264316 335400 267378
rect 336568 264330 336596 274314
rect 336752 269074 336780 277766
rect 337752 271040 337804 271046
rect 337752 270982 337804 270988
rect 337200 269816 337252 269822
rect 337200 269758 337252 269764
rect 336740 269068 336792 269074
rect 336740 269010 336792 269016
rect 337212 264330 337240 269758
rect 337764 264330 337792 270982
rect 338132 269686 338160 277766
rect 340156 276010 340184 277780
rect 340892 277766 341366 277794
rect 340144 276004 340196 276010
rect 340144 275946 340196 275952
rect 340236 275324 340288 275330
rect 340236 275266 340288 275272
rect 338856 274780 338908 274786
rect 338856 274722 338908 274728
rect 338868 269958 338896 274722
rect 338856 269952 338908 269958
rect 338856 269894 338908 269900
rect 339040 269952 339092 269958
rect 339040 269894 339092 269900
rect 338120 269680 338172 269686
rect 338120 269622 338172 269628
rect 338304 266892 338356 266898
rect 338304 266834 338356 266840
rect 336122 264302 336596 264330
rect 336858 264302 337240 264330
rect 337594 264302 337792 264330
rect 338316 264316 338344 266834
rect 339052 264316 339080 269894
rect 339408 269068 339460 269074
rect 339408 269010 339460 269016
rect 339420 266762 339448 269010
rect 340052 267028 340104 267034
rect 340052 266970 340104 266976
rect 340064 266762 340092 266970
rect 339408 266756 339460 266762
rect 339408 266698 339460 266704
rect 340052 266756 340104 266762
rect 340052 266698 340104 266704
rect 340248 264330 340276 275266
rect 340696 272128 340748 272134
rect 340696 272070 340748 272076
rect 340708 264330 340736 272070
rect 340892 268666 340920 277766
rect 342260 276004 342312 276010
rect 342260 275946 342312 275952
rect 342272 273970 342300 275946
rect 342260 273964 342312 273970
rect 342260 273906 342312 273912
rect 342456 271726 342484 277780
rect 343652 275738 343680 277780
rect 343824 275868 343876 275874
rect 343824 275810 343876 275816
rect 343640 275732 343692 275738
rect 343640 275674 343692 275680
rect 343548 274236 343600 274242
rect 343548 274178 343600 274184
rect 342444 271720 342496 271726
rect 342444 271662 342496 271668
rect 343364 270632 343416 270638
rect 343364 270574 343416 270580
rect 341248 269680 341300 269686
rect 341248 269622 341300 269628
rect 340880 268660 340932 268666
rect 340880 268602 340932 268608
rect 339802 264302 340276 264330
rect 340538 264302 340736 264330
rect 341260 264316 341288 269622
rect 342168 268388 342220 268394
rect 342168 268330 342220 268336
rect 342180 267442 342208 268330
rect 342720 267572 342772 267578
rect 342720 267514 342772 267520
rect 342168 267436 342220 267442
rect 342168 267378 342220 267384
rect 341800 267300 341852 267306
rect 341800 267242 341852 267248
rect 341984 267300 342036 267306
rect 341984 267242 342036 267248
rect 341812 267034 341840 267242
rect 341800 267028 341852 267034
rect 341800 266970 341852 266976
rect 341996 264316 342024 267242
rect 342732 264316 342760 267514
rect 343376 267170 343404 270574
rect 343560 267578 343588 274178
rect 343836 273086 343864 275810
rect 344848 274786 344876 277780
rect 345216 277766 346058 277794
rect 346780 277766 347254 277794
rect 348160 277766 348450 277794
rect 344836 274780 344888 274786
rect 344836 274722 344888 274728
rect 344652 273964 344704 273970
rect 344652 273906 344704 273912
rect 343824 273080 343876 273086
rect 343824 273022 343876 273028
rect 344192 270904 344244 270910
rect 344192 270846 344244 270852
rect 343548 267572 343600 267578
rect 343548 267514 343600 267520
rect 343364 267164 343416 267170
rect 343364 267106 343416 267112
rect 343456 266756 343508 266762
rect 343456 266698 343508 266704
rect 343468 264316 343496 266698
rect 344204 264316 344232 270846
rect 344664 264330 344692 273906
rect 345216 268938 345244 277766
rect 345388 275732 345440 275738
rect 345388 275674 345440 275680
rect 345400 273222 345428 275674
rect 345388 273216 345440 273222
rect 345388 273158 345440 273164
rect 345480 273080 345532 273086
rect 345480 273022 345532 273028
rect 345204 268932 345256 268938
rect 345204 268874 345256 268880
rect 345492 266490 345520 273022
rect 345664 271584 345716 271590
rect 345664 271526 345716 271532
rect 346584 271584 346636 271590
rect 346584 271526 346636 271532
rect 345676 270774 345704 271526
rect 345664 270768 345716 270774
rect 345664 270710 345716 270716
rect 346400 267572 346452 267578
rect 346400 267514 346452 267520
rect 345480 266484 345532 266490
rect 345480 266426 345532 266432
rect 345664 266416 345716 266422
rect 345664 266358 345716 266364
rect 344664 264302 344954 264330
rect 345676 264316 345704 266358
rect 346412 264316 346440 267514
rect 346596 266626 346624 271526
rect 346780 271454 346808 277766
rect 347780 271720 347832 271726
rect 347780 271662 347832 271668
rect 346768 271448 346820 271454
rect 346768 271390 346820 271396
rect 347136 267844 347188 267850
rect 347136 267786 347188 267792
rect 346584 266620 346636 266626
rect 346584 266562 346636 266568
rect 347148 264316 347176 267786
rect 347792 267034 347820 271662
rect 348160 270638 348188 277766
rect 349632 271862 349660 277780
rect 350736 276010 350764 277780
rect 351946 277766 352236 277794
rect 350724 276004 350776 276010
rect 350724 275946 350776 275952
rect 350540 275188 350592 275194
rect 350540 275130 350592 275136
rect 350552 274514 350580 275130
rect 350540 274508 350592 274514
rect 350540 274450 350592 274456
rect 351828 274508 351880 274514
rect 351828 274450 351880 274456
rect 349620 271856 349672 271862
rect 349620 271798 349672 271804
rect 350080 271448 350132 271454
rect 350080 271390 350132 271396
rect 348148 270632 348200 270638
rect 348148 270574 348200 270580
rect 349344 268932 349396 268938
rect 349344 268874 349396 268880
rect 347780 267028 347832 267034
rect 347780 266970 347832 266976
rect 348608 267028 348660 267034
rect 348608 266970 348660 266976
rect 347872 266620 347924 266626
rect 347872 266562 347924 266568
rect 347884 264316 347912 266562
rect 348620 264316 348648 266970
rect 349356 264316 349384 268874
rect 350092 264316 350120 271390
rect 351644 270224 351696 270230
rect 351644 270166 351696 270172
rect 350816 267164 350868 267170
rect 350816 267106 350868 267112
rect 350828 264316 350856 267106
rect 351656 266762 351684 270166
rect 351644 266756 351696 266762
rect 351644 266698 351696 266704
rect 351840 264330 351868 274450
rect 352208 271658 352236 277766
rect 352196 271652 352248 271658
rect 352196 271594 352248 271600
rect 353128 270774 353156 277780
rect 354324 275874 354352 277780
rect 355324 276004 355376 276010
rect 355324 275946 355376 275952
rect 354312 275868 354364 275874
rect 354312 275810 354364 275816
rect 353392 274780 353444 274786
rect 353392 274722 353444 274728
rect 353116 270768 353168 270774
rect 353116 270710 353168 270716
rect 353208 270632 353260 270638
rect 353208 270574 353260 270580
rect 353024 266756 353076 266762
rect 353024 266698 353076 266704
rect 352288 266416 352340 266422
rect 352288 266358 352340 266364
rect 351578 264302 351868 264330
rect 352300 264316 352328 266358
rect 353036 264316 353064 266698
rect 353220 266422 353248 270574
rect 353404 268802 353432 274722
rect 353944 273284 353996 273290
rect 353944 273226 353996 273232
rect 353392 268796 353444 268802
rect 353392 268738 353444 268744
rect 353760 268660 353812 268666
rect 353760 268602 353812 268608
rect 353208 266416 353260 266422
rect 353208 266358 353260 266364
rect 353772 264316 353800 268602
rect 353956 267714 353984 273226
rect 354588 270768 354640 270774
rect 354588 270710 354640 270716
rect 354600 267734 354628 270710
rect 355336 270502 355364 275946
rect 355520 274786 355548 277780
rect 356072 277766 356730 277794
rect 355508 274780 355560 274786
rect 355508 274722 355560 274728
rect 355876 271992 355928 271998
rect 355876 271934 355928 271940
rect 355324 270496 355376 270502
rect 355324 270438 355376 270444
rect 354772 269408 354824 269414
rect 354772 269350 354824 269356
rect 353944 267708 353996 267714
rect 353944 267650 353996 267656
rect 354508 267706 354628 267734
rect 354508 264316 354536 267706
rect 354784 266422 354812 269350
rect 355232 267300 355284 267306
rect 355232 267242 355284 267248
rect 354772 266416 354824 266422
rect 354772 266358 354824 266364
rect 355244 264316 355272 267242
rect 355888 264330 355916 271934
rect 356072 268258 356100 277766
rect 356888 275868 356940 275874
rect 356888 275810 356940 275816
rect 356900 270910 356928 275810
rect 357912 275194 357940 277780
rect 359016 277394 359044 277780
rect 358924 277366 359044 277394
rect 357900 275188 357952 275194
rect 357900 275130 357952 275136
rect 358728 274780 358780 274786
rect 358728 274722 358780 274728
rect 358740 273834 358768 274722
rect 358728 273828 358780 273834
rect 358728 273770 358780 273776
rect 358084 273556 358136 273562
rect 358084 273498 358136 273504
rect 356888 270904 356940 270910
rect 356888 270846 356940 270852
rect 357164 270904 357216 270910
rect 357164 270846 357216 270852
rect 356060 268252 356112 268258
rect 356060 268194 356112 268200
rect 357176 264330 357204 270846
rect 357440 267708 357492 267714
rect 357440 267650 357492 267656
rect 355888 264302 355994 264330
rect 356730 264302 357204 264330
rect 357452 264316 357480 267650
rect 358096 266898 358124 273498
rect 358924 269074 358952 277366
rect 359464 271584 359516 271590
rect 359464 271526 359516 271532
rect 359476 271046 359504 271526
rect 360212 271318 360240 277780
rect 361408 272950 361436 277780
rect 361396 272944 361448 272950
rect 361396 272886 361448 272892
rect 361304 271856 361356 271862
rect 361304 271798 361356 271804
rect 360200 271312 360252 271318
rect 360200 271254 360252 271260
rect 359464 271040 359516 271046
rect 359464 270982 359516 270988
rect 360108 271040 360160 271046
rect 360108 270982 360160 270988
rect 359292 270286 359872 270314
rect 359292 269686 359320 270286
rect 359844 270230 359872 270286
rect 359648 270224 359700 270230
rect 359648 270166 359700 270172
rect 359832 270224 359884 270230
rect 359832 270166 359884 270172
rect 359660 269958 359688 270166
rect 359464 269952 359516 269958
rect 359464 269894 359516 269900
rect 359648 269952 359700 269958
rect 359648 269894 359700 269900
rect 359476 269686 359504 269894
rect 359280 269680 359332 269686
rect 359280 269622 359332 269628
rect 359464 269680 359516 269686
rect 359464 269622 359516 269628
rect 358912 269068 358964 269074
rect 358912 269010 358964 269016
rect 358544 268932 358596 268938
rect 358544 268874 358596 268880
rect 358084 266892 358136 266898
rect 358084 266834 358136 266840
rect 358556 264330 358584 268874
rect 359280 268524 359332 268530
rect 359280 268466 359332 268472
rect 359292 268258 359320 268466
rect 359280 268252 359332 268258
rect 359280 268194 359332 268200
rect 359648 266892 359700 266898
rect 359648 266834 359700 266840
rect 358912 266416 358964 266422
rect 358912 266358 358964 266364
rect 358202 264302 358584 264330
rect 358924 264316 358952 266358
rect 359660 264316 359688 266834
rect 360120 266422 360148 270982
rect 360384 268116 360436 268122
rect 360384 268058 360436 268064
rect 360108 266416 360160 266422
rect 360108 266358 360160 266364
rect 360396 264316 360424 268058
rect 361316 264330 361344 271798
rect 362604 271182 362632 277780
rect 363616 277766 363814 277794
rect 362776 272264 362828 272270
rect 362776 272206 362828 272212
rect 362592 271176 362644 271182
rect 362592 271118 362644 271124
rect 362788 266422 362816 272206
rect 363616 271726 363644 277766
rect 364996 274786 365024 277780
rect 365628 275188 365680 275194
rect 365628 275130 365680 275136
rect 364984 274780 365036 274786
rect 364984 274722 365036 274728
rect 365444 274780 365496 274786
rect 365444 274722 365496 274728
rect 364248 272400 364300 272406
rect 364248 272342 364300 272348
rect 363604 271720 363656 271726
rect 363604 271662 363656 271668
rect 363788 271720 363840 271726
rect 363788 271662 363840 271668
rect 362960 266892 363012 266898
rect 362960 266834 363012 266840
rect 362972 266490 363000 266834
rect 362960 266484 363012 266490
rect 362960 266426 363012 266432
rect 361856 266416 361908 266422
rect 361856 266358 361908 266364
rect 362776 266416 362828 266422
rect 362776 266358 362828 266364
rect 361146 264302 361344 264330
rect 361868 264316 361896 266358
rect 362592 266076 362644 266082
rect 362592 266018 362644 266024
rect 362604 264316 362632 266018
rect 363800 264330 363828 271662
rect 364260 264330 364288 272342
rect 365456 271590 365484 274722
rect 365640 274650 365668 275130
rect 365628 274644 365680 274650
rect 365628 274586 365680 274592
rect 366100 272814 366128 277780
rect 367296 277394 367324 277780
rect 367204 277366 367324 277394
rect 367008 273828 367060 273834
rect 367008 273770 367060 273776
rect 366088 272808 366140 272814
rect 366088 272750 366140 272756
rect 365444 271584 365496 271590
rect 365444 271526 365496 271532
rect 365628 271176 365680 271182
rect 365628 271118 365680 271124
rect 364800 268796 364852 268802
rect 364800 268738 364852 268744
rect 363354 264302 363828 264330
rect 364090 264302 364288 264330
rect 364812 264316 364840 268738
rect 365640 267734 365668 271118
rect 365812 267980 365864 267986
rect 365812 267922 365864 267928
rect 365548 267706 365668 267734
rect 365548 264316 365576 267706
rect 365824 266626 365852 267922
rect 365996 267708 366048 267714
rect 365996 267650 366048 267656
rect 366008 267034 366036 267650
rect 366638 267336 366694 267345
rect 366638 267271 366694 267280
rect 365996 267028 366048 267034
rect 365996 266970 366048 266976
rect 365812 266620 365864 266626
rect 365812 266562 365864 266568
rect 366652 264330 366680 267271
rect 366298 264302 366680 264330
rect 367020 264316 367048 273770
rect 367204 268258 367232 277366
rect 368492 272678 368520 277780
rect 369688 276010 369716 277780
rect 369676 276004 369728 276010
rect 369676 275946 369728 275952
rect 369952 276004 370004 276010
rect 369952 275946 370004 275952
rect 368480 272672 368532 272678
rect 368480 272614 368532 272620
rect 369768 272672 369820 272678
rect 369768 272614 369820 272620
rect 367744 270496 367796 270502
rect 367744 270438 367796 270444
rect 367192 268252 367244 268258
rect 367192 268194 367244 268200
rect 367756 264316 367784 270438
rect 369122 270192 369178 270201
rect 369122 270127 369178 270136
rect 369136 266898 369164 270127
rect 369308 268932 369360 268938
rect 369308 268874 369360 268880
rect 369492 268932 369544 268938
rect 369492 268874 369544 268880
rect 369320 268122 369348 268874
rect 369308 268116 369360 268122
rect 369308 268058 369360 268064
rect 369124 266892 369176 266898
rect 369124 266834 369176 266840
rect 369306 266792 369362 266801
rect 369306 266727 369308 266736
rect 369360 266727 369362 266736
rect 369308 266698 369360 266704
rect 368480 265804 368532 265810
rect 368480 265746 368532 265752
rect 368492 264316 368520 265746
rect 369504 264330 369532 268874
rect 369780 265810 369808 272614
rect 369964 268666 369992 275946
rect 370884 275738 370912 277780
rect 370872 275732 370924 275738
rect 370872 275674 370924 275680
rect 371884 274100 371936 274106
rect 371884 274042 371936 274048
rect 371896 273254 371924 274042
rect 371620 273226 371924 273254
rect 370320 271312 370372 271318
rect 370320 271254 370372 271260
rect 369952 268660 370004 268666
rect 369952 268602 370004 268608
rect 369768 265804 369820 265810
rect 369768 265746 369820 265752
rect 370332 264330 370360 271254
rect 371620 267578 371648 273226
rect 372080 273086 372108 277780
rect 372632 277766 373290 277794
rect 372068 273080 372120 273086
rect 372068 273022 372120 273028
rect 372436 273080 372488 273086
rect 372436 273022 372488 273028
rect 371792 272808 371844 272814
rect 371792 272750 371844 272756
rect 371804 272542 371832 272750
rect 371792 272536 371844 272542
rect 371792 272478 371844 272484
rect 371976 272536 372028 272542
rect 371976 272478 372028 272484
rect 371988 272134 372016 272478
rect 371976 272128 372028 272134
rect 371976 272070 372028 272076
rect 371608 267572 371660 267578
rect 371608 267514 371660 267520
rect 371792 267572 371844 267578
rect 371792 267514 371844 267520
rect 370502 267336 370558 267345
rect 370502 267271 370504 267280
rect 370556 267271 370558 267280
rect 370504 267242 370556 267248
rect 371424 267164 371476 267170
rect 371424 267106 371476 267112
rect 370688 266892 370740 266898
rect 370688 266834 370740 266840
rect 369242 264302 369532 264330
rect 369978 264302 370360 264330
rect 370700 264316 370728 266834
rect 371436 264316 371464 267106
rect 371804 266801 371832 267514
rect 371790 266792 371846 266801
rect 371790 266727 371846 266736
rect 372448 264330 372476 273022
rect 372632 269278 372660 277766
rect 374184 275732 374236 275738
rect 374184 275674 374236 275680
rect 374196 272542 374224 275674
rect 374380 275602 374408 277780
rect 374368 275596 374420 275602
rect 374368 275538 374420 275544
rect 374644 275596 374696 275602
rect 374644 275538 374696 275544
rect 374368 273692 374420 273698
rect 374368 273634 374420 273640
rect 374184 272536 374236 272542
rect 374184 272478 374236 272484
rect 374380 270314 374408 273634
rect 374656 273426 374684 275538
rect 375576 275194 375604 277780
rect 375564 275188 375616 275194
rect 375564 275130 375616 275136
rect 376116 274916 376168 274922
rect 376116 274858 376168 274864
rect 374644 273420 374696 273426
rect 374644 273362 374696 273368
rect 375012 272536 375064 272542
rect 375012 272478 375064 272484
rect 374104 270286 374408 270314
rect 373724 269680 373776 269686
rect 373724 269622 373776 269628
rect 372988 269544 373040 269550
rect 372988 269486 373040 269492
rect 373448 269544 373500 269550
rect 373736 269521 373764 269622
rect 373448 269486 373500 269492
rect 373722 269512 373778 269521
rect 373000 269278 373028 269486
rect 372620 269272 372672 269278
rect 372620 269214 372672 269220
rect 372988 269272 373040 269278
rect 372988 269214 373040 269220
rect 373460 267714 373488 269486
rect 373722 269447 373778 269456
rect 373448 267708 373500 267714
rect 373448 267650 373500 267656
rect 373632 267708 373684 267714
rect 373632 267650 373684 267656
rect 372896 266620 372948 266626
rect 372896 266562 372948 266568
rect 372186 264302 372476 264330
rect 372908 264316 372936 266562
rect 373644 264316 373672 267650
rect 374104 266762 374132 270286
rect 374828 270224 374880 270230
rect 374288 270172 374828 270178
rect 374288 270166 374880 270172
rect 374288 270150 374868 270166
rect 374288 269278 374316 270150
rect 374460 270088 374512 270094
rect 374460 270030 374512 270036
rect 374276 269272 374328 269278
rect 374276 269214 374328 269220
rect 374472 269210 374500 270030
rect 374460 269204 374512 269210
rect 374460 269146 374512 269152
rect 374644 268660 374696 268666
rect 374644 268602 374696 268608
rect 374656 268394 374684 268602
rect 374644 268388 374696 268394
rect 374644 268330 374696 268336
rect 375024 266914 375052 272478
rect 375196 269544 375248 269550
rect 375194 269512 375196 269521
rect 375248 269512 375250 269521
rect 375194 269447 375250 269456
rect 375840 269068 375892 269074
rect 375840 269010 375892 269016
rect 374840 266886 375052 266914
rect 374092 266756 374144 266762
rect 374092 266698 374144 266704
rect 374840 264330 374868 266886
rect 375104 266756 375156 266762
rect 375104 266698 375156 266704
rect 374394 264302 374868 264330
rect 375116 264316 375144 266698
rect 375852 264316 375880 269010
rect 376128 267850 376156 274858
rect 376576 272944 376628 272950
rect 376576 272886 376628 272892
rect 376116 267844 376168 267850
rect 376116 267786 376168 267792
rect 376588 264316 376616 272886
rect 376772 270230 376800 277780
rect 377968 272814 377996 277780
rect 379164 275602 379192 277780
rect 379532 277766 380374 277794
rect 379152 275596 379204 275602
rect 379152 275538 379204 275544
rect 378784 275120 378836 275126
rect 378784 275062 378836 275068
rect 378796 274378 378824 275062
rect 378784 274372 378836 274378
rect 378784 274314 378836 274320
rect 378968 273420 379020 273426
rect 378968 273362 379020 273368
rect 377956 272808 378008 272814
rect 377956 272750 378008 272756
rect 378140 272808 378192 272814
rect 378140 272750 378192 272756
rect 378152 272542 378180 272750
rect 378140 272536 378192 272542
rect 378140 272478 378192 272484
rect 378784 271992 378836 271998
rect 378784 271934 378836 271940
rect 376760 270224 376812 270230
rect 376944 270224 376996 270230
rect 376760 270166 376812 270172
rect 376942 270192 376944 270201
rect 376996 270192 376998 270201
rect 376942 270127 376998 270136
rect 377126 270056 377182 270065
rect 377126 269991 377182 270000
rect 377140 267578 377168 269991
rect 378048 267844 378100 267850
rect 378048 267786 378100 267792
rect 377128 267572 377180 267578
rect 377128 267514 377180 267520
rect 377312 267572 377364 267578
rect 377312 267514 377364 267520
rect 377324 264316 377352 267514
rect 378060 264316 378088 267786
rect 378796 264316 378824 271934
rect 378980 267034 379008 273362
rect 379152 270360 379204 270366
rect 379150 270328 379152 270337
rect 379336 270360 379388 270366
rect 379204 270328 379206 270337
rect 379532 270337 379560 277766
rect 380716 276956 380768 276962
rect 380716 276898 380768 276904
rect 379336 270302 379388 270308
rect 379518 270328 379574 270337
rect 379150 270263 379206 270272
rect 379348 270065 379376 270302
rect 379518 270263 379574 270272
rect 380530 270328 380586 270337
rect 380530 270263 380586 270272
rect 379334 270056 379390 270065
rect 379334 269991 379390 270000
rect 379334 267608 379390 267617
rect 379334 267543 379336 267552
rect 379388 267543 379390 267552
rect 379520 267572 379572 267578
rect 379336 267514 379388 267520
rect 379520 267514 379572 267520
rect 378968 267028 379020 267034
rect 378968 266970 379020 266976
rect 379532 264316 379560 267514
rect 380544 267442 380572 270263
rect 380532 267436 380584 267442
rect 380532 267378 380584 267384
rect 379704 267028 379756 267034
rect 379704 266970 379756 266976
rect 379716 266762 379744 266970
rect 379704 266756 379756 266762
rect 379704 266698 379756 266704
rect 380728 264330 380756 276898
rect 380900 275596 380952 275602
rect 380900 275538 380952 275544
rect 380912 272134 380940 275538
rect 381556 275466 381584 277780
rect 382384 277766 382674 277794
rect 381544 275460 381596 275466
rect 381544 275402 381596 275408
rect 382384 273290 382412 277766
rect 382648 275460 382700 275466
rect 382648 275402 382700 275408
rect 382660 274786 382688 275402
rect 382648 274780 382700 274786
rect 382648 274722 382700 274728
rect 382832 274780 382884 274786
rect 382832 274722 382884 274728
rect 382372 273284 382424 273290
rect 382372 273226 382424 273232
rect 380900 272128 380952 272134
rect 380900 272070 380952 272076
rect 382188 272128 382240 272134
rect 382188 272070 382240 272076
rect 381358 267608 381414 267617
rect 381358 267543 381360 267552
rect 381412 267543 381414 267552
rect 381360 267514 381412 267520
rect 382200 266762 382228 272070
rect 382464 268524 382516 268530
rect 382464 268466 382516 268472
rect 380992 266756 381044 266762
rect 380992 266698 381044 266704
rect 382188 266756 382240 266762
rect 382188 266698 382240 266704
rect 380282 264302 380756 264330
rect 381004 264316 381032 266698
rect 382096 266212 382148 266218
rect 382096 266154 382148 266160
rect 382108 264330 382136 266154
rect 381754 264302 382136 264330
rect 382476 264316 382504 268466
rect 382844 268394 382872 274722
rect 383856 273254 383884 277780
rect 383856 273226 383976 273254
rect 383200 271584 383252 271590
rect 383200 271526 383252 271532
rect 382832 268388 382884 268394
rect 382832 268330 382884 268336
rect 383212 264316 383240 271526
rect 383384 270360 383436 270366
rect 383568 270360 383620 270366
rect 383384 270302 383436 270308
rect 383566 270328 383568 270337
rect 383620 270328 383622 270337
rect 383396 269657 383424 270302
rect 383566 270263 383622 270272
rect 383658 270056 383714 270065
rect 383658 269991 383714 270000
rect 383672 269906 383700 269991
rect 383580 269878 383700 269906
rect 383580 269822 383608 269878
rect 383568 269816 383620 269822
rect 383568 269758 383620 269764
rect 383752 269816 383804 269822
rect 383752 269758 383804 269764
rect 383764 269657 383792 269758
rect 383382 269648 383438 269657
rect 383382 269583 383438 269592
rect 383750 269648 383806 269657
rect 383750 269583 383806 269592
rect 383948 269278 383976 273226
rect 384304 272536 384356 272542
rect 384304 272478 384356 272484
rect 384120 269544 384172 269550
rect 384118 269512 384120 269521
rect 384172 269512 384174 269521
rect 384118 269447 384174 269456
rect 383936 269272 383988 269278
rect 383936 269214 383988 269220
rect 384120 269204 384172 269210
rect 384120 269146 384172 269152
rect 384132 266218 384160 269146
rect 384316 267578 384344 272478
rect 384488 269544 384540 269550
rect 384488 269486 384540 269492
rect 384500 269210 384528 269486
rect 384488 269204 384540 269210
rect 384488 269146 384540 269152
rect 385052 268666 385080 277780
rect 386248 275126 386276 277780
rect 386984 277766 387458 277794
rect 386420 275596 386472 275602
rect 386420 275538 386472 275544
rect 386432 275194 386460 275538
rect 386420 275188 386472 275194
rect 386420 275130 386472 275136
rect 386236 275120 386288 275126
rect 386236 275062 386288 275068
rect 386420 275052 386472 275058
rect 386420 274994 386472 275000
rect 386432 274786 386460 274994
rect 386420 274780 386472 274786
rect 386420 274722 386472 274728
rect 385960 273284 386012 273290
rect 385960 273226 386012 273232
rect 385040 268660 385092 268666
rect 385040 268602 385092 268608
rect 384304 267572 384356 267578
rect 384304 267514 384356 267520
rect 384488 267572 384540 267578
rect 384488 267514 384540 267520
rect 384120 266212 384172 266218
rect 384120 266154 384172 266160
rect 384500 264330 384528 267514
rect 385408 266756 385460 266762
rect 385408 266698 385460 266704
rect 384672 265940 384724 265946
rect 384672 265882 384724 265888
rect 383962 264302 384528 264330
rect 384684 264316 384712 265882
rect 385420 264316 385448 266698
rect 385972 264330 386000 273226
rect 386984 270065 387012 277766
rect 387340 276820 387392 276826
rect 387340 276762 387392 276768
rect 386970 270056 387026 270065
rect 386970 269991 387026 270000
rect 387352 264330 387380 276762
rect 388640 275466 388668 277780
rect 388628 275460 388680 275466
rect 388628 275402 388680 275408
rect 388076 274780 388128 274786
rect 388076 274722 388128 274728
rect 388088 271454 388116 274722
rect 389744 273562 389772 277780
rect 390572 277766 390954 277794
rect 390284 274644 390336 274650
rect 390284 274586 390336 274592
rect 389732 273556 389784 273562
rect 389732 273498 389784 273504
rect 388272 272598 388668 272626
rect 388272 272542 388300 272598
rect 388260 272536 388312 272542
rect 388260 272478 388312 272484
rect 388444 272536 388496 272542
rect 388444 272478 388496 272484
rect 388456 271998 388484 272478
rect 388640 271998 388668 272598
rect 388444 271992 388496 271998
rect 388444 271934 388496 271940
rect 388628 271992 388680 271998
rect 388628 271934 388680 271940
rect 388628 271584 388680 271590
rect 388628 271526 388680 271532
rect 388812 271584 388864 271590
rect 388812 271526 388864 271532
rect 388076 271448 388128 271454
rect 388076 271390 388128 271396
rect 388640 271318 388668 271526
rect 388628 271312 388680 271318
rect 388628 271254 388680 271260
rect 388444 270360 388496 270366
rect 388444 270302 388496 270308
rect 388628 270360 388680 270366
rect 388628 270302 388680 270308
rect 388456 269278 388484 270302
rect 388640 269550 388668 270302
rect 388628 269544 388680 269550
rect 388628 269486 388680 269492
rect 388444 269272 388496 269278
rect 388444 269214 388496 269220
rect 388352 268660 388404 268666
rect 388352 268602 388404 268608
rect 387616 268388 387668 268394
rect 387616 268330 387668 268336
rect 385972 264302 386170 264330
rect 386906 264302 387380 264330
rect 387628 264316 387656 268330
rect 388364 267850 388392 268602
rect 388352 267844 388404 267850
rect 388352 267786 388404 267792
rect 388168 267572 388220 267578
rect 388168 267514 388220 267520
rect 388352 267572 388404 267578
rect 388352 267514 388404 267520
rect 388180 267345 388208 267514
rect 388166 267336 388222 267345
rect 388166 267271 388222 267280
rect 388364 264316 388392 267514
rect 388824 266762 388852 271526
rect 388996 269544 389048 269550
rect 388994 269512 388996 269521
rect 389048 269512 389050 269521
rect 388994 269447 389050 269456
rect 390100 267844 390152 267850
rect 390100 267786 390152 267792
rect 390112 267306 390140 267786
rect 390100 267300 390152 267306
rect 390100 267242 390152 267248
rect 388812 266756 388864 266762
rect 388812 266698 388864 266704
rect 389088 265804 389140 265810
rect 389088 265746 389140 265752
rect 389100 264316 389128 265746
rect 390296 264330 390324 274586
rect 390572 269550 390600 277766
rect 391572 275596 391624 275602
rect 391572 275538 391624 275544
rect 390560 269544 390612 269550
rect 390560 269486 390612 269492
rect 391296 269544 391348 269550
rect 391296 269486 391348 269492
rect 390466 267336 390522 267345
rect 390466 267271 390468 267280
rect 390520 267271 390522 267280
rect 390468 267242 390520 267248
rect 390560 266756 390612 266762
rect 390560 266698 390612 266704
rect 389850 264302 390324 264330
rect 390572 264316 390600 266698
rect 391308 264316 391336 269486
rect 391584 266762 391612 275538
rect 392136 275466 392164 277780
rect 393332 275738 393360 277780
rect 393700 277766 394542 277794
rect 393320 275732 393372 275738
rect 393320 275674 393372 275680
rect 392124 275460 392176 275466
rect 392124 275402 392176 275408
rect 391940 275324 391992 275330
rect 391940 275266 391992 275272
rect 391952 274242 391980 275266
rect 393228 274372 393280 274378
rect 393228 274314 393280 274320
rect 391940 274236 391992 274242
rect 391940 274178 391992 274184
rect 391756 271584 391808 271590
rect 391754 271552 391756 271561
rect 391940 271584 391992 271590
rect 391808 271552 391810 271561
rect 391940 271526 391992 271532
rect 391754 271487 391810 271496
rect 391952 267850 391980 271526
rect 391940 267844 391992 267850
rect 391940 267786 391992 267792
rect 392582 267608 392638 267617
rect 392582 267543 392584 267552
rect 392636 267543 392638 267552
rect 392768 267572 392820 267578
rect 392584 267514 392636 267520
rect 392768 267514 392820 267520
rect 391756 267436 391808 267442
rect 391756 267378 391808 267384
rect 392032 267436 392084 267442
rect 392032 267378 392084 267384
rect 391768 266762 391796 267378
rect 391572 266756 391624 266762
rect 391572 266698 391624 266704
rect 391756 266756 391808 266762
rect 391756 266698 391808 266704
rect 392044 264316 392072 267378
rect 392780 264316 392808 267514
rect 393240 267442 393268 274314
rect 393700 270094 393728 277766
rect 395436 275732 395488 275738
rect 395436 275674 395488 275680
rect 394332 274236 394384 274242
rect 394332 274178 394384 274184
rect 393688 270088 393740 270094
rect 393688 270030 393740 270036
rect 393688 269408 393740 269414
rect 393686 269376 393688 269385
rect 393872 269408 393924 269414
rect 393740 269376 393742 269385
rect 393872 269350 393924 269356
rect 393686 269311 393742 269320
rect 393410 267608 393466 267617
rect 393410 267543 393466 267552
rect 393424 267442 393452 267543
rect 393228 267436 393280 267442
rect 393228 267378 393280 267384
rect 393412 267436 393464 267442
rect 393412 267378 393464 267384
rect 393884 264330 393912 269350
rect 394344 267734 394372 274178
rect 394792 273556 394844 273562
rect 394792 273498 394844 273504
rect 394804 273290 394832 273498
rect 394792 273284 394844 273290
rect 394792 273226 394844 273232
rect 394976 273216 395028 273222
rect 394976 273158 395028 273164
rect 394988 271998 395016 273158
rect 394976 271992 395028 271998
rect 394976 271934 395028 271940
rect 393530 264302 393912 264330
rect 394252 267706 394372 267734
rect 394252 264316 394280 267706
rect 395448 264330 395476 275674
rect 395724 274106 395752 277780
rect 396724 275460 396776 275466
rect 396724 275402 396776 275408
rect 395712 274100 395764 274106
rect 395712 274042 395764 274048
rect 396736 273970 396764 275402
rect 396920 275330 396948 277780
rect 397656 277766 398038 277794
rect 396908 275324 396960 275330
rect 396908 275266 396960 275272
rect 397460 275324 397512 275330
rect 397460 275266 397512 275272
rect 397276 274100 397328 274106
rect 397276 274042 397328 274048
rect 396724 273964 396776 273970
rect 396724 273906 396776 273912
rect 395896 269952 395948 269958
rect 395896 269894 395948 269900
rect 395908 264330 395936 269894
rect 396172 267980 396224 267986
rect 396172 267922 396224 267928
rect 396184 267170 396212 267922
rect 396172 267164 396224 267170
rect 396172 267106 396224 267112
rect 396262 266520 396318 266529
rect 396262 266455 396264 266464
rect 396316 266455 396318 266464
rect 396264 266426 396316 266432
rect 397288 266422 397316 274042
rect 397472 273562 397500 275266
rect 397460 273556 397512 273562
rect 397460 273498 397512 273504
rect 397656 270094 397684 277766
rect 399220 275874 399248 277780
rect 399208 275868 399260 275874
rect 399208 275810 399260 275816
rect 400220 275868 400272 275874
rect 400220 275810 400272 275816
rect 399666 275768 399722 275777
rect 399666 275703 399668 275712
rect 399720 275703 399722 275712
rect 399852 275732 399904 275738
rect 399668 275674 399720 275680
rect 399852 275674 399904 275680
rect 398748 273964 398800 273970
rect 398748 273906 398800 273912
rect 397644 270088 397696 270094
rect 397644 270030 397696 270036
rect 398288 270088 398340 270094
rect 398288 270030 398340 270036
rect 397920 269680 397972 269686
rect 397918 269648 397920 269657
rect 397972 269648 397974 269657
rect 397918 269583 397974 269592
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 395002 264302 395476 264330
rect 395738 264302 395936 264330
rect 396460 264316 396488 266358
rect 397184 266280 397236 266286
rect 397184 266222 397236 266228
rect 397196 264316 397224 266222
rect 398300 264330 398328 270030
rect 398472 269816 398524 269822
rect 398472 269758 398524 269764
rect 398484 269414 398512 269758
rect 398472 269408 398524 269414
rect 398472 269350 398524 269356
rect 398760 267734 398788 273906
rect 398930 269648 398986 269657
rect 398930 269583 398986 269592
rect 398944 269414 398972 269583
rect 398932 269408 398984 269414
rect 398932 269350 398984 269356
rect 398668 267706 398788 267734
rect 398472 267300 398524 267306
rect 398472 267242 398524 267248
rect 398484 266529 398512 267242
rect 398470 266520 398526 266529
rect 398470 266455 398526 266464
rect 397946 264302 398328 264330
rect 398668 264316 398696 267706
rect 399864 264330 399892 275674
rect 400232 274514 400260 275810
rect 400416 275466 400444 277780
rect 400770 275768 400826 275777
rect 400588 275732 400640 275738
rect 400770 275703 400772 275712
rect 400588 275674 400640 275680
rect 400824 275703 400826 275712
rect 400772 275674 400824 275680
rect 400600 275466 400628 275674
rect 400404 275460 400456 275466
rect 400404 275402 400456 275408
rect 400588 275460 400640 275466
rect 400588 275402 400640 275408
rect 400220 274508 400272 274514
rect 400220 274450 400272 274456
rect 401324 274508 401376 274514
rect 401324 274450 401376 274456
rect 400126 269784 400182 269793
rect 400126 269719 400182 269728
rect 399418 264302 399892 264330
rect 400140 264316 400168 269719
rect 401336 264330 401364 274450
rect 401612 269385 401640 277780
rect 402072 277766 402822 277794
rect 402072 269498 402100 277766
rect 402428 276548 402480 276554
rect 402428 276490 402480 276496
rect 401796 269470 402100 269498
rect 401796 269414 401824 269470
rect 401784 269408 401836 269414
rect 401598 269376 401654 269385
rect 401784 269350 401836 269356
rect 401968 269408 402020 269414
rect 401968 269350 402020 269356
rect 401598 269311 401654 269320
rect 401980 267306 402008 269350
rect 402440 267734 402468 276490
rect 404004 274922 404032 277780
rect 404372 277766 405214 277794
rect 405752 277766 406318 277794
rect 403992 274916 404044 274922
rect 403992 274858 404044 274864
rect 404176 274916 404228 274922
rect 404176 274858 404228 274864
rect 402610 271552 402666 271561
rect 402610 271487 402666 271496
rect 402624 270450 402652 271487
rect 402978 271008 403034 271017
rect 402978 270943 403034 270952
rect 402992 270858 403020 270943
rect 404188 270858 404216 274858
rect 402900 270830 403020 270858
rect 404004 270830 404216 270858
rect 402900 270774 402928 270830
rect 404004 270774 404032 270830
rect 402888 270768 402940 270774
rect 402888 270710 402940 270716
rect 403072 270768 403124 270774
rect 403072 270710 403124 270716
rect 403992 270768 404044 270774
rect 403992 270710 404044 270716
rect 402796 270632 402848 270638
rect 402794 270600 402796 270609
rect 402934 270632 402986 270638
rect 402848 270600 402850 270609
rect 403084 270609 403112 270710
rect 402934 270574 402986 270580
rect 403070 270600 403126 270609
rect 402794 270535 402850 270544
rect 402946 270450 402974 270574
rect 403070 270535 403126 270544
rect 404174 270600 404230 270609
rect 404174 270535 404230 270544
rect 402624 270422 402974 270450
rect 402348 267706 402468 267734
rect 401968 267300 402020 267306
rect 401968 267242 402020 267248
rect 401600 266416 401652 266422
rect 401600 266358 401652 266364
rect 400890 264302 401364 264330
rect 401612 264316 401640 266358
rect 402348 264316 402376 267706
rect 402980 267300 403032 267306
rect 402980 267242 403032 267248
rect 402992 266506 403020 267242
rect 402900 266478 403020 266506
rect 402900 266422 402928 266478
rect 404188 266422 404216 270535
rect 404372 267850 404400 277766
rect 405188 273556 405240 273562
rect 405188 273498 405240 273504
rect 404360 267844 404412 267850
rect 404360 267786 404412 267792
rect 402888 266416 402940 266422
rect 402888 266358 402940 266364
rect 403072 266416 403124 266422
rect 403072 266358 403124 266364
rect 404176 266416 404228 266422
rect 404176 266358 404228 266364
rect 403084 264316 403112 266358
rect 404544 265668 404596 265674
rect 404544 265610 404596 265616
rect 403808 265532 403860 265538
rect 403808 265474 403860 265480
rect 403820 264316 403848 265474
rect 404556 264316 404584 265610
rect 405200 264330 405228 273498
rect 405372 272264 405424 272270
rect 405372 272206 405424 272212
rect 405384 271998 405412 272206
rect 405372 271992 405424 271998
rect 405372 271934 405424 271940
rect 405752 270230 405780 277766
rect 405924 270632 405976 270638
rect 405922 270600 405924 270609
rect 405976 270600 405978 270609
rect 405922 270535 405978 270544
rect 405740 270224 405792 270230
rect 405740 270166 405792 270172
rect 405924 270224 405976 270230
rect 406752 270224 406804 270230
rect 405924 270166 405976 270172
rect 406750 270192 406752 270201
rect 406804 270192 406806 270201
rect 405936 266626 405964 270166
rect 406750 270127 406806 270136
rect 405924 266620 405976 266626
rect 405924 266562 405976 266568
rect 406384 266552 406436 266558
rect 406384 266494 406436 266500
rect 406396 264330 406424 266494
rect 406948 264330 406976 278666
rect 546696 278594 547078 278610
rect 437204 278588 437256 278594
rect 437204 278530 437256 278536
rect 546684 278588 547078 278594
rect 546736 278582 547078 278588
rect 546684 278530 546736 278536
rect 424692 277840 424744 277846
rect 407500 276010 407528 277780
rect 407488 276004 407540 276010
rect 407488 275946 407540 275952
rect 408224 276004 408276 276010
rect 408224 275946 408276 275952
rect 407396 270224 407448 270230
rect 408040 270224 408092 270230
rect 407396 270166 407448 270172
rect 407776 270184 408040 270212
rect 407408 269686 407436 270166
rect 407580 269952 407632 269958
rect 407580 269894 407632 269900
rect 407592 269686 407620 269894
rect 407396 269680 407448 269686
rect 407396 269622 407448 269628
rect 407580 269680 407632 269686
rect 407580 269622 407632 269628
rect 407776 269226 407804 270184
rect 408040 270166 408092 270172
rect 407500 269198 407804 269226
rect 407304 268116 407356 268122
rect 407304 268058 407356 268064
rect 407316 267850 407344 268058
rect 407304 267844 407356 267850
rect 407304 267786 407356 267792
rect 405200 264302 405306 264330
rect 406042 264302 406424 264330
rect 406778 264302 406976 264330
rect 407500 264316 407528 269198
rect 407764 269068 407816 269074
rect 407764 269010 407816 269016
rect 407948 269068 408000 269074
rect 407948 269010 408000 269016
rect 407776 268122 407804 269010
rect 407764 268116 407816 268122
rect 407764 268058 407816 268064
rect 407960 267986 407988 269010
rect 407948 267980 408000 267986
rect 407948 267922 408000 267928
rect 408236 264316 408264 275946
rect 408696 274786 408724 277780
rect 409420 277092 409472 277098
rect 409420 277034 409472 277040
rect 408684 274780 408736 274786
rect 408684 274722 408736 274728
rect 408512 270286 409000 270314
rect 408512 270230 408540 270286
rect 408500 270224 408552 270230
rect 408776 270224 408828 270230
rect 408500 270166 408552 270172
rect 408774 270192 408776 270201
rect 408828 270192 408830 270201
rect 408774 270127 408830 270136
rect 408972 270094 409000 270286
rect 408592 270088 408644 270094
rect 408960 270088 409012 270094
rect 408644 270036 408724 270042
rect 408592 270030 408724 270036
rect 408960 270030 409012 270036
rect 408604 270014 408724 270030
rect 408696 269278 408724 270014
rect 408454 269272 408506 269278
rect 408684 269272 408736 269278
rect 408506 269220 408540 269226
rect 408454 269214 408540 269220
rect 408684 269214 408736 269220
rect 408466 269198 408540 269214
rect 408512 269113 408540 269198
rect 408498 269104 408554 269113
rect 408498 269039 408554 269048
rect 409432 264330 409460 277034
rect 409892 273426 409920 277780
rect 410892 276140 410944 276146
rect 410892 276082 410944 276088
rect 409880 273420 409932 273426
rect 409880 273362 409932 273368
rect 409694 271688 409750 271697
rect 409694 271623 409750 271632
rect 408986 264302 409460 264330
rect 409708 264316 409736 271623
rect 410904 267850 410932 276082
rect 411088 275874 411116 277780
rect 411076 275868 411128 275874
rect 411076 275810 411128 275816
rect 412284 274922 412312 277780
rect 412652 277766 413402 277794
rect 412272 274916 412324 274922
rect 412272 274858 412324 274864
rect 411260 274780 411312 274786
rect 411260 274722 411312 274728
rect 411272 271017 411300 274722
rect 411904 272128 411956 272134
rect 411904 272070 411956 272076
rect 411258 271008 411314 271017
rect 411258 270943 411314 270952
rect 411168 267980 411220 267986
rect 411168 267922 411220 267928
rect 410892 267844 410944 267850
rect 410892 267786 410944 267792
rect 410798 266384 410854 266393
rect 410798 266319 410854 266328
rect 410812 264330 410840 266319
rect 410458 264302 410840 264330
rect 411180 264316 411208 267922
rect 411916 264316 411944 272070
rect 412652 269278 412680 277766
rect 413744 277704 413796 277710
rect 413744 277646 413796 277652
rect 413468 271448 413520 271454
rect 413468 271390 413520 271396
rect 412914 271144 412970 271153
rect 412914 271079 412970 271088
rect 412928 270774 412956 271079
rect 413480 271046 413508 271390
rect 413284 271040 413336 271046
rect 413284 270982 413336 270988
rect 413468 271040 413520 271046
rect 413468 270982 413520 270988
rect 413296 270774 413324 270982
rect 412916 270768 412968 270774
rect 412916 270710 412968 270716
rect 413284 270768 413336 270774
rect 413284 270710 413336 270716
rect 413468 269680 413520 269686
rect 413468 269622 413520 269628
rect 413480 269414 413508 269622
rect 413468 269408 413520 269414
rect 413468 269350 413520 269356
rect 412640 269272 412692 269278
rect 412640 269214 412692 269220
rect 413100 268252 413152 268258
rect 413100 268194 413152 268200
rect 413112 267986 413140 268194
rect 413468 268116 413520 268122
rect 413468 268058 413520 268064
rect 412916 267980 412968 267986
rect 412916 267922 412968 267928
rect 413100 267980 413152 267986
rect 413100 267922 413152 267928
rect 412928 267866 412956 267922
rect 413480 267866 413508 268058
rect 412640 267844 412692 267850
rect 412928 267838 413508 267866
rect 412640 267786 412692 267792
rect 412652 264316 412680 267786
rect 413468 267232 413520 267238
rect 413468 267174 413520 267180
rect 413480 267050 413508 267174
rect 413020 267034 413508 267050
rect 413008 267028 413508 267034
rect 413060 267022 413508 267028
rect 413008 266970 413060 266976
rect 412822 266928 412878 266937
rect 412822 266863 412824 266872
rect 412876 266863 412878 266872
rect 412824 266834 412876 266840
rect 413756 264330 413784 277646
rect 414388 275188 414440 275194
rect 414388 275130 414440 275136
rect 414400 274922 414428 275130
rect 414584 275058 414612 277780
rect 415216 275324 415268 275330
rect 415216 275266 415268 275272
rect 414572 275052 414624 275058
rect 414572 274994 414624 275000
rect 414388 274916 414440 274922
rect 414388 274858 414440 274864
rect 414664 273352 414716 273358
rect 414664 273294 414716 273300
rect 413928 271448 413980 271454
rect 413928 271390 413980 271396
rect 413940 271153 413968 271390
rect 413926 271144 413982 271153
rect 413926 271079 413982 271088
rect 414112 269680 414164 269686
rect 414112 269622 414164 269628
rect 413402 264302 413784 264330
rect 414124 264316 414152 269622
rect 414676 266937 414704 273294
rect 415228 271998 415256 275266
rect 415492 275052 415544 275058
rect 415492 274994 415544 275000
rect 415216 271992 415268 271998
rect 415216 271934 415268 271940
rect 415504 267850 415532 274994
rect 415780 274786 415808 277780
rect 416792 277766 416990 277794
rect 415768 274780 415820 274786
rect 415768 274722 415820 274728
rect 416412 273420 416464 273426
rect 416412 273362 416464 273368
rect 416424 273254 416452 273362
rect 416332 273226 416452 273254
rect 415676 273216 415728 273222
rect 415676 273158 415728 273164
rect 415688 271998 415716 273158
rect 415676 271992 415728 271998
rect 415676 271934 415728 271940
rect 415858 269512 415914 269521
rect 415858 269447 415914 269456
rect 415492 267844 415544 267850
rect 415492 267786 415544 267792
rect 415676 267844 415728 267850
rect 415676 267786 415728 267792
rect 414662 266928 414718 266937
rect 414662 266863 414718 266872
rect 414848 266416 414900 266422
rect 414848 266358 414900 266364
rect 414860 264316 414888 266358
rect 415688 266286 415716 267786
rect 415676 266280 415728 266286
rect 415676 266222 415728 266228
rect 415872 264330 415900 269447
rect 415610 264302 415900 264330
rect 416332 264316 416360 273226
rect 416792 269113 416820 277766
rect 418172 274922 418200 277780
rect 419000 277766 419382 277794
rect 418344 275324 418396 275330
rect 418344 275266 418396 275272
rect 418528 275324 418580 275330
rect 418528 275266 418580 275272
rect 418356 274922 418384 275266
rect 418160 274916 418212 274922
rect 418160 274858 418212 274864
rect 418344 274916 418396 274922
rect 418344 274858 418396 274864
rect 417976 274780 418028 274786
rect 417976 274722 418028 274728
rect 417988 273254 418016 274722
rect 417896 273226 418016 273254
rect 417700 270904 417752 270910
rect 417698 270872 417700 270881
rect 417752 270872 417754 270881
rect 417698 270807 417754 270816
rect 416778 269104 416834 269113
rect 416778 269039 416834 269048
rect 416686 268152 416742 268161
rect 416686 268087 416688 268096
rect 416740 268087 416742 268096
rect 416872 268116 416924 268122
rect 416688 268058 416740 268064
rect 416872 268058 416924 268064
rect 416884 267238 416912 268058
rect 417698 267880 417754 267889
rect 417698 267815 417754 267824
rect 417712 267714 417740 267815
rect 417700 267708 417752 267714
rect 417700 267650 417752 267656
rect 417896 267306 417924 273226
rect 418160 270904 418212 270910
rect 418158 270872 418160 270881
rect 418212 270872 418214 270881
rect 418158 270807 418214 270816
rect 418066 268152 418122 268161
rect 418066 268087 418122 268096
rect 418080 267850 418108 268087
rect 418540 267986 418568 275266
rect 419000 270910 419028 277766
rect 420368 276412 420420 276418
rect 420368 276354 420420 276360
rect 418988 270904 419040 270910
rect 418988 270846 419040 270852
rect 419448 270904 419500 270910
rect 419448 270846 419500 270852
rect 418528 267980 418580 267986
rect 418528 267922 418580 267928
rect 418068 267844 418120 267850
rect 418068 267786 418120 267792
rect 417056 267300 417108 267306
rect 417056 267242 417108 267248
rect 417884 267300 417936 267306
rect 417884 267242 417936 267248
rect 418068 267300 418120 267306
rect 418068 267242 418120 267248
rect 416872 267232 416924 267238
rect 416872 267174 416924 267180
rect 417068 264316 417096 267242
rect 418080 267186 418108 267242
rect 417620 267158 418108 267186
rect 417240 267028 417292 267034
rect 417240 266970 417292 266976
rect 417252 266422 417280 266970
rect 417620 266558 417648 267158
rect 417608 266552 417660 266558
rect 417608 266494 417660 266500
rect 419460 266422 419488 270846
rect 417240 266416 417292 266422
rect 417424 266416 417476 266422
rect 417240 266358 417292 266364
rect 417422 266384 417424 266393
rect 418528 266416 418580 266422
rect 417476 266384 417478 266393
rect 418528 266358 418580 266364
rect 419448 266416 419500 266422
rect 419448 266358 419500 266364
rect 417422 266319 417478 266328
rect 417792 265260 417844 265266
rect 417792 265202 417844 265208
rect 417804 264316 417832 265202
rect 418540 264316 418568 266358
rect 419448 266280 419500 266286
rect 419448 266222 419500 266228
rect 419460 264330 419488 266222
rect 420380 264330 420408 276354
rect 420564 273698 420592 277780
rect 421668 276010 421696 277780
rect 422496 277766 422878 277794
rect 423692 277766 424074 277794
rect 424692 277782 424744 277788
rect 422208 277568 422260 277574
rect 422208 277510 422260 277516
rect 421656 276004 421708 276010
rect 421656 275946 421708 275952
rect 421840 276004 421892 276010
rect 421840 275946 421892 275952
rect 421852 275330 421880 275946
rect 421840 275324 421892 275330
rect 421840 275266 421892 275272
rect 422024 275324 422076 275330
rect 422024 275266 422076 275272
rect 422036 274938 422064 275266
rect 422220 275074 422248 277510
rect 421944 274922 422064 274938
rect 421932 274916 422064 274922
rect 421984 274910 422064 274916
rect 422128 275046 422248 275074
rect 421932 274858 421984 274864
rect 420552 273692 420604 273698
rect 420552 273634 420604 273640
rect 422128 273254 422156 275046
rect 422300 274916 422352 274922
rect 422300 274858 422352 274864
rect 422312 274802 422340 274858
rect 422036 273226 422156 273254
rect 422220 274774 422340 274802
rect 422036 267734 422064 273226
rect 422036 267706 422156 267734
rect 421748 267028 421800 267034
rect 421748 266970 421800 266976
rect 420734 266656 420790 266665
rect 420734 266591 420790 266600
rect 419290 264302 419488 264330
rect 420026 264302 420408 264330
rect 420748 264316 420776 266591
rect 421760 266506 421788 266970
rect 421760 266490 421972 266506
rect 421760 266484 421984 266490
rect 421760 266478 421932 266484
rect 421932 266426 421984 266432
rect 422128 266336 422156 267706
rect 422036 266308 422156 266336
rect 421840 266212 421892 266218
rect 421840 266154 421892 266160
rect 421852 264330 421880 266154
rect 421498 264302 421880 264330
rect 422036 264330 422064 266308
rect 422220 266218 422248 274774
rect 422496 270774 422524 277766
rect 422944 275324 422996 275330
rect 422944 275266 422996 275272
rect 422956 275210 422984 275266
rect 422956 275194 423352 275210
rect 422956 275188 423364 275194
rect 422956 275182 423312 275188
rect 423312 275130 423364 275136
rect 423220 274916 423272 274922
rect 423220 274858 423272 274864
rect 423232 274802 423260 274858
rect 422680 274786 423260 274802
rect 422668 274780 423260 274786
rect 422720 274774 423260 274780
rect 422668 274722 422720 274728
rect 422668 273692 422720 273698
rect 422668 273634 422720 273640
rect 422484 270768 422536 270774
rect 422484 270710 422536 270716
rect 422680 267889 422708 273634
rect 423692 269278 423720 277766
rect 424508 272400 424560 272406
rect 424506 272368 424508 272377
rect 424560 272368 424562 272377
rect 424506 272303 424562 272312
rect 424508 271176 424560 271182
rect 424508 271118 424560 271124
rect 424520 270774 424548 271118
rect 424508 270768 424560 270774
rect 424508 270710 424560 270716
rect 423680 269272 423732 269278
rect 423680 269214 423732 269220
rect 423864 269272 423916 269278
rect 423864 269214 423916 269220
rect 422944 267980 422996 267986
rect 422944 267922 422996 267928
rect 422666 267880 422722 267889
rect 422666 267815 422722 267824
rect 422392 266892 422444 266898
rect 422392 266834 422444 266840
rect 422404 266354 422432 266834
rect 422392 266348 422444 266354
rect 422392 266290 422444 266296
rect 422208 266212 422260 266218
rect 422208 266154 422260 266160
rect 422036 264302 422234 264330
rect 422956 264316 422984 267922
rect 423876 266665 423904 269214
rect 423862 266656 423918 266665
rect 423862 266591 423918 266600
rect 424048 266348 424100 266354
rect 424048 266290 424100 266296
rect 424060 264330 424088 266290
rect 424704 264330 424732 277782
rect 425256 276010 425284 277780
rect 425244 276004 425296 276010
rect 425244 275946 425296 275952
rect 426072 276004 426124 276010
rect 426072 275946 426124 275952
rect 425242 268288 425298 268297
rect 425242 268223 425298 268232
rect 424874 268016 424930 268025
rect 424874 267951 424876 267960
rect 424928 267951 424930 267960
rect 424876 267922 424928 267928
rect 425256 266914 425284 268223
rect 424980 266886 425284 266914
rect 424980 266762 425008 266886
rect 424968 266756 425020 266762
rect 424968 266698 425020 266704
rect 425152 266756 425204 266762
rect 425152 266698 425204 266704
rect 423706 264302 424088 264330
rect 424442 264302 424732 264330
rect 425164 264316 425192 266698
rect 426084 264330 426112 275946
rect 426254 273592 426310 273601
rect 426254 273527 426310 273536
rect 426268 266762 426296 273527
rect 426452 271862 426480 277780
rect 427096 277766 427662 277794
rect 428292 277766 428858 277794
rect 429764 277766 429962 277794
rect 427096 275194 427124 277766
rect 427084 275188 427136 275194
rect 427084 275130 427136 275136
rect 427268 275188 427320 275194
rect 427268 275130 427320 275136
rect 427280 272377 427308 275130
rect 427266 272368 427322 272377
rect 427266 272303 427322 272312
rect 427084 272264 427136 272270
rect 427084 272206 427136 272212
rect 427096 271998 427124 272206
rect 427084 271992 427136 271998
rect 427084 271934 427136 271940
rect 427728 271992 427780 271998
rect 427728 271934 427780 271940
rect 426440 271856 426492 271862
rect 426440 271798 426492 271804
rect 427544 271856 427596 271862
rect 427544 271798 427596 271804
rect 427084 271448 427136 271454
rect 427084 271390 427136 271396
rect 427096 271046 427124 271390
rect 427084 271040 427136 271046
rect 427084 270982 427136 270988
rect 427084 267708 427136 267714
rect 427084 267650 427136 267656
rect 426898 267064 426954 267073
rect 427096 267034 427124 267650
rect 427358 267608 427414 267617
rect 427358 267543 427360 267552
rect 427412 267543 427414 267552
rect 427360 267514 427412 267520
rect 426898 266999 426900 267008
rect 426952 266999 426954 267008
rect 427084 267028 427136 267034
rect 426900 266970 426952 266976
rect 427084 266970 427136 266976
rect 427556 266762 427584 271798
rect 427740 270494 427768 271934
rect 427648 270466 427768 270494
rect 427648 266914 427676 270466
rect 428002 267608 428058 267617
rect 428002 267543 428004 267552
rect 428056 267543 428058 267552
rect 428004 267514 428056 267520
rect 428094 267336 428150 267345
rect 428094 267271 428150 267280
rect 427648 266886 427768 266914
rect 426256 266756 426308 266762
rect 426256 266698 426308 266704
rect 426624 266756 426676 266762
rect 426624 266698 426676 266704
rect 427544 266756 427596 266762
rect 427544 266698 427596 266704
rect 425914 264302 426112 264330
rect 426636 264316 426664 266698
rect 427740 264330 427768 266886
rect 427912 266756 427964 266762
rect 427912 266698 427964 266704
rect 427924 266354 427952 266698
rect 427912 266348 427964 266354
rect 427912 266290 427964 266296
rect 427386 264302 427768 264330
rect 428108 264316 428136 267271
rect 428292 266082 428320 277766
rect 429290 272232 429346 272241
rect 429290 272167 429346 272176
rect 429106 270736 429162 270745
rect 429106 270671 429162 270680
rect 428462 268016 428518 268025
rect 428462 267951 428464 267960
rect 428516 267951 428518 267960
rect 428464 267922 428516 267928
rect 428280 266076 428332 266082
rect 428280 266018 428332 266024
rect 429120 264330 429148 270671
rect 429304 268297 429332 272167
rect 429764 271726 429792 277766
rect 431144 275194 431172 277780
rect 432340 277394 432368 277780
rect 433536 277394 433564 277780
rect 434746 277766 435220 277794
rect 432340 277366 432460 277394
rect 431132 275188 431184 275194
rect 431132 275130 431184 275136
rect 431316 275188 431368 275194
rect 431316 275130 431368 275136
rect 429752 271720 429804 271726
rect 429752 271662 429804 271668
rect 430212 271584 430264 271590
rect 430212 271526 430264 271532
rect 430028 271448 430080 271454
rect 430028 271390 430080 271396
rect 430040 270774 430068 271390
rect 430224 271182 430252 271526
rect 430212 271176 430264 271182
rect 430212 271118 430264 271124
rect 431328 270774 431356 275130
rect 432050 273592 432106 273601
rect 432050 273527 432106 273536
rect 432064 273290 432092 273527
rect 432052 273284 432104 273290
rect 432432 273254 432460 277366
rect 432052 273226 432104 273232
rect 432248 273226 432460 273254
rect 433444 277366 433564 277394
rect 431868 273216 431920 273222
rect 431868 273158 431920 273164
rect 431880 272513 431908 273158
rect 431866 272504 431922 272513
rect 431866 272439 431922 272448
rect 431498 271144 431554 271153
rect 431498 271079 431554 271088
rect 430028 270768 430080 270774
rect 430028 270710 430080 270716
rect 430304 270768 430356 270774
rect 430304 270710 430356 270716
rect 431316 270768 431368 270774
rect 431316 270710 431368 270716
rect 429934 269240 429990 269249
rect 429934 269175 429990 269184
rect 429290 268288 429346 268297
rect 429290 268223 429346 268232
rect 429948 264330 429976 269175
rect 428858 264302 429148 264330
rect 429594 264302 429976 264330
rect 430316 264316 430344 270710
rect 431512 264330 431540 271079
rect 431776 271040 431828 271046
rect 431776 270982 431828 270988
rect 431066 264302 431540 264330
rect 431788 264316 431816 270982
rect 432248 268802 432276 273226
rect 433444 271454 433472 277366
rect 434350 274136 434406 274145
rect 434350 274071 434406 274080
rect 433432 271448 433484 271454
rect 432970 271416 433026 271425
rect 433432 271390 433484 271396
rect 433616 271448 433668 271454
rect 433616 271390 433668 271396
rect 432970 271351 433026 271360
rect 432420 270768 432472 270774
rect 432420 270710 432472 270716
rect 432432 270502 432460 270710
rect 432420 270496 432472 270502
rect 432420 270438 432472 270444
rect 432604 270496 432656 270502
rect 432604 270438 432656 270444
rect 432616 269414 432644 270438
rect 432604 269408 432656 269414
rect 432604 269350 432656 269356
rect 432788 269408 432840 269414
rect 432788 269350 432840 269356
rect 432800 269249 432828 269350
rect 432786 269240 432842 269249
rect 432786 269175 432842 269184
rect 432788 269068 432840 269074
rect 432788 269010 432840 269016
rect 432236 268796 432288 268802
rect 432236 268738 432288 268744
rect 432800 268546 432828 269010
rect 432432 268518 432828 268546
rect 432432 268258 432460 268518
rect 432420 268252 432472 268258
rect 432420 268194 432472 268200
rect 432604 268252 432656 268258
rect 432604 268194 432656 268200
rect 432616 267073 432644 268194
rect 432788 267708 432840 267714
rect 432788 267650 432840 267656
rect 432602 267064 432658 267073
rect 432602 266999 432658 267008
rect 432800 266762 432828 267650
rect 432788 266756 432840 266762
rect 432788 266698 432840 266704
rect 432984 264330 433012 271351
rect 433628 271153 433656 271390
rect 433614 271144 433670 271153
rect 433614 271079 433670 271088
rect 433248 266756 433300 266762
rect 433248 266698 433300 266704
rect 432538 264302 433012 264330
rect 433260 264316 433288 266698
rect 434364 264330 434392 274071
rect 435192 271726 435220 277766
rect 435928 273834 435956 277780
rect 436112 277766 437046 277794
rect 435916 273828 435968 273834
rect 435916 273770 435968 273776
rect 435180 271720 435232 271726
rect 435180 271662 435232 271668
rect 435364 271720 435416 271726
rect 435364 271662 435416 271668
rect 435376 271454 435404 271662
rect 435364 271448 435416 271454
rect 435364 271390 435416 271396
rect 436112 270774 436140 277766
rect 436560 276140 436612 276146
rect 436560 276082 436612 276088
rect 436572 275194 436600 276082
rect 436744 276004 436796 276010
rect 436744 275946 436796 275952
rect 436756 275194 436784 275946
rect 436560 275188 436612 275194
rect 436560 275130 436612 275136
rect 436744 275188 436796 275194
rect 436744 275130 436796 275136
rect 437216 273254 437244 278530
rect 644664 278452 644716 278458
rect 644664 278394 644716 278400
rect 641994 278080 642050 278089
rect 641994 278015 642050 278024
rect 527732 277840 527784 277846
rect 436664 273226 437244 273254
rect 437952 277766 438242 277794
rect 438872 277766 439438 277794
rect 436100 270768 436152 270774
rect 436284 270768 436336 270774
rect 436100 270710 436152 270716
rect 436282 270736 436284 270745
rect 436336 270736 436338 270745
rect 436282 270671 436338 270680
rect 436006 267744 436062 267753
rect 436006 267679 436008 267688
rect 436060 267679 436062 267688
rect 436008 267650 436060 267656
rect 435088 266348 435140 266354
rect 435088 266290 435140 266296
rect 435100 264330 435128 266290
rect 435456 264784 435508 264790
rect 435456 264726 435508 264732
rect 434010 264302 434392 264330
rect 434746 264302 435128 264330
rect 435468 264316 435496 264726
rect 436664 264330 436692 273226
rect 437952 272921 437980 277766
rect 436926 272912 436982 272921
rect 436926 272847 436982 272856
rect 437938 272912 437994 272921
rect 437938 272847 437994 272856
rect 436940 272678 436968 272847
rect 437388 272808 437440 272814
rect 437388 272750 437440 272756
rect 437572 272808 437624 272814
rect 437572 272750 437624 272756
rect 436928 272672 436980 272678
rect 436928 272614 436980 272620
rect 437112 272672 437164 272678
rect 437112 272614 437164 272620
rect 437124 272241 437152 272614
rect 437400 272354 437428 272750
rect 437584 272513 437612 272750
rect 437570 272504 437626 272513
rect 437570 272439 437626 272448
rect 437400 272326 437612 272354
rect 437584 272270 437612 272326
rect 437388 272264 437440 272270
rect 437110 272232 437166 272241
rect 437110 272167 437166 272176
rect 437386 272232 437388 272241
rect 437572 272264 437624 272270
rect 437440 272232 437442 272241
rect 437572 272206 437624 272212
rect 437386 272167 437442 272176
rect 438674 270056 438730 270065
rect 438674 269991 438730 270000
rect 437018 269104 437074 269113
rect 437018 269039 437074 269048
rect 437032 268802 437060 269039
rect 437020 268796 437072 268802
rect 437020 268738 437072 268744
rect 437388 268796 437440 268802
rect 437388 268738 437440 268744
rect 437400 268274 437428 268738
rect 437032 268246 437428 268274
rect 437032 268122 437060 268246
rect 437020 268116 437072 268122
rect 437020 268058 437072 268064
rect 437204 268116 437256 268122
rect 437204 268058 437256 268064
rect 436218 264302 436692 264330
rect 437216 264194 437244 268058
rect 437386 267744 437442 267753
rect 437386 267679 437388 267688
rect 437440 267679 437442 267688
rect 437388 267650 437440 267656
rect 437386 266792 437442 266801
rect 437386 266727 437388 266736
rect 437440 266727 437442 266736
rect 437664 266756 437716 266762
rect 437388 266698 437440 266704
rect 437664 266698 437716 266704
rect 437676 266354 437704 266698
rect 437664 266348 437716 266354
rect 437664 266290 437716 266296
rect 437664 264988 437716 264994
rect 437664 264930 437716 264936
rect 437676 264316 437704 264930
rect 438688 264330 438716 269991
rect 438872 269113 438900 277766
rect 440620 271590 440648 277780
rect 441632 277766 441830 277794
rect 443026 277766 443224 277794
rect 441632 272814 441660 277766
rect 442908 276276 442960 276282
rect 442908 276218 442960 276224
rect 442920 273254 442948 276218
rect 442828 273226 442948 273254
rect 441620 272808 441672 272814
rect 441620 272750 441672 272756
rect 442264 272808 442316 272814
rect 442264 272750 442316 272756
rect 442276 272406 442304 272750
rect 442264 272400 442316 272406
rect 442264 272342 442316 272348
rect 442448 272400 442500 272406
rect 442448 272342 442500 272348
rect 442460 272241 442488 272342
rect 442446 272232 442502 272241
rect 442446 272167 442502 272176
rect 441526 271960 441582 271969
rect 441526 271895 441582 271904
rect 440608 271584 440660 271590
rect 440608 271526 440660 271532
rect 440976 271584 441028 271590
rect 440976 271526 441028 271532
rect 439136 271448 439188 271454
rect 439136 271390 439188 271396
rect 438858 269104 438914 269113
rect 438858 269039 438914 269048
rect 438426 264302 438716 264330
rect 439148 264316 439176 271390
rect 439872 265124 439924 265130
rect 439872 265066 439924 265072
rect 439884 264316 439912 265066
rect 440988 264330 441016 271526
rect 441342 268968 441398 268977
rect 441342 268903 441344 268912
rect 441396 268903 441398 268912
rect 441344 268874 441396 268880
rect 441540 264330 441568 271895
rect 442092 270558 442488 270586
rect 442092 270230 442120 270558
rect 442460 270502 442488 270558
rect 442264 270496 442316 270502
rect 442264 270438 442316 270444
rect 442448 270496 442500 270502
rect 442448 270438 442500 270444
rect 442276 270230 442304 270438
rect 442080 270224 442132 270230
rect 442080 270166 442132 270172
rect 442264 270224 442316 270230
rect 442264 270166 442316 270172
rect 442080 268660 442132 268666
rect 442080 268602 442132 268608
rect 442092 268258 442120 268602
rect 442080 268252 442132 268258
rect 442080 268194 442132 268200
rect 442448 268116 442500 268122
rect 442448 268058 442500 268064
rect 442460 266801 442488 268058
rect 442446 266792 442502 266801
rect 442446 266727 442502 266736
rect 442080 266212 442132 266218
rect 442080 266154 442132 266160
rect 440634 264302 441016 264330
rect 441370 264302 441568 264330
rect 442092 264316 442120 266154
rect 442828 264316 442856 273226
rect 443196 268977 443224 277766
rect 443840 277766 444222 277794
rect 444944 277766 445326 277794
rect 443840 273086 443868 277766
rect 443828 273080 443880 273086
rect 443828 273022 443880 273028
rect 444012 273080 444064 273086
rect 444012 273022 444064 273028
rect 444024 272406 444052 273022
rect 444012 272400 444064 272406
rect 444012 272342 444064 272348
rect 444196 272400 444248 272406
rect 444196 272342 444248 272348
rect 444208 271969 444236 272342
rect 444194 271960 444250 271969
rect 444194 271895 444250 271904
rect 444944 270502 444972 277766
rect 446218 275496 446274 275505
rect 446218 275431 446274 275440
rect 446232 273254 446260 275431
rect 446508 273834 446536 277780
rect 446496 273828 446548 273834
rect 446496 273770 446548 273776
rect 446404 273692 446456 273698
rect 446404 273634 446456 273640
rect 446416 273290 446444 273634
rect 446048 273226 446260 273254
rect 446404 273284 446456 273290
rect 446404 273226 446456 273232
rect 445390 272232 445446 272241
rect 445390 272167 445446 272176
rect 444932 270496 444984 270502
rect 444932 270438 444984 270444
rect 445116 270496 445168 270502
rect 445116 270438 445168 270444
rect 443550 270328 443606 270337
rect 443550 270263 443606 270272
rect 443182 268968 443238 268977
rect 443182 268903 443238 268912
rect 443564 264316 443592 270263
rect 445128 270065 445156 270438
rect 445114 270056 445170 270065
rect 445114 269991 445170 270000
rect 444288 265396 444340 265402
rect 444288 265338 444340 265344
rect 444300 264316 444328 265338
rect 445404 264330 445432 272167
rect 446048 271425 446076 273226
rect 447704 272270 447732 277780
rect 448532 277766 448914 277794
rect 449912 277766 450110 277794
rect 448152 273828 448204 273834
rect 448152 273770 448204 273776
rect 447692 272264 447744 272270
rect 447876 272264 447928 272270
rect 447692 272206 447744 272212
rect 447874 272232 447876 272241
rect 447928 272232 447930 272241
rect 447874 272167 447930 272176
rect 447094 271584 447146 271590
rect 446692 271532 447094 271538
rect 446692 271526 447146 271532
rect 446692 271510 447134 271526
rect 446692 271454 446720 271510
rect 446680 271448 446732 271454
rect 446034 271416 446090 271425
rect 446034 271351 446090 271360
rect 446310 271416 446366 271425
rect 446680 271390 446732 271396
rect 446310 271351 446366 271360
rect 446324 267734 446352 271351
rect 447048 268932 447100 268938
rect 447048 268874 447100 268880
rect 447060 268569 447088 268874
rect 447046 268560 447102 268569
rect 447046 268495 447102 268504
rect 446140 267706 446352 267734
rect 446140 264330 446168 267706
rect 446862 266248 446918 266257
rect 446862 266183 446918 266192
rect 446876 264330 446904 266183
rect 447600 266076 447652 266082
rect 447600 266018 447652 266024
rect 447612 264330 447640 266018
rect 448164 264330 448192 273770
rect 448334 271960 448390 271969
rect 448334 271895 448390 271904
rect 448348 266082 448376 271895
rect 448532 268569 448560 277766
rect 449714 273184 449770 273193
rect 449714 273119 449770 273128
rect 448518 268560 448574 268569
rect 448518 268495 448574 268504
rect 448704 266348 448756 266354
rect 448704 266290 448756 266296
rect 448336 266076 448388 266082
rect 448336 266018 448388 266024
rect 448520 266076 448572 266082
rect 448520 266018 448572 266024
rect 448532 265538 448560 266018
rect 448520 265532 448572 265538
rect 448520 265474 448572 265480
rect 445050 264302 445432 264330
rect 445786 264302 446168 264330
rect 446522 264302 446904 264330
rect 447258 264302 447640 264330
rect 447994 264302 448192 264330
rect 448716 264316 448744 266290
rect 449070 266248 449126 266257
rect 448888 266212 448940 266218
rect 449070 266183 449072 266192
rect 448888 266154 448940 266160
rect 449124 266183 449126 266192
rect 449072 266154 449124 266160
rect 448900 265402 448928 266154
rect 448888 265396 448940 265402
rect 448888 265338 448940 265344
rect 449728 264330 449756 273119
rect 449912 269074 449940 277766
rect 450728 276140 450780 276146
rect 450728 276082 450780 276088
rect 450544 273080 450596 273086
rect 450544 273022 450596 273028
rect 450556 272921 450584 273022
rect 450542 272912 450598 272921
rect 450542 272847 450598 272856
rect 449900 269068 449952 269074
rect 449900 269010 449952 269016
rect 450174 267064 450230 267073
rect 450174 266999 450230 267008
rect 449466 264302 449756 264330
rect 450188 264316 450216 266999
rect 450740 264330 450768 276082
rect 451004 273216 451056 273222
rect 451002 273184 451004 273193
rect 451056 273184 451058 273193
rect 451002 273119 451058 273128
rect 451292 273086 451320 277780
rect 452120 277766 452502 277794
rect 452672 277766 453606 277794
rect 454236 277766 454802 277794
rect 451280 273080 451332 273086
rect 451280 273022 451332 273028
rect 451096 272944 451148 272950
rect 452120 272921 452148 277766
rect 451096 272886 451148 272892
rect 452106 272912 452162 272921
rect 451108 271969 451136 272886
rect 452106 272847 452162 272856
rect 452106 272504 452162 272513
rect 452106 272439 452162 272448
rect 451094 271960 451150 271969
rect 451094 271895 451150 271904
rect 451246 271646 451596 271674
rect 451246 271590 451274 271646
rect 451234 271584 451286 271590
rect 451234 271526 451286 271532
rect 451372 271584 451424 271590
rect 451372 271526 451424 271532
rect 451384 271425 451412 271526
rect 451568 271425 451596 271646
rect 451370 271416 451426 271425
rect 451370 271351 451426 271360
rect 451554 271416 451610 271425
rect 451554 271351 451610 271360
rect 452120 264330 452148 272439
rect 452384 268932 452436 268938
rect 452384 268874 452436 268880
rect 450740 264302 450938 264330
rect 451674 264302 452148 264330
rect 452396 264316 452424 268874
rect 452672 268802 452700 277766
rect 454040 273080 454092 273086
rect 454040 273022 454092 273028
rect 453762 272912 453818 272921
rect 453762 272847 453818 272856
rect 453120 269068 453172 269074
rect 453120 269010 453172 269016
rect 452660 268796 452712 268802
rect 452660 268738 452712 268744
rect 453132 264316 453160 269010
rect 453776 264330 453804 272847
rect 454052 272814 454080 273022
rect 454040 272808 454092 272814
rect 454040 272750 454092 272756
rect 454236 272542 454264 277766
rect 454866 273864 454922 273873
rect 454866 273799 454922 273808
rect 454684 272944 454736 272950
rect 454682 272912 454684 272921
rect 454736 272912 454738 272921
rect 454682 272847 454738 272856
rect 454224 272536 454276 272542
rect 454408 272536 454460 272542
rect 454224 272478 454276 272484
rect 454406 272504 454408 272513
rect 454460 272504 454462 272513
rect 454406 272439 454462 272448
rect 454880 267073 454908 273799
rect 455984 272678 456012 277780
rect 457180 276962 457208 277780
rect 458192 277766 458390 277794
rect 459586 277766 459876 277794
rect 457444 277228 457496 277234
rect 457444 277170 457496 277176
rect 457168 276956 457220 276962
rect 457168 276898 457220 276904
rect 457456 273254 457484 277170
rect 457088 273226 457484 273254
rect 455972 272672 456024 272678
rect 455972 272614 456024 272620
rect 456524 272536 456576 272542
rect 456524 272478 456576 272484
rect 455142 269240 455198 269249
rect 455142 269175 455198 269184
rect 455156 268530 455184 269175
rect 455604 268932 455656 268938
rect 455604 268874 455656 268880
rect 455616 268666 455644 268874
rect 455604 268660 455656 268666
rect 455604 268602 455656 268608
rect 455144 268524 455196 268530
rect 455144 268466 455196 268472
rect 455328 268524 455380 268530
rect 455328 268466 455380 268472
rect 454866 267064 454922 267073
rect 454866 266999 454922 267008
rect 454958 266384 455014 266393
rect 454958 266319 455014 266328
rect 454972 264330 455000 266319
rect 453776 264302 453882 264330
rect 454618 264302 455000 264330
rect 455340 264316 455368 268466
rect 456536 264330 456564 272478
rect 456890 271416 456946 271425
rect 456890 271351 456946 271360
rect 456904 271182 456932 271351
rect 456754 271176 456806 271182
rect 456752 271144 456754 271153
rect 456892 271176 456944 271182
rect 456806 271144 456808 271153
rect 456892 271118 456944 271124
rect 456752 271079 456808 271088
rect 456798 269240 456854 269249
rect 456798 269175 456854 269184
rect 456812 268938 456840 269175
rect 456800 268932 456852 268938
rect 456800 268874 456852 268880
rect 457088 266506 457116 273226
rect 458192 273086 458220 277766
rect 458180 273080 458232 273086
rect 458180 273022 458232 273028
rect 458638 272232 458694 272241
rect 458638 272167 458694 272176
rect 457902 268152 457958 268161
rect 457902 268087 457958 268096
rect 456766 266478 457116 266506
rect 456766 266218 456794 266478
rect 456890 266384 456946 266393
rect 456890 266319 456946 266328
rect 457166 266384 457222 266393
rect 457166 266319 457222 266328
rect 456904 266218 456932 266319
rect 456754 266212 456806 266218
rect 456754 266154 456806 266160
rect 456892 266212 456944 266218
rect 456892 266154 456944 266160
rect 457180 264330 457208 266319
rect 457916 264330 457944 268087
rect 458652 264330 458680 272167
rect 459848 270366 459876 277766
rect 460032 277766 460690 277794
rect 461504 277766 461886 277794
rect 462332 277766 463082 277794
rect 464080 277766 464278 277794
rect 465184 277766 465474 277794
rect 459836 270360 459888 270366
rect 459836 270302 459888 270308
rect 459374 270056 459430 270065
rect 459374 269991 459430 270000
rect 459388 264330 459416 269991
rect 460032 268938 460060 277766
rect 460938 274408 460994 274417
rect 460938 274343 460994 274352
rect 460952 273986 460980 274343
rect 460768 273958 460980 273986
rect 460768 273698 460796 273958
rect 461030 273864 461086 273873
rect 461030 273799 461032 273808
rect 461084 273799 461086 273808
rect 461032 273770 461084 273776
rect 460756 273692 460808 273698
rect 460756 273634 460808 273640
rect 461504 273254 461532 277766
rect 461504 273226 461624 273254
rect 461400 273080 461452 273086
rect 461400 273022 461452 273028
rect 461412 272678 461440 273022
rect 461400 272672 461452 272678
rect 461400 272614 461452 272620
rect 460846 272504 460902 272513
rect 460846 272439 460902 272448
rect 460020 268932 460072 268938
rect 460020 268874 460072 268880
rect 460110 268424 460166 268433
rect 460110 268359 460166 268368
rect 460124 264330 460152 268359
rect 460860 264330 460888 272439
rect 461596 271318 461624 273226
rect 461768 272536 461820 272542
rect 461766 272504 461768 272513
rect 461820 272504 461822 272513
rect 461766 272439 461822 272448
rect 461584 271312 461636 271318
rect 461584 271254 461636 271260
rect 461768 271312 461820 271318
rect 461768 271254 461820 271260
rect 461780 271153 461808 271254
rect 461766 271144 461822 271153
rect 461766 271079 461822 271088
rect 461768 270224 461820 270230
rect 461768 270166 461820 270172
rect 461780 270065 461808 270166
rect 461766 270056 461822 270065
rect 461766 269991 461822 270000
rect 462332 269226 462360 277766
rect 464080 273254 464108 277766
rect 463988 273226 464108 273254
rect 462502 271280 462558 271289
rect 462502 271215 462558 271224
rect 461412 269198 462360 269226
rect 461412 268938 461440 269198
rect 461596 269074 461808 269090
rect 461596 269068 461820 269074
rect 461596 269062 461768 269068
rect 461400 268932 461452 268938
rect 461400 268874 461452 268880
rect 461596 268818 461624 269062
rect 461768 269010 461820 269016
rect 461860 268932 461912 268938
rect 461860 268874 461912 268880
rect 461412 268790 461624 268818
rect 461412 268666 461440 268790
rect 461582 268696 461638 268705
rect 461400 268660 461452 268666
rect 461872 268682 461900 268874
rect 462136 268796 462188 268802
rect 462136 268738 462188 268744
rect 461582 268631 461638 268640
rect 461780 268654 461900 268682
rect 461400 268602 461452 268608
rect 461030 266112 461086 266121
rect 461030 266047 461086 266056
rect 461044 265946 461072 266047
rect 461032 265940 461084 265946
rect 461032 265882 461084 265888
rect 461216 264648 461268 264654
rect 461216 264590 461268 264596
rect 456090 264302 456564 264330
rect 456826 264302 457208 264330
rect 457562 264302 457944 264330
rect 458298 264302 458680 264330
rect 459034 264302 459416 264330
rect 459770 264302 460152 264330
rect 460506 264302 460888 264330
rect 461228 264316 461256 264590
rect 461596 264330 461624 268631
rect 461780 268530 461808 268654
rect 461768 268524 461820 268530
rect 461768 268466 461820 268472
rect 461952 268524 462004 268530
rect 461952 268466 462004 268472
rect 461964 268161 461992 268466
rect 462148 268394 462176 268738
rect 462318 268424 462374 268433
rect 462136 268388 462188 268394
rect 462318 268359 462320 268368
rect 462136 268330 462188 268336
rect 462372 268359 462374 268368
rect 462320 268330 462372 268336
rect 461950 268152 462006 268161
rect 461950 268087 462006 268096
rect 462516 266393 462544 271215
rect 463606 266792 463662 266801
rect 463606 266727 463662 266736
rect 462502 266384 462558 266393
rect 462502 266319 462558 266328
rect 461766 266112 461822 266121
rect 461766 266047 461768 266056
rect 461820 266047 461822 266056
rect 461768 266018 461820 266024
rect 462686 265840 462742 265849
rect 462686 265775 462742 265784
rect 461596 264302 461978 264330
rect 462700 264316 462728 265775
rect 463620 264330 463648 266727
rect 463988 266082 464016 273226
rect 464894 272504 464950 272513
rect 464894 272439 464950 272448
rect 464710 268152 464766 268161
rect 464710 268087 464766 268096
rect 464724 267442 464752 268087
rect 464712 267436 464764 267442
rect 464712 267378 464764 267384
rect 463976 266076 464028 266082
rect 463976 266018 464028 266024
rect 464160 266076 464212 266082
rect 464160 266018 464212 266024
rect 463450 264302 463648 264330
rect 464172 264316 464200 266018
rect 464908 264316 464936 272439
rect 465184 271318 465212 277766
rect 466656 276010 466684 277780
rect 467656 277432 467708 277438
rect 467656 277374 467708 277380
rect 465724 276004 465776 276010
rect 465724 275946 465776 275952
rect 465908 276004 465960 276010
rect 465908 275946 465960 275952
rect 466644 276004 466696 276010
rect 466644 275946 466696 275952
rect 467104 276004 467156 276010
rect 467104 275946 467156 275952
rect 465736 275330 465764 275946
rect 465540 275324 465592 275330
rect 465540 275266 465592 275272
rect 465724 275324 465776 275330
rect 465724 275266 465776 275272
rect 465552 275210 465580 275266
rect 465920 275210 465948 275946
rect 465552 275182 465948 275210
rect 467116 273254 467144 275946
rect 467668 273254 467696 277374
rect 467852 276826 467880 277780
rect 468036 277766 468970 277794
rect 469232 277766 470166 277794
rect 470612 277766 471362 277794
rect 472176 277766 472558 277794
rect 473464 277766 473754 277794
rect 474752 277766 474950 277794
rect 467840 276820 467892 276826
rect 467840 276762 467892 276768
rect 467116 273226 467512 273254
rect 466274 272776 466330 272785
rect 466274 272711 466330 272720
rect 466288 272542 466316 272711
rect 466276 272536 466328 272542
rect 466276 272478 466328 272484
rect 466460 272536 466512 272542
rect 466460 272478 466512 272484
rect 466472 272354 466500 272478
rect 466288 272326 466500 272354
rect 466288 272241 466316 272326
rect 466274 272232 466330 272241
rect 466274 272167 466330 272176
rect 466458 271416 466514 271425
rect 466458 271351 466514 271360
rect 465172 271312 465224 271318
rect 465356 271312 465408 271318
rect 465172 271254 465224 271260
rect 465354 271280 465356 271289
rect 465408 271280 465410 271289
rect 466472 271266 466500 271351
rect 465354 271215 465410 271224
rect 466426 271238 466500 271266
rect 466426 271182 466454 271238
rect 466414 271176 466466 271182
rect 465998 271144 466054 271153
rect 466552 271176 466604 271182
rect 466414 271118 466466 271124
rect 466550 271144 466552 271153
rect 466604 271144 466606 271153
rect 465998 271079 466054 271088
rect 466550 271079 466606 271088
rect 465816 266484 465868 266490
rect 465816 266426 465868 266432
rect 465828 265305 465856 266426
rect 465814 265296 465870 265305
rect 465814 265231 465870 265240
rect 466012 264330 466040 271079
rect 466458 268968 466514 268977
rect 466458 268903 466514 268912
rect 466472 268818 466500 268903
rect 466426 268802 466500 268818
rect 466414 268796 466500 268802
rect 466466 268790 466500 268796
rect 467012 268796 467064 268802
rect 466414 268738 466466 268744
rect 467012 268738 467064 268744
rect 466288 268666 466868 268682
rect 466276 268660 466880 268666
rect 466328 268654 466828 268660
rect 466276 268602 466328 268608
rect 466828 268602 466880 268608
rect 467024 268546 467052 268738
rect 466564 268518 467052 268546
rect 466366 268424 466422 268433
rect 466564 268394 466592 268518
rect 466734 268424 466790 268433
rect 466366 268359 466422 268368
rect 466552 268388 466604 268394
rect 466182 267608 466238 267617
rect 466182 267543 466238 267552
rect 466196 267170 466224 267543
rect 466184 267164 466236 267170
rect 466184 267106 466236 267112
rect 466184 267028 466236 267034
rect 466184 266970 466236 266976
rect 466196 266529 466224 266970
rect 466182 266520 466238 266529
rect 466182 266455 466238 266464
rect 465658 264302 466040 264330
rect 466380 264316 466408 268359
rect 466734 268359 466736 268368
rect 466552 268330 466604 268336
rect 466788 268359 466790 268368
rect 466736 268330 466788 268336
rect 467010 267608 467066 267617
rect 467010 267543 467066 267552
rect 466828 267436 466880 267442
rect 466828 267378 466880 267384
rect 466840 267073 466868 267378
rect 467024 267170 467052 267543
rect 467012 267164 467064 267170
rect 467012 267106 467064 267112
rect 466826 267064 466882 267073
rect 466826 266999 466882 267008
rect 466920 266484 466972 266490
rect 466920 266426 466972 266432
rect 466932 265305 466960 266426
rect 467484 265962 467512 273226
rect 467392 265946 467512 265962
rect 467380 265940 467512 265946
rect 467432 265934 467512 265940
rect 467576 273226 467696 273254
rect 467380 265882 467432 265888
rect 466918 265296 466974 265305
rect 466918 265231 466974 265240
rect 467576 264330 467604 273226
rect 468036 268977 468064 277766
rect 469036 276820 469088 276826
rect 469036 276762 469088 276768
rect 469048 273254 469076 276762
rect 468956 273226 469076 273254
rect 468022 268968 468078 268977
rect 468022 268903 468078 268912
rect 468206 267744 468262 267753
rect 468206 267679 468262 267688
rect 468220 264330 468248 267679
rect 467130 264302 467604 264330
rect 467866 264302 468248 264330
rect 468956 264194 468984 273226
rect 469232 268161 469260 277766
rect 470230 274680 470286 274689
rect 470230 274615 470232 274624
rect 470284 274615 470286 274624
rect 470416 274644 470468 274650
rect 470232 274586 470284 274592
rect 470416 274586 470468 274592
rect 470428 274417 470456 274586
rect 470414 274408 470470 274417
rect 470414 274343 470470 274352
rect 470612 273254 470640 277766
rect 472176 274689 472204 277766
rect 472992 276956 473044 276962
rect 472992 276898 473044 276904
rect 472162 274680 472218 274689
rect 472162 274615 472218 274624
rect 470612 273226 470732 273254
rect 469600 270422 469996 270450
rect 469600 269550 469628 270422
rect 469968 270366 469996 270422
rect 469772 270360 469824 270366
rect 469772 270302 469824 270308
rect 469956 270360 470008 270366
rect 469956 270302 470008 270308
rect 469784 269550 469812 270302
rect 470506 270056 470562 270065
rect 470506 269991 470562 270000
rect 469588 269544 469640 269550
rect 469588 269486 469640 269492
rect 469772 269544 469824 269550
rect 469772 269486 469824 269492
rect 469218 268152 469274 268161
rect 469218 268087 469274 268096
rect 470520 267306 470548 269991
rect 469680 267300 469732 267306
rect 469680 267242 469732 267248
rect 470508 267300 470560 267306
rect 470508 267242 470560 267248
rect 469692 264330 469720 267242
rect 470046 267064 470102 267073
rect 470046 266999 470102 267008
rect 469338 264302 469720 264330
rect 470060 264316 470088 266999
rect 470704 266098 470732 273226
rect 472254 270600 472310 270609
rect 472254 270535 472310 270544
rect 471426 267744 471482 267753
rect 471426 267679 471428 267688
rect 471480 267679 471482 267688
rect 471428 267650 471480 267656
rect 471060 267572 471112 267578
rect 471060 267514 471112 267520
rect 471072 267306 471100 267514
rect 471060 267300 471112 267306
rect 471060 267242 471112 267248
rect 470612 266070 470732 266098
rect 470612 265810 470640 266070
rect 470784 265940 470836 265946
rect 470784 265882 470836 265888
rect 470600 265804 470652 265810
rect 470600 265746 470652 265752
rect 470796 264316 470824 265882
rect 471888 264512 471940 264518
rect 471888 264454 471940 264460
rect 471900 264330 471928 264454
rect 471546 264302 471928 264330
rect 472268 264316 472296 270535
rect 473004 264316 473032 276898
rect 473464 275602 473492 277766
rect 473452 275596 473504 275602
rect 473452 275538 473504 275544
rect 474004 275596 474056 275602
rect 474004 275538 474056 275544
rect 473726 268152 473782 268161
rect 473726 268087 473782 268096
rect 473740 264316 473768 268087
rect 474016 266801 474044 275538
rect 474752 270366 474780 277766
rect 475212 276134 475792 276162
rect 475212 275602 475240 276134
rect 475764 276010 475792 276134
rect 475568 276004 475620 276010
rect 475568 275946 475620 275952
rect 475752 276004 475804 276010
rect 475752 275946 475804 275952
rect 475200 275596 475252 275602
rect 475200 275538 475252 275544
rect 475384 275596 475436 275602
rect 475384 275538 475436 275544
rect 475396 275330 475424 275538
rect 475580 275330 475608 275946
rect 475384 275324 475436 275330
rect 475384 275266 475436 275272
rect 475568 275324 475620 275330
rect 475568 275266 475620 275272
rect 475384 274644 475436 274650
rect 475384 274586 475436 274592
rect 475568 274644 475620 274650
rect 475568 274586 475620 274592
rect 475396 274242 475424 274586
rect 475200 274236 475252 274242
rect 475200 274178 475252 274184
rect 475384 274236 475436 274242
rect 475384 274178 475436 274184
rect 475212 274122 475240 274178
rect 475580 274122 475608 274586
rect 475842 274408 475898 274417
rect 476132 274378 476160 277780
rect 476316 277766 477250 277794
rect 477512 277766 478446 277794
rect 475842 274343 475898 274352
rect 476120 274372 476172 274378
rect 475212 274094 475608 274122
rect 475660 272400 475712 272406
rect 475660 272342 475712 272348
rect 475672 272241 475700 272342
rect 475658 272232 475714 272241
rect 475658 272167 475714 272176
rect 474740 270360 474792 270366
rect 474740 270302 474792 270308
rect 474924 270360 474976 270366
rect 474924 270302 474976 270308
rect 474936 270065 474964 270302
rect 474922 270056 474978 270065
rect 474922 269991 474978 270000
rect 475566 268424 475622 268433
rect 475566 268359 475622 268368
rect 474002 266792 474058 266801
rect 474002 266727 474058 266736
rect 474646 266792 474702 266801
rect 474646 266727 474702 266736
rect 474660 264330 474688 266727
rect 475580 264330 475608 268359
rect 474490 264302 474688 264330
rect 475226 264302 475608 264330
rect 475856 264330 475884 274343
rect 476120 274314 476172 274320
rect 476026 272776 476082 272785
rect 476026 272711 476082 272720
rect 476040 272406 476068 272711
rect 476028 272400 476080 272406
rect 476028 272342 476080 272348
rect 476028 269816 476080 269822
rect 476028 269758 476080 269764
rect 476040 269249 476068 269758
rect 476026 269240 476082 269249
rect 476026 269175 476082 269184
rect 476316 267306 476344 277766
rect 477040 269816 477092 269822
rect 477040 269758 477092 269764
rect 476304 267300 476356 267306
rect 476304 267242 476356 267248
rect 476488 267300 476540 267306
rect 476488 267242 476540 267248
rect 476500 266762 476528 267242
rect 476488 266756 476540 266762
rect 476488 266698 476540 266704
rect 477052 264330 477080 269758
rect 477512 269249 477540 277766
rect 479628 274650 479656 277780
rect 480168 276004 480220 276010
rect 480168 275946 480220 275952
rect 480352 276004 480404 276010
rect 480352 275946 480404 275952
rect 480180 275777 480208 275946
rect 480364 275777 480392 275946
rect 480166 275768 480222 275777
rect 480166 275703 480222 275712
rect 480350 275768 480406 275777
rect 480824 275738 480852 277780
rect 481652 277766 482034 277794
rect 480350 275703 480406 275712
rect 480812 275732 480864 275738
rect 480812 275674 480864 275680
rect 480996 275732 481048 275738
rect 480996 275674 481048 275680
rect 479996 275590 480392 275618
rect 479616 274644 479668 274650
rect 479616 274586 479668 274592
rect 479800 274644 479852 274650
rect 479800 274586 479852 274592
rect 479812 274417 479840 274586
rect 479798 274408 479854 274417
rect 478604 274372 478656 274378
rect 479798 274343 479854 274352
rect 478604 274314 478656 274320
rect 477498 269240 477554 269249
rect 477498 269175 477554 269184
rect 477408 265804 477460 265810
rect 477408 265746 477460 265752
rect 475856 264302 475962 264330
rect 476698 264302 477080 264330
rect 477420 264316 477448 265746
rect 478616 264330 478644 274314
rect 479996 272898 480024 275590
rect 480364 275466 480392 275590
rect 481008 275482 481036 275674
rect 480168 275460 480220 275466
rect 480168 275402 480220 275408
rect 480352 275460 480404 275466
rect 480352 275402 480404 275408
rect 480548 275454 481036 275482
rect 480180 275346 480208 275402
rect 480548 275346 480576 275454
rect 480180 275318 480576 275346
rect 481454 275224 481510 275233
rect 481454 275159 481510 275168
rect 479536 272870 480024 272898
rect 479536 267034 479564 272870
rect 480074 272776 480130 272785
rect 480074 272711 480130 272720
rect 480994 272776 481050 272785
rect 480994 272711 481050 272720
rect 480088 272406 480116 272711
rect 480076 272400 480128 272406
rect 480076 272342 480128 272348
rect 480214 272400 480266 272406
rect 480214 272342 480266 272348
rect 480074 272232 480130 272241
rect 480226 272218 480254 272342
rect 481008 272241 481036 272711
rect 480130 272190 480254 272218
rect 480994 272232 481050 272241
rect 480074 272167 480130 272176
rect 480994 272167 481050 272176
rect 480260 271584 480312 271590
rect 480260 271526 480312 271532
rect 480536 271584 480588 271590
rect 480536 271526 480588 271532
rect 480272 271266 480300 271526
rect 480548 271425 480576 271526
rect 480534 271416 480590 271425
rect 480534 271351 480590 271360
rect 480720 271312 480772 271318
rect 480272 271260 480720 271266
rect 480272 271254 480772 271260
rect 480272 271238 480760 271254
rect 480260 271176 480312 271182
rect 480442 271144 480498 271153
rect 480312 271124 480442 271130
rect 480260 271118 480442 271124
rect 480272 271102 480442 271118
rect 480442 271079 480498 271088
rect 480074 270056 480130 270065
rect 480074 269991 480130 270000
rect 480088 269822 480116 269991
rect 480536 269952 480588 269958
rect 480536 269894 480588 269900
rect 480076 269816 480128 269822
rect 480076 269758 480128 269764
rect 480258 268968 480314 268977
rect 480258 268903 480314 268912
rect 480272 268546 480300 268903
rect 480088 268530 480300 268546
rect 480076 268524 480300 268530
rect 480128 268518 480300 268524
rect 480076 268466 480128 268472
rect 480350 268424 480406 268433
rect 480350 268359 480352 268368
rect 480404 268359 480406 268368
rect 480352 268330 480404 268336
rect 480548 267734 480576 269894
rect 480272 267706 480576 267734
rect 480272 267594 480300 267706
rect 480180 267566 480300 267594
rect 480180 267442 480208 267566
rect 480168 267436 480220 267442
rect 480168 267378 480220 267384
rect 480352 267436 480404 267442
rect 480352 267378 480404 267384
rect 479524 267028 479576 267034
rect 479524 266970 479576 266976
rect 479708 267028 479760 267034
rect 479708 266970 479760 266976
rect 479720 266762 479748 266970
rect 479890 266792 479946 266801
rect 478880 266756 478932 266762
rect 478880 266698 478932 266704
rect 479708 266756 479760 266762
rect 479890 266727 479892 266736
rect 479708 266698 479760 266704
rect 479944 266727 479946 266736
rect 479892 266698 479944 266704
rect 478170 264302 478644 264330
rect 478892 264316 478920 266698
rect 479614 265840 479670 265849
rect 479614 265775 479670 265784
rect 479628 264316 479656 265775
rect 480364 264316 480392 267378
rect 481468 264330 481496 275159
rect 481652 269550 481680 277766
rect 483018 276040 483074 276049
rect 483018 275975 483074 275984
rect 482558 274408 482614 274417
rect 482558 274343 482614 274352
rect 481640 269544 481692 269550
rect 481640 269486 481692 269492
rect 482192 264376 482244 264382
rect 481114 264302 481496 264330
rect 481850 264324 482192 264330
rect 481850 264318 482244 264324
rect 481850 264302 482232 264318
rect 482572 264316 482600 274343
rect 483032 270065 483060 275975
rect 483216 274106 483244 277780
rect 484320 276010 484348 277780
rect 484504 277766 485530 277794
rect 484308 276004 484360 276010
rect 484308 275946 484360 275952
rect 483204 274100 483256 274106
rect 483204 274042 483256 274048
rect 483018 270056 483074 270065
rect 483018 269991 483074 270000
rect 484504 269822 484532 277766
rect 485780 276004 485832 276010
rect 485780 275946 485832 275952
rect 484860 275460 484912 275466
rect 484860 275402 484912 275408
rect 485044 275460 485096 275466
rect 485044 275402 485096 275408
rect 484872 275074 484900 275402
rect 485056 275194 485084 275402
rect 485044 275188 485096 275194
rect 485044 275130 485096 275136
rect 485228 275188 485280 275194
rect 485228 275130 485280 275136
rect 485240 275074 485268 275130
rect 484872 275046 485268 275074
rect 485044 274236 485096 274242
rect 485044 274178 485096 274184
rect 485228 274236 485280 274242
rect 485228 274178 485280 274184
rect 485056 273970 485084 274178
rect 485044 273964 485096 273970
rect 485044 273906 485096 273912
rect 484492 269816 484544 269822
rect 484492 269758 484544 269764
rect 484308 269544 484360 269550
rect 484308 269486 484360 269492
rect 483110 267608 483166 267617
rect 483110 267543 483166 267552
rect 483124 267442 483152 267543
rect 483112 267436 483164 267442
rect 483112 267378 483164 267384
rect 483296 267436 483348 267442
rect 483296 267378 483348 267384
rect 483308 264316 483336 267378
rect 484320 264330 484348 269486
rect 485240 264330 485268 274178
rect 485594 270872 485650 270881
rect 485594 270807 485650 270816
rect 485608 267734 485636 270807
rect 485792 270609 485820 275946
rect 486712 274106 486740 277780
rect 487908 275738 487936 277780
rect 488552 277766 489118 277794
rect 487896 275732 487948 275738
rect 487896 275674 487948 275680
rect 488080 275732 488132 275738
rect 488080 275674 488132 275680
rect 486700 274100 486752 274106
rect 486700 274042 486752 274048
rect 487068 274100 487120 274106
rect 487068 274042 487120 274048
rect 485778 270600 485834 270609
rect 485778 270535 485834 270544
rect 486240 269816 486292 269822
rect 486240 269758 486292 269764
rect 484058 264302 484348 264330
rect 484794 264302 485268 264330
rect 485516 267706 485636 267734
rect 485516 264316 485544 267706
rect 486252 264316 486280 269758
rect 487080 267734 487108 274042
rect 487802 273048 487858 273057
rect 487802 272983 487858 272992
rect 487618 272776 487674 272785
rect 487618 272711 487674 272720
rect 487632 272406 487660 272711
rect 487620 272400 487672 272406
rect 487620 272342 487672 272348
rect 487816 272134 487844 272983
rect 487804 272128 487856 272134
rect 487804 272070 487856 272076
rect 487618 271960 487674 271969
rect 487618 271895 487674 271904
rect 487632 271318 487660 271895
rect 488092 271674 488120 275674
rect 487816 271646 488120 271674
rect 487620 271312 487672 271318
rect 487620 271254 487672 271260
rect 486988 267706 487108 267734
rect 486988 264316 487016 267706
rect 487816 267170 487844 271646
rect 488552 270042 488580 277766
rect 489918 276040 489974 276049
rect 489736 276004 489788 276010
rect 489918 275975 489920 275984
rect 489736 275946 489788 275952
rect 489972 275975 489974 275984
rect 490102 276040 490158 276049
rect 490102 275975 490158 275984
rect 489920 275946 489972 275952
rect 489748 275777 489776 275946
rect 490116 275890 490144 275975
rect 489886 275862 490144 275890
rect 489734 275768 489790 275777
rect 489886 275738 489914 275862
rect 490010 275768 490066 275777
rect 489734 275703 489790 275712
rect 489874 275732 489926 275738
rect 490010 275703 490012 275712
rect 489874 275674 489926 275680
rect 490064 275703 490066 275712
rect 490012 275674 490064 275680
rect 490300 275482 490328 277780
rect 491496 276049 491524 277780
rect 492232 277766 492614 277794
rect 493060 277766 493810 277794
rect 494532 277766 495006 277794
rect 495820 277766 496202 277794
rect 497016 277766 497398 277794
rect 492232 276554 492260 277766
rect 492220 276548 492272 276554
rect 492220 276490 492272 276496
rect 491850 276176 491906 276185
rect 491850 276111 491906 276120
rect 491482 276040 491538 276049
rect 491482 275975 491538 275984
rect 490116 275454 490328 275482
rect 489874 275188 489926 275194
rect 489874 275130 489926 275136
rect 489886 275074 489914 275130
rect 489886 275046 489960 275074
rect 489932 274961 489960 275046
rect 489918 274952 489974 274961
rect 489918 274887 489974 274896
rect 490116 274666 490144 275454
rect 489932 274638 490144 274666
rect 489932 274514 489960 274638
rect 490470 274544 490526 274553
rect 489920 274508 489972 274514
rect 489920 274450 489972 274456
rect 490104 274508 490156 274514
rect 490470 274479 490526 274488
rect 490104 274450 490156 274456
rect 489734 274408 489790 274417
rect 489790 274366 489960 274394
rect 489734 274343 489790 274352
rect 489932 274242 489960 274366
rect 489736 274236 489788 274242
rect 489736 274178 489788 274184
rect 489920 274236 489972 274242
rect 489920 274178 489972 274184
rect 489458 273864 489514 273873
rect 489458 273799 489514 273808
rect 489276 271584 489328 271590
rect 489276 271526 489328 271532
rect 489288 271425 489316 271526
rect 489274 271416 489330 271425
rect 489274 271351 489330 271360
rect 488000 270014 488580 270042
rect 488000 269793 488028 270014
rect 488172 269952 488224 269958
rect 488170 269920 488172 269929
rect 488356 269952 488408 269958
rect 488224 269920 488226 269929
rect 488356 269894 488408 269900
rect 488170 269855 488226 269864
rect 487986 269784 488042 269793
rect 487986 269719 488042 269728
rect 487804 267164 487856 267170
rect 487804 267106 487856 267112
rect 488078 266792 488134 266801
rect 488078 266727 488134 266736
rect 488092 264330 488120 266727
rect 487738 264302 488120 264330
rect 488368 264330 488396 269894
rect 489472 264330 489500 273799
rect 489748 273601 489776 274178
rect 490116 273601 490144 274450
rect 489734 273592 489790 273601
rect 489734 273527 489790 273536
rect 490102 273592 490158 273601
rect 490102 273527 490158 273536
rect 489748 272870 490236 272898
rect 489748 272270 489776 272870
rect 490208 272270 490236 272870
rect 489736 272264 489788 272270
rect 490196 272264 490248 272270
rect 489736 272206 489788 272212
rect 490010 272232 490066 272241
rect 490196 272206 490248 272212
rect 490010 272167 490066 272176
rect 490024 272066 490052 272167
rect 490012 272060 490064 272066
rect 490012 272002 490064 272008
rect 489874 271992 489926 271998
rect 489642 271960 489698 271969
rect 489926 271940 490052 271946
rect 489874 271934 490052 271940
rect 489886 271918 490052 271934
rect 489642 271895 489698 271904
rect 489656 271590 489684 271895
rect 490024 271833 490052 271918
rect 490010 271824 490066 271833
rect 490010 271759 490066 271768
rect 489644 271584 489696 271590
rect 489644 271526 489696 271532
rect 490102 271416 490158 271425
rect 490102 271351 490158 271360
rect 489920 271176 489972 271182
rect 489642 271144 489698 271153
rect 489698 271124 489920 271130
rect 489698 271118 489972 271124
rect 489698 271102 489960 271118
rect 489642 271079 489698 271088
rect 490116 270638 490144 271351
rect 490286 271144 490342 271153
rect 490286 271079 490342 271088
rect 489920 270632 489972 270638
rect 489920 270574 489972 270580
rect 490104 270632 490156 270638
rect 490104 270574 490156 270580
rect 489932 270450 489960 270574
rect 490300 270450 490328 271079
rect 489932 270422 490328 270450
rect 489734 269920 489790 269929
rect 489734 269855 489790 269864
rect 489748 269634 489776 269855
rect 489748 269606 489960 269634
rect 489932 269550 489960 269606
rect 489736 269544 489788 269550
rect 489736 269486 489788 269492
rect 489920 269544 489972 269550
rect 489920 269486 489972 269492
rect 489748 269249 489776 269486
rect 489734 269240 489790 269249
rect 489734 269175 489790 269184
rect 490484 267734 490512 274479
rect 490654 273048 490710 273057
rect 490654 272983 490710 272992
rect 491206 273048 491262 273057
rect 491206 272983 491262 272992
rect 490668 272406 490696 272983
rect 490656 272400 490708 272406
rect 490656 272342 490708 272348
rect 489932 267730 490512 267734
rect 489886 267706 490512 267730
rect 489886 267702 489960 267706
rect 489734 267608 489790 267617
rect 489886 267594 489914 267702
rect 489790 267566 489914 267594
rect 490470 267608 490526 267617
rect 489734 267543 489790 267552
rect 490470 267543 490472 267552
rect 490524 267543 490526 267552
rect 490656 267572 490708 267578
rect 490472 267514 490524 267520
rect 490656 267514 490708 267520
rect 489736 267436 489788 267442
rect 489736 267378 489788 267384
rect 490196 267436 490248 267442
rect 490196 267378 490248 267384
rect 489748 266529 489776 267378
rect 489920 267164 489972 267170
rect 489920 267106 489972 267112
rect 489734 266520 489790 266529
rect 489734 266455 489790 266464
rect 488368 264302 488474 264330
rect 489210 264302 489500 264330
rect 489932 264316 489960 267106
rect 490208 266801 490236 267378
rect 490194 266792 490250 266801
rect 490194 266727 490250 266736
rect 490470 266792 490526 266801
rect 490470 266727 490526 266736
rect 490104 266620 490156 266626
rect 490104 266562 490156 266568
rect 490116 266506 490144 266562
rect 490484 266506 490512 266727
rect 490116 266478 490512 266506
rect 490668 264316 490696 267514
rect 491220 267170 491248 272983
rect 491390 267608 491446 267617
rect 491390 267543 491446 267552
rect 491404 267170 491432 267543
rect 491208 267164 491260 267170
rect 491208 267106 491260 267112
rect 491392 267164 491444 267170
rect 491392 267106 491444 267112
rect 491864 264330 491892 276111
rect 493060 271153 493088 277766
rect 493324 276548 493376 276554
rect 493324 276490 493376 276496
rect 493046 271144 493102 271153
rect 493046 271079 493102 271088
rect 492126 267608 492182 267617
rect 492126 267543 492182 267552
rect 491418 264302 491892 264330
rect 492140 264316 492168 267543
rect 493336 266626 493364 276490
rect 494532 275194 494560 277766
rect 494980 276004 495032 276010
rect 494980 275946 495032 275952
rect 495348 276004 495400 276010
rect 495348 275946 495400 275952
rect 494992 275602 495020 275946
rect 494980 275596 495032 275602
rect 494980 275538 495032 275544
rect 494980 275460 495032 275466
rect 494980 275402 495032 275408
rect 494520 275188 494572 275194
rect 494520 275130 494572 275136
rect 494992 274961 495020 275402
rect 494978 274952 495034 274961
rect 494978 274887 495034 274896
rect 494888 274508 494940 274514
rect 494888 274450 494940 274456
rect 495072 274508 495124 274514
rect 495072 274450 495124 274456
rect 494900 274106 494928 274450
rect 494888 274100 494940 274106
rect 494888 274042 494940 274048
rect 495084 273986 495112 274450
rect 494520 273964 494572 273970
rect 494520 273906 494572 273912
rect 494716 273958 495112 273986
rect 494532 273562 494560 273906
rect 494336 273556 494388 273562
rect 494336 273498 494388 273504
rect 494520 273556 494572 273562
rect 494520 273498 494572 273504
rect 494348 273442 494376 273498
rect 494716 273442 494744 273958
rect 494348 273414 494744 273442
rect 495070 270600 495126 270609
rect 493980 270558 495070 270586
rect 493690 270056 493746 270065
rect 493690 269991 493746 270000
rect 493324 266620 493376 266626
rect 493324 266562 493376 266568
rect 493704 266490 493732 269991
rect 492864 266484 492916 266490
rect 492864 266426 492916 266432
rect 493692 266484 493744 266490
rect 493692 266426 493744 266432
rect 492876 264316 492904 266426
rect 493980 264330 494008 270558
rect 495070 270535 495126 270544
rect 494520 269952 494572 269958
rect 494572 269900 494928 269906
rect 494520 269894 494928 269900
rect 494532 269878 494928 269894
rect 494900 269822 494928 269878
rect 494888 269816 494940 269822
rect 494888 269758 494940 269764
rect 494150 267880 494206 267889
rect 494150 267815 494206 267824
rect 494164 267578 494192 267815
rect 494152 267572 494204 267578
rect 494152 267514 494204 267520
rect 494520 267572 494572 267578
rect 494520 267514 494572 267520
rect 494532 266529 494560 267514
rect 494704 267164 494756 267170
rect 494704 267106 494756 267112
rect 494888 267164 494940 267170
rect 494888 267106 494940 267112
rect 494716 266626 494744 267106
rect 494900 266801 494928 267106
rect 494886 266792 494942 266801
rect 494886 266727 494942 266736
rect 494704 266620 494756 266626
rect 494704 266562 494756 266568
rect 494518 266520 494574 266529
rect 494336 266484 494388 266490
rect 495360 266490 495388 275946
rect 495820 267734 495848 277766
rect 497016 274514 497044 277766
rect 497462 276448 497518 276457
rect 497462 276383 497518 276392
rect 497186 274544 497242 274553
rect 497004 274508 497056 274514
rect 497186 274479 497188 274488
rect 497004 274450 497056 274456
rect 497240 274479 497242 274488
rect 497188 274450 497240 274456
rect 496726 271144 496782 271153
rect 496726 271079 496782 271088
rect 495636 267706 495848 267734
rect 494518 266455 494574 266464
rect 495348 266484 495400 266490
rect 494336 266426 494388 266432
rect 495348 266426 495400 266432
rect 493626 264302 494008 264330
rect 494348 264316 494376 266426
rect 495636 265674 495664 267706
rect 496542 266792 496598 266801
rect 496542 266727 496598 266736
rect 495808 266484 495860 266490
rect 495808 266426 495860 266432
rect 495624 265668 495676 265674
rect 495624 265610 495676 265616
rect 495438 264344 495494 264353
rect 495098 264302 495438 264330
rect 495820 264316 495848 266426
rect 496556 264316 496584 266727
rect 496740 266490 496768 271079
rect 497476 267073 497504 276383
rect 498580 275466 498608 277780
rect 500052 277766 500894 277794
rect 501800 277766 502090 277794
rect 502352 277766 503286 277794
rect 499578 277400 499634 277409
rect 499578 277335 499634 277344
rect 499592 277114 499620 277335
rect 499500 277098 499620 277114
rect 499488 277092 499620 277098
rect 499540 277086 499620 277092
rect 499764 277092 499816 277098
rect 499488 277034 499540 277040
rect 499764 277034 499816 277040
rect 499224 276678 499574 276706
rect 499224 276185 499252 276678
rect 499546 276554 499574 276678
rect 499396 276548 499448 276554
rect 499396 276490 499448 276496
rect 499534 276548 499586 276554
rect 499534 276490 499586 276496
rect 499210 276176 499266 276185
rect 499210 276111 499266 276120
rect 499408 276049 499436 276490
rect 499776 276049 499804 277034
rect 499394 276040 499450 276049
rect 499394 275975 499450 275984
rect 499762 276040 499818 276049
rect 499762 275975 499818 275984
rect 498568 275460 498620 275466
rect 498568 275402 498620 275408
rect 498752 275460 498804 275466
rect 498752 275402 498804 275408
rect 497646 273592 497702 273601
rect 497646 273527 497702 273536
rect 497660 267170 497688 273527
rect 498764 272354 498792 275402
rect 499210 272776 499266 272785
rect 499266 272734 499436 272762
rect 499210 272711 499266 272720
rect 499408 272406 499436 272734
rect 498672 272326 498792 272354
rect 499028 272400 499080 272406
rect 499028 272342 499080 272348
rect 499396 272400 499448 272406
rect 499396 272342 499448 272348
rect 497648 267164 497700 267170
rect 497648 267106 497700 267112
rect 497462 267064 497518 267073
rect 497462 266999 497518 267008
rect 498014 266520 498070 266529
rect 496728 266484 496780 266490
rect 498672 266490 498700 272326
rect 498842 272232 498898 272241
rect 498842 272167 498898 272176
rect 498856 272066 498884 272167
rect 499040 272134 499068 272342
rect 499854 272232 499910 272241
rect 499684 272190 499854 272218
rect 499684 272134 499712 272190
rect 499854 272167 499910 272176
rect 499028 272128 499080 272134
rect 499028 272070 499080 272076
rect 499672 272128 499724 272134
rect 499672 272070 499724 272076
rect 498844 272060 498896 272066
rect 498844 272002 498896 272008
rect 499534 271992 499586 271998
rect 499408 271940 499534 271946
rect 499408 271934 499586 271940
rect 499408 271918 499574 271934
rect 499408 271833 499436 271918
rect 499394 271824 499450 271833
rect 499394 271759 499450 271768
rect 499762 271688 499818 271697
rect 499592 271646 499762 271674
rect 499592 270722 499620 271646
rect 499762 271623 499818 271632
rect 499500 270694 499620 270722
rect 499500 270638 499528 270694
rect 499488 270632 499540 270638
rect 499672 270632 499724 270638
rect 499488 270574 499540 270580
rect 499670 270600 499672 270609
rect 499724 270600 499726 270609
rect 499670 270535 499726 270544
rect 499396 270088 499448 270094
rect 499394 270056 499396 270065
rect 499534 270088 499586 270094
rect 499448 270056 499450 270065
rect 500052 270065 500080 277766
rect 501800 275874 501828 277766
rect 502352 277409 502380 277766
rect 502338 277400 502394 277409
rect 504468 277394 504496 277780
rect 505296 277766 505678 277794
rect 506492 277766 506874 277794
rect 504468 277366 504588 277394
rect 502338 277335 502394 277344
rect 504364 276004 504416 276010
rect 504364 275946 504416 275952
rect 501788 275868 501840 275874
rect 501788 275810 501840 275816
rect 501972 275868 502024 275874
rect 501972 275810 502024 275816
rect 501142 275768 501198 275777
rect 501142 275703 501198 275712
rect 500224 272128 500276 272134
rect 500224 272070 500276 272076
rect 500236 271969 500264 272070
rect 500222 271960 500278 271969
rect 500222 271895 500278 271904
rect 499534 270030 499586 270036
rect 500038 270056 500094 270065
rect 499394 269991 499450 270000
rect 499546 269906 499574 270030
rect 500038 269991 500094 270000
rect 499316 269878 499574 269906
rect 499316 269822 499344 269878
rect 499304 269816 499356 269822
rect 499304 269758 499356 269764
rect 499580 269816 499632 269822
rect 499580 269758 499632 269764
rect 499210 269240 499266 269249
rect 499210 269175 499266 269184
rect 499224 269090 499252 269175
rect 499592 269090 499620 269758
rect 499762 269240 499818 269249
rect 499762 269175 499818 269184
rect 499224 269062 499620 269090
rect 499210 268968 499266 268977
rect 499210 268903 499266 268912
rect 499394 268968 499450 268977
rect 499394 268903 499450 268912
rect 499224 268546 499252 268903
rect 499408 268666 499436 268903
rect 499396 268660 499448 268666
rect 499396 268602 499448 268608
rect 499534 268660 499586 268666
rect 499534 268602 499586 268608
rect 499546 268546 499574 268602
rect 499224 268518 499574 268546
rect 499534 267164 499586 267170
rect 499534 267106 499586 267112
rect 499026 267064 499082 267073
rect 499546 267050 499574 267106
rect 499026 266999 499082 267008
rect 499224 267022 499574 267050
rect 498014 266455 498070 266464
rect 498660 266484 498712 266490
rect 496728 266426 496780 266432
rect 497280 265668 497332 265674
rect 497280 265610 497332 265616
rect 497292 264316 497320 265610
rect 498028 264316 498056 266455
rect 498660 266426 498712 266432
rect 499040 264330 499068 266999
rect 499224 266801 499252 267022
rect 499210 266792 499266 266801
rect 499210 266727 499266 266736
rect 499394 266520 499450 266529
rect 499212 266484 499264 266490
rect 499394 266455 499396 266464
rect 499212 266426 499264 266432
rect 499448 266455 499450 266464
rect 499396 266426 499448 266432
rect 498778 264302 499068 264330
rect 499224 264330 499252 266426
rect 499776 264353 499804 269175
rect 501156 268977 501184 275703
rect 501984 275448 502012 275810
rect 504376 275466 504404 275946
rect 501800 275420 502012 275448
rect 504364 275460 504416 275466
rect 501800 275058 501828 275420
rect 504364 275402 504416 275408
rect 501972 275324 502024 275330
rect 501972 275266 502024 275272
rect 501984 275058 502012 275266
rect 501788 275052 501840 275058
rect 501788 274994 501840 275000
rect 501972 275052 502024 275058
rect 501972 274994 502024 275000
rect 503626 274680 503682 274689
rect 503626 274615 503682 274624
rect 503640 269521 503668 274615
rect 504560 270881 504588 277366
rect 504732 276004 504784 276010
rect 504732 275946 504784 275952
rect 504744 275777 504772 275946
rect 504730 275768 504786 275777
rect 504730 275703 504786 275712
rect 505296 273601 505324 277766
rect 505282 273592 505338 273601
rect 505282 273527 505338 273536
rect 504546 270872 504602 270881
rect 504546 270807 504602 270816
rect 503626 269512 503682 269521
rect 503626 269447 503682 269456
rect 501142 268968 501198 268977
rect 501142 268903 501198 268912
rect 506492 267850 506520 277766
rect 507964 277394 507992 277780
rect 507872 277366 507992 277394
rect 508700 277766 509174 277794
rect 510080 277766 510370 277794
rect 510632 277766 511566 277794
rect 512012 277766 512762 277794
rect 507872 272241 507900 277366
rect 508700 275874 508728 277766
rect 510080 277710 510108 277766
rect 510068 277704 510120 277710
rect 510068 277646 510120 277652
rect 508884 277222 509280 277250
rect 508884 276457 508912 277222
rect 509252 277098 509280 277222
rect 509056 277092 509108 277098
rect 509056 277034 509108 277040
rect 509240 277092 509292 277098
rect 509240 277034 509292 277040
rect 508870 276448 508926 276457
rect 508870 276383 508926 276392
rect 509068 276010 509096 277034
rect 509056 276004 509108 276010
rect 509056 275946 509108 275952
rect 508688 275868 508740 275874
rect 508688 275810 508740 275816
rect 509238 275768 509294 275777
rect 509238 275703 509294 275712
rect 509252 275074 509280 275703
rect 509206 275046 509280 275074
rect 509206 274922 509234 275046
rect 509194 274916 509246 274922
rect 509194 274858 509246 274864
rect 509332 274916 509384 274922
rect 509332 274858 509384 274864
rect 509344 274689 509372 274858
rect 509330 274680 509386 274689
rect 509330 274615 509386 274624
rect 507858 272232 507914 272241
rect 507858 272167 507914 272176
rect 509422 271688 509478 271697
rect 509422 271623 509478 271632
rect 509436 270910 509464 271623
rect 509194 270904 509246 270910
rect 509424 270904 509476 270910
rect 509246 270852 509280 270858
rect 509194 270846 509280 270852
rect 509424 270846 509476 270852
rect 509206 270830 509280 270846
rect 509252 270745 509280 270830
rect 509238 270736 509294 270745
rect 509238 270671 509294 270680
rect 508884 269742 509280 269770
rect 508884 267889 508912 269742
rect 509252 269686 509280 269742
rect 509056 269680 509108 269686
rect 509056 269622 509108 269628
rect 509240 269680 509292 269686
rect 509240 269622 509292 269628
rect 509068 269249 509096 269622
rect 510632 269249 510660 277766
rect 512012 276010 512040 277766
rect 512000 276004 512052 276010
rect 512000 275946 512052 275952
rect 512184 276004 512236 276010
rect 512184 275946 512236 275952
rect 512196 275777 512224 275946
rect 512182 275768 512238 275777
rect 512182 275703 512238 275712
rect 513944 274922 513972 277780
rect 513932 274916 513984 274922
rect 513932 274858 513984 274864
rect 514116 274916 514168 274922
rect 514116 274858 514168 274864
rect 514128 272785 514156 274858
rect 515140 273426 515168 277780
rect 516244 276010 516272 277780
rect 516428 277766 517454 277794
rect 518360 277766 518650 277794
rect 518912 277766 519846 277794
rect 516232 276004 516284 276010
rect 516232 275946 516284 275952
rect 515128 273420 515180 273426
rect 515128 273362 515180 273368
rect 514114 272776 514170 272785
rect 514114 272711 514170 272720
rect 509054 269240 509110 269249
rect 509054 269175 509110 269184
rect 510618 269240 510674 269249
rect 510618 269175 510674 269184
rect 508870 267880 508926 267889
rect 506480 267844 506532 267850
rect 508870 267815 508926 267824
rect 506480 267786 506532 267792
rect 514024 266892 514076 266898
rect 514024 266834 514076 266840
rect 514208 266892 514260 266898
rect 514208 266834 514260 266840
rect 514036 266626 514064 266834
rect 513840 266620 513892 266626
rect 513840 266562 513892 266568
rect 514024 266620 514076 266626
rect 514024 266562 514076 266568
rect 513852 266506 513880 266562
rect 514220 266506 514248 266834
rect 513852 266478 514248 266506
rect 516428 265266 516456 277766
rect 518360 270745 518388 277766
rect 518346 270736 518402 270745
rect 518346 270671 518402 270680
rect 518912 266626 518940 277766
rect 521028 276418 521056 277780
rect 521672 277766 522238 277794
rect 521016 276412 521068 276418
rect 521016 276354 521068 276360
rect 521672 269278 521700 277766
rect 523420 277394 523448 277780
rect 524524 277574 524552 277780
rect 524708 277766 525734 277794
rect 525904 277766 526930 277794
rect 527784 277788 528126 277794
rect 527732 277782 528126 277788
rect 527744 277766 528126 277782
rect 524512 277568 524564 277574
rect 524512 277510 524564 277516
rect 523328 277366 523448 277394
rect 523328 274786 523356 277366
rect 523684 276004 523736 276010
rect 523684 275946 523736 275952
rect 523500 275188 523552 275194
rect 523500 275130 523552 275136
rect 523512 274786 523540 275130
rect 523316 274780 523368 274786
rect 523316 274722 523368 274728
rect 523500 274780 523552 274786
rect 523500 274722 523552 274728
rect 521660 269272 521712 269278
rect 521660 269214 521712 269220
rect 518900 266620 518952 266626
rect 518900 266562 518952 266568
rect 516416 265260 516468 265266
rect 516416 265202 516468 265208
rect 523696 264994 523724 275946
rect 524708 267986 524736 277766
rect 524696 267980 524748 267986
rect 524696 267922 524748 267928
rect 525904 266898 525932 277766
rect 529308 273562 529336 277780
rect 530504 274786 530532 277780
rect 531228 276140 531280 276146
rect 531228 276082 531280 276088
rect 531240 274922 531268 276082
rect 531228 274916 531280 274922
rect 531228 274858 531280 274864
rect 530492 274780 530544 274786
rect 530492 274722 530544 274728
rect 529296 273556 529348 273562
rect 529296 273498 529348 273504
rect 531608 271862 531636 277780
rect 532804 271998 532832 277780
rect 532988 277766 534014 277794
rect 532792 271992 532844 271998
rect 532792 271934 532844 271940
rect 531596 271856 531648 271862
rect 531596 271798 531648 271804
rect 532988 267345 533016 277766
rect 533344 276004 533396 276010
rect 533344 275946 533396 275952
rect 533356 274786 533384 275946
rect 533344 274780 533396 274786
rect 533344 274722 533396 274728
rect 533528 271720 533580 271726
rect 533528 271662 533580 271668
rect 533540 270910 533568 271662
rect 533528 270904 533580 270910
rect 533528 270846 533580 270852
rect 535196 270774 535224 277780
rect 535472 277766 536406 277794
rect 535184 270768 535236 270774
rect 535184 270710 535236 270716
rect 535472 269414 535500 277766
rect 537588 275194 537616 277780
rect 537576 275188 537628 275194
rect 537576 275130 537628 275136
rect 537760 275188 537812 275194
rect 537760 275130 537812 275136
rect 535460 269408 535512 269414
rect 535460 269350 535512 269356
rect 532974 267336 533030 267345
rect 532974 267271 533030 267280
rect 525892 266892 525944 266898
rect 525892 266834 525944 266840
rect 537772 265130 537800 275130
rect 538784 271862 538812 277780
rect 538772 271856 538824 271862
rect 538772 271798 538824 271804
rect 539888 271046 539916 277780
rect 541084 275505 541112 277780
rect 541268 277766 542294 277794
rect 541070 275496 541126 275505
rect 541070 275431 541126 275440
rect 539876 271040 539928 271046
rect 539876 270982 539928 270988
rect 538864 270904 538916 270910
rect 538864 270846 538916 270852
rect 538876 267714 538904 270846
rect 541268 268122 541296 277766
rect 543476 274145 543504 277780
rect 543752 277766 544686 277794
rect 545132 277766 545882 277794
rect 547892 277766 548182 277794
rect 543462 274136 543518 274145
rect 543462 274071 543518 274080
rect 541256 268116 541308 268122
rect 541256 268058 541308 268064
rect 538864 267708 538916 267714
rect 538864 267650 538916 267656
rect 543752 267306 543780 277766
rect 543740 267300 543792 267306
rect 543740 267242 543792 267248
rect 537760 265124 537812 265130
rect 537760 265066 537812 265072
rect 523684 264988 523736 264994
rect 523684 264930 523736 264936
rect 545132 264790 545160 277766
rect 547892 268258 547920 277766
rect 549364 274786 549392 277780
rect 549548 277766 550574 277794
rect 549352 274780 549404 274786
rect 549352 274722 549404 274728
rect 549548 270502 549576 277766
rect 551560 272400 551612 272406
rect 551560 272342 551612 272348
rect 551572 271998 551600 272342
rect 551560 271992 551612 271998
rect 551560 271934 551612 271940
rect 551756 271726 551784 277780
rect 552952 275194 552980 277780
rect 553872 277766 554162 277794
rect 552940 275188 552992 275194
rect 552940 275130 552992 275136
rect 552848 274780 552900 274786
rect 552848 274722 552900 274728
rect 552664 272400 552716 272406
rect 552664 272342 552716 272348
rect 552676 272134 552704 272342
rect 552664 272128 552716 272134
rect 552664 272070 552716 272076
rect 551744 271720 551796 271726
rect 551744 271662 551796 271668
rect 549536 270496 549588 270502
rect 549536 270438 549588 270444
rect 547880 268252 547932 268258
rect 547880 268194 547932 268200
rect 552860 265402 552888 274722
rect 553872 271454 553900 277766
rect 555252 271998 555280 277780
rect 556160 275188 556212 275194
rect 556160 275130 556212 275136
rect 556172 273698 556200 275130
rect 556448 274786 556476 277780
rect 557644 276282 557672 277780
rect 557920 277766 558854 277794
rect 559300 277766 560050 277794
rect 557632 276276 557684 276282
rect 557632 276218 557684 276224
rect 556436 274780 556488 274786
rect 556436 274722 556488 274728
rect 556160 273692 556212 273698
rect 556160 273634 556212 273640
rect 555240 271992 555292 271998
rect 555240 271934 555292 271940
rect 554044 271720 554096 271726
rect 554044 271662 554096 271668
rect 553860 271448 553912 271454
rect 553860 271390 553912 271396
rect 554056 267034 554084 271662
rect 557920 270337 557948 277766
rect 557906 270328 557962 270337
rect 557906 270263 557962 270272
rect 554044 267028 554096 267034
rect 554044 266970 554096 266976
rect 559300 265538 559328 277766
rect 561232 272270 561260 277780
rect 561220 272264 561272 272270
rect 561220 272206 561272 272212
rect 562428 271590 562456 277780
rect 563532 277234 563560 277780
rect 563520 277228 563572 277234
rect 563520 277170 563572 277176
rect 564728 272814 564756 277780
rect 565924 275194 565952 277780
rect 566108 277766 567134 277794
rect 565912 275188 565964 275194
rect 565912 275130 565964 275136
rect 564716 272808 564768 272814
rect 564716 272750 564768 272756
rect 562416 271584 562468 271590
rect 562416 271526 562468 271532
rect 566108 266354 566136 277766
rect 568316 273222 568344 277780
rect 569512 273834 569540 277780
rect 570708 274922 570736 277780
rect 570972 277432 571024 277438
rect 570972 277374 571024 277380
rect 570984 275194 571012 277374
rect 570972 275188 571024 275194
rect 570972 275130 571024 275136
rect 570696 274916 570748 274922
rect 570696 274858 570748 274864
rect 569500 273828 569552 273834
rect 569500 273770 569552 273776
rect 568304 273216 568356 273222
rect 568304 273158 568356 273164
rect 571812 273086 571840 277780
rect 572732 277766 573022 277794
rect 571800 273080 571852 273086
rect 571800 273022 571852 273028
rect 571984 273080 572036 273086
rect 571984 273022 572036 273028
rect 571996 266762 572024 273022
rect 572732 269074 572760 277766
rect 574204 275874 574232 277780
rect 574192 275868 574244 275874
rect 574192 275810 574244 275816
rect 575400 272950 575428 277780
rect 575676 277766 576610 277794
rect 576872 277766 577806 277794
rect 578528 277766 578910 277794
rect 575388 272944 575440 272950
rect 575388 272886 575440 272892
rect 572720 269068 572772 269074
rect 572720 269010 572772 269016
rect 571984 266756 572036 266762
rect 571984 266698 572036 266704
rect 566096 266348 566148 266354
rect 566096 266290 566148 266296
rect 575676 266218 575704 277766
rect 576872 268938 576900 277766
rect 578528 272678 578556 277766
rect 578884 272808 578936 272814
rect 578884 272750 578936 272756
rect 578516 272672 578568 272678
rect 578516 272614 578568 272620
rect 576860 268932 576912 268938
rect 576860 268874 576912 268880
rect 578896 267617 578924 272750
rect 580092 271318 580120 277780
rect 581012 277766 581302 277794
rect 580080 271312 580132 271318
rect 580080 271254 580132 271260
rect 581012 268666 581040 277766
rect 582484 272542 582512 277780
rect 582760 277766 583694 277794
rect 583864 277766 584890 277794
rect 582472 272536 582524 272542
rect 582472 272478 582524 272484
rect 582760 270230 582788 277766
rect 582748 270224 582800 270230
rect 582748 270166 582800 270172
rect 583864 268802 583892 277766
rect 585784 272536 585836 272542
rect 585784 272478 585836 272484
rect 583852 268796 583904 268802
rect 583852 268738 583904 268744
rect 581000 268660 581052 268666
rect 581000 268602 581052 268608
rect 578882 267608 578938 267617
rect 585796 267578 585824 272478
rect 586072 272406 586100 277780
rect 586532 277766 587190 277794
rect 587912 277766 588386 277794
rect 589292 277766 589582 277794
rect 586060 272400 586112 272406
rect 586060 272342 586112 272348
rect 578882 267543 578938 267552
rect 585784 267572 585836 267578
rect 585784 267514 585836 267520
rect 575664 266212 575716 266218
rect 575664 266154 575716 266160
rect 559288 265532 559340 265538
rect 559288 265474 559340 265480
rect 552848 265396 552900 265402
rect 552848 265338 552900 265344
rect 545120 264784 545172 264790
rect 545120 264726 545172 264732
rect 586532 264654 586560 277766
rect 587912 268705 587940 277766
rect 587898 268696 587954 268705
rect 587898 268631 587954 268640
rect 589292 266121 589320 277766
rect 590764 277394 590792 277780
rect 590672 277366 590792 277394
rect 591040 277766 591974 277794
rect 590672 269550 590700 277366
rect 590660 269544 590712 269550
rect 590660 269486 590712 269492
rect 589278 266112 589334 266121
rect 591040 266082 591068 277766
rect 593156 272513 593184 277780
rect 593142 272504 593198 272513
rect 593142 272439 593198 272448
rect 594352 271182 594380 277780
rect 594812 277766 595470 277794
rect 596192 277766 596666 277794
rect 594340 271176 594392 271182
rect 594340 271118 594392 271124
rect 594812 268530 594840 277766
rect 596192 275346 596220 277766
rect 596100 275318 596220 275346
rect 596100 275194 596128 275318
rect 596088 275188 596140 275194
rect 596088 275130 596140 275136
rect 597468 275188 597520 275194
rect 597468 275130 597520 275136
rect 597480 274650 597508 275130
rect 597468 274644 597520 274650
rect 597468 274586 597520 274592
rect 597848 270910 597876 277780
rect 599044 276826 599072 277780
rect 599320 277766 600254 277794
rect 599032 276820 599084 276826
rect 599032 276762 599084 276768
rect 597836 270904 597888 270910
rect 597836 270846 597888 270852
rect 599320 270366 599348 277766
rect 601436 277098 601464 277780
rect 601804 277766 602554 277794
rect 603092 277766 603750 277794
rect 601424 277092 601476 277098
rect 601424 277034 601476 277040
rect 599308 270360 599360 270366
rect 599308 270302 599360 270308
rect 594800 268524 594852 268530
rect 594800 268466 594852 268472
rect 601608 268524 601660 268530
rect 601608 268466 601660 268472
rect 601620 266490 601648 268466
rect 601608 266484 601660 266490
rect 601608 266426 601660 266432
rect 589278 266047 589334 266056
rect 591028 266076 591080 266082
rect 591028 266018 591080 266024
rect 601804 265946 601832 277766
rect 601792 265940 601844 265946
rect 601792 265882 601844 265888
rect 586520 264648 586572 264654
rect 586520 264590 586572 264596
rect 603092 264518 603120 277766
rect 604932 275738 604960 277780
rect 606128 276962 606156 277780
rect 607324 277394 607352 277780
rect 607232 277366 607352 277394
rect 606116 276956 606168 276962
rect 606116 276898 606168 276904
rect 604920 275732 604972 275738
rect 604920 275674 604972 275680
rect 607232 268433 607260 277366
rect 608520 273086 608548 277780
rect 608888 277766 609730 277794
rect 608508 273080 608560 273086
rect 608508 273022 608560 273028
rect 607218 268424 607274 268433
rect 608888 268394 608916 277766
rect 610072 275732 610124 275738
rect 610072 275674 610124 275680
rect 610084 274378 610112 275674
rect 610820 275194 610848 277780
rect 612016 275602 612044 277780
rect 612752 277766 613226 277794
rect 612004 275596 612056 275602
rect 612004 275538 612056 275544
rect 610808 275188 610860 275194
rect 610808 275130 610860 275136
rect 610072 274372 610124 274378
rect 610072 274314 610124 274320
rect 607218 268359 607274 268368
rect 608876 268388 608928 268394
rect 608876 268330 608928 268336
rect 612752 265810 612780 277766
rect 614408 275738 614436 277780
rect 615604 277394 615632 277780
rect 616616 277766 616814 277794
rect 615604 277366 615724 277394
rect 614396 275732 614448 275738
rect 614396 275674 614448 275680
rect 614764 274712 614816 274718
rect 614764 274654 614816 274660
rect 614776 265849 614804 274654
rect 615696 271726 615724 277366
rect 616616 274718 616644 277766
rect 616788 276548 616840 276554
rect 616788 276490 616840 276496
rect 616800 276010 616828 276490
rect 616788 276004 616840 276010
rect 616788 275946 616840 275952
rect 616604 274712 616656 274718
rect 616604 274654 616656 274660
rect 617996 274514 618024 277780
rect 619100 275233 619128 277780
rect 619086 275224 619142 275233
rect 619086 275159 619142 275168
rect 619640 274848 619692 274854
rect 619640 274790 619692 274796
rect 618904 274712 618956 274718
rect 618904 274654 618956 274660
rect 617984 274508 618036 274514
rect 617984 274450 618036 274456
rect 615684 271720 615736 271726
rect 615684 271662 615736 271668
rect 614762 265840 614818 265849
rect 612740 265804 612792 265810
rect 614762 265775 614818 265784
rect 612740 265746 612792 265752
rect 603080 264512 603132 264518
rect 603080 264454 603132 264460
rect 618916 264382 618944 274654
rect 619652 269822 619680 274790
rect 620296 274718 620324 277780
rect 620284 274712 620336 274718
rect 620284 274654 620336 274660
rect 621492 274242 621520 277780
rect 621480 274236 621532 274242
rect 621480 274178 621532 274184
rect 622688 272542 622716 277780
rect 623884 274854 623912 277780
rect 623872 274848 623924 274854
rect 623872 274790 623924 274796
rect 625080 274106 625108 277780
rect 625068 274100 625120 274106
rect 625068 274042 625120 274048
rect 622676 272536 622728 272542
rect 622676 272478 622728 272484
rect 625804 271584 625856 271590
rect 625804 271526 625856 271532
rect 620284 270224 620336 270230
rect 620284 270166 620336 270172
rect 620296 269958 620324 270166
rect 620284 269952 620336 269958
rect 620284 269894 620336 269900
rect 619640 269816 619692 269822
rect 619640 269758 619692 269764
rect 625816 267442 625844 271526
rect 626184 271425 626212 277780
rect 626552 277766 627394 277794
rect 626170 271416 626226 271425
rect 626170 271351 626226 271360
rect 626552 270094 626580 277766
rect 628576 273970 628604 277780
rect 628564 273964 628616 273970
rect 628564 273906 628616 273912
rect 629772 271590 629800 277780
rect 630692 277766 630982 277794
rect 629760 271584 629812 271590
rect 629760 271526 629812 271532
rect 626540 270088 626592 270094
rect 626540 270030 626592 270036
rect 630692 269958 630720 277766
rect 632164 273873 632192 277780
rect 633360 275058 633388 277780
rect 633636 277766 634478 277794
rect 633348 275052 633400 275058
rect 633348 274994 633400 275000
rect 632704 273964 632756 273970
rect 632704 273906 632756 273912
rect 632150 273864 632206 273873
rect 632150 273799 632206 273808
rect 630680 269952 630732 269958
rect 630680 269894 630732 269900
rect 625804 267436 625856 267442
rect 625804 267378 625856 267384
rect 632716 267170 632744 273906
rect 633636 269686 633664 277766
rect 635660 276010 635688 277780
rect 635648 276004 635700 276010
rect 635648 275946 635700 275952
rect 636856 272814 636884 277780
rect 637592 277766 638066 277794
rect 636844 272808 636896 272814
rect 636844 272750 636896 272756
rect 637592 270065 637620 277766
rect 639248 270638 639276 277780
rect 640444 275466 640472 277780
rect 640720 277766 641654 277794
rect 640432 275460 640484 275466
rect 640432 275402 640484 275408
rect 639236 270632 639288 270638
rect 639236 270574 639288 270580
rect 637578 270056 637634 270065
rect 637578 269991 637634 270000
rect 636200 269816 636252 269822
rect 640720 269793 640748 277766
rect 636200 269758 636252 269764
rect 640706 269784 640762 269793
rect 633624 269680 633676 269686
rect 633624 269622 633676 269628
rect 632704 267164 632756 267170
rect 632704 267106 632756 267112
rect 636212 267073 636240 269758
rect 640706 269719 640762 269728
rect 636198 267064 636254 267073
rect 636198 266999 636254 267008
rect 618904 264376 618956 264382
rect 499762 264344 499818 264353
rect 499224 264302 499514 264330
rect 495438 264279 495494 264288
rect 618904 264318 618956 264324
rect 499762 264279 499818 264288
rect 436954 264166 437244 264194
rect 468602 264166 468984 264194
rect 511538 262712 511594 262721
rect 511538 262647 511594 262656
rect 511552 261526 511580 262647
rect 511540 261520 511592 261526
rect 511540 261462 511592 261468
rect 568580 261520 568632 261526
rect 568580 261462 568632 261468
rect 511354 260264 511410 260273
rect 511354 260199 511410 260208
rect 511368 260030 511396 260199
rect 511356 260024 511408 260030
rect 511356 259966 511408 259972
rect 514024 260024 514076 260030
rect 514024 259966 514076 259972
rect 511446 257816 511502 257825
rect 511446 257751 511502 257760
rect 511460 256766 511488 257751
rect 511448 256760 511500 256766
rect 511448 256702 511500 256708
rect 511170 255368 511226 255377
rect 511170 255303 511226 255312
rect 510618 250472 510674 250481
rect 510618 250407 510674 250416
rect 510632 249830 510660 250407
rect 510620 249824 510672 249830
rect 510620 249766 510672 249772
rect 511184 249082 511212 255303
rect 511906 252920 511962 252929
rect 511906 252855 511962 252864
rect 511920 252618 511948 252855
rect 511908 252612 511960 252618
rect 511908 252554 511960 252560
rect 513288 249824 513340 249830
rect 513288 249766 513340 249772
rect 511172 249076 511224 249082
rect 511172 249018 511224 249024
rect 511078 248024 511134 248033
rect 511078 247959 511134 247968
rect 128832 247302 129228 247330
rect 128832 247110 128860 247302
rect 129004 247240 129056 247246
rect 129004 247182 129056 247188
rect 128820 247104 128872 247110
rect 128820 247046 128872 247052
rect 116872 230846 117268 230874
rect 108948 230784 109000 230790
rect 108948 230726 109000 230732
rect 89628 230648 89680 230654
rect 89628 230590 89680 230596
rect 79968 230512 80020 230518
rect 79968 230454 80020 230460
rect 69664 229900 69716 229906
rect 69664 229842 69716 229848
rect 66904 229764 66956 229770
rect 66904 229706 66956 229712
rect 65984 227996 66036 228002
rect 65984 227938 66036 227944
rect 63592 227044 63644 227050
rect 63592 226986 63644 226992
rect 63408 220652 63460 220658
rect 63408 220594 63460 220600
rect 63420 217410 63448 220594
rect 63604 220250 63632 226986
rect 63960 220856 64012 220862
rect 63960 220798 64012 220804
rect 63592 220244 63644 220250
rect 63592 220186 63644 220192
rect 63972 217410 64000 220798
rect 64788 220108 64840 220114
rect 64788 220050 64840 220056
rect 64800 217410 64828 220050
rect 65996 217410 66024 227938
rect 66718 222048 66774 222057
rect 66718 221983 66774 221992
rect 66732 217410 66760 221983
rect 66916 220862 66944 229706
rect 68928 228404 68980 228410
rect 68928 228346 68980 228352
rect 68468 224256 68520 224262
rect 68468 224198 68520 224204
rect 66904 220856 66956 220862
rect 66904 220798 66956 220804
rect 67364 220788 67416 220794
rect 67364 220730 67416 220736
rect 67376 217410 67404 220730
rect 68480 217410 68508 224198
rect 68940 217410 68968 228346
rect 69676 220794 69704 229842
rect 75828 228540 75880 228546
rect 75828 228482 75880 228488
rect 72516 227180 72568 227186
rect 72516 227122 72568 227128
rect 71686 224224 71742 224233
rect 71686 224159 71742 224168
rect 70032 221468 70084 221474
rect 70032 221410 70084 221416
rect 69664 220788 69716 220794
rect 69664 220730 69716 220736
rect 70044 217410 70072 221410
rect 70860 219700 70912 219706
rect 70860 219642 70912 219648
rect 70872 217410 70900 219642
rect 71700 217410 71728 224159
rect 72528 217410 72556 227122
rect 75000 224528 75052 224534
rect 75000 224470 75052 224476
rect 74264 223168 74316 223174
rect 74264 223110 74316 223116
rect 72882 221232 72938 221241
rect 72882 221167 72938 221176
rect 63112 217382 63448 217410
rect 63940 217382 64000 217410
rect 64768 217382 64828 217410
rect 65596 217382 66024 217410
rect 66424 217382 66760 217410
rect 67252 217382 67404 217410
rect 68080 217382 68508 217410
rect 68908 217382 68968 217410
rect 69736 217382 70072 217410
rect 70564 217382 70900 217410
rect 71392 217382 71728 217410
rect 72220 217382 72556 217410
rect 72896 217410 72924 221167
rect 74276 217410 74304 223110
rect 75012 217410 75040 224470
rect 75840 217410 75868 228482
rect 78404 225752 78456 225758
rect 78404 225694 78456 225700
rect 77024 224800 77076 224806
rect 77024 224742 77076 224748
rect 76656 220516 76708 220522
rect 76656 220458 76708 220464
rect 76668 217410 76696 220458
rect 77036 220114 77064 224742
rect 77208 220244 77260 220250
rect 77208 220186 77260 220192
rect 77024 220108 77076 220114
rect 77024 220050 77076 220056
rect 77220 217410 77248 220186
rect 78416 217410 78444 225694
rect 79784 223032 79836 223038
rect 79784 222974 79836 222980
rect 79140 220788 79192 220794
rect 79140 220730 79192 220736
rect 79152 217410 79180 220730
rect 79796 217410 79824 222974
rect 79980 220794 80008 230454
rect 82912 230172 82964 230178
rect 82912 230114 82964 230120
rect 82544 227316 82596 227322
rect 82544 227258 82596 227264
rect 81348 225480 81400 225486
rect 81348 225422 81400 225428
rect 80796 221876 80848 221882
rect 80796 221818 80848 221824
rect 79968 220788 80020 220794
rect 79968 220730 80020 220736
rect 80152 220788 80204 220794
rect 80152 220730 80204 220736
rect 80164 220522 80192 220730
rect 80152 220516 80204 220522
rect 80152 220458 80204 220464
rect 80808 217410 80836 221818
rect 81360 217410 81388 225422
rect 82556 217410 82584 227258
rect 82924 223174 82952 230114
rect 88248 230036 88300 230042
rect 88248 229978 88300 229984
rect 84936 226160 84988 226166
rect 84936 226102 84988 226108
rect 82912 223168 82964 223174
rect 82912 223110 82964 223116
rect 83280 223168 83332 223174
rect 83280 223110 83332 223116
rect 83292 217410 83320 223110
rect 83924 219836 83976 219842
rect 83924 219778 83976 219784
rect 83936 217410 83964 219778
rect 84948 217410 84976 226102
rect 88064 225888 88116 225894
rect 88064 225830 88116 225836
rect 86684 223304 86736 223310
rect 86684 223246 86736 223252
rect 86696 217410 86724 223246
rect 87420 220516 87472 220522
rect 87420 220458 87472 220464
rect 87432 217410 87460 220458
rect 88076 217410 88104 225830
rect 88260 220522 88288 229978
rect 89640 220522 89668 230590
rect 107568 230308 107620 230314
rect 107568 230250 107620 230256
rect 99840 228948 99892 228954
rect 99840 228890 99892 228896
rect 96528 228812 96580 228818
rect 96528 228754 96580 228760
rect 93216 228676 93268 228682
rect 93216 228618 93268 228624
rect 92388 226024 92440 226030
rect 92388 225966 92440 225972
rect 91560 223440 91612 223446
rect 91560 223382 91612 223388
rect 88248 220516 88300 220522
rect 88248 220458 88300 220464
rect 89076 220516 89128 220522
rect 89076 220458 89128 220464
rect 89628 220516 89680 220522
rect 89628 220458 89680 220464
rect 88892 219836 88944 219842
rect 88892 219778 88944 219784
rect 88904 219570 88932 219778
rect 88892 219564 88944 219570
rect 88892 219506 88944 219512
rect 89088 217410 89116 220458
rect 89444 220380 89496 220386
rect 89444 220322 89496 220328
rect 72896 217382 73048 217410
rect 73876 217382 74304 217410
rect 74704 217382 75040 217410
rect 75532 217382 75868 217410
rect 76360 217382 76696 217410
rect 77188 217382 77248 217410
rect 78016 217382 78444 217410
rect 78844 217382 79180 217410
rect 79672 217382 79824 217410
rect 80500 217382 80836 217410
rect 81328 217382 81388 217410
rect 82156 217382 82584 217410
rect 82984 217382 83320 217410
rect 83812 217382 83964 217410
rect 84640 217382 84976 217410
rect 86296 217382 86724 217410
rect 87124 217382 87460 217410
rect 87952 217382 88104 217410
rect 88780 217382 89116 217410
rect 89456 217410 89484 220322
rect 91572 217410 91600 223382
rect 92400 217410 92428 225966
rect 93228 217410 93256 228618
rect 94964 223576 95016 223582
rect 94964 223518 95016 223524
rect 94976 217410 95004 223518
rect 95700 220516 95752 220522
rect 95700 220458 95752 220464
rect 95712 217410 95740 220458
rect 96540 217410 96568 228754
rect 97356 227452 97408 227458
rect 97356 227394 97408 227400
rect 97368 217410 97396 227394
rect 97908 226296 97960 226302
rect 97908 226238 97960 226244
rect 97724 221740 97776 221746
rect 97724 221682 97776 221688
rect 89456 217382 89608 217410
rect 91264 217382 91600 217410
rect 92092 217382 92428 217410
rect 92920 217382 93256 217410
rect 94576 217382 95004 217410
rect 95404 217382 95740 217410
rect 96232 217382 96568 217410
rect 97060 217382 97396 217410
rect 97736 217410 97764 221682
rect 97920 220522 97948 226238
rect 99104 224664 99156 224670
rect 99104 224606 99156 224612
rect 97908 220516 97960 220522
rect 97908 220458 97960 220464
rect 99116 217410 99144 224606
rect 99852 217410 99880 228890
rect 104808 225344 104860 225350
rect 104808 225286 104860 225292
rect 102140 222624 102192 222630
rect 102140 222566 102192 222572
rect 101496 222488 101548 222494
rect 101496 222430 101548 222436
rect 101508 217410 101536 222430
rect 102152 220794 102180 222566
rect 102140 220788 102192 220794
rect 102140 220730 102192 220736
rect 103980 220108 104032 220114
rect 103980 220050 104032 220056
rect 101864 219972 101916 219978
rect 101864 219914 101916 219920
rect 97736 217382 97888 217410
rect 98716 217382 99144 217410
rect 99544 217382 99880 217410
rect 101200 217382 101536 217410
rect 101876 217410 101904 219914
rect 103152 219836 103204 219842
rect 103152 219778 103204 219784
rect 103164 217410 103192 219778
rect 103992 217410 104020 220050
rect 104820 219978 104848 225286
rect 104808 219972 104860 219978
rect 104808 219914 104860 219920
rect 107580 219434 107608 230250
rect 108120 220788 108172 220794
rect 108120 220730 108172 220736
rect 107396 219406 107608 219434
rect 104808 219020 104860 219026
rect 104808 218962 104860 218968
rect 104820 217410 104848 218962
rect 106188 218884 106240 218890
rect 106188 218826 106240 218832
rect 105636 218748 105688 218754
rect 105636 218690 105688 218696
rect 105648 217410 105676 218690
rect 106200 217410 106228 218826
rect 107396 217410 107424 219406
rect 108132 217410 108160 220730
rect 108960 217410 108988 230726
rect 116872 230518 116900 230846
rect 117240 230790 117268 230846
rect 117044 230784 117096 230790
rect 117044 230726 117096 230732
rect 117228 230784 117280 230790
rect 117228 230726 117280 230732
rect 117056 230518 117084 230726
rect 116860 230512 116912 230518
rect 116860 230454 116912 230460
rect 117044 230512 117096 230518
rect 117044 230454 117096 230460
rect 117228 229628 117280 229634
rect 117228 229570 117280 229576
rect 111062 229528 111118 229537
rect 111062 229463 111118 229472
rect 109776 229084 109828 229090
rect 109776 229026 109828 229032
rect 109788 217410 109816 229026
rect 111076 221882 111104 229463
rect 115664 227452 115716 227458
rect 115664 227394 115716 227400
rect 114468 222760 114520 222766
rect 114468 222702 114520 222708
rect 111064 221876 111116 221882
rect 111064 221818 111116 221824
rect 111432 221876 111484 221882
rect 111432 221818 111484 221824
rect 111444 217410 111472 221818
rect 113916 219972 113968 219978
rect 113916 219914 113968 219920
rect 112904 219292 112956 219298
rect 112904 219234 112956 219240
rect 112260 219156 112312 219162
rect 112260 219098 112312 219104
rect 112272 217410 112300 219098
rect 112916 217410 112944 219234
rect 113928 217410 113956 219914
rect 114480 217410 114508 222702
rect 115676 217410 115704 227394
rect 116400 222012 116452 222018
rect 116400 221954 116452 221960
rect 116412 217410 116440 221954
rect 117240 217410 117268 229570
rect 126888 229492 126940 229498
rect 126888 229434 126940 229440
rect 118792 228268 118844 228274
rect 118792 228210 118844 228216
rect 118608 227724 118660 227730
rect 118608 227666 118660 227672
rect 118056 219428 118108 219434
rect 118056 219370 118108 219376
rect 118068 217410 118096 219370
rect 118620 217410 118648 227666
rect 118804 219842 118832 228210
rect 122196 226908 122248 226914
rect 122196 226850 122248 226856
rect 120080 225072 120132 225078
rect 120080 225014 120132 225020
rect 119712 222148 119764 222154
rect 119712 222090 119764 222096
rect 118792 219836 118844 219842
rect 118792 219778 118844 219784
rect 119724 217410 119752 222090
rect 120092 220658 120120 225014
rect 121368 224936 121420 224942
rect 121368 224878 121420 224884
rect 120080 220652 120132 220658
rect 120080 220594 120132 220600
rect 120540 220516 120592 220522
rect 120540 220458 120592 220464
rect 120552 217410 120580 220458
rect 121380 217410 121408 224878
rect 122208 217410 122236 226850
rect 124680 224120 124732 224126
rect 124680 224062 124732 224068
rect 122564 221332 122616 221338
rect 122564 221274 122616 221280
rect 101876 217382 102028 217410
rect 102856 217382 103192 217410
rect 103684 217382 104020 217410
rect 104512 217382 104848 217410
rect 105340 217382 105676 217410
rect 106168 217382 106228 217410
rect 106996 217382 107424 217410
rect 107824 217382 108160 217410
rect 108652 217382 108988 217410
rect 109480 217382 109816 217410
rect 111136 217382 111472 217410
rect 111964 217382 112300 217410
rect 112792 217382 112944 217410
rect 113620 217382 113956 217410
rect 114448 217382 114508 217410
rect 115276 217382 115704 217410
rect 116104 217382 116440 217410
rect 116932 217382 117268 217410
rect 117760 217382 118096 217410
rect 118588 217382 118648 217410
rect 119416 217382 119752 217410
rect 120244 217382 120580 217410
rect 121072 217382 121408 217410
rect 121900 217382 122236 217410
rect 122576 217410 122604 221274
rect 123852 220788 123904 220794
rect 123852 220730 123904 220736
rect 123864 217410 123892 220730
rect 124692 217410 124720 224062
rect 125324 222488 125376 222494
rect 125324 222430 125376 222436
rect 125336 217410 125364 222430
rect 126152 220924 126204 220930
rect 126152 220866 126204 220872
rect 126164 220658 126192 220866
rect 126152 220652 126204 220658
rect 126152 220594 126204 220600
rect 126336 220652 126388 220658
rect 126336 220594 126388 220600
rect 126348 217410 126376 220594
rect 126900 217410 126928 229434
rect 127072 227860 127124 227866
rect 127072 227802 127124 227808
rect 127084 220930 127112 227802
rect 127808 227724 127860 227730
rect 127808 227666 127860 227672
rect 127820 227610 127848 227666
rect 127268 227594 127848 227610
rect 127256 227588 127848 227594
rect 127308 227582 127848 227588
rect 127256 227530 127308 227536
rect 128820 226772 128872 226778
rect 128820 226714 128872 226720
rect 127072 220924 127124 220930
rect 127072 220866 127124 220872
rect 127808 220788 127860 220794
rect 127808 220730 127860 220736
rect 127992 220788 128044 220794
rect 127992 220730 128044 220736
rect 127820 220522 127848 220730
rect 127624 220516 127676 220522
rect 127624 220458 127676 220464
rect 127808 220516 127860 220522
rect 127808 220458 127860 220464
rect 127636 219978 127664 220458
rect 127624 219972 127676 219978
rect 127624 219914 127676 219920
rect 128004 217410 128032 220730
rect 128832 217410 128860 226714
rect 129016 225593 129044 247182
rect 129200 230897 129228 247302
rect 130382 245712 130438 245721
rect 130382 245647 130438 245656
rect 129186 230888 129242 230897
rect 129186 230823 129242 230832
rect 130396 225865 130424 245647
rect 510710 240680 510766 240689
rect 510710 240615 510766 240624
rect 507490 237960 507546 237969
rect 507490 237895 507546 237904
rect 132590 230888 132646 230897
rect 132590 230823 132592 230832
rect 132644 230823 132646 230832
rect 144642 230888 144698 230897
rect 144642 230823 144698 230832
rect 132592 230794 132644 230800
rect 132408 230784 132460 230790
rect 132460 230732 132540 230738
rect 132408 230726 132540 230732
rect 132420 230710 132540 230726
rect 132512 230625 132540 230710
rect 132498 230616 132554 230625
rect 132498 230551 132554 230560
rect 144656 229770 144684 230823
rect 145838 230344 145894 230353
rect 145838 230279 145894 230288
rect 146022 230344 146078 230353
rect 146022 230279 146078 230288
rect 144644 229764 144696 229770
rect 144644 229706 144696 229712
rect 144828 229764 144880 229770
rect 144828 229706 144880 229712
rect 133788 229356 133840 229362
rect 133788 229298 133840 229304
rect 132224 226636 132276 226642
rect 132224 226578 132276 226584
rect 130382 225856 130438 225865
rect 130382 225791 130438 225800
rect 129002 225584 129058 225593
rect 129002 225519 129058 225528
rect 131028 223984 131080 223990
rect 131028 223926 131080 223932
rect 129464 221196 129516 221202
rect 129464 221138 129516 221144
rect 129476 217410 129504 221138
rect 130198 220416 130254 220425
rect 130198 220351 130254 220360
rect 130212 217410 130240 220351
rect 131040 217410 131068 223926
rect 132236 217410 132264 226578
rect 132960 218612 133012 218618
rect 132960 218554 133012 218560
rect 132972 217410 133000 218554
rect 133800 217410 133828 229298
rect 140688 229220 140740 229226
rect 140688 229162 140740 229168
rect 137100 227724 137152 227730
rect 137100 227666 137152 227672
rect 137284 227724 137336 227730
rect 137284 227666 137336 227672
rect 137112 226658 137140 227666
rect 137296 226778 137324 227666
rect 137284 226772 137336 226778
rect 137284 226714 137336 226720
rect 137468 226772 137520 226778
rect 137468 226714 137520 226720
rect 137480 226658 137508 226714
rect 137112 226630 137508 226658
rect 138756 226432 138808 226438
rect 138756 226374 138808 226380
rect 134984 225208 135036 225214
rect 134984 225150 135036 225156
rect 134708 223848 134760 223854
rect 134708 223790 134760 223796
rect 134720 217410 134748 223790
rect 122576 217382 122728 217410
rect 123556 217382 123892 217410
rect 124384 217382 124720 217410
rect 125212 217382 125364 217410
rect 126040 217382 126376 217410
rect 126868 217382 126928 217410
rect 127696 217382 128032 217410
rect 128524 217382 128860 217410
rect 129352 217382 129504 217410
rect 130180 217382 130240 217410
rect 131008 217382 131068 217410
rect 131836 217382 132264 217410
rect 132664 217382 133000 217410
rect 133492 217382 133828 217410
rect 134320 217382 134748 217410
rect 134996 217410 135024 225150
rect 136546 222864 136602 222873
rect 136546 222799 136602 222808
rect 136560 220794 136588 222799
rect 137928 220924 137980 220930
rect 137928 220866 137980 220872
rect 136548 220788 136600 220794
rect 136548 220730 136600 220736
rect 136916 220788 136968 220794
rect 136916 220730 136968 220736
rect 136928 219842 136956 220730
rect 136916 219836 136968 219842
rect 136916 219778 136968 219784
rect 137100 219836 137152 219842
rect 137100 219778 137152 219784
rect 136272 218476 136324 218482
rect 136272 218418 136324 218424
rect 136284 217410 136312 218418
rect 137112 217410 137140 219778
rect 137940 217410 137968 220866
rect 138768 217410 138796 226374
rect 139124 221060 139176 221066
rect 139124 221002 139176 221008
rect 134996 217382 135148 217410
rect 135976 217382 136312 217410
rect 136804 217382 137140 217410
rect 137632 217382 137968 217410
rect 138460 217382 138796 217410
rect 139136 217410 139164 221002
rect 140700 219434 140728 229162
rect 144840 229094 144868 229706
rect 145852 229265 145880 230279
rect 145838 229256 145894 229265
rect 145838 229191 145894 229200
rect 144380 229066 144868 229094
rect 142894 228032 142950 228041
rect 142894 227967 142950 227976
rect 142158 227760 142214 227769
rect 142158 227695 142214 227704
rect 142172 227202 142200 227695
rect 142126 227174 142200 227202
rect 142126 227050 142154 227174
rect 142114 227044 142166 227050
rect 142114 226986 142166 226992
rect 142252 227044 142304 227050
rect 142252 226986 142304 226992
rect 142264 226930 142292 226986
rect 142126 226902 142292 226930
rect 142126 226778 142154 226902
rect 142114 226772 142166 226778
rect 142114 226714 142166 226720
rect 142252 226772 142304 226778
rect 142252 226714 142304 226720
rect 142264 226658 142292 226714
rect 142172 226630 142292 226658
rect 142172 226506 142200 226630
rect 141884 226500 141936 226506
rect 141884 226442 141936 226448
rect 142160 226500 142212 226506
rect 142160 226442 142212 226448
rect 142342 226502 142398 226511
rect 141700 226432 141752 226438
rect 141698 226400 141700 226409
rect 141752 226400 141754 226409
rect 141698 226335 141754 226344
rect 141240 223712 141292 223718
rect 141240 223654 141292 223660
rect 140516 219406 140728 219434
rect 140516 217410 140544 219406
rect 141252 217410 141280 223654
rect 141896 219434 141924 226442
rect 142342 226437 142398 226446
rect 142158 223136 142214 223145
rect 142158 223071 142214 223080
rect 142172 222986 142200 223071
rect 142126 222958 142200 222986
rect 142126 222902 142154 222958
rect 142114 222896 142166 222902
rect 142114 222838 142166 222844
rect 142436 222896 142488 222902
rect 142436 222838 142488 222844
rect 142618 222864 142674 222873
rect 142448 222714 142476 222838
rect 142618 222799 142674 222808
rect 142172 222686 142476 222714
rect 142172 222442 142200 222686
rect 142126 222414 142200 222442
rect 142126 222358 142154 222414
rect 142632 222358 142660 222799
rect 142114 222352 142166 222358
rect 142114 222294 142166 222300
rect 142620 222352 142672 222358
rect 142620 222294 142672 222300
rect 142068 219836 142120 219842
rect 142068 219778 142120 219784
rect 142252 219836 142304 219842
rect 142252 219778 142304 219784
rect 142080 219609 142108 219778
rect 142264 219609 142292 219778
rect 142066 219600 142122 219609
rect 142066 219535 142122 219544
rect 142250 219600 142306 219609
rect 142250 219535 142306 219544
rect 141896 219406 142108 219434
rect 142080 217410 142108 219406
rect 142908 217410 142936 227967
rect 144380 221610 144408 229066
rect 146036 224398 146064 230279
rect 147034 224496 147090 224505
rect 147034 224431 147090 224440
rect 146024 224392 146076 224398
rect 146024 224334 146076 224340
rect 146208 224392 146260 224398
rect 146208 224334 146260 224340
rect 144368 221604 144420 221610
rect 144368 221546 144420 221552
rect 144552 221604 144604 221610
rect 144552 221546 144604 221552
rect 143078 219736 143134 219745
rect 143078 219671 143080 219680
rect 143132 219671 143134 219680
rect 143264 219700 143316 219706
rect 143080 219642 143132 219648
rect 143264 219642 143316 219648
rect 139136 217382 139288 217410
rect 140116 217382 140544 217410
rect 140944 217382 141280 217410
rect 141772 217382 142108 217410
rect 142600 217382 142936 217410
rect 143276 217410 143304 219642
rect 144564 217410 144592 221546
rect 146220 219434 146248 224334
rect 145392 219406 146248 219434
rect 145392 217410 145420 219406
rect 146208 218340 146260 218346
rect 146208 218282 146260 218288
rect 146220 217410 146248 218282
rect 147048 217410 147076 224431
rect 147678 220688 147734 220697
rect 147678 220623 147734 220632
rect 147692 220266 147720 220623
rect 147646 220238 147720 220266
rect 147646 220114 147674 220238
rect 147634 220108 147686 220114
rect 147634 220050 147686 220056
rect 147772 220108 147824 220114
rect 147772 220050 147824 220056
rect 147784 219745 147812 220050
rect 148060 220017 148088 231676
rect 148336 231662 148626 231690
rect 148336 223145 148364 231662
rect 149164 226137 149192 231676
rect 149520 228132 149572 228138
rect 149520 228074 149572 228080
rect 149150 226128 149206 226137
rect 149150 226063 149206 226072
rect 148322 223136 148378 223145
rect 148322 223071 148378 223080
rect 148966 222864 149022 222873
rect 148966 222799 149022 222808
rect 148980 220114 149008 222799
rect 148968 220108 149020 220114
rect 148968 220050 149020 220056
rect 149152 220108 149204 220114
rect 149152 220050 149204 220056
rect 148046 220008 148102 220017
rect 148046 219943 148102 219952
rect 147770 219736 147826 219745
rect 147770 219671 147826 219680
rect 149164 219450 149192 220050
rect 148796 219422 149192 219450
rect 147588 218204 147640 218210
rect 147588 218146 147640 218152
rect 147600 217410 147628 218146
rect 148796 217410 148824 219422
rect 149532 217410 149560 228074
rect 149716 225622 149744 231676
rect 150268 229770 150296 231676
rect 150544 231662 150834 231690
rect 150544 230353 150572 231662
rect 150530 230344 150586 230353
rect 150530 230279 150586 230288
rect 150256 229764 150308 229770
rect 150256 229706 150308 229712
rect 150440 229764 150492 229770
rect 150440 229706 150492 229712
rect 150452 228682 150480 229706
rect 150440 228676 150492 228682
rect 150440 228618 150492 228624
rect 150624 228676 150676 228682
rect 150624 228618 150676 228624
rect 150636 228274 150664 228618
rect 150624 228268 150676 228274
rect 150624 228210 150676 228216
rect 150808 228268 150860 228274
rect 150808 228210 150860 228216
rect 150820 228041 150848 228210
rect 150806 228032 150862 228041
rect 150806 227967 150862 227976
rect 151372 226681 151400 231676
rect 151924 229265 151952 231676
rect 152200 231662 152490 231690
rect 152752 231662 153042 231690
rect 153304 231662 153594 231690
rect 153856 231662 154146 231690
rect 151910 229256 151966 229265
rect 151910 229191 151966 229200
rect 151358 226672 151414 226681
rect 151358 226607 151414 226616
rect 149704 225616 149756 225622
rect 149704 225558 149756 225564
rect 151176 225616 151228 225622
rect 151176 225558 151228 225564
rect 151188 224954 151216 225558
rect 151450 225312 151506 225321
rect 151450 225247 151506 225256
rect 151188 224926 151308 224954
rect 150162 223408 150218 223417
rect 150162 223343 150218 223352
rect 150176 220114 150204 223343
rect 150346 220144 150402 220153
rect 150164 220108 150216 220114
rect 150346 220079 150402 220088
rect 151084 220108 151136 220114
rect 150164 220050 150216 220056
rect 150360 217410 150388 220079
rect 151084 220050 151136 220056
rect 151096 217410 151124 220050
rect 143276 217382 143428 217410
rect 144256 217382 144592 217410
rect 145084 217382 145420 217410
rect 145912 217382 146248 217410
rect 146740 217382 147076 217410
rect 147568 217382 147628 217410
rect 148396 217382 148824 217410
rect 149224 217382 149560 217410
rect 150052 217382 150388 217410
rect 150880 217382 151124 217410
rect 151280 217410 151308 224926
rect 151464 224806 151492 225247
rect 151636 225072 151688 225078
rect 151634 225040 151636 225049
rect 151774 225072 151826 225078
rect 151688 225040 151690 225049
rect 152200 225049 152228 231662
rect 152752 225321 152780 231662
rect 153304 227769 153332 231662
rect 153856 230897 153884 231662
rect 153842 230888 153898 230897
rect 153842 230823 153898 230832
rect 153750 230344 153806 230353
rect 153750 230279 153806 230288
rect 153764 230178 153792 230279
rect 153752 230172 153804 230178
rect 153752 230114 153804 230120
rect 153936 230172 153988 230178
rect 153936 230114 153988 230120
rect 153948 229906 153976 230114
rect 153936 229900 153988 229906
rect 153936 229842 153988 229848
rect 154120 229900 154172 229906
rect 154120 229842 154172 229848
rect 153290 227760 153346 227769
rect 153290 227695 153346 227704
rect 152738 225312 152794 225321
rect 152738 225247 152794 225256
rect 151774 225014 151826 225020
rect 152186 225040 152242 225049
rect 151634 224975 151690 224984
rect 151786 224954 151814 225014
rect 152186 224975 152242 224984
rect 151786 224926 151952 224954
rect 151452 224800 151504 224806
rect 151452 224742 151504 224748
rect 151728 224800 151780 224806
rect 151728 224742 151780 224748
rect 151740 224534 151768 224742
rect 151728 224528 151780 224534
rect 151924 224505 151952 224926
rect 152096 224528 152148 224534
rect 151728 224470 151780 224476
rect 151910 224496 151966 224505
rect 152096 224470 152148 224476
rect 151910 224431 151966 224440
rect 151636 221468 151688 221474
rect 151636 221410 151688 221416
rect 151820 221468 151872 221474
rect 151820 221410 151872 221416
rect 151648 221241 151676 221410
rect 151634 221232 151690 221241
rect 151634 221167 151690 221176
rect 151832 220114 151860 221410
rect 152108 220697 152136 224470
rect 152292 222958 152688 222986
rect 152292 222630 152320 222958
rect 152660 222902 152688 222958
rect 152464 222896 152516 222902
rect 152464 222838 152516 222844
rect 152648 222896 152700 222902
rect 152648 222838 152700 222844
rect 152476 222630 152504 222838
rect 152280 222624 152332 222630
rect 152280 222566 152332 222572
rect 152464 222624 152516 222630
rect 152464 222566 152516 222572
rect 154132 220794 154160 229842
rect 154684 229094 154712 231676
rect 154684 229066 154804 229094
rect 154302 226672 154358 226681
rect 154302 226607 154358 226616
rect 152464 220788 152516 220794
rect 152464 220730 152516 220736
rect 153660 220788 153712 220794
rect 153660 220730 153712 220736
rect 154120 220788 154172 220794
rect 154120 220730 154172 220736
rect 152094 220688 152150 220697
rect 152094 220623 152150 220632
rect 152476 220114 152504 220730
rect 151820 220108 151872 220114
rect 151820 220050 151872 220056
rect 152464 220108 152516 220114
rect 152464 220050 152516 220056
rect 152830 219736 152886 219745
rect 152830 219671 152886 219680
rect 152844 217410 152872 219671
rect 153672 217410 153700 220730
rect 154316 217410 154344 226607
rect 154776 222057 154804 229066
rect 155040 224528 155092 224534
rect 155038 224496 155040 224505
rect 155092 224496 155094 224505
rect 155038 224431 155094 224440
rect 155236 224262 155264 231676
rect 155788 228002 155816 231676
rect 156340 230178 156368 231676
rect 156524 231662 156906 231690
rect 157458 231662 157840 231690
rect 156328 230172 156380 230178
rect 156328 230114 156380 230120
rect 156524 229094 156552 231662
rect 156248 229066 156552 229094
rect 155776 227996 155828 228002
rect 155776 227938 155828 227944
rect 155960 227996 156012 228002
rect 155960 227938 156012 227944
rect 155972 227882 156000 227938
rect 155880 227854 156000 227882
rect 155408 224528 155460 224534
rect 155408 224470 155460 224476
rect 155224 224256 155276 224262
rect 155224 224198 155276 224204
rect 154762 222048 154818 222057
rect 154762 221983 154818 221992
rect 154488 220788 154540 220794
rect 154488 220730 154540 220736
rect 154500 219706 154528 220730
rect 154670 219736 154726 219745
rect 154488 219700 154540 219706
rect 154670 219671 154672 219680
rect 154488 219642 154540 219648
rect 154724 219671 154726 219680
rect 154672 219642 154724 219648
rect 155420 217410 155448 224470
rect 155592 224256 155644 224262
rect 155592 224198 155644 224204
rect 155604 223417 155632 224198
rect 155590 223408 155646 223417
rect 155590 223343 155646 223352
rect 155880 217410 155908 227854
rect 156248 221241 156276 229066
rect 156602 228032 156658 228041
rect 156602 227967 156658 227976
rect 156616 227186 156644 227967
rect 157430 227760 157486 227769
rect 157430 227695 157486 227704
rect 157444 227322 157472 227695
rect 157812 227338 157840 231662
rect 157996 228410 158024 231676
rect 158180 231662 158562 231690
rect 158916 231662 159114 231690
rect 159376 231662 159666 231690
rect 157984 228404 158036 228410
rect 157984 228346 158036 228352
rect 157432 227316 157484 227322
rect 157812 227310 158024 227338
rect 157432 227258 157484 227264
rect 157708 227248 157760 227254
rect 157536 227196 157708 227202
rect 157536 227190 157760 227196
rect 156604 227180 156656 227186
rect 156604 227122 156656 227128
rect 157536 227174 157748 227190
rect 157536 227050 157564 227174
rect 157524 227044 157576 227050
rect 157524 226986 157576 226992
rect 157800 227044 157852 227050
rect 157800 226986 157852 226992
rect 157812 226681 157840 226986
rect 157798 226672 157854 226681
rect 157798 226607 157854 226616
rect 157338 224768 157394 224777
rect 157338 224703 157394 224712
rect 157352 224618 157380 224703
rect 157306 224590 157380 224618
rect 157306 224534 157334 224590
rect 157294 224528 157346 224534
rect 157432 224528 157484 224534
rect 157294 224470 157346 224476
rect 157430 224496 157432 224505
rect 157484 224496 157486 224505
rect 157430 224431 157486 224440
rect 157798 224496 157854 224505
rect 157798 224431 157854 224440
rect 157294 223168 157346 223174
rect 157154 223136 157210 223145
rect 157432 223168 157484 223174
rect 157294 223110 157346 223116
rect 157430 223136 157432 223145
rect 157484 223136 157486 223145
rect 157154 223071 157210 223080
rect 157168 222902 157196 223071
rect 157306 222986 157334 223110
rect 157430 223071 157486 223080
rect 157306 222958 157564 222986
rect 157156 222896 157208 222902
rect 157340 222896 157392 222902
rect 157156 222838 157208 222844
rect 157338 222864 157340 222873
rect 157536 222873 157564 222958
rect 157392 222864 157394 222873
rect 157338 222799 157394 222808
rect 157522 222864 157578 222873
rect 157522 222799 157578 222808
rect 156234 221232 156290 221241
rect 156234 221167 156290 221176
rect 157812 220697 157840 224431
rect 157996 224233 158024 227310
rect 157982 224224 158038 224233
rect 157982 224159 158038 224168
rect 157982 223136 158038 223145
rect 157982 223071 158038 223080
rect 156878 220688 156934 220697
rect 156878 220623 156934 220632
rect 157798 220688 157854 220697
rect 157798 220623 157854 220632
rect 156892 220250 156920 220623
rect 156880 220244 156932 220250
rect 156880 220186 156932 220192
rect 156800 220114 157380 220130
rect 156800 220108 157392 220114
rect 156800 220102 157340 220108
rect 156800 219706 156828 220102
rect 157340 220050 157392 220056
rect 156788 219700 156840 219706
rect 156788 219642 156840 219648
rect 156972 219700 157024 219706
rect 156972 219642 157024 219648
rect 156984 217410 157012 219642
rect 157996 217410 158024 223071
rect 158180 222902 158208 231662
rect 158442 229120 158498 229129
rect 158442 229055 158498 229064
rect 158456 225486 158484 229055
rect 158444 225480 158496 225486
rect 158444 225422 158496 225428
rect 158628 225480 158680 225486
rect 158628 225422 158680 225428
rect 158168 222896 158220 222902
rect 158352 222896 158404 222902
rect 158168 222838 158220 222844
rect 158350 222864 158352 222873
rect 158404 222864 158406 222873
rect 158350 222799 158406 222808
rect 158640 217410 158668 225422
rect 158916 220969 158944 231662
rect 159376 224806 159404 231662
rect 159732 230036 159784 230042
rect 159732 229978 159784 229984
rect 159744 229770 159772 229978
rect 159732 229764 159784 229770
rect 159732 229706 159784 229712
rect 159732 228404 159784 228410
rect 159732 228346 159784 228352
rect 159744 224954 159772 228346
rect 160204 228041 160232 231676
rect 160480 231662 160770 231690
rect 161124 231662 161322 231690
rect 160480 230353 160508 231662
rect 160466 230344 160522 230353
rect 160466 230279 160522 230288
rect 160744 229900 160796 229906
rect 160744 229842 160796 229848
rect 160190 228032 160246 228041
rect 160190 227967 160246 227976
rect 159560 224926 159772 224954
rect 159364 224800 159416 224806
rect 159364 224742 159416 224748
rect 158902 220960 158958 220969
rect 158902 220895 158958 220904
rect 159560 217410 159588 224926
rect 159732 224800 159784 224806
rect 159732 224742 159784 224748
rect 159744 224534 159772 224742
rect 159732 224528 159784 224534
rect 159916 224528 159968 224534
rect 159732 224470 159784 224476
rect 159914 224496 159916 224505
rect 159968 224496 159970 224505
rect 159914 224431 159970 224440
rect 160756 221474 160784 229842
rect 161124 223174 161152 231662
rect 161478 230344 161534 230353
rect 161478 230279 161534 230288
rect 161492 225162 161520 230279
rect 161860 225758 161888 231676
rect 162412 228546 162440 231676
rect 162400 228540 162452 228546
rect 162400 228482 162452 228488
rect 162400 226160 162452 226166
rect 162400 226102 162452 226108
rect 161848 225752 161900 225758
rect 161848 225694 161900 225700
rect 161308 225134 161520 225162
rect 161308 225078 161336 225134
rect 161296 225072 161348 225078
rect 161296 225014 161348 225020
rect 161480 225072 161532 225078
rect 161480 225014 161532 225020
rect 161492 224777 161520 225014
rect 161478 224768 161534 224777
rect 161478 224703 161534 224712
rect 161940 223440 161992 223446
rect 161940 223382 161992 223388
rect 161952 223174 161980 223382
rect 161112 223168 161164 223174
rect 161112 223110 161164 223116
rect 161940 223168 161992 223174
rect 161940 223110 161992 223116
rect 159824 221468 159876 221474
rect 159824 221410 159876 221416
rect 160008 221468 160060 221474
rect 160008 221410 160060 221416
rect 160744 221468 160796 221474
rect 160744 221410 160796 221416
rect 160928 221468 160980 221474
rect 160928 221410 160980 221416
rect 159836 221241 159864 221410
rect 159822 221232 159878 221241
rect 159822 221167 159878 221176
rect 160020 217410 160048 221410
rect 160940 221241 160968 221410
rect 160926 221232 160982 221241
rect 160926 221167 160982 221176
rect 161110 221232 161166 221241
rect 161110 221167 161166 221176
rect 160926 219600 160982 219609
rect 160926 219535 160928 219544
rect 160980 219535 160982 219544
rect 160928 219506 160980 219512
rect 161124 217410 161152 221167
rect 162412 220522 162440 226102
rect 162964 224534 162992 231676
rect 162952 224528 163004 224534
rect 162952 224470 163004 224476
rect 163136 224528 163188 224534
rect 163136 224470 163188 224476
rect 163148 224346 163176 224470
rect 162780 224318 163176 224346
rect 161756 220516 161808 220522
rect 161756 220458 161808 220464
rect 161940 220516 161992 220522
rect 161940 220458 161992 220464
rect 162400 220516 162452 220522
rect 162400 220458 162452 220464
rect 162584 220516 162636 220522
rect 162584 220458 162636 220464
rect 161768 220250 161796 220458
rect 161296 220244 161348 220250
rect 161296 220186 161348 220192
rect 161756 220244 161808 220250
rect 161756 220186 161808 220192
rect 161308 219570 161336 220186
rect 161296 219564 161348 219570
rect 161296 219506 161348 219512
rect 161952 217410 161980 220458
rect 162596 219570 162624 220458
rect 162584 219564 162636 219570
rect 162584 219506 162636 219512
rect 162780 217410 162808 224318
rect 163516 223038 163544 231676
rect 163792 231662 164082 231690
rect 164344 231662 164634 231690
rect 163792 229129 163820 231662
rect 164344 230625 164372 231662
rect 164330 230616 164386 230625
rect 164330 230551 164386 230560
rect 165172 229537 165200 231676
rect 165632 231662 165738 231690
rect 166000 231662 166290 231690
rect 166552 231662 166842 231690
rect 165158 229528 165214 229537
rect 165158 229463 165214 229472
rect 163778 229120 163834 229129
rect 165632 229106 165660 231662
rect 163778 229055 163834 229064
rect 165540 229078 165660 229106
rect 165160 227180 165212 227186
rect 165160 227122 165212 227128
rect 165172 224954 165200 227122
rect 165080 224926 165200 224954
rect 163504 223032 163556 223038
rect 163504 222974 163556 222980
rect 164148 223032 164200 223038
rect 164148 222974 164200 222980
rect 163596 219564 163648 219570
rect 163596 219506 163648 219512
rect 163608 217410 163636 219506
rect 164160 217410 164188 222974
rect 165080 220522 165108 224926
rect 165252 223168 165304 223174
rect 165252 223110 165304 223116
rect 165068 220516 165120 220522
rect 165068 220458 165120 220464
rect 165264 217410 165292 223110
rect 165540 222902 165568 229078
rect 166000 226030 166028 231662
rect 166264 228540 166316 228546
rect 166264 228482 166316 228488
rect 165988 226024 166040 226030
rect 165988 225966 166040 225972
rect 166276 224954 166304 228482
rect 166552 227769 166580 231662
rect 166814 230888 166870 230897
rect 166814 230823 166870 230832
rect 166828 230178 166856 230823
rect 166998 230344 167054 230353
rect 166998 230279 167054 230288
rect 167012 230178 167040 230279
rect 166816 230172 166868 230178
rect 166816 230114 166868 230120
rect 167000 230172 167052 230178
rect 167000 230114 167052 230120
rect 166538 227760 166594 227769
rect 166538 227695 166594 227704
rect 167000 226296 167052 226302
rect 166998 226264 167000 226273
rect 167184 226296 167236 226302
rect 167052 226264 167054 226273
rect 167184 226238 167236 226244
rect 166998 226199 167054 226208
rect 166448 226024 166500 226030
rect 166448 225966 166500 225972
rect 166184 224926 166304 224954
rect 165710 223136 165766 223145
rect 165710 223071 165766 223080
rect 165724 222902 165752 223071
rect 165528 222896 165580 222902
rect 165528 222838 165580 222844
rect 165712 222896 165764 222902
rect 165712 222838 165764 222844
rect 165620 220516 165672 220522
rect 165620 220458 165672 220464
rect 165632 219609 165660 220458
rect 165986 220416 166042 220425
rect 165986 220351 165988 220360
rect 166040 220351 166042 220360
rect 165988 220322 166040 220328
rect 165618 219600 165674 219609
rect 165618 219535 165674 219544
rect 166184 217410 166212 224926
rect 166460 220522 166488 225966
rect 167196 225894 167224 226238
rect 167380 226030 167408 231676
rect 167656 231662 167946 231690
rect 167368 226024 167420 226030
rect 167368 225966 167420 225972
rect 167184 225888 167236 225894
rect 167184 225830 167236 225836
rect 167656 223446 167684 231662
rect 168484 226030 168512 231676
rect 168668 231662 169050 231690
rect 169312 231662 169602 231690
rect 168472 226024 168524 226030
rect 168472 225966 168524 225972
rect 168288 225888 168340 225894
rect 168288 225830 168340 225836
rect 167828 225752 167880 225758
rect 167828 225694 167880 225700
rect 167644 223440 167696 223446
rect 167644 223382 167696 223388
rect 166644 221598 166994 221626
rect 166644 221241 166672 221598
rect 166966 221474 166994 221598
rect 166816 221468 166868 221474
rect 166816 221410 166868 221416
rect 166954 221468 167006 221474
rect 166954 221410 167006 221416
rect 166630 221232 166686 221241
rect 166630 221167 166686 221176
rect 166828 221105 166856 221410
rect 166814 221096 166870 221105
rect 166814 221031 166870 221040
rect 166448 220516 166500 220522
rect 166448 220458 166500 220464
rect 166632 220516 166684 220522
rect 166632 220458 166684 220464
rect 166644 217410 166672 220458
rect 166954 220244 167006 220250
rect 166828 220204 166954 220232
rect 166828 219978 166856 220204
rect 166954 220186 167006 220192
rect 166816 219972 166868 219978
rect 166816 219914 166868 219920
rect 166954 219972 167006 219978
rect 166954 219914 167006 219920
rect 166966 219858 166994 219914
rect 166920 219830 166994 219858
rect 166920 219570 166948 219830
rect 166908 219564 166960 219570
rect 166908 219506 166960 219512
rect 167840 217410 167868 225694
rect 168300 217410 168328 225830
rect 151280 217382 151708 217410
rect 152536 217382 152872 217410
rect 153364 217382 153700 217410
rect 154192 217382 154344 217410
rect 155020 217382 155448 217410
rect 155848 217382 155908 217410
rect 156676 217382 157012 217410
rect 157504 217382 158024 217410
rect 158332 217382 158668 217410
rect 159160 217382 159588 217410
rect 159988 217382 160048 217410
rect 160816 217382 161152 217410
rect 161644 217382 161980 217410
rect 162472 217382 162808 217410
rect 163300 217382 163636 217410
rect 164128 217382 164188 217410
rect 164956 217382 165292 217410
rect 165784 217382 166212 217410
rect 166612 217382 166672 217410
rect 167440 217382 167868 217410
rect 168268 217382 168328 217410
rect 62764 217320 62816 217326
rect 62764 217262 62816 217268
rect 110308 217258 110460 217274
rect 110308 217252 110472 217258
rect 110308 217246 110420 217252
rect 110420 217194 110472 217200
rect 100372 217122 100708 217138
rect 100372 217116 100720 217122
rect 100372 217110 100668 217116
rect 100668 217058 100720 217064
rect 93748 216986 93900 217002
rect 93748 216980 93912 216986
rect 93748 216974 93860 216980
rect 93860 216922 93912 216928
rect 90436 216850 90772 216866
rect 90436 216844 90784 216850
rect 90436 216838 90732 216844
rect 90732 216786 90784 216792
rect 85468 216714 85620 216730
rect 168668 216714 168696 231662
rect 169312 230897 169340 231662
rect 169298 230888 169354 230897
rect 169298 230823 169354 230832
rect 168838 230344 168894 230353
rect 168838 230279 168894 230288
rect 168852 230042 168880 230279
rect 170140 230042 170168 231676
rect 168840 230036 168892 230042
rect 168840 229978 168892 229984
rect 169024 230036 169076 230042
rect 169024 229978 169076 229984
rect 170128 230036 170180 230042
rect 170128 229978 170180 229984
rect 169036 220425 169064 229978
rect 170034 229528 170090 229537
rect 170034 229463 170090 229472
rect 169022 220416 169078 220425
rect 170048 220386 170076 229463
rect 170692 223310 170720 231676
rect 171244 230654 171272 231676
rect 171428 231662 171810 231690
rect 172072 231662 172362 231690
rect 172624 231662 172914 231690
rect 171232 230648 171284 230654
rect 171232 230590 171284 230596
rect 171140 230036 171192 230042
rect 171140 229978 171192 229984
rect 171152 228818 171180 229978
rect 171140 228812 171192 228818
rect 171140 228754 171192 228760
rect 170680 223304 170732 223310
rect 170680 223246 170732 223252
rect 170864 223304 170916 223310
rect 170864 223246 170916 223252
rect 169022 220351 169078 220360
rect 170036 220380 170088 220386
rect 170036 220322 170088 220328
rect 170220 220380 170272 220386
rect 170220 220322 170272 220328
rect 169392 219564 169444 219570
rect 169392 219506 169444 219512
rect 169404 217410 169432 219506
rect 170232 217410 170260 220322
rect 170876 219434 170904 223246
rect 171138 222048 171194 222057
rect 171138 221983 171194 221992
rect 171152 221898 171180 221983
rect 171060 221870 171180 221898
rect 171060 221746 171088 221870
rect 171048 221740 171100 221746
rect 171048 221682 171100 221688
rect 171232 221740 171284 221746
rect 171232 221682 171284 221688
rect 171244 221218 171272 221682
rect 171060 221190 171272 221218
rect 171060 221066 171088 221190
rect 171230 221096 171286 221105
rect 171048 221060 171100 221066
rect 171230 221031 171232 221040
rect 171048 221002 171100 221008
rect 171284 221031 171286 221040
rect 171232 221002 171284 221008
rect 171048 220244 171100 220250
rect 171048 220186 171100 220192
rect 171060 219881 171088 220186
rect 171046 219872 171102 219881
rect 171046 219807 171102 219816
rect 171428 219434 171456 231662
rect 172072 230353 172100 231662
rect 172058 230344 172114 230353
rect 172058 230279 172114 230288
rect 172334 228032 172390 228041
rect 172334 227967 172390 227976
rect 171876 220244 171928 220250
rect 171876 220186 171928 220192
rect 170876 219406 170996 219434
rect 170968 217410 170996 219406
rect 169096 217382 169432 217410
rect 169924 217382 170260 217410
rect 170752 217382 170996 217410
rect 171152 219406 171456 219434
rect 171152 216850 171180 219406
rect 171888 217410 171916 220186
rect 171580 217382 171916 217410
rect 172348 217410 172376 227967
rect 172624 223446 172652 231662
rect 173452 226302 173480 231676
rect 174018 231662 174400 231690
rect 173440 226296 173492 226302
rect 173624 226296 173676 226302
rect 173440 226238 173492 226244
rect 173622 226264 173624 226273
rect 173676 226264 173678 226273
rect 173622 226199 173678 226208
rect 173256 226160 173308 226166
rect 173256 226102 173308 226108
rect 172612 223440 172664 223446
rect 172612 223382 172664 223388
rect 173072 223168 173124 223174
rect 173072 223110 173124 223116
rect 173084 223009 173112 223110
rect 173070 223000 173126 223009
rect 173070 222935 173126 222944
rect 173268 219881 173296 226102
rect 173808 223576 173860 223582
rect 173808 223518 173860 223524
rect 173532 223440 173584 223446
rect 173532 223382 173584 223388
rect 173544 222630 173572 223382
rect 173532 222624 173584 222630
rect 173532 222566 173584 222572
rect 173438 220416 173494 220425
rect 173438 220351 173494 220360
rect 173452 220250 173480 220351
rect 173440 220244 173492 220250
rect 173440 220186 173492 220192
rect 173624 220244 173676 220250
rect 173624 220186 173676 220192
rect 173254 219872 173310 219881
rect 173254 219807 173310 219816
rect 173636 217410 173664 220186
rect 173820 219570 173848 223518
rect 174084 223032 174136 223038
rect 174082 223000 174084 223009
rect 174136 223000 174138 223009
rect 174082 222935 174138 222944
rect 173808 219564 173860 219570
rect 173808 219506 173860 219512
rect 174176 219564 174228 219570
rect 174176 219506 174228 219512
rect 174188 217410 174216 219506
rect 172348 217382 172408 217410
rect 173236 217382 173664 217410
rect 174064 217382 174216 217410
rect 174372 216986 174400 231662
rect 174556 230042 174584 231676
rect 174832 231662 175122 231690
rect 174544 230036 174596 230042
rect 174544 229978 174596 229984
rect 174832 222057 174860 231662
rect 175004 230036 175056 230042
rect 175004 229978 175056 229984
rect 175016 229537 175044 229978
rect 175002 229528 175058 229537
rect 175002 229463 175058 229472
rect 175660 226302 175688 231676
rect 175844 231662 176226 231690
rect 176672 231662 176778 231690
rect 177040 231662 177330 231690
rect 175844 227322 175872 231662
rect 176028 229066 176516 229094
rect 175832 227316 175884 227322
rect 175832 227258 175884 227264
rect 175648 226296 175700 226302
rect 175648 226238 175700 226244
rect 175832 226296 175884 226302
rect 175832 226238 175884 226244
rect 175188 222624 175240 222630
rect 175188 222566 175240 222572
rect 174818 222048 174874 222057
rect 174818 221983 174874 221992
rect 175200 217410 175228 222566
rect 175844 220425 175872 226238
rect 175830 220416 175886 220425
rect 175830 220351 175886 220360
rect 175832 218748 175884 218754
rect 175832 218690 175884 218696
rect 175844 218074 175872 218690
rect 175832 218068 175884 218074
rect 175832 218010 175884 218016
rect 176028 217410 176056 229066
rect 176488 228954 176516 229066
rect 176476 228948 176528 228954
rect 176672 228936 176700 231662
rect 176844 230444 176896 230450
rect 176844 230386 176896 230392
rect 176856 229090 176884 230386
rect 176844 229084 176896 229090
rect 176844 229026 176896 229032
rect 176476 228890 176528 228896
rect 176626 228908 176700 228936
rect 176626 228818 176654 228908
rect 176614 228812 176666 228818
rect 176614 228754 176666 228760
rect 176752 226296 176804 226302
rect 176752 226238 176804 226244
rect 176476 226160 176528 226166
rect 176474 226128 176476 226137
rect 176764 226137 176792 226238
rect 176528 226128 176530 226137
rect 176474 226063 176530 226072
rect 176750 226128 176806 226137
rect 176750 226063 176806 226072
rect 177040 223446 177068 231662
rect 177868 224670 177896 231676
rect 178328 231662 178434 231690
rect 178132 225344 178184 225350
rect 178130 225312 178132 225321
rect 178184 225312 178186 225321
rect 178130 225247 178186 225256
rect 177856 224664 177908 224670
rect 177856 224606 177908 224612
rect 178040 224664 178092 224670
rect 178040 224606 178092 224612
rect 178052 224482 178080 224606
rect 177868 224454 178080 224482
rect 177028 223440 177080 223446
rect 177028 223382 177080 223388
rect 176566 220824 176622 220833
rect 176566 220759 176622 220768
rect 176580 219570 176608 220759
rect 177868 220561 177896 224454
rect 177854 220552 177910 220561
rect 177854 220487 177910 220496
rect 176568 219564 176620 219570
rect 176568 219506 176620 219512
rect 177672 219564 177724 219570
rect 177672 219506 177724 219512
rect 176200 219020 176252 219026
rect 176200 218962 176252 218968
rect 176568 219020 176620 219026
rect 176568 218962 176620 218968
rect 176212 218754 176240 218962
rect 176200 218748 176252 218754
rect 176200 218690 176252 218696
rect 176580 217410 176608 218962
rect 177684 217410 177712 219506
rect 178328 219434 178356 231662
rect 178972 228682 179000 231676
rect 179538 231662 179736 231690
rect 179236 228812 179288 228818
rect 179236 228754 179288 228760
rect 178960 228676 179012 228682
rect 178960 228618 179012 228624
rect 179052 227316 179104 227322
rect 179052 227258 179104 227264
rect 179064 226914 179092 227258
rect 179052 226908 179104 226914
rect 179052 226850 179104 226856
rect 178500 225344 178552 225350
rect 178500 225286 178552 225292
rect 174892 217382 175228 217410
rect 175720 217382 176056 217410
rect 176548 217382 176608 217410
rect 177376 217382 177712 217410
rect 178052 219406 178356 219434
rect 178052 217122 178080 219406
rect 178512 217410 178540 225286
rect 179248 222194 179276 228754
rect 179156 222166 179276 222194
rect 179156 219434 179184 222166
rect 179064 219406 179184 219434
rect 179064 217410 179092 219406
rect 179708 218754 179736 231662
rect 179892 231662 180090 231690
rect 179892 225321 179920 231662
rect 179878 225312 179934 225321
rect 179878 225247 179934 225256
rect 180628 224806 180656 231676
rect 180996 231662 181194 231690
rect 180798 226128 180854 226137
rect 180798 226063 180854 226072
rect 180812 225894 180840 226063
rect 180800 225888 180852 225894
rect 180800 225830 180852 225836
rect 180616 224800 180668 224806
rect 180616 224742 180668 224748
rect 180800 224800 180852 224806
rect 180800 224742 180852 224748
rect 180812 224618 180840 224742
rect 180168 224590 180840 224618
rect 179696 218748 179748 218754
rect 179696 218690 179748 218696
rect 180168 217410 180196 224590
rect 180708 223576 180760 223582
rect 180708 223518 180760 223524
rect 180522 219600 180578 219609
rect 180522 219535 180524 219544
rect 180576 219535 180578 219544
rect 180524 219506 180576 219512
rect 180720 219434 180748 223518
rect 180996 220402 181024 231662
rect 181260 230716 181312 230722
rect 181260 230658 181312 230664
rect 181272 230450 181300 230658
rect 181260 230444 181312 230450
rect 181260 230386 181312 230392
rect 181444 230444 181496 230450
rect 181444 230386 181496 230392
rect 181456 229634 181484 230386
rect 181444 229628 181496 229634
rect 181444 229570 181496 229576
rect 181732 227866 181760 231676
rect 182298 231662 182680 231690
rect 182088 229628 182140 229634
rect 182088 229570 182140 229576
rect 182100 228834 182128 229570
rect 182008 228806 182128 228834
rect 182364 228812 182416 228818
rect 181720 227860 181772 227866
rect 181720 227802 181772 227808
rect 181352 226160 181404 226166
rect 181350 226128 181352 226137
rect 181404 226128 181406 226137
rect 181350 226063 181406 226072
rect 182008 224954 182036 228806
rect 182364 228754 182416 228760
rect 182180 228676 182232 228682
rect 182180 228618 182232 228624
rect 182192 228562 182220 228618
rect 181916 224926 182036 224954
rect 182100 228534 182220 228562
rect 181916 224806 181944 224926
rect 181904 224800 181956 224806
rect 181904 224742 181956 224748
rect 182100 224074 182128 228534
rect 182376 228041 182404 228754
rect 182362 228032 182418 228041
rect 182362 227967 182418 227976
rect 181824 224046 182128 224074
rect 181166 223000 181222 223009
rect 181166 222935 181222 222944
rect 181180 222222 181208 222935
rect 181168 222216 181220 222222
rect 181168 222158 181220 222164
rect 181444 222148 181496 222154
rect 181444 222090 181496 222096
rect 181456 221898 181484 222090
rect 181272 221870 181484 221898
rect 181272 221746 181300 221870
rect 181260 221740 181312 221746
rect 181260 221682 181312 221688
rect 181444 221740 181496 221746
rect 181444 221682 181496 221688
rect 181456 220833 181484 221682
rect 181442 220824 181498 220833
rect 181442 220759 181498 220768
rect 178204 217382 178540 217410
rect 179032 217382 179092 217410
rect 179860 217382 180196 217410
rect 180536 219406 180748 219434
rect 180904 220374 181024 220402
rect 181166 220416 181222 220425
rect 180904 219434 180932 220374
rect 181166 220351 181222 220360
rect 181180 220266 181208 220351
rect 181088 220250 181208 220266
rect 181076 220244 181208 220250
rect 181128 220238 181208 220244
rect 181076 220186 181128 220192
rect 181168 219564 181220 219570
rect 181168 219506 181220 219512
rect 180904 219406 181024 219434
rect 180536 217410 180564 219406
rect 180996 218890 181024 219406
rect 181180 219026 181208 219506
rect 181824 219434 181852 224046
rect 181994 222048 182050 222057
rect 181994 221983 181996 221992
rect 182048 221983 182050 221992
rect 182180 222012 182232 222018
rect 181996 221954 182048 221960
rect 182180 221954 182232 221960
rect 182192 219609 182220 221954
rect 182178 219600 182234 219609
rect 182178 219535 182234 219544
rect 182652 219434 182680 231662
rect 182836 230314 182864 231676
rect 183112 231662 183402 231690
rect 183848 231662 183954 231690
rect 183112 230722 183140 231662
rect 183100 230716 183152 230722
rect 183100 230658 183152 230664
rect 182824 230308 182876 230314
rect 182824 230250 182876 230256
rect 183468 230308 183520 230314
rect 183468 230250 183520 230256
rect 182824 227044 182876 227050
rect 182824 226986 182876 226992
rect 182836 219434 182864 226986
rect 183480 222154 183508 230250
rect 183468 222148 183520 222154
rect 183468 222090 183520 222096
rect 183848 221882 183876 231662
rect 184492 230586 184520 231676
rect 185058 231662 185256 231690
rect 184480 230580 184532 230586
rect 184480 230522 184532 230528
rect 184848 224936 184900 224942
rect 184848 224878 184900 224884
rect 184296 222148 184348 222154
rect 184296 222090 184348 222096
rect 183836 221876 183888 221882
rect 183836 221818 183888 221824
rect 183282 219600 183338 219609
rect 183282 219535 183284 219544
rect 183336 219535 183338 219544
rect 183468 219564 183520 219570
rect 183284 219506 183336 219512
rect 183468 219506 183520 219512
rect 181824 219406 181944 219434
rect 181168 219020 181220 219026
rect 181168 218962 181220 218968
rect 180984 218884 181036 218890
rect 180984 218826 181036 218832
rect 181916 217410 181944 219406
rect 182560 219406 182680 219434
rect 182744 219406 182864 219434
rect 182560 218074 182588 219406
rect 182548 218068 182600 218074
rect 182548 218010 182600 218016
rect 182744 217410 182772 219406
rect 183480 217410 183508 219506
rect 184308 217410 184336 222090
rect 184860 217410 184888 224878
rect 185030 223408 185086 223417
rect 185030 223343 185086 223352
rect 185044 222766 185072 223343
rect 185032 222760 185084 222766
rect 185032 222702 185084 222708
rect 180536 217382 180688 217410
rect 181516 217382 181944 217410
rect 182344 217382 182772 217410
rect 183172 217382 183508 217410
rect 184000 217382 184336 217410
rect 184828 217382 184888 217410
rect 185228 217258 185256 231662
rect 185412 231662 185610 231690
rect 185780 231662 186162 231690
rect 186608 231662 186714 231690
rect 185412 219298 185440 231662
rect 185780 224954 185808 231662
rect 185952 227044 186004 227050
rect 185952 226986 186004 226992
rect 186136 227044 186188 227050
rect 186136 226986 186188 226992
rect 185964 226681 185992 226986
rect 185950 226672 186006 226681
rect 185950 226607 186006 226616
rect 185596 224926 185808 224954
rect 185596 223417 185624 224926
rect 185582 223408 185638 223417
rect 185582 223343 185638 223352
rect 185584 223168 185636 223174
rect 185584 223110 185636 223116
rect 185768 223168 185820 223174
rect 185768 223110 185820 223116
rect 185596 222630 185624 223110
rect 185780 222766 185808 223110
rect 185768 222760 185820 222766
rect 185768 222702 185820 222708
rect 185584 222624 185636 222630
rect 185584 222566 185636 222572
rect 185768 222012 185820 222018
rect 185768 221954 185820 221960
rect 185584 221876 185636 221882
rect 185584 221818 185636 221824
rect 185596 221338 185624 221818
rect 185780 221338 185808 221954
rect 185584 221332 185636 221338
rect 185584 221274 185636 221280
rect 185768 221332 185820 221338
rect 185768 221274 185820 221280
rect 186148 219434 186176 226986
rect 186056 219406 186176 219434
rect 185400 219292 185452 219298
rect 185400 219234 185452 219240
rect 186056 217410 186084 219406
rect 186608 219162 186636 231662
rect 187252 227186 187280 231676
rect 187424 230444 187476 230450
rect 187424 230386 187476 230392
rect 187240 227180 187292 227186
rect 187240 227122 187292 227128
rect 187054 225040 187110 225049
rect 187054 224975 187110 224984
rect 187068 224806 187096 224975
rect 187056 224800 187108 224806
rect 187056 224742 187108 224748
rect 187240 224800 187292 224806
rect 187240 224742 187292 224748
rect 186872 220244 186924 220250
rect 186872 220186 186924 220192
rect 186596 219156 186648 219162
rect 186596 219098 186648 219104
rect 186884 217410 186912 220186
rect 187252 219434 187280 224742
rect 187436 220250 187464 230386
rect 187804 222057 187832 231676
rect 187988 231662 188370 231690
rect 187988 229094 188016 231662
rect 187988 229066 188200 229094
rect 187976 227044 188028 227050
rect 187976 226986 188028 226992
rect 187988 226681 188016 226986
rect 187974 226672 188030 226681
rect 187974 226607 188030 226616
rect 187790 222048 187846 222057
rect 187790 221983 187846 221992
rect 187424 220244 187476 220250
rect 187424 220186 187476 220192
rect 187608 220244 187660 220250
rect 187608 220186 187660 220192
rect 187620 219978 187648 220186
rect 187608 219972 187660 219978
rect 187608 219914 187660 219920
rect 187792 219972 187844 219978
rect 187792 219914 187844 219920
rect 187804 219570 187832 219914
rect 187974 219600 188030 219609
rect 187792 219564 187844 219570
rect 187974 219535 187976 219544
rect 187792 219506 187844 219512
rect 188028 219535 188030 219544
rect 187976 219506 188028 219512
rect 188172 219434 188200 229066
rect 188908 227458 188936 231676
rect 189184 231662 189474 231690
rect 189644 231662 190026 231690
rect 189184 230586 189212 231662
rect 189172 230580 189224 230586
rect 189172 230522 189224 230528
rect 188896 227452 188948 227458
rect 188896 227394 188948 227400
rect 189080 227452 189132 227458
rect 189080 227394 189132 227400
rect 189092 227338 189120 227394
rect 188816 227310 189120 227338
rect 187252 219406 187556 219434
rect 187528 217410 187556 219406
rect 188160 219428 188212 219434
rect 188160 219370 188212 219376
rect 188436 217864 188488 217870
rect 188436 217806 188488 217812
rect 188448 217410 188476 217806
rect 185656 217382 186084 217410
rect 186484 217382 186912 217410
rect 187312 217382 187556 217410
rect 188140 217382 188476 217410
rect 188816 217410 188844 227310
rect 189644 223009 189672 231662
rect 190564 230602 190592 231676
rect 190564 230574 190684 230602
rect 190274 230480 190330 230489
rect 190274 230415 190276 230424
rect 190328 230415 190330 230424
rect 190458 230480 190514 230489
rect 190458 230415 190460 230424
rect 190276 230386 190328 230392
rect 190512 230415 190514 230424
rect 190460 230386 190512 230392
rect 190656 229650 190684 230574
rect 190380 229622 190684 229650
rect 190380 229378 190408 229622
rect 190918 229528 190974 229537
rect 190918 229463 190920 229472
rect 190972 229463 190974 229472
rect 190920 229434 190972 229440
rect 190380 229350 190500 229378
rect 190472 229106 190500 229350
rect 190642 229256 190698 229265
rect 190642 229191 190698 229200
rect 190380 229094 190500 229106
rect 190012 229078 190500 229094
rect 190012 229066 190408 229078
rect 190012 225049 190040 229066
rect 190276 226296 190328 226302
rect 190274 226264 190276 226273
rect 190414 226296 190466 226302
rect 190328 226264 190330 226273
rect 190414 226238 190466 226244
rect 190274 226199 190330 226208
rect 190426 226114 190454 226238
rect 190196 226086 190454 226114
rect 189998 225040 190054 225049
rect 189998 224975 190054 224984
rect 190196 224890 190224 226086
rect 189920 224862 190224 224890
rect 189630 223000 189686 223009
rect 189630 222935 189686 222944
rect 188988 222148 189040 222154
rect 188988 222090 189040 222096
rect 189000 217870 189028 222090
rect 189920 220425 189948 224862
rect 190656 224777 190684 229191
rect 191116 227594 191144 231676
rect 191392 231662 191682 231690
rect 191944 231662 192234 231690
rect 191104 227588 191156 227594
rect 191104 227530 191156 227536
rect 191392 226273 191420 231662
rect 191748 230580 191800 230586
rect 191748 230522 191800 230528
rect 191760 230042 191788 230522
rect 191748 230036 191800 230042
rect 191748 229978 191800 229984
rect 191564 229628 191616 229634
rect 191564 229570 191616 229576
rect 191576 229265 191604 229570
rect 191562 229256 191618 229265
rect 191562 229191 191618 229200
rect 191378 226264 191434 226273
rect 191378 226199 191434 226208
rect 190366 224768 190422 224777
rect 190366 224703 190422 224712
rect 190642 224768 190698 224777
rect 190642 224703 190698 224712
rect 190380 224126 190408 224703
rect 190368 224120 190420 224126
rect 190368 224062 190420 224068
rect 191748 224120 191800 224126
rect 191748 224062 191800 224068
rect 191564 222760 191616 222766
rect 191564 222702 191616 222708
rect 189906 220416 189962 220425
rect 189906 220351 189962 220360
rect 190092 219428 190144 219434
rect 190092 219370 190144 219376
rect 188988 217864 189040 217870
rect 188988 217806 189040 217812
rect 190104 217410 190132 219370
rect 190920 217864 190972 217870
rect 190920 217806 190972 217812
rect 190932 217410 190960 217806
rect 191576 217410 191604 222702
rect 191760 217870 191788 224062
rect 191944 221882 191972 231662
rect 192116 230036 192168 230042
rect 192116 229978 192168 229984
rect 192128 227322 192156 229978
rect 192772 229634 192800 231676
rect 193324 230042 193352 231676
rect 193600 231662 193890 231690
rect 194060 231662 194442 231690
rect 194704 231662 194994 231690
rect 193600 230586 193628 231662
rect 193588 230580 193640 230586
rect 193588 230522 193640 230528
rect 193312 230036 193364 230042
rect 193312 229978 193364 229984
rect 192760 229628 192812 229634
rect 192760 229570 192812 229576
rect 192668 227588 192720 227594
rect 192668 227530 192720 227536
rect 192116 227316 192168 227322
rect 192116 227258 192168 227264
rect 192484 222012 192536 222018
rect 192484 221954 192536 221960
rect 191932 221876 191984 221882
rect 191932 221818 191984 221824
rect 192298 221232 192354 221241
rect 192496 221202 192524 221954
rect 192298 221167 192300 221176
rect 192352 221167 192354 221176
rect 192484 221196 192536 221202
rect 192300 221138 192352 221144
rect 192484 221138 192536 221144
rect 192482 220688 192538 220697
rect 192482 220623 192484 220632
rect 192536 220623 192538 220632
rect 192484 220594 192536 220600
rect 191748 217864 191800 217870
rect 191748 217806 191800 217812
rect 192680 217410 192708 227530
rect 193494 224224 193550 224233
rect 193494 224159 193550 224168
rect 193508 223854 193536 224159
rect 193496 223848 193548 223854
rect 193496 223790 193548 223796
rect 192852 222080 192904 222086
rect 192852 222022 192904 222028
rect 188816 217382 188968 217410
rect 189796 217382 190132 217410
rect 190624 217382 190960 217410
rect 191452 217382 191604 217410
rect 192280 217382 192708 217410
rect 192864 217410 192892 222022
rect 194060 220697 194088 231662
rect 194232 229628 194284 229634
rect 194232 229570 194284 229576
rect 194244 222086 194272 229570
rect 194704 229094 194732 231662
rect 195244 230036 195296 230042
rect 195244 229978 195296 229984
rect 195256 229498 195284 229978
rect 195244 229492 195296 229498
rect 195244 229434 195296 229440
rect 194612 229066 194732 229094
rect 195532 229094 195560 231676
rect 195888 229628 195940 229634
rect 195888 229570 195940 229576
rect 195532 229066 195652 229094
rect 194416 224936 194468 224942
rect 194416 224878 194468 224884
rect 194428 223990 194456 224878
rect 194416 223984 194468 223990
rect 194416 223926 194468 223932
rect 194612 222358 194640 229066
rect 195072 226358 195468 226386
rect 195072 226302 195100 226358
rect 195060 226296 195112 226302
rect 195060 226238 195112 226244
rect 195244 226296 195296 226302
rect 195244 226238 195296 226244
rect 195256 225214 195284 226238
rect 195440 225214 195468 226358
rect 195244 225208 195296 225214
rect 195244 225150 195296 225156
rect 195428 225208 195480 225214
rect 195428 225150 195480 225156
rect 194876 224936 194928 224942
rect 194876 224878 194928 224884
rect 194888 224670 194916 224878
rect 194876 224664 194928 224670
rect 194876 224606 194928 224612
rect 194968 222488 195020 222494
rect 194968 222430 195020 222436
rect 194600 222352 194652 222358
rect 194600 222294 194652 222300
rect 194232 222080 194284 222086
rect 194232 222022 194284 222028
rect 194416 222012 194468 222018
rect 194416 221954 194468 221960
rect 194046 220688 194102 220697
rect 193036 220652 193088 220658
rect 194046 220623 194102 220632
rect 193036 220594 193088 220600
rect 193048 219570 193076 220594
rect 193036 219564 193088 219570
rect 193036 219506 193088 219512
rect 194428 219434 194456 221954
rect 194980 220794 195008 222430
rect 195624 222358 195652 229066
rect 195900 228274 195928 229570
rect 196084 229537 196112 231676
rect 196360 231662 196650 231690
rect 196912 231662 197202 231690
rect 196070 229528 196126 229537
rect 196070 229463 196126 229472
rect 195888 228268 195940 228274
rect 195888 228210 195940 228216
rect 195612 222352 195664 222358
rect 195612 222294 195664 222300
rect 195152 222148 195204 222154
rect 195152 222090 195204 222096
rect 195164 220930 195192 222090
rect 196360 221241 196388 231662
rect 196912 223854 196940 231662
rect 197740 227730 197768 231676
rect 197728 227724 197780 227730
rect 197728 227666 197780 227672
rect 197452 227180 197504 227186
rect 197452 227122 197504 227128
rect 197268 224664 197320 224670
rect 197268 224606 197320 224612
rect 196900 223848 196952 223854
rect 196900 223790 196952 223796
rect 196346 221232 196402 221241
rect 196346 221167 196402 221176
rect 195152 220924 195204 220930
rect 195152 220866 195204 220872
rect 195336 220924 195388 220930
rect 195336 220866 195388 220872
rect 194968 220788 195020 220794
rect 194968 220730 195020 220736
rect 195152 220788 195204 220794
rect 195152 220730 195204 220736
rect 194244 219406 194456 219434
rect 194244 217410 194272 219406
rect 195164 217410 195192 220730
rect 195348 219842 195376 220866
rect 195336 219836 195388 219842
rect 195336 219778 195388 219784
rect 195888 219836 195940 219842
rect 195888 219778 195940 219784
rect 195900 217410 195928 219778
rect 196716 219428 196768 219434
rect 196716 219370 196768 219376
rect 196728 217410 196756 219370
rect 197280 217410 197308 224606
rect 197464 219842 197492 227122
rect 198292 224942 198320 231676
rect 198858 231662 199056 231690
rect 198280 224936 198332 224942
rect 198280 224878 198332 224884
rect 198464 224936 198516 224942
rect 198464 224878 198516 224884
rect 197452 219836 197504 219842
rect 197452 219778 197504 219784
rect 198476 217410 198504 224878
rect 199028 218618 199056 231662
rect 199212 231662 199410 231690
rect 199672 231662 199962 231690
rect 199212 224233 199240 231662
rect 199384 227724 199436 227730
rect 199384 227666 199436 227672
rect 199198 224224 199254 224233
rect 199198 224159 199254 224168
rect 199396 223530 199424 227666
rect 199672 226642 199700 231662
rect 200500 229362 200528 231676
rect 200684 231662 201066 231690
rect 200488 229356 200540 229362
rect 200488 229298 200540 229304
rect 199660 226636 199712 226642
rect 199660 226578 199712 226584
rect 199212 223502 199424 223530
rect 199016 218612 199068 218618
rect 199016 218554 199068 218560
rect 199212 217410 199240 223502
rect 200118 222048 200174 222057
rect 200118 221983 200174 221992
rect 200132 221626 200160 221983
rect 200086 221610 200160 221626
rect 200074 221604 200160 221610
rect 200126 221598 200160 221604
rect 200304 221604 200356 221610
rect 200074 221546 200126 221552
rect 200304 221546 200356 221552
rect 200316 221105 200344 221546
rect 199474 221096 199530 221105
rect 199474 221031 199530 221040
rect 200302 221096 200358 221105
rect 200302 221031 200358 221040
rect 199488 220930 199516 221031
rect 199476 220924 199528 220930
rect 199476 220866 199528 220872
rect 199844 220856 199896 220862
rect 199658 220824 199714 220833
rect 199844 220798 199896 220804
rect 199658 220759 199660 220768
rect 199712 220759 199714 220768
rect 199660 220730 199712 220736
rect 199856 217410 199884 220798
rect 200684 219434 200712 231662
rect 200856 229220 200908 229226
rect 200856 229162 200908 229168
rect 200868 229094 200896 229162
rect 200868 229066 201080 229094
rect 200856 223848 200908 223854
rect 200856 223790 200908 223796
rect 200408 219406 200712 219434
rect 200408 218482 200436 219406
rect 200396 218476 200448 218482
rect 200396 218418 200448 218424
rect 200868 217410 200896 223790
rect 201052 220862 201080 229066
rect 201604 222290 201632 231676
rect 201788 231662 202170 231690
rect 202340 231662 202722 231690
rect 201788 226302 201816 231662
rect 201960 226364 202012 226370
rect 201960 226306 202012 226312
rect 201776 226296 201828 226302
rect 201776 226238 201828 226244
rect 201592 222284 201644 222290
rect 201592 222226 201644 222232
rect 201224 222148 201276 222154
rect 201224 222090 201276 222096
rect 201040 220856 201092 220862
rect 201040 220798 201092 220804
rect 192864 217382 193108 217410
rect 193936 217382 194272 217410
rect 194764 217382 195192 217410
rect 195592 217382 195928 217410
rect 196420 217382 196756 217410
rect 197248 217382 197308 217410
rect 198076 217382 198504 217410
rect 198904 217382 199240 217410
rect 199732 217382 199884 217410
rect 200560 217382 200896 217410
rect 201236 217410 201264 222090
rect 201972 220833 202000 226306
rect 202340 221610 202368 231662
rect 203260 230314 203288 231676
rect 203248 230308 203300 230314
rect 203248 230250 203300 230256
rect 202788 229628 202840 229634
rect 202788 229570 202840 229576
rect 202602 229392 202658 229401
rect 202800 229362 202828 229570
rect 203524 229492 203576 229498
rect 203524 229434 203576 229440
rect 202602 229327 202604 229336
rect 202656 229327 202658 229336
rect 202788 229356 202840 229362
rect 202604 229298 202656 229304
rect 202788 229298 202840 229304
rect 203536 229094 203564 229434
rect 203536 229066 203656 229094
rect 202328 221604 202380 221610
rect 202328 221546 202380 221552
rect 201958 220824 202014 220833
rect 201958 220759 202014 220768
rect 203432 220788 203484 220794
rect 203432 220730 203484 220736
rect 201592 219836 201644 219842
rect 201592 219778 201644 219784
rect 201604 219434 201632 219778
rect 202326 219736 202382 219745
rect 202326 219671 202328 219680
rect 202380 219671 202382 219680
rect 202512 219700 202564 219706
rect 202328 219642 202380 219648
rect 202512 219642 202564 219648
rect 201592 219428 201644 219434
rect 201592 219370 201644 219376
rect 202524 217410 202552 219642
rect 203444 217410 203472 220730
rect 203628 220522 203656 229066
rect 203812 223718 203840 231676
rect 204364 226506 204392 231676
rect 204548 231662 204930 231690
rect 205284 231662 205482 231690
rect 205836 231662 206034 231690
rect 204548 229401 204576 231662
rect 204720 230580 204772 230586
rect 204720 230522 204772 230528
rect 204732 230178 204760 230522
rect 205088 230308 205140 230314
rect 205088 230250 205140 230256
rect 204720 230172 204772 230178
rect 204720 230114 204772 230120
rect 205100 229634 205128 230250
rect 205088 229628 205140 229634
rect 205088 229570 205140 229576
rect 204534 229392 204590 229401
rect 205284 229362 205312 231662
rect 205456 230444 205508 230450
rect 205456 230386 205508 230392
rect 205468 229634 205496 230386
rect 205456 229628 205508 229634
rect 205456 229570 205508 229576
rect 204534 229327 204590 229336
rect 205272 229356 205324 229362
rect 205272 229298 205324 229304
rect 205548 229356 205600 229362
rect 205548 229298 205600 229304
rect 205560 228002 205588 229298
rect 205836 229094 205864 231662
rect 206008 230444 206060 230450
rect 206008 230386 206060 230392
rect 206020 229226 206048 230386
rect 206008 229220 206060 229226
rect 206008 229162 206060 229168
rect 205836 229066 205956 229094
rect 205548 227996 205600 228002
rect 205548 227938 205600 227944
rect 204536 227860 204588 227866
rect 204536 227802 204588 227808
rect 204352 226500 204404 226506
rect 204352 226442 204404 226448
rect 204548 224754 204576 227802
rect 204904 227180 204956 227186
rect 204904 227122 204956 227128
rect 205088 227180 205140 227186
rect 205088 227122 205140 227128
rect 204916 226914 204944 227122
rect 204904 226908 204956 226914
rect 204904 226850 204956 226856
rect 205100 226778 205128 227122
rect 205088 226772 205140 226778
rect 205088 226714 205140 226720
rect 205640 226772 205692 226778
rect 205640 226714 205692 226720
rect 205456 226296 205508 226302
rect 205456 226238 205508 226244
rect 204364 224726 204576 224754
rect 203800 223712 203852 223718
rect 203800 223654 203852 223660
rect 204168 220924 204220 220930
rect 204168 220866 204220 220872
rect 203616 220516 203668 220522
rect 203616 220458 203668 220464
rect 204180 217410 204208 220866
rect 204364 220153 204392 224726
rect 204536 224664 204588 224670
rect 204536 224606 204588 224612
rect 204720 224664 204772 224670
rect 204720 224606 204772 224612
rect 204548 223854 204576 224606
rect 204732 224262 204760 224606
rect 204720 224256 204772 224262
rect 204720 224198 204772 224204
rect 204904 224256 204956 224262
rect 204904 224198 204956 224204
rect 204916 223990 204944 224198
rect 204904 223984 204956 223990
rect 204904 223926 204956 223932
rect 204536 223848 204588 223854
rect 204536 223790 204588 223796
rect 204720 221604 204772 221610
rect 204720 221546 204772 221552
rect 204732 221338 204760 221546
rect 204720 221332 204772 221338
rect 204720 221274 204772 221280
rect 205272 220788 205324 220794
rect 205272 220730 205324 220736
rect 205088 220244 205140 220250
rect 205088 220186 205140 220192
rect 204350 220144 204406 220153
rect 204350 220079 204406 220088
rect 204628 220108 204680 220114
rect 204628 220050 204680 220056
rect 204640 219434 204668 220050
rect 205100 219842 205128 220186
rect 205088 219836 205140 219842
rect 205088 219778 205140 219784
rect 205284 219706 205312 220730
rect 205272 219700 205324 219706
rect 205272 219642 205324 219648
rect 204994 219464 205050 219473
rect 204628 219428 204680 219434
rect 204994 219399 205050 219408
rect 204628 219370 204680 219376
rect 205008 217410 205036 219399
rect 201236 217382 201388 217410
rect 202216 217382 202552 217410
rect 203044 217382 203472 217410
rect 203872 217382 204208 217410
rect 204700 217382 205036 217410
rect 205468 217410 205496 226238
rect 205652 219473 205680 226714
rect 205928 222057 205956 229066
rect 206572 226642 206600 231676
rect 207124 229094 207152 231676
rect 207676 229094 207704 231676
rect 207952 231662 208242 231690
rect 207124 229066 207428 229094
rect 207676 229066 207796 229094
rect 206560 226636 206612 226642
rect 206560 226578 206612 226584
rect 206836 224392 206888 224398
rect 206834 224360 206836 224369
rect 207020 224392 207072 224398
rect 206888 224360 206890 224369
rect 207020 224334 207072 224340
rect 206834 224295 206890 224304
rect 205914 222048 205970 222057
rect 205914 221983 205970 221992
rect 206652 219836 206704 219842
rect 206652 219778 206704 219784
rect 205914 219736 205970 219745
rect 205914 219671 205916 219680
rect 205968 219671 205970 219680
rect 205916 219642 205968 219648
rect 205638 219464 205694 219473
rect 205638 219399 205694 219408
rect 206664 217410 206692 219778
rect 207032 218210 207060 224334
rect 207204 222488 207256 222494
rect 207204 222430 207256 222436
rect 207216 219706 207244 222430
rect 207400 222358 207428 229066
rect 207388 222352 207440 222358
rect 207388 222294 207440 222300
rect 207480 221196 207532 221202
rect 207480 221138 207532 221144
rect 207204 219700 207256 219706
rect 207204 219642 207256 219648
rect 207020 218204 207072 218210
rect 207020 218146 207072 218152
rect 207492 217410 207520 221138
rect 207768 218346 207796 229066
rect 207952 224398 207980 231662
rect 207940 224392 207992 224398
rect 208780 224369 208808 231676
rect 209332 229634 209360 231676
rect 209792 231662 209898 231690
rect 210160 231662 210450 231690
rect 210712 231662 211002 231690
rect 209320 229628 209372 229634
rect 209320 229570 209372 229576
rect 209792 229106 209820 231662
rect 209700 229078 209820 229106
rect 209700 228138 209728 229078
rect 209688 228132 209740 228138
rect 209688 228074 209740 228080
rect 208952 227996 209004 228002
rect 208952 227938 209004 227944
rect 207940 224334 207992 224340
rect 208766 224360 208822 224369
rect 208766 224295 208822 224304
rect 208400 223712 208452 223718
rect 208400 223654 208452 223660
rect 208412 219434 208440 223654
rect 208964 219434 208992 227938
rect 210160 221066 210188 231662
rect 210712 224670 210740 231662
rect 211160 229220 211212 229226
rect 211160 229162 211212 229168
rect 211172 228546 211200 229162
rect 211160 228540 211212 228546
rect 211160 228482 211212 228488
rect 211540 227866 211568 231676
rect 211712 229628 211764 229634
rect 211712 229570 211764 229576
rect 211528 227860 211580 227866
rect 211528 227802 211580 227808
rect 210700 224664 210752 224670
rect 210700 224606 210752 224612
rect 210884 224664 210936 224670
rect 210884 224606 210936 224612
rect 210424 224392 210476 224398
rect 210424 224334 210476 224340
rect 210148 221060 210200 221066
rect 210148 221002 210200 221008
rect 209686 219872 209742 219881
rect 209686 219807 209688 219816
rect 209740 219807 209742 219816
rect 209870 219872 209926 219881
rect 209870 219807 209872 219816
rect 209688 219778 209740 219784
rect 209924 219807 209926 219816
rect 209872 219778 209924 219784
rect 209688 219700 209740 219706
rect 209688 219642 209740 219648
rect 208320 219406 208440 219434
rect 208872 219406 208992 219434
rect 207756 218340 207808 218346
rect 207756 218282 207808 218288
rect 208320 217410 208348 219406
rect 208872 217410 208900 219406
rect 209700 217410 209728 219642
rect 210436 219434 210464 224334
rect 210424 219428 210476 219434
rect 210424 219370 210476 219376
rect 210896 217410 210924 224606
rect 211724 219994 211752 229570
rect 212092 224398 212120 231676
rect 212264 228540 212316 228546
rect 212264 228482 212316 228488
rect 212276 225570 212304 228482
rect 212644 227186 212672 231676
rect 212632 227180 212684 227186
rect 212632 227122 212684 227128
rect 213196 225622 213224 231676
rect 213380 231662 213762 231690
rect 213380 229770 213408 231662
rect 214104 229900 214156 229906
rect 214104 229842 214156 229848
rect 213368 229764 213420 229770
rect 213368 229706 213420 229712
rect 213552 229764 213604 229770
rect 213552 229706 213604 229712
rect 212184 225542 212304 225570
rect 213184 225616 213236 225622
rect 213184 225558 213236 225564
rect 212184 224482 212212 225542
rect 212356 225480 212408 225486
rect 212356 225422 212408 225428
rect 212540 225480 212592 225486
rect 212540 225422 212592 225428
rect 212368 225321 212396 225422
rect 212354 225312 212410 225321
rect 212354 225247 212410 225256
rect 212552 225078 212580 225422
rect 212540 225072 212592 225078
rect 212540 225014 212592 225020
rect 212184 224454 212488 224482
rect 212080 224392 212132 224398
rect 212080 224334 212132 224340
rect 211448 219966 211752 219994
rect 211448 219842 211476 219966
rect 211436 219836 211488 219842
rect 211436 219778 211488 219784
rect 211620 219836 211672 219842
rect 211620 219778 211672 219784
rect 211632 217410 211660 219778
rect 212460 217410 212488 224454
rect 213366 222864 213422 222873
rect 213366 222799 213422 222808
rect 213380 222630 213408 222799
rect 213368 222624 213420 222630
rect 213368 222566 213420 222572
rect 213276 221468 213328 221474
rect 213276 221410 213328 221416
rect 213288 221066 213316 221410
rect 213276 221060 213328 221066
rect 213276 221002 213328 221008
rect 213564 219434 213592 229706
rect 214116 229537 214144 229842
rect 214102 229528 214158 229537
rect 214102 229463 214158 229472
rect 214300 229362 214328 231676
rect 214472 229900 214524 229906
rect 214472 229842 214524 229848
rect 214288 229356 214340 229362
rect 214288 229298 214340 229304
rect 214484 228410 214512 229842
rect 214654 229528 214710 229537
rect 214654 229463 214710 229472
rect 214668 229362 214696 229463
rect 214656 229356 214708 229362
rect 214656 229298 214708 229304
rect 214852 229094 214880 231676
rect 214852 229066 215248 229094
rect 214472 228404 214524 228410
rect 214472 228346 214524 228352
rect 214932 228404 214984 228410
rect 214932 228346 214984 228352
rect 214380 225752 214432 225758
rect 214380 225694 214432 225700
rect 214564 225752 214616 225758
rect 214564 225694 214616 225700
rect 214196 225616 214248 225622
rect 214196 225558 214248 225564
rect 214208 225350 214236 225558
rect 214196 225344 214248 225350
rect 214196 225286 214248 225292
rect 214392 225078 214420 225694
rect 214576 225214 214604 225694
rect 214748 225344 214800 225350
rect 214746 225312 214748 225321
rect 214800 225312 214802 225321
rect 214944 225298 214972 228346
rect 214944 225270 215064 225298
rect 214746 225247 214802 225256
rect 214564 225208 214616 225214
rect 214564 225150 214616 225156
rect 214380 225072 214432 225078
rect 214380 225014 214432 225020
rect 214378 224904 214434 224913
rect 214378 224839 214434 224848
rect 213736 222624 213788 222630
rect 213736 222566 213788 222572
rect 213380 219406 213592 219434
rect 213380 217410 213408 219406
rect 205468 217382 205528 217410
rect 206356 217382 206692 217410
rect 207184 217382 207520 217410
rect 208012 217382 208348 217410
rect 208840 217382 208900 217410
rect 209668 217382 209728 217410
rect 210496 217382 210924 217410
rect 211324 217382 211660 217410
rect 212152 217382 212488 217410
rect 212980 217382 213408 217410
rect 213748 217410 213776 222566
rect 214392 219842 214420 224839
rect 214564 224392 214616 224398
rect 214564 224334 214616 224340
rect 214576 223718 214604 224334
rect 214564 223712 214616 223718
rect 214564 223654 214616 223660
rect 214564 223032 214616 223038
rect 214564 222974 214616 222980
rect 214748 223032 214800 223038
rect 214748 222974 214800 222980
rect 214576 222358 214604 222974
rect 214760 222873 214788 222974
rect 214746 222864 214802 222873
rect 214746 222799 214802 222808
rect 214564 222352 214616 222358
rect 214564 222294 214616 222300
rect 214748 221332 214800 221338
rect 214748 221274 214800 221280
rect 214760 220930 214788 221274
rect 214748 220924 214800 220930
rect 214748 220866 214800 220872
rect 214564 220652 214616 220658
rect 214564 220594 214616 220600
rect 214576 219842 214604 220594
rect 214380 219836 214432 219842
rect 214380 219778 214432 219784
rect 214564 219836 214616 219842
rect 214564 219778 214616 219784
rect 215036 217410 215064 225270
rect 215220 222902 215248 229066
rect 215404 225486 215432 231676
rect 215392 225480 215444 225486
rect 215392 225422 215444 225428
rect 215576 225480 215628 225486
rect 215576 225422 215628 225428
rect 215588 224913 215616 225422
rect 215760 225208 215812 225214
rect 215760 225150 215812 225156
rect 215574 224904 215630 224913
rect 215574 224839 215630 224848
rect 215208 222896 215260 222902
rect 215208 222838 215260 222844
rect 215772 217410 215800 225150
rect 215956 222494 215984 231676
rect 216508 229906 216536 231676
rect 216876 231662 217074 231690
rect 216496 229900 216548 229906
rect 216496 229842 216548 229848
rect 215944 222488 215996 222494
rect 215944 222430 215996 222436
rect 216876 221066 216904 231662
rect 217612 225350 217640 231676
rect 218164 229362 218192 231676
rect 218152 229356 218204 229362
rect 218152 229298 218204 229304
rect 217600 225344 217652 225350
rect 217600 225286 217652 225292
rect 218716 224534 218744 231676
rect 218992 231662 219282 231690
rect 218704 224528 218756 224534
rect 218704 224470 218756 224476
rect 218992 223038 219020 231662
rect 219820 225894 219848 231676
rect 220004 231662 220386 231690
rect 220004 229094 220032 231662
rect 220452 229900 220504 229906
rect 220452 229842 220504 229848
rect 220004 229066 220124 229094
rect 219808 225888 219860 225894
rect 219808 225830 219860 225836
rect 219164 225480 219216 225486
rect 219164 225422 219216 225428
rect 218980 223032 219032 223038
rect 218980 222974 219032 222980
rect 218060 222896 218112 222902
rect 218060 222838 218112 222844
rect 216864 221060 216916 221066
rect 216864 221002 216916 221008
rect 217416 221060 217468 221066
rect 217416 221002 217468 221008
rect 216312 220652 216364 220658
rect 216312 220594 216364 220600
rect 216324 217410 216352 220594
rect 217428 217410 217456 221002
rect 218072 219434 218100 222838
rect 217980 219406 218100 219434
rect 217980 217410 218008 219406
rect 219176 217410 219204 225422
rect 219716 220652 219768 220658
rect 219716 220594 219768 220600
rect 219900 220652 219952 220658
rect 219900 220594 219952 220600
rect 219728 220386 219756 220594
rect 219532 220380 219584 220386
rect 219532 220322 219584 220328
rect 219716 220380 219768 220386
rect 219716 220322 219768 220328
rect 219346 220144 219402 220153
rect 219544 220114 219572 220322
rect 219346 220079 219348 220088
rect 219400 220079 219402 220088
rect 219532 220108 219584 220114
rect 219348 220050 219400 220056
rect 219532 220050 219584 220056
rect 219912 217410 219940 220594
rect 220096 220153 220124 229066
rect 220464 220658 220492 229842
rect 220924 229362 220952 231676
rect 220912 229356 220964 229362
rect 220912 229298 220964 229304
rect 220820 229220 220872 229226
rect 220820 229162 220872 229168
rect 220832 228818 220860 229162
rect 220820 228812 220872 228818
rect 220820 228754 220872 228760
rect 221476 225078 221504 231676
rect 221752 231662 222042 231690
rect 221464 225072 221516 225078
rect 221464 225014 221516 225020
rect 220636 222488 220688 222494
rect 220636 222430 220688 222436
rect 220452 220652 220504 220658
rect 220452 220594 220504 220600
rect 220082 220144 220138 220153
rect 220082 220079 220138 220088
rect 220648 217410 220676 222430
rect 221752 222358 221780 231662
rect 222580 229498 222608 231676
rect 222568 229492 222620 229498
rect 222568 229434 222620 229440
rect 222200 229356 222252 229362
rect 222200 229298 222252 229304
rect 222212 229090 222240 229298
rect 222200 229084 222252 229090
rect 222200 229026 222252 229032
rect 222108 228812 222160 228818
rect 222108 228754 222160 228760
rect 221740 222352 221792 222358
rect 221740 222294 221792 222300
rect 221556 220652 221608 220658
rect 221556 220594 221608 220600
rect 221568 217410 221596 220594
rect 222120 217410 222148 228754
rect 222292 225072 222344 225078
rect 222292 225014 222344 225020
rect 222304 220658 222332 225014
rect 223132 223446 223160 231676
rect 223120 223440 223172 223446
rect 223120 223382 223172 223388
rect 223684 223310 223712 231676
rect 224236 226166 224264 231676
rect 224420 231662 224802 231690
rect 224224 226160 224276 226166
rect 224224 226102 224276 226108
rect 224224 225888 224276 225894
rect 224224 225830 224276 225836
rect 224236 225622 224264 225830
rect 224224 225616 224276 225622
rect 224224 225558 224276 225564
rect 224420 224652 224448 231662
rect 225340 229226 225368 231676
rect 225524 231662 225906 231690
rect 225328 229220 225380 229226
rect 225328 229162 225380 229168
rect 223868 224624 224448 224652
rect 223672 223304 223724 223310
rect 223672 223246 223724 223252
rect 223868 220658 223896 224624
rect 224224 223168 224276 223174
rect 224224 223110 224276 223116
rect 222292 220652 222344 220658
rect 222292 220594 222344 220600
rect 222476 220652 222528 220658
rect 222476 220594 222528 220600
rect 223856 220652 223908 220658
rect 223856 220594 223908 220600
rect 224040 220652 224092 220658
rect 224040 220594 224092 220600
rect 222488 220114 222516 220594
rect 224052 220386 224080 220594
rect 224040 220380 224092 220386
rect 224040 220322 224092 220328
rect 222476 220108 222528 220114
rect 222476 220050 222528 220056
rect 223212 220108 223264 220114
rect 223212 220050 223264 220056
rect 223224 217410 223252 220050
rect 224236 219434 224264 223110
rect 225524 221746 225552 231662
rect 225696 226160 225748 226166
rect 225696 226102 225748 226108
rect 225512 221740 225564 221746
rect 225512 221682 225564 221688
rect 224500 220652 224552 220658
rect 224500 220594 224552 220600
rect 224512 220114 224540 220594
rect 224500 220108 224552 220114
rect 224500 220050 224552 220056
rect 224684 220108 224736 220114
rect 224684 220050 224736 220056
rect 224052 219406 224264 219434
rect 224052 217410 224080 219406
rect 224696 217410 224724 220050
rect 225708 217410 225736 226102
rect 226444 226030 226472 231676
rect 226616 228132 226668 228138
rect 226616 228074 226668 228080
rect 226432 226024 226484 226030
rect 226432 225966 226484 225972
rect 226064 223440 226116 223446
rect 226064 223382 226116 223388
rect 213748 217382 213808 217410
rect 214636 217382 215064 217410
rect 215464 217382 215800 217410
rect 216292 217382 216352 217410
rect 217120 217382 217456 217410
rect 217948 217382 218008 217410
rect 218776 217382 219204 217410
rect 219604 217382 219940 217410
rect 220432 217382 220676 217410
rect 221260 217382 221596 217410
rect 222088 217382 222148 217410
rect 222916 217382 223252 217410
rect 223744 217382 224080 217410
rect 224572 217382 224724 217410
rect 225400 217382 225736 217410
rect 226076 217410 226104 223382
rect 226628 220114 226656 228074
rect 226996 225758 227024 231676
rect 227352 229492 227404 229498
rect 227352 229434 227404 229440
rect 226984 225752 227036 225758
rect 226984 225694 227036 225700
rect 227168 225752 227220 225758
rect 227168 225694 227220 225700
rect 227180 225078 227208 225694
rect 227168 225072 227220 225078
rect 227168 225014 227220 225020
rect 227364 223446 227392 229434
rect 227548 229362 227576 231676
rect 227916 231662 228114 231690
rect 227536 229356 227588 229362
rect 227536 229298 227588 229304
rect 227352 223440 227404 223446
rect 227352 223382 227404 223388
rect 227628 223440 227680 223446
rect 227628 223382 227680 223388
rect 227444 223304 227496 223310
rect 227444 223246 227496 223252
rect 226616 220108 226668 220114
rect 226616 220050 226668 220056
rect 227456 217410 227484 223246
rect 227640 223174 227668 223382
rect 227628 223168 227680 223174
rect 227628 223110 227680 223116
rect 227916 221610 227944 231662
rect 228652 223174 228680 231676
rect 229218 231662 229508 231690
rect 229192 229356 229244 229362
rect 229192 229298 229244 229304
rect 229008 228948 229060 228954
rect 229008 228890 229060 228896
rect 228640 223168 228692 223174
rect 228640 223110 228692 223116
rect 228180 223032 228232 223038
rect 228180 222974 228232 222980
rect 227904 221604 227956 221610
rect 227904 221546 227956 221552
rect 228192 217410 228220 222974
rect 229020 217410 229048 228890
rect 229204 224670 229232 229298
rect 229192 224664 229244 224670
rect 229192 224606 229244 224612
rect 229480 220386 229508 231662
rect 229756 229158 229784 231676
rect 229744 229152 229796 229158
rect 229744 229094 229796 229100
rect 230308 223582 230336 231676
rect 230860 225894 230888 231676
rect 231412 230042 231440 231676
rect 231400 230036 231452 230042
rect 231400 229978 231452 229984
rect 231964 227050 231992 231676
rect 232240 231662 232530 231690
rect 232240 229094 232268 231662
rect 232148 229066 232268 229094
rect 231952 227044 232004 227050
rect 231952 226986 232004 226992
rect 230848 225888 230900 225894
rect 230848 225830 230900 225836
rect 231676 225072 231728 225078
rect 231676 225014 231728 225020
rect 230296 223576 230348 223582
rect 230296 223518 230348 223524
rect 230388 221604 230440 221610
rect 230388 221546 230440 221552
rect 229468 220380 229520 220386
rect 229468 220322 229520 220328
rect 229836 219972 229888 219978
rect 229836 219914 229888 219920
rect 229848 217410 229876 219914
rect 230400 217410 230428 221546
rect 231492 220380 231544 220386
rect 231492 220322 231544 220328
rect 231504 217410 231532 220322
rect 231688 219502 231716 225014
rect 231860 224664 231912 224670
rect 231860 224606 231912 224612
rect 231872 224126 231900 224606
rect 231860 224120 231912 224126
rect 231860 224062 231912 224068
rect 231860 221740 231912 221746
rect 231860 221682 231912 221688
rect 231872 220114 231900 221682
rect 232148 221474 232176 229066
rect 233068 228682 233096 231676
rect 233436 231662 233634 231690
rect 233056 228676 233108 228682
rect 233056 228618 233108 228624
rect 232320 224528 232372 224534
rect 232320 224470 232372 224476
rect 232136 221468 232188 221474
rect 232136 221410 232188 221416
rect 231860 220108 231912 220114
rect 231860 220050 231912 220056
rect 231676 219496 231728 219502
rect 231676 219438 231728 219444
rect 232332 217410 232360 224470
rect 233436 221746 233464 231662
rect 233884 229220 233936 229226
rect 233884 229162 233936 229168
rect 233700 229084 233752 229090
rect 233700 229026 233752 229032
rect 233712 228138 233740 229026
rect 233700 228132 233752 228138
rect 233700 228074 233752 228080
rect 233424 221740 233476 221746
rect 233424 221682 233476 221688
rect 233700 221740 233752 221746
rect 233700 221682 233752 221688
rect 232688 220652 232740 220658
rect 232688 220594 232740 220600
rect 232872 220652 232924 220658
rect 232872 220594 232924 220600
rect 232700 220114 232728 220594
rect 232688 220108 232740 220114
rect 232688 220050 232740 220056
rect 232884 217410 232912 220594
rect 233712 217410 233740 221682
rect 233896 220658 233924 229162
rect 234172 227322 234200 231676
rect 234160 227316 234212 227322
rect 234160 227258 234212 227264
rect 234724 224806 234752 231676
rect 235000 231662 235290 231690
rect 234712 224800 234764 224806
rect 234712 224742 234764 224748
rect 234620 224256 234672 224262
rect 234620 224198 234672 224204
rect 233884 220652 233936 220658
rect 233884 220594 233936 220600
rect 234632 219434 234660 224198
rect 235000 224126 235028 231662
rect 235828 230178 235856 231676
rect 235816 230172 235868 230178
rect 235816 230114 235868 230120
rect 236000 230172 236052 230178
rect 236000 230114 236052 230120
rect 236012 227594 236040 230114
rect 236000 227588 236052 227594
rect 236000 227530 236052 227536
rect 236380 227458 236408 231676
rect 236368 227452 236420 227458
rect 236368 227394 236420 227400
rect 236000 227316 236052 227322
rect 236000 227258 236052 227264
rect 235724 227180 235776 227186
rect 235724 227122 235776 227128
rect 234988 224120 235040 224126
rect 234988 224062 235040 224068
rect 234540 219406 234660 219434
rect 234540 217410 234568 219406
rect 235736 217410 235764 227122
rect 236012 220386 236040 227258
rect 236932 224670 236960 231676
rect 237288 227044 237340 227050
rect 237288 226986 237340 226992
rect 236920 224664 236972 224670
rect 236920 224606 236972 224612
rect 236460 220652 236512 220658
rect 236460 220594 236512 220600
rect 236000 220380 236052 220386
rect 236000 220322 236052 220328
rect 236472 217410 236500 220594
rect 237300 217410 237328 226986
rect 237484 221882 237512 231676
rect 238036 225078 238064 231676
rect 238588 230178 238616 231676
rect 238956 231662 239154 231690
rect 238576 230172 238628 230178
rect 238576 230114 238628 230120
rect 238024 225072 238076 225078
rect 238024 225014 238076 225020
rect 238576 224664 238628 224670
rect 238576 224606 238628 224612
rect 237472 221876 237524 221882
rect 237472 221818 237524 221824
rect 238116 219496 238168 219502
rect 238116 219438 238168 219444
rect 238128 217410 238156 219438
rect 226076 217382 226228 217410
rect 227056 217382 227484 217410
rect 227884 217382 228220 217410
rect 228712 217382 229048 217410
rect 229540 217382 229876 217410
rect 230368 217382 230428 217410
rect 231196 217382 231532 217410
rect 232024 217382 232360 217410
rect 232852 217382 232912 217410
rect 233680 217382 233740 217410
rect 234508 217382 234568 217410
rect 235336 217382 235764 217410
rect 236164 217382 236500 217410
rect 236992 217382 237328 217410
rect 237820 217382 238156 217410
rect 238588 217410 238616 224606
rect 238956 222018 238984 231662
rect 239692 222766 239720 231676
rect 240244 230314 240272 231676
rect 240232 230308 240284 230314
rect 240232 230250 240284 230256
rect 240796 226914 240824 231676
rect 241164 231662 241362 231690
rect 240968 230172 241020 230178
rect 240968 230114 241020 230120
rect 240784 226908 240836 226914
rect 240784 226850 240836 226856
rect 240600 224800 240652 224806
rect 240600 224742 240652 224748
rect 239680 222760 239732 222766
rect 239680 222702 239732 222708
rect 238944 222012 238996 222018
rect 238944 221954 238996 221960
rect 240048 221468 240100 221474
rect 240048 221410 240100 221416
rect 239588 220788 239640 220794
rect 239588 220730 239640 220736
rect 239772 220788 239824 220794
rect 239772 220730 239824 220736
rect 239600 220386 239628 220730
rect 239588 220380 239640 220386
rect 239588 220322 239640 220328
rect 239784 217410 239812 220730
rect 240060 219502 240088 221410
rect 240048 219496 240100 219502
rect 240048 219438 240100 219444
rect 240612 217410 240640 224742
rect 240980 220794 241008 230114
rect 241164 223990 241192 231662
rect 241900 226642 241928 231676
rect 242084 231662 242466 231690
rect 241888 226636 241940 226642
rect 241888 226578 241940 226584
rect 241152 223984 241204 223990
rect 241152 223926 241204 223932
rect 240968 220788 241020 220794
rect 240968 220730 241020 220736
rect 241244 220788 241296 220794
rect 241244 220730 241296 220736
rect 241256 217410 241284 220730
rect 242084 220250 242112 231662
rect 243004 227730 243032 231676
rect 243188 231662 243570 231690
rect 243740 231662 244122 231690
rect 242992 227724 243044 227730
rect 242992 227666 243044 227672
rect 242256 227452 242308 227458
rect 242256 227394 242308 227400
rect 242072 220244 242124 220250
rect 242072 220186 242124 220192
rect 242268 217410 242296 227394
rect 243188 223854 243216 231662
rect 243544 230036 243596 230042
rect 243544 229978 243596 229984
rect 243556 229226 243584 229978
rect 243544 229220 243596 229226
rect 243544 229162 243596 229168
rect 243360 226432 243412 226438
rect 243360 226374 243412 226380
rect 243176 223848 243228 223854
rect 243176 223790 243228 223796
rect 242900 223644 242952 223650
rect 242900 223586 242952 223592
rect 242624 220380 242676 220386
rect 242624 220322 242676 220328
rect 238588 217382 238648 217410
rect 239476 217382 239812 217410
rect 240304 217382 240640 217410
rect 241132 217382 241284 217410
rect 241960 217382 242296 217410
rect 242636 217410 242664 220322
rect 242912 220250 242940 223586
rect 242900 220244 242952 220250
rect 242900 220186 242952 220192
rect 243372 219842 243400 226374
rect 243740 224942 243768 231662
rect 244660 230450 244688 231676
rect 244648 230444 244700 230450
rect 244648 230386 244700 230392
rect 243728 224936 243780 224942
rect 243728 224878 243780 224884
rect 244556 224936 244608 224942
rect 244556 224878 244608 224884
rect 243912 221876 243964 221882
rect 243912 221818 243964 221824
rect 243728 220652 243780 220658
rect 243728 220594 243780 220600
rect 243544 220244 243596 220250
rect 243544 220186 243596 220192
rect 243556 219978 243584 220186
rect 243740 219978 243768 220594
rect 243544 219972 243596 219978
rect 243544 219914 243596 219920
rect 243728 219972 243780 219978
rect 243728 219914 243780 219920
rect 243360 219836 243412 219842
rect 243360 219778 243412 219784
rect 243924 217410 243952 221818
rect 244568 220794 244596 224878
rect 245212 223650 245240 231676
rect 245476 228676 245528 228682
rect 245476 228618 245528 228624
rect 245200 223644 245252 223650
rect 245200 223586 245252 223592
rect 244556 220788 244608 220794
rect 244556 220730 244608 220736
rect 244740 220720 244792 220726
rect 244740 220662 244792 220668
rect 244752 217410 244780 220662
rect 245488 217410 245516 228618
rect 245764 221338 245792 231676
rect 245948 231662 246330 231690
rect 245948 222154 245976 231662
rect 246868 226438 246896 231676
rect 246856 226432 246908 226438
rect 246856 226374 246908 226380
rect 247420 226302 247448 231676
rect 247604 231662 247986 231690
rect 247408 226296 247460 226302
rect 247408 226238 247460 226244
rect 246764 225616 246816 225622
rect 246764 225558 246816 225564
rect 245936 222148 245988 222154
rect 245936 222090 245988 222096
rect 246396 222080 246448 222086
rect 246396 222022 246448 222028
rect 245752 221332 245804 221338
rect 245752 221274 245804 221280
rect 246408 217410 246436 222022
rect 242636 217382 242788 217410
rect 243616 217382 243952 217410
rect 244444 217382 244780 217410
rect 245272 217382 245516 217410
rect 246100 217382 246436 217410
rect 246776 217410 246804 225558
rect 247604 221202 247632 231662
rect 247776 230308 247828 230314
rect 247776 230250 247828 230256
rect 247788 222086 247816 230250
rect 248524 226846 248552 231676
rect 249076 229634 249104 231676
rect 249352 231662 249642 231690
rect 249064 229628 249116 229634
rect 249064 229570 249116 229576
rect 249352 228274 249380 231662
rect 250180 229362 250208 231676
rect 250168 229356 250220 229362
rect 250168 229298 250220 229304
rect 250444 229288 250496 229294
rect 250444 229230 250496 229236
rect 250456 229094 250484 229230
rect 250364 229066 250484 229094
rect 249340 228268 249392 228274
rect 249340 228210 249392 228216
rect 248880 228132 248932 228138
rect 248880 228074 248932 228080
rect 248512 226840 248564 226846
rect 248512 226782 248564 226788
rect 248144 222148 248196 222154
rect 248144 222090 248196 222096
rect 247776 222080 247828 222086
rect 247776 222022 247828 222028
rect 247960 222012 248012 222018
rect 247960 221954 248012 221960
rect 247592 221196 247644 221202
rect 247592 221138 247644 221144
rect 247972 220726 248000 221954
rect 247960 220720 248012 220726
rect 247960 220662 248012 220668
rect 248156 219706 248184 222090
rect 248144 219700 248196 219706
rect 248144 219642 248196 219648
rect 248052 219496 248104 219502
rect 248052 219438 248104 219444
rect 248064 217410 248092 219438
rect 248892 217410 248920 228074
rect 249708 227588 249760 227594
rect 249708 227530 249760 227536
rect 249524 220652 249576 220658
rect 249524 220594 249576 220600
rect 249536 217410 249564 220594
rect 249720 219502 249748 227530
rect 250364 220522 250392 229066
rect 250732 224398 250760 231676
rect 250720 224392 250772 224398
rect 250720 224334 250772 224340
rect 250536 223576 250588 223582
rect 250536 223518 250588 223524
rect 250352 220516 250404 220522
rect 250352 220458 250404 220464
rect 249708 219496 249760 219502
rect 249708 219438 249760 219444
rect 250548 217410 250576 223518
rect 251284 222154 251312 231676
rect 251836 228546 251864 231676
rect 252112 231662 252402 231690
rect 251824 228540 251876 228546
rect 251824 228482 251876 228488
rect 252112 222630 252140 231662
rect 252744 225888 252796 225894
rect 252744 225830 252796 225836
rect 252284 223168 252336 223174
rect 252284 223110 252336 223116
rect 252100 222624 252152 222630
rect 252100 222566 252152 222572
rect 251272 222148 251324 222154
rect 251272 222090 251324 222096
rect 251088 220788 251140 220794
rect 251088 220730 251140 220736
rect 251100 217410 251128 220730
rect 252296 217410 252324 223110
rect 252756 220794 252784 225830
rect 252940 225350 252968 231676
rect 253492 229770 253520 231676
rect 253480 229764 253532 229770
rect 253480 229706 253532 229712
rect 253756 228540 253808 228546
rect 253756 228482 253808 228488
rect 252928 225344 252980 225350
rect 252928 225286 252980 225292
rect 252744 220788 252796 220794
rect 252744 220730 252796 220736
rect 253020 220788 253072 220794
rect 253020 220730 253072 220736
rect 252836 220516 252888 220522
rect 252836 220458 252888 220464
rect 252848 220250 252876 220458
rect 252836 220244 252888 220250
rect 252836 220186 252888 220192
rect 253032 217410 253060 220730
rect 253572 220516 253624 220522
rect 253572 220458 253624 220464
rect 253584 220114 253612 220458
rect 253572 220108 253624 220114
rect 253572 220050 253624 220056
rect 253768 217410 253796 228482
rect 254044 225214 254072 231676
rect 254320 231662 254610 231690
rect 254032 225208 254084 225214
rect 254032 225150 254084 225156
rect 254320 221066 254348 231662
rect 255148 228410 255176 231676
rect 255700 229294 255728 231676
rect 255976 231662 256266 231690
rect 255688 229288 255740 229294
rect 255688 229230 255740 229236
rect 255136 228404 255188 228410
rect 255136 228346 255188 228352
rect 255228 226024 255280 226030
rect 255228 225966 255280 225972
rect 254308 221060 254360 221066
rect 254308 221002 254360 221008
rect 254676 219700 254728 219706
rect 254676 219642 254728 219648
rect 254688 217410 254716 219642
rect 255240 217410 255268 225966
rect 255976 225486 256004 231662
rect 256332 230444 256384 230450
rect 256332 230386 256384 230392
rect 255964 225480 256016 225486
rect 255964 225422 256016 225428
rect 256344 220794 256372 230386
rect 256516 228404 256568 228410
rect 256516 228346 256568 228352
rect 256332 220788 256384 220794
rect 256332 220730 256384 220736
rect 256332 220516 256384 220522
rect 256332 220458 256384 220464
rect 256344 217410 256372 220458
rect 256528 219706 256556 228346
rect 256804 222494 256832 231676
rect 257356 222902 257384 231676
rect 257908 229906 257936 231676
rect 257896 229900 257948 229906
rect 257896 229842 257948 229848
rect 258460 228818 258488 231676
rect 258736 231662 259026 231690
rect 258736 229094 258764 231662
rect 259092 229764 259144 229770
rect 259092 229706 259144 229712
rect 258644 229066 258764 229094
rect 258448 228812 258500 228818
rect 258448 228754 258500 228760
rect 258644 223446 258672 229066
rect 258632 223440 258684 223446
rect 258632 223382 258684 223388
rect 258816 223440 258868 223446
rect 258816 223382 258868 223388
rect 257344 222896 257396 222902
rect 257344 222838 257396 222844
rect 257988 222896 258040 222902
rect 257988 222838 258040 222844
rect 256792 222488 256844 222494
rect 256792 222430 256844 222436
rect 257160 221332 257212 221338
rect 257160 221274 257212 221280
rect 256516 219700 256568 219706
rect 256516 219642 256568 219648
rect 257172 217410 257200 221274
rect 258000 217410 258028 222838
rect 258828 217410 258856 223382
rect 246776 217382 246928 217410
rect 247756 217382 248092 217410
rect 248584 217382 248920 217410
rect 249412 217382 249564 217410
rect 250240 217382 250576 217410
rect 251068 217382 251128 217410
rect 251896 217382 252324 217410
rect 252724 217382 253060 217410
rect 253552 217382 253796 217410
rect 254380 217382 254716 217410
rect 255208 217382 255268 217410
rect 256036 217382 256372 217410
rect 256864 217382 257200 217410
rect 257692 217382 258028 217410
rect 258520 217382 258856 217410
rect 259104 217410 259132 229706
rect 259564 225758 259592 231676
rect 259840 231662 260130 231690
rect 259552 225752 259604 225758
rect 259552 225694 259604 225700
rect 259840 220250 259868 231662
rect 260668 226166 260696 231676
rect 261220 229094 261248 231676
rect 261128 229066 261248 229094
rect 261772 229090 261800 231676
rect 262324 229498 262352 231676
rect 262312 229492 262364 229498
rect 262312 229434 262364 229440
rect 261760 229084 261812 229090
rect 260656 226160 260708 226166
rect 260656 226102 260708 226108
rect 260564 225752 260616 225758
rect 260564 225694 260616 225700
rect 259828 220244 259880 220250
rect 259828 220186 259880 220192
rect 260576 217410 260604 225694
rect 261128 223310 261156 229066
rect 261760 229026 261812 229032
rect 262876 228954 262904 231676
rect 263152 231662 263442 231690
rect 262864 228948 262916 228954
rect 262864 228890 262916 228896
rect 262128 227792 262180 227798
rect 262128 227734 262180 227740
rect 261116 223304 261168 223310
rect 261116 223246 261168 223252
rect 261300 223304 261352 223310
rect 261300 223246 261352 223252
rect 261312 217410 261340 223246
rect 261668 222148 261720 222154
rect 261668 222090 261720 222096
rect 261680 221746 261708 222090
rect 261668 221740 261720 221746
rect 261668 221682 261720 221688
rect 261944 221740 261996 221746
rect 261944 221682 261996 221688
rect 261956 217410 261984 221682
rect 262140 219978 262168 227734
rect 263152 221610 263180 231662
rect 263416 227044 263468 227050
rect 263416 226986 263468 226992
rect 263140 221604 263192 221610
rect 263140 221546 263192 221552
rect 262956 220244 263008 220250
rect 262956 220186 263008 220192
rect 262128 219972 262180 219978
rect 262128 219914 262180 219920
rect 262968 217410 262996 220186
rect 259104 217382 259348 217410
rect 260176 217382 260604 217410
rect 261004 217382 261340 217410
rect 261832 217382 261984 217410
rect 262660 217382 262996 217410
rect 263428 217410 263456 226986
rect 263980 223038 264008 231676
rect 264256 231662 264546 231690
rect 263968 223032 264020 223038
rect 263968 222974 264020 222980
rect 264256 220114 264284 231662
rect 265084 224534 265112 231676
rect 265360 231662 265650 231690
rect 265360 229094 265388 231662
rect 265268 229066 265388 229094
rect 265072 224528 265124 224534
rect 265072 224470 265124 224476
rect 265268 222154 265296 229066
rect 265440 228812 265492 228818
rect 265440 228754 265492 228760
rect 265256 222148 265308 222154
rect 265256 222090 265308 222096
rect 264244 220108 264296 220114
rect 264244 220050 264296 220056
rect 264612 219632 264664 219638
rect 264612 219574 264664 219580
rect 264624 217410 264652 219574
rect 265452 217410 265480 228754
rect 266188 227322 266216 231676
rect 266740 230042 266768 231676
rect 267200 231662 267306 231690
rect 266728 230036 266780 230042
rect 266728 229978 266780 229984
rect 267004 229900 267056 229906
rect 267004 229842 267056 229848
rect 266176 227316 266228 227322
rect 266176 227258 266228 227264
rect 267016 222154 267044 229842
rect 267200 227186 267228 231662
rect 267556 227316 267608 227322
rect 267556 227258 267608 227264
rect 267188 227180 267240 227186
rect 267188 227122 267240 227128
rect 267372 227180 267424 227186
rect 267372 227122 267424 227128
rect 266268 222148 266320 222154
rect 266268 222090 266320 222096
rect 267004 222148 267056 222154
rect 267004 222090 267056 222096
rect 267188 222148 267240 222154
rect 267188 222090 267240 222096
rect 266280 217410 266308 222090
rect 267200 221746 267228 222090
rect 267188 221740 267240 221746
rect 267188 221682 267240 221688
rect 267096 220788 267148 220794
rect 267096 220730 267148 220736
rect 267108 217410 267136 220730
rect 263428 217382 263488 217410
rect 264316 217382 264652 217410
rect 265144 217382 265480 217410
rect 265972 217382 266308 217410
rect 266800 217382 267136 217410
rect 267384 217410 267412 227122
rect 267568 220794 267596 227258
rect 267844 226914 267872 231676
rect 267832 226908 267884 226914
rect 267832 226850 267884 226856
rect 268396 224262 268424 231676
rect 268948 227798 268976 231676
rect 268936 227792 268988 227798
rect 268936 227734 268988 227740
rect 269500 224670 269528 231676
rect 270052 224806 270080 231676
rect 270040 224800 270092 224806
rect 270040 224742 270092 224748
rect 269488 224664 269540 224670
rect 269488 224606 269540 224612
rect 270224 224528 270276 224534
rect 270224 224470 270276 224476
rect 268384 224256 268436 224262
rect 268384 224198 268436 224204
rect 268752 221604 268804 221610
rect 268752 221546 268804 221552
rect 267556 220788 267608 220794
rect 267556 220730 267608 220736
rect 268764 217410 268792 221546
rect 269580 220108 269632 220114
rect 269580 220050 269632 220056
rect 269592 217410 269620 220050
rect 270236 219638 270264 224470
rect 270408 224256 270460 224262
rect 270408 224198 270460 224204
rect 270224 219632 270276 219638
rect 270224 219574 270276 219580
rect 270420 217410 270448 224198
rect 270604 221474 270632 231676
rect 271156 230178 271184 231676
rect 271144 230172 271196 230178
rect 271144 230114 271196 230120
rect 271708 227458 271736 231676
rect 272076 231662 272274 231690
rect 271696 227452 271748 227458
rect 271696 227394 271748 227400
rect 271604 224392 271656 224398
rect 271604 224334 271656 224340
rect 270592 221468 270644 221474
rect 270592 221410 270644 221416
rect 271236 221468 271288 221474
rect 271236 221410 271288 221416
rect 271248 217410 271276 221410
rect 267384 217382 267628 217410
rect 268456 217382 268792 217410
rect 269284 217382 269620 217410
rect 270112 217382 270448 217410
rect 270940 217382 271276 217410
rect 271616 217410 271644 224334
rect 272076 221882 272104 231662
rect 272524 227724 272576 227730
rect 272524 227666 272576 227672
rect 272536 227050 272564 227666
rect 272524 227044 272576 227050
rect 272524 226986 272576 226992
rect 272812 224942 272840 231676
rect 273378 231662 273760 231690
rect 273732 229094 273760 231662
rect 273548 229066 273760 229094
rect 272800 224936 272852 224942
rect 272800 224878 272852 224884
rect 272984 223984 273036 223990
rect 272984 223926 273036 223932
rect 272064 221876 272116 221882
rect 272064 221818 272116 221824
rect 272996 217410 273024 223926
rect 273548 220386 273576 229066
rect 273916 228682 273944 231676
rect 274192 231662 274482 231690
rect 274744 231662 275034 231690
rect 273904 228676 273956 228682
rect 273904 228618 273956 228624
rect 273720 226160 273772 226166
rect 273720 226102 273772 226108
rect 273536 220380 273588 220386
rect 273536 220322 273588 220328
rect 273732 217410 273760 226102
rect 274192 225622 274220 231662
rect 274180 225616 274232 225622
rect 274180 225558 274232 225564
rect 274744 222018 274772 231662
rect 275572 230314 275600 231676
rect 275560 230308 275612 230314
rect 275560 230250 275612 230256
rect 275652 230036 275704 230042
rect 275652 229978 275704 229984
rect 275376 228948 275428 228954
rect 275376 228890 275428 228896
rect 274732 222012 274784 222018
rect 274732 221954 274784 221960
rect 274364 220380 274416 220386
rect 274364 220322 274416 220328
rect 274376 217410 274404 220322
rect 275388 217410 275416 228890
rect 275664 223990 275692 229978
rect 276124 228274 276152 231676
rect 276400 231662 276690 231690
rect 276400 229094 276428 231662
rect 276400 229066 276520 229094
rect 276296 228676 276348 228682
rect 276296 228618 276348 228624
rect 276112 228268 276164 228274
rect 276112 228210 276164 228216
rect 275652 223984 275704 223990
rect 275652 223926 275704 223932
rect 275652 220788 275704 220794
rect 275652 220730 275704 220736
rect 271616 217382 271768 217410
rect 272596 217382 273024 217410
rect 273424 217382 273760 217410
rect 274252 217382 274404 217410
rect 275080 217382 275416 217410
rect 275664 217410 275692 220730
rect 276308 220386 276336 228618
rect 276492 223582 276520 229066
rect 277228 227594 277256 231676
rect 277596 231662 277794 231690
rect 277216 227588 277268 227594
rect 277216 227530 277268 227536
rect 276480 223576 276532 223582
rect 276480 223518 276532 223524
rect 277124 223576 277176 223582
rect 277124 223518 277176 223524
rect 276296 220380 276348 220386
rect 276296 220322 276348 220328
rect 277136 217410 277164 223518
rect 277596 220930 277624 231662
rect 278332 223174 278360 231676
rect 278884 228546 278912 231676
rect 278872 228540 278924 228546
rect 278872 228482 278924 228488
rect 279436 225894 279464 231676
rect 279988 230450 280016 231676
rect 279976 230444 280028 230450
rect 279976 230386 280028 230392
rect 279884 230172 279936 230178
rect 279884 230114 279936 230120
rect 279424 225888 279476 225894
rect 279424 225830 279476 225836
rect 279608 225616 279660 225622
rect 279608 225558 279660 225564
rect 278320 223168 278372 223174
rect 278320 223110 278372 223116
rect 278688 223032 278740 223038
rect 278688 222974 278740 222980
rect 277584 220924 277636 220930
rect 277584 220866 277636 220872
rect 277860 220652 277912 220658
rect 277860 220594 277912 220600
rect 277872 217410 277900 220594
rect 278700 217410 278728 222974
rect 279620 220658 279648 225558
rect 279608 220652 279660 220658
rect 279608 220594 279660 220600
rect 279896 219434 279924 230114
rect 280540 226030 280568 231676
rect 280724 231662 281106 231690
rect 280528 226024 280580 226030
rect 280528 225966 280580 225972
rect 280068 221740 280120 221746
rect 280068 221682 280120 221688
rect 279620 219406 279924 219434
rect 279620 217410 279648 219406
rect 280080 217410 280108 221682
rect 280724 221338 280752 231662
rect 281644 228410 281672 231676
rect 281920 231662 282210 231690
rect 282472 231662 282762 231690
rect 281920 229094 281948 231662
rect 281828 229066 281948 229094
rect 281632 228404 281684 228410
rect 281632 228346 281684 228352
rect 281264 224664 281316 224670
rect 281264 224606 281316 224612
rect 280712 221332 280764 221338
rect 280712 221274 280764 221280
rect 281276 217410 281304 224606
rect 281828 220522 281856 229066
rect 282000 228404 282052 228410
rect 282000 228346 282052 228352
rect 281816 220516 281868 220522
rect 281816 220458 281868 220464
rect 282012 217410 282040 228346
rect 282472 223446 282500 231662
rect 283300 225758 283328 231676
rect 283656 227044 283708 227050
rect 283656 226986 283708 226992
rect 283288 225752 283340 225758
rect 283288 225694 283340 225700
rect 282460 223440 282512 223446
rect 282460 223382 282512 223388
rect 282552 220380 282604 220386
rect 282552 220322 282604 220328
rect 282564 217410 282592 220322
rect 283668 217410 283696 226986
rect 283852 222902 283880 231676
rect 284404 229770 284432 231676
rect 284588 231662 284970 231690
rect 284392 229764 284444 229770
rect 284392 229706 284444 229712
rect 283840 222896 283892 222902
rect 283840 222838 283892 222844
rect 284024 222896 284076 222902
rect 284024 222838 284076 222844
rect 275664 217382 275908 217410
rect 276736 217382 277164 217410
rect 277564 217382 277900 217410
rect 278392 217382 278728 217410
rect 279220 217382 279648 217410
rect 280048 217382 280108 217410
rect 280876 217382 281304 217410
rect 281704 217382 282040 217410
rect 282532 217382 282592 217410
rect 283360 217382 283696 217410
rect 284036 217410 284064 222838
rect 284588 222154 284616 231662
rect 284944 230376 284996 230382
rect 284944 230318 284996 230324
rect 284576 222148 284628 222154
rect 284576 222090 284628 222096
rect 284956 220250 284984 230318
rect 285508 227730 285536 231676
rect 285496 227724 285548 227730
rect 285496 227666 285548 227672
rect 286060 223310 286088 231676
rect 286612 230382 286640 231676
rect 286600 230376 286652 230382
rect 286600 230318 286652 230324
rect 287164 228818 287192 231676
rect 287440 231662 287730 231690
rect 287152 228812 287204 228818
rect 287152 228754 287204 228760
rect 286968 228540 287020 228546
rect 286968 228482 287020 228488
rect 286048 223304 286100 223310
rect 286048 223246 286100 223252
rect 285312 221876 285364 221882
rect 285312 221818 285364 221824
rect 284944 220244 284996 220250
rect 284944 220186 284996 220192
rect 285324 217410 285352 221818
rect 286140 220244 286192 220250
rect 286140 220186 286192 220192
rect 286152 217410 286180 220186
rect 286980 217410 287008 228482
rect 287440 227322 287468 231662
rect 287704 229560 287756 229566
rect 287704 229502 287756 229508
rect 287716 229094 287744 229502
rect 287624 229066 287744 229094
rect 287428 227316 287480 227322
rect 287428 227258 287480 227264
rect 287624 220114 287652 229066
rect 288268 224534 288296 231676
rect 288820 229906 288848 231676
rect 289004 231662 289386 231690
rect 288808 229900 288860 229906
rect 288808 229842 288860 229848
rect 288256 224528 288308 224534
rect 288256 224470 288308 224476
rect 288348 223168 288400 223174
rect 288348 223110 288400 223116
rect 287612 220108 287664 220114
rect 287612 220050 287664 220056
rect 287796 220108 287848 220114
rect 287796 220050 287848 220056
rect 287808 217410 287836 220050
rect 288360 217410 288388 223110
rect 289004 222018 289032 231662
rect 289544 226364 289596 226370
rect 289544 226306 289596 226312
rect 288992 222012 289044 222018
rect 288992 221954 289044 221960
rect 288624 221604 288676 221610
rect 288624 221546 288676 221552
rect 288636 220114 288664 221546
rect 288624 220108 288676 220114
rect 288624 220050 288676 220056
rect 289556 217410 289584 226306
rect 289924 224262 289952 231676
rect 290200 231662 290490 231690
rect 290200 227186 290228 231662
rect 290464 230444 290516 230450
rect 290464 230386 290516 230392
rect 290188 227180 290240 227186
rect 290188 227122 290240 227128
rect 290280 225752 290332 225758
rect 290280 225694 290332 225700
rect 289912 224256 289964 224262
rect 289912 224198 289964 224204
rect 290292 217410 290320 225694
rect 290476 220794 290504 230386
rect 291028 229566 291056 231676
rect 291016 229560 291068 229566
rect 291016 229502 291068 229508
rect 291580 224398 291608 231676
rect 291936 228812 291988 228818
rect 291936 228754 291988 228760
rect 291568 224392 291620 224398
rect 291568 224334 291620 224340
rect 291200 224256 291252 224262
rect 291200 224198 291252 224204
rect 290464 220788 290516 220794
rect 290464 220730 290516 220736
rect 291212 219434 291240 224198
rect 290844 219406 291240 219434
rect 290844 217410 290872 219406
rect 291948 217410 291976 228754
rect 292132 226166 292160 231676
rect 292120 226160 292172 226166
rect 292120 226102 292172 226108
rect 292684 221474 292712 231676
rect 293236 230042 293264 231676
rect 293512 231662 293802 231690
rect 293224 230036 293276 230042
rect 293224 229978 293276 229984
rect 293512 228954 293540 231662
rect 293868 229764 293920 229770
rect 293868 229706 293920 229712
rect 293500 228948 293552 228954
rect 293500 228890 293552 228896
rect 293684 227180 293736 227186
rect 293684 227122 293736 227128
rect 292672 221468 292724 221474
rect 292672 221410 292724 221416
rect 292304 220108 292356 220114
rect 292304 220050 292356 220056
rect 284036 217382 284188 217410
rect 285016 217382 285352 217410
rect 285844 217382 286180 217410
rect 286672 217382 287008 217410
rect 287500 217382 287836 217410
rect 288328 217382 288388 217410
rect 289156 217382 289584 217410
rect 289984 217382 290320 217410
rect 290812 217382 290872 217410
rect 291640 217382 291976 217410
rect 292316 217410 292344 220050
rect 293696 217410 293724 227122
rect 293880 226370 293908 229706
rect 293868 226364 293920 226370
rect 293868 226306 293920 226312
rect 294340 223582 294368 231676
rect 294892 228682 294920 231676
rect 295444 230450 295472 231676
rect 295432 230444 295484 230450
rect 295432 230386 295484 230392
rect 294880 228676 294932 228682
rect 294880 228618 294932 228624
rect 295248 228676 295300 228682
rect 295248 228618 295300 228624
rect 294328 223576 294380 223582
rect 294328 223518 294380 223524
rect 293960 223304 294012 223310
rect 293960 223246 294012 223252
rect 293972 220250 294000 223246
rect 293960 220244 294012 220250
rect 293960 220186 294012 220192
rect 294420 219496 294472 219502
rect 294420 219438 294472 219444
rect 294432 217410 294460 219438
rect 295260 217410 295288 228618
rect 295996 223038 296024 231676
rect 296180 231662 296562 231690
rect 295984 223032 296036 223038
rect 295984 222974 296036 222980
rect 296180 221746 296208 231662
rect 296720 230376 296772 230382
rect 296720 230318 296772 230324
rect 296732 224670 296760 230318
rect 297100 225622 297128 231676
rect 297652 230178 297680 231676
rect 297640 230172 297692 230178
rect 297640 230114 297692 230120
rect 297364 229900 297416 229906
rect 297364 229842 297416 229848
rect 297088 225616 297140 225622
rect 297088 225558 297140 225564
rect 296720 224664 296772 224670
rect 296720 224606 296772 224612
rect 296628 224392 296680 224398
rect 296628 224334 296680 224340
rect 296168 221740 296220 221746
rect 296168 221682 296220 221688
rect 296076 220856 296128 220862
rect 296076 220798 296128 220804
rect 296088 217410 296116 220798
rect 296640 217410 296668 224334
rect 297376 220862 297404 229842
rect 298204 228410 298232 231676
rect 298480 231662 298770 231690
rect 298192 228404 298244 228410
rect 298192 228346 298244 228352
rect 298480 227050 298508 231662
rect 299308 230382 299336 231676
rect 299296 230376 299348 230382
rect 299296 230318 299348 230324
rect 299860 230110 299888 231676
rect 300136 231662 300426 231690
rect 298744 230104 298796 230110
rect 298744 230046 298796 230052
rect 299848 230104 299900 230110
rect 299848 230046 299900 230052
rect 298468 227044 298520 227050
rect 298468 226986 298520 226992
rect 298008 225616 298060 225622
rect 298008 225558 298060 225564
rect 297364 220856 297416 220862
rect 297364 220798 297416 220804
rect 297732 220516 297784 220522
rect 297732 220458 297784 220464
rect 297744 217410 297772 220458
rect 298020 219502 298048 225558
rect 298560 221468 298612 221474
rect 298560 221410 298612 221416
rect 298008 219496 298060 219502
rect 298008 219438 298060 219444
rect 298572 217410 298600 221410
rect 298756 220386 298784 230046
rect 299388 227044 299440 227050
rect 299388 226986 299440 226992
rect 299400 220522 299428 226986
rect 299756 222624 299808 222630
rect 299756 222566 299808 222572
rect 299388 220516 299440 220522
rect 299388 220458 299440 220464
rect 298744 220380 298796 220386
rect 298744 220322 298796 220328
rect 299204 220244 299256 220250
rect 299204 220186 299256 220192
rect 299216 217410 299244 220186
rect 299768 220114 299796 222566
rect 300136 221882 300164 231662
rect 300492 230376 300544 230382
rect 300492 230318 300544 230324
rect 300504 222902 300532 230318
rect 300964 228546 300992 231676
rect 301516 230382 301544 231676
rect 301504 230376 301556 230382
rect 301504 230318 301556 230324
rect 300952 228540 301004 228546
rect 300952 228482 301004 228488
rect 302068 223310 302096 231676
rect 302056 223304 302108 223310
rect 302056 223246 302108 223252
rect 302620 223174 302648 231676
rect 303172 225758 303200 231676
rect 303160 225752 303212 225758
rect 303160 225694 303212 225700
rect 303344 225752 303396 225758
rect 303344 225694 303396 225700
rect 302608 223168 302660 223174
rect 302608 223110 302660 223116
rect 302240 223032 302292 223038
rect 302240 222974 302292 222980
rect 300492 222896 300544 222902
rect 300492 222838 300544 222844
rect 300124 221876 300176 221882
rect 300124 221818 300176 221824
rect 300124 221740 300176 221746
rect 300124 221682 300176 221688
rect 299756 220108 299808 220114
rect 299756 220050 299808 220056
rect 300136 217410 300164 221682
rect 300768 220380 300820 220386
rect 300768 220322 300820 220328
rect 300780 217410 300808 220322
rect 302252 219434 302280 222974
rect 302700 220788 302752 220794
rect 302700 220730 302752 220736
rect 301884 219406 302280 219434
rect 301884 217410 301912 219406
rect 302712 217410 302740 220730
rect 303356 220250 303384 225694
rect 303528 222896 303580 222902
rect 303528 222838 303580 222844
rect 303344 220244 303396 220250
rect 303344 220186 303396 220192
rect 303540 217410 303568 222838
rect 303724 221610 303752 231676
rect 304276 229770 304304 231676
rect 304264 229764 304316 229770
rect 304264 229706 304316 229712
rect 304828 228818 304856 231676
rect 304816 228812 304868 228818
rect 304816 228754 304868 228760
rect 304356 228404 304408 228410
rect 304356 228346 304408 228352
rect 303712 221604 303764 221610
rect 303712 221546 303764 221552
rect 304368 217410 304396 228346
rect 305380 227186 305408 231676
rect 305644 230036 305696 230042
rect 305644 229978 305696 229984
rect 305368 227180 305420 227186
rect 305368 227122 305420 227128
rect 305000 224528 305052 224534
rect 305000 224470 305052 224476
rect 304632 220652 304684 220658
rect 304632 220594 304684 220600
rect 292316 217382 292468 217410
rect 293296 217382 293724 217410
rect 294124 217382 294460 217410
rect 294952 217382 295288 217410
rect 295780 217382 296116 217410
rect 296608 217382 296668 217410
rect 297436 217382 297772 217410
rect 298264 217382 298600 217410
rect 299092 217382 299244 217410
rect 299920 217382 300164 217410
rect 300748 217382 300808 217410
rect 301576 217382 301912 217410
rect 302404 217382 302740 217410
rect 303232 217382 303568 217410
rect 304060 217382 304396 217410
rect 304644 217410 304672 220594
rect 305012 220386 305040 224470
rect 305656 220794 305684 229978
rect 305932 224262 305960 231676
rect 305920 224256 305972 224262
rect 305920 224198 305972 224204
rect 306484 222630 306512 231676
rect 307036 228682 307064 231676
rect 307024 228676 307076 228682
rect 307024 228618 307076 228624
rect 307588 224398 307616 231676
rect 308140 225622 308168 231676
rect 308692 229906 308720 231676
rect 308680 229900 308732 229906
rect 308680 229842 308732 229848
rect 308864 229900 308916 229906
rect 308864 229842 308916 229848
rect 308496 227792 308548 227798
rect 308496 227734 308548 227740
rect 308128 225616 308180 225622
rect 308128 225558 308180 225564
rect 307576 224392 307628 224398
rect 307576 224334 307628 224340
rect 307484 224256 307536 224262
rect 307484 224198 307536 224204
rect 306472 222624 306524 222630
rect 306472 222566 306524 222572
rect 305644 220788 305696 220794
rect 305644 220730 305696 220736
rect 306840 220516 306892 220522
rect 306840 220458 306892 220464
rect 305000 220380 305052 220386
rect 305000 220322 305052 220328
rect 306012 219496 306064 219502
rect 306012 219438 306064 219444
rect 306024 217410 306052 219438
rect 306852 217410 306880 220458
rect 307496 219502 307524 224198
rect 307668 220312 307720 220318
rect 307668 220254 307720 220260
rect 307484 219496 307536 219502
rect 307484 219438 307536 219444
rect 307680 217410 307708 220254
rect 308508 217410 308536 227734
rect 308876 219434 308904 229842
rect 309244 221474 309272 231676
rect 309520 231662 309810 231690
rect 309520 221746 309548 231662
rect 310348 227050 310376 231676
rect 310336 227044 310388 227050
rect 310336 226986 310388 226992
rect 310900 225758 310928 231676
rect 311072 227044 311124 227050
rect 311072 226986 311124 226992
rect 310888 225752 310940 225758
rect 310888 225694 310940 225700
rect 310612 223440 310664 223446
rect 310612 223382 310664 223388
rect 309508 221740 309560 221746
rect 309508 221682 309560 221688
rect 310060 221740 310112 221746
rect 310060 221682 310112 221688
rect 309232 221468 309284 221474
rect 309232 221410 309284 221416
rect 304644 217382 304888 217410
rect 305716 217382 306052 217410
rect 306544 217382 306880 217410
rect 307372 217382 307708 217410
rect 308200 217382 308536 217410
rect 308784 219406 308904 219434
rect 308784 217410 308812 219406
rect 310072 217410 310100 221682
rect 310624 220522 310652 223382
rect 310612 220516 310664 220522
rect 310612 220458 310664 220464
rect 311084 219434 311112 226986
rect 311452 223038 311480 231676
rect 311440 223032 311492 223038
rect 311440 222974 311492 222980
rect 312004 222902 312032 231676
rect 312556 224534 312584 231676
rect 313108 230042 313136 231676
rect 313476 231662 313674 231690
rect 313096 230036 313148 230042
rect 313096 229978 313148 229984
rect 312728 225752 312780 225758
rect 312728 225694 312780 225700
rect 312544 224528 312596 224534
rect 312544 224470 312596 224476
rect 311992 222896 312044 222902
rect 311992 222838 312044 222844
rect 311624 219632 311676 219638
rect 311624 219574 311676 219580
rect 310992 219406 311112 219434
rect 310992 217410 311020 219406
rect 311636 217410 311664 219574
rect 312740 217410 312768 225694
rect 313096 223576 313148 223582
rect 313096 223518 313148 223524
rect 308784 217382 309028 217410
rect 309856 217382 310100 217410
rect 310684 217382 311020 217410
rect 311512 217382 311664 217410
rect 312340 217382 312768 217410
rect 313108 217410 313136 223518
rect 313476 220862 313504 231662
rect 314212 223446 314240 231676
rect 314764 228410 314792 231676
rect 315040 231662 315330 231690
rect 314752 228404 314804 228410
rect 314752 228346 314804 228352
rect 315040 224262 315068 231662
rect 315868 227798 315896 231676
rect 316144 231662 316434 231690
rect 315856 227792 315908 227798
rect 315856 227734 315908 227740
rect 315856 227656 315908 227662
rect 315856 227598 315908 227604
rect 315028 224256 315080 224262
rect 315028 224198 315080 224204
rect 314200 223440 314252 223446
rect 314200 223382 314252 223388
rect 314384 222896 314436 222902
rect 314384 222838 314436 222844
rect 313464 220856 313516 220862
rect 313464 220798 313516 220804
rect 314396 217410 314424 222838
rect 315120 221604 315172 221610
rect 315120 221546 315172 221552
rect 315132 217410 315160 221546
rect 315868 220318 315896 227598
rect 316144 221746 316172 231662
rect 316972 227798 317000 231676
rect 317524 229906 317552 231676
rect 317800 231662 318090 231690
rect 317512 229900 317564 229906
rect 317512 229842 317564 229848
rect 317512 229492 317564 229498
rect 317512 229434 317564 229440
rect 316960 227792 317012 227798
rect 316960 227734 317012 227740
rect 317328 227792 317380 227798
rect 317328 227734 317380 227740
rect 316132 221740 316184 221746
rect 316132 221682 316184 221688
rect 316040 221468 316092 221474
rect 316040 221410 316092 221416
rect 315856 220312 315908 220318
rect 315856 220254 315908 220260
rect 316052 219450 316080 221410
rect 316776 220788 316828 220794
rect 316776 220730 316828 220736
rect 315960 219422 316080 219450
rect 315960 217410 315988 219422
rect 316788 217410 316816 220730
rect 317340 217410 317368 227734
rect 317524 225758 317552 229434
rect 317512 225752 317564 225758
rect 317512 225694 317564 225700
rect 317800 219638 317828 231662
rect 318628 223582 318656 231676
rect 319180 227050 319208 231676
rect 319444 230376 319496 230382
rect 319444 230318 319496 230324
rect 319168 227044 319220 227050
rect 319168 226986 319220 226992
rect 318616 223576 318668 223582
rect 318616 223518 318668 223524
rect 319456 221610 319484 230318
rect 319732 229498 319760 231676
rect 320284 230382 320312 231676
rect 320560 231662 320850 231690
rect 320272 230376 320324 230382
rect 320272 230318 320324 230324
rect 319720 229492 319772 229498
rect 319720 229434 319772 229440
rect 320088 229356 320140 229362
rect 320088 229298 320140 229304
rect 320100 222902 320128 229298
rect 320088 222896 320140 222902
rect 320088 222838 320140 222844
rect 319444 221604 319496 221610
rect 319444 221546 319496 221552
rect 320560 220794 320588 231662
rect 321388 229362 321416 231676
rect 321664 231662 321954 231690
rect 322216 231662 322506 231690
rect 323058 231662 323440 231690
rect 321376 229356 321428 229362
rect 321376 229298 321428 229304
rect 321376 229152 321428 229158
rect 321376 229094 321428 229100
rect 321388 220794 321416 229094
rect 321664 221474 321692 231662
rect 321836 229696 321888 229702
rect 321836 229638 321888 229644
rect 321848 227798 321876 229638
rect 321836 227792 321888 227798
rect 321836 227734 321888 227740
rect 321652 221468 321704 221474
rect 321652 221410 321704 221416
rect 320548 220788 320600 220794
rect 320548 220730 320600 220736
rect 320916 220788 320968 220794
rect 320916 220730 320968 220736
rect 321376 220788 321428 220794
rect 321376 220730 321428 220736
rect 320088 220516 320140 220522
rect 320088 220458 320140 220464
rect 318432 220380 318484 220386
rect 318432 220322 318484 220328
rect 317788 219632 317840 219638
rect 317788 219574 317840 219580
rect 318444 217410 318472 220322
rect 319260 220108 319312 220114
rect 319260 220050 319312 220056
rect 319272 217410 319300 220050
rect 320100 217410 320128 220458
rect 320928 217410 320956 220730
rect 321192 220652 321244 220658
rect 321192 220594 321244 220600
rect 313108 217382 313168 217410
rect 313996 217382 314424 217410
rect 314824 217382 315160 217410
rect 315652 217382 315988 217410
rect 316480 217382 316816 217410
rect 317308 217382 317368 217410
rect 318136 217382 318472 217410
rect 318964 217382 319300 217410
rect 319792 217382 320128 217410
rect 320620 217382 320956 217410
rect 321204 217410 321232 220594
rect 322216 220386 322244 231662
rect 323412 229094 323440 231662
rect 323596 229702 323624 231676
rect 323872 231662 324162 231690
rect 323584 229696 323636 229702
rect 323584 229638 323636 229644
rect 323228 229066 323440 229094
rect 323228 220522 323256 229066
rect 323400 220788 323452 220794
rect 323400 220730 323452 220736
rect 323216 220516 323268 220522
rect 323216 220458 323268 220464
rect 322204 220380 322256 220386
rect 322204 220322 322256 220328
rect 322572 219768 322624 219774
rect 322572 219710 322624 219716
rect 322584 217410 322612 219710
rect 323412 217410 323440 220730
rect 323872 220114 323900 231662
rect 324700 220658 324728 231676
rect 324976 231662 325266 231690
rect 324976 220794 325004 231662
rect 325804 229158 325832 231676
rect 325988 231662 326370 231690
rect 326632 231662 326922 231690
rect 327368 231662 327474 231690
rect 327736 231662 328026 231690
rect 328578 231662 328868 231690
rect 325792 229152 325844 229158
rect 325792 229094 325844 229100
rect 324964 220788 325016 220794
rect 324964 220730 325016 220736
rect 324688 220652 324740 220658
rect 324688 220594 324740 220600
rect 325608 220380 325660 220386
rect 325608 220322 325660 220328
rect 323860 220108 323912 220114
rect 323860 220050 323912 220056
rect 324228 219632 324280 219638
rect 324228 219574 324280 219580
rect 324240 217410 324268 219574
rect 325056 219496 325108 219502
rect 325056 219438 325108 219444
rect 325068 217410 325096 219438
rect 325620 217410 325648 220322
rect 325988 219774 326016 231662
rect 326632 229094 326660 231662
rect 326540 229066 326660 229094
rect 325976 219768 326028 219774
rect 325976 219710 326028 219716
rect 326540 219502 326568 229066
rect 327368 220794 327396 231662
rect 326712 220788 326764 220794
rect 326712 220730 326764 220736
rect 327356 220788 327408 220794
rect 327356 220730 327408 220736
rect 326528 219496 326580 219502
rect 326528 219438 326580 219444
rect 326724 217410 326752 220730
rect 327540 220652 327592 220658
rect 327540 220594 327592 220600
rect 327552 217410 327580 220594
rect 327736 219638 327764 231662
rect 328840 229094 328868 231662
rect 328748 229066 328868 229094
rect 328932 231662 329130 231690
rect 329300 231662 329682 231690
rect 328184 220788 328236 220794
rect 328184 220730 328236 220736
rect 327724 219632 327776 219638
rect 327724 219574 327776 219580
rect 328196 217410 328224 220730
rect 328748 220386 328776 229066
rect 328932 220794 328960 231662
rect 328920 220788 328972 220794
rect 328920 220730 328972 220736
rect 329104 220788 329156 220794
rect 329104 220730 329156 220736
rect 328736 220380 328788 220386
rect 328736 220322 328788 220328
rect 329116 217410 329144 220730
rect 321204 217382 321448 217410
rect 322276 217382 322612 217410
rect 323104 217382 323440 217410
rect 323932 217382 324268 217410
rect 324760 217382 325096 217410
rect 325588 217382 325648 217410
rect 326416 217382 326752 217410
rect 327244 217382 327580 217410
rect 328072 217382 328224 217410
rect 328900 217382 329144 217410
rect 329300 217410 329328 231662
rect 330220 220658 330248 231676
rect 330496 231662 330786 231690
rect 331338 231662 331628 231690
rect 330496 220794 330524 231662
rect 330484 220788 330536 220794
rect 330484 220730 330536 220736
rect 330852 220788 330904 220794
rect 330852 220730 330904 220736
rect 330208 220652 330260 220658
rect 330208 220594 330260 220600
rect 330864 217410 330892 220730
rect 331600 217410 331628 231662
rect 331876 230382 331904 231676
rect 332152 231662 332442 231690
rect 332704 231662 332994 231690
rect 331864 230376 331916 230382
rect 331864 230318 331916 230324
rect 332152 220794 332180 231662
rect 332140 220788 332192 220794
rect 332140 220730 332192 220736
rect 332704 219434 332732 231662
rect 333532 230382 333560 231676
rect 333060 230376 333112 230382
rect 333060 230318 333112 230324
rect 333520 230376 333572 230382
rect 333520 230318 333572 230324
rect 332520 219406 332732 219434
rect 332520 217410 332548 219406
rect 333072 217410 333100 230318
rect 334084 229294 334112 231676
rect 334360 231662 334650 231690
rect 334072 229288 334124 229294
rect 334072 229230 334124 229236
rect 334360 220794 334388 231662
rect 334532 230376 334584 230382
rect 334532 230318 334584 230324
rect 333888 220788 333940 220794
rect 333888 220730 333940 220736
rect 334348 220788 334400 220794
rect 334348 220730 334400 220736
rect 333900 217410 333928 220730
rect 334544 219434 334572 230318
rect 335188 229106 335216 231676
rect 335740 230178 335768 231676
rect 335728 230172 335780 230178
rect 335728 230114 335780 230120
rect 336292 229838 336320 231676
rect 336280 229832 336332 229838
rect 336280 229774 336332 229780
rect 335544 229288 335596 229294
rect 335544 229230 335596 229236
rect 335188 229078 335400 229106
rect 329300 217382 329728 217410
rect 330556 217382 330892 217410
rect 331384 217382 331628 217410
rect 332212 217382 332548 217410
rect 333040 217382 333100 217410
rect 333868 217382 333928 217410
rect 334452 219406 334572 219434
rect 334452 217410 334480 219406
rect 335372 217410 335400 229078
rect 335556 229094 335584 229230
rect 335556 229066 335952 229094
rect 335924 217410 335952 229066
rect 336844 217410 336872 231676
rect 337410 231662 337884 231690
rect 337292 230172 337344 230178
rect 337292 230114 337344 230120
rect 337304 229094 337332 230114
rect 337856 229094 337884 231662
rect 337948 230330 337976 231676
rect 337948 230302 338068 230330
rect 338040 230246 338068 230302
rect 338028 230240 338080 230246
rect 338028 230182 338080 230188
rect 338500 230110 338528 231676
rect 338488 230104 338540 230110
rect 338488 230046 338540 230052
rect 339052 229974 339080 231676
rect 339604 230382 339632 231676
rect 340170 231662 340552 231690
rect 339592 230376 339644 230382
rect 339592 230318 339644 230324
rect 339040 229968 339092 229974
rect 339040 229910 339092 229916
rect 340144 229968 340196 229974
rect 340144 229910 340196 229916
rect 339776 229832 339828 229838
rect 339776 229774 339828 229780
rect 337304 229066 337608 229094
rect 337856 229066 338436 229094
rect 337580 217410 337608 229066
rect 338408 217410 338436 229066
rect 339788 219434 339816 229774
rect 339696 219406 339816 219434
rect 339696 217410 339724 219406
rect 334452 217382 334696 217410
rect 335372 217382 335524 217410
rect 335924 217382 336352 217410
rect 336844 217382 337180 217410
rect 337580 217382 338008 217410
rect 338408 217382 338836 217410
rect 339664 217382 339724 217410
rect 340156 217410 340184 229910
rect 340524 229770 340552 231662
rect 340512 229764 340564 229770
rect 340512 229706 340564 229712
rect 340708 219502 340736 231676
rect 340972 230376 341024 230382
rect 340972 230318 341024 230324
rect 340696 219496 340748 219502
rect 340696 219438 340748 219444
rect 340984 217870 341012 230318
rect 341260 229906 341288 231676
rect 341812 230246 341840 231676
rect 341432 230240 341484 230246
rect 341432 230182 341484 230188
rect 341800 230240 341852 230246
rect 341800 230182 341852 230188
rect 341248 229900 341300 229906
rect 341248 229842 341300 229848
rect 341444 219434 341472 230182
rect 342364 229634 342392 231676
rect 342720 230104 342772 230110
rect 342720 230046 342772 230052
rect 342352 229628 342404 229634
rect 342352 229570 342404 229576
rect 341352 219406 341472 219434
rect 340972 217864 341024 217870
rect 340972 217806 341024 217812
rect 341352 217410 341380 219406
rect 341800 217864 341852 217870
rect 341800 217806 341852 217812
rect 340156 217382 340492 217410
rect 341320 217382 341380 217410
rect 341812 217410 341840 217806
rect 342732 217410 342760 230046
rect 342916 222902 342944 231676
rect 343376 231662 343482 231690
rect 343376 229430 343404 231662
rect 343732 230240 343784 230246
rect 343732 230182 343784 230188
rect 343548 229628 343600 229634
rect 343548 229570 343600 229576
rect 343364 229424 343416 229430
rect 343364 229366 343416 229372
rect 342904 222896 342956 222902
rect 342904 222838 342956 222844
rect 343560 221746 343588 229570
rect 343744 229566 343772 230182
rect 344020 230042 344048 231676
rect 344586 231662 344876 231690
rect 344008 230036 344060 230042
rect 344008 229978 344060 229984
rect 344100 229900 344152 229906
rect 344100 229842 344152 229848
rect 343916 229764 343968 229770
rect 343916 229706 343968 229712
rect 343732 229560 343784 229566
rect 343732 229502 343784 229508
rect 343548 221740 343600 221746
rect 343548 221682 343600 221688
rect 343928 217870 343956 229706
rect 343916 217864 343968 217870
rect 343916 217806 343968 217812
rect 344112 217410 344140 229842
rect 344848 221610 344876 231662
rect 345124 223446 345152 231676
rect 345676 230246 345704 231676
rect 345664 230240 345716 230246
rect 345664 230182 345716 230188
rect 345388 229560 345440 229566
rect 345388 229502 345440 229508
rect 345112 223440 345164 223446
rect 345112 223382 345164 223388
rect 344836 221604 344888 221610
rect 344836 221546 344888 221552
rect 344284 217864 344336 217870
rect 344284 217806 344336 217812
rect 341812 217382 342148 217410
rect 342732 217382 342976 217410
rect 343804 217382 344140 217410
rect 344296 217410 344324 217806
rect 345400 217410 345428 229502
rect 346228 220794 346256 231676
rect 346794 231662 347176 231690
rect 346676 229424 346728 229430
rect 346676 229366 346728 229372
rect 346216 220788 346268 220794
rect 346216 220730 346268 220736
rect 345940 219496 345992 219502
rect 345940 219438 345992 219444
rect 345952 217410 345980 219438
rect 346688 217410 346716 229366
rect 347148 222154 347176 231662
rect 347332 228546 347360 231676
rect 347320 228540 347372 228546
rect 347320 228482 347372 228488
rect 347884 224806 347912 231676
rect 348450 231662 348924 231690
rect 348240 230036 348292 230042
rect 348240 229978 348292 229984
rect 348252 229094 348280 229978
rect 348252 229066 348372 229094
rect 347872 224800 347924 224806
rect 347872 224742 347924 224748
rect 347136 222148 347188 222154
rect 347136 222090 347188 222096
rect 347872 221740 347924 221746
rect 347872 221682 347924 221688
rect 347884 217410 347912 221682
rect 348344 217410 348372 229066
rect 348896 219502 348924 231662
rect 348988 229650 349016 231676
rect 349540 230042 349568 231676
rect 349712 230240 349764 230246
rect 349712 230182 349764 230188
rect 349528 230036 349580 230042
rect 349528 229978 349580 229984
rect 348988 229634 349108 229650
rect 348988 229628 349120 229634
rect 348988 229622 349068 229628
rect 349068 229570 349120 229576
rect 349724 229094 349752 230182
rect 350092 229094 350120 231676
rect 350644 229294 350672 231676
rect 350632 229288 350684 229294
rect 350632 229230 350684 229236
rect 349724 229066 350028 229094
rect 350092 229066 350212 229094
rect 349252 222896 349304 222902
rect 349252 222838 349304 222844
rect 348884 219496 348936 219502
rect 348884 219438 348936 219444
rect 349264 217410 349292 222838
rect 350000 217410 350028 229066
rect 350184 223582 350212 229066
rect 351196 228410 351224 231676
rect 351184 228404 351236 228410
rect 351184 228346 351236 228352
rect 350172 223576 350224 223582
rect 350172 223518 350224 223524
rect 351748 221746 351776 231676
rect 352300 225758 352328 231676
rect 352866 231662 353248 231690
rect 353024 229628 353076 229634
rect 353024 229570 353076 229576
rect 352288 225752 352340 225758
rect 352288 225694 352340 225700
rect 352472 223440 352524 223446
rect 352472 223382 352524 223388
rect 351736 221740 351788 221746
rect 351736 221682 351788 221688
rect 350908 221604 350960 221610
rect 350908 221546 350960 221552
rect 350920 217410 350948 221546
rect 351920 220788 351972 220794
rect 351920 220730 351972 220736
rect 351932 217410 351960 220730
rect 352484 217410 352512 223382
rect 353036 223174 353064 229570
rect 353024 223168 353076 223174
rect 353024 223110 353076 223116
rect 353220 220114 353248 231662
rect 353404 230382 353432 231676
rect 353392 230376 353444 230382
rect 353392 230318 353444 230324
rect 353956 227050 353984 231676
rect 354416 231662 354522 231690
rect 353944 227044 353996 227050
rect 353944 226986 353996 226992
rect 353484 224800 353536 224806
rect 353484 224742 353536 224748
rect 353208 220108 353260 220114
rect 353208 220050 353260 220056
rect 353496 217410 353524 224742
rect 354416 223038 354444 231662
rect 355060 230382 355088 231676
rect 355626 231662 356008 231690
rect 354588 230376 354640 230382
rect 354588 230318 354640 230324
rect 355048 230376 355100 230382
rect 355048 230318 355100 230324
rect 354404 223032 354456 223038
rect 354404 222974 354456 222980
rect 354220 222148 354272 222154
rect 354220 222090 354272 222096
rect 354232 217410 354260 222090
rect 354600 221610 354628 230318
rect 355324 229288 355376 229294
rect 355324 229230 355376 229236
rect 354588 221604 354640 221610
rect 354588 221546 354640 221552
rect 355336 220794 355364 229230
rect 355692 223576 355744 223582
rect 355692 223518 355744 223524
rect 355324 220788 355376 220794
rect 355324 220730 355376 220736
rect 355704 220658 355732 223518
rect 355980 222902 356008 231662
rect 356164 229634 356192 231676
rect 356730 231662 357112 231690
rect 356704 230376 356756 230382
rect 356704 230318 356756 230324
rect 356336 230036 356388 230042
rect 356336 229978 356388 229984
rect 356152 229628 356204 229634
rect 356152 229570 356204 229576
rect 356152 228540 356204 228546
rect 356152 228482 356204 228488
rect 355968 222896 356020 222902
rect 355968 222838 356020 222844
rect 355692 220652 355744 220658
rect 355692 220594 355744 220600
rect 355048 219496 355100 219502
rect 355048 219438 355100 219444
rect 355060 217410 355088 219438
rect 356164 217410 356192 228482
rect 356348 228002 356376 229978
rect 356716 229094 356744 230318
rect 356716 229066 356928 229094
rect 356336 227996 356388 228002
rect 356336 227938 356388 227944
rect 356704 220652 356756 220658
rect 356704 220594 356756 220600
rect 356716 217410 356744 220594
rect 356900 220250 356928 229066
rect 357084 225622 357112 231662
rect 357268 230246 357296 231676
rect 357834 231662 358216 231690
rect 357256 230240 357308 230246
rect 357256 230182 357308 230188
rect 357624 225752 357676 225758
rect 357624 225694 357676 225700
rect 357072 225616 357124 225622
rect 357072 225558 357124 225564
rect 357440 223168 357492 223174
rect 357440 223110 357492 223116
rect 356888 220244 356940 220250
rect 356888 220186 356940 220192
rect 357452 217410 357480 223110
rect 357636 220658 357664 225694
rect 358188 221474 358216 231662
rect 358372 224262 358400 231676
rect 358924 229906 358952 231676
rect 359476 230382 359504 231676
rect 359464 230376 359516 230382
rect 359464 230318 359516 230324
rect 359740 230240 359792 230246
rect 359740 230182 359792 230188
rect 358912 229900 358964 229906
rect 358912 229842 358964 229848
rect 359096 227996 359148 228002
rect 359096 227938 359148 227944
rect 358360 224256 358412 224262
rect 358360 224198 358412 224204
rect 358176 221468 358228 221474
rect 358176 221410 358228 221416
rect 358360 220788 358412 220794
rect 358360 220730 358412 220736
rect 357624 220652 357676 220658
rect 357624 220594 357676 220600
rect 358372 217410 358400 220730
rect 359108 217410 359136 227938
rect 359752 224398 359780 230182
rect 360028 228682 360056 231676
rect 360580 228818 360608 231676
rect 361132 230178 361160 231676
rect 361488 230376 361540 230382
rect 361488 230318 361540 230324
rect 361120 230172 361172 230178
rect 361120 230114 361172 230120
rect 360568 228812 360620 228818
rect 360568 228754 360620 228760
rect 360016 228676 360068 228682
rect 360016 228618 360068 228624
rect 360752 228404 360804 228410
rect 360752 228346 360804 228352
rect 359740 224392 359792 224398
rect 359740 224334 359792 224340
rect 360200 220652 360252 220658
rect 360200 220594 360252 220600
rect 360212 217410 360240 220594
rect 360764 217410 360792 228346
rect 361500 227186 361528 230318
rect 361684 229770 361712 231676
rect 362250 231662 362632 231690
rect 362408 229900 362460 229906
rect 362408 229842 362460 229848
rect 361672 229764 361724 229770
rect 361672 229706 361724 229712
rect 361488 227180 361540 227186
rect 361488 227122 361540 227128
rect 362420 223310 362448 229842
rect 362408 223304 362460 223310
rect 362408 223246 362460 223252
rect 362604 221882 362632 231662
rect 362788 225758 362816 231676
rect 363340 230042 363368 231676
rect 363906 231662 364196 231690
rect 363972 230172 364024 230178
rect 363972 230114 364024 230120
rect 363328 230036 363380 230042
rect 363328 229978 363380 229984
rect 363144 229628 363196 229634
rect 363144 229570 363196 229576
rect 362776 225752 362828 225758
rect 362776 225694 362828 225700
rect 363156 223174 363184 229570
rect 363984 228410 364012 230114
rect 363972 228404 364024 228410
rect 363972 228346 364024 228352
rect 363144 223168 363196 223174
rect 363144 223110 363196 223116
rect 363236 223032 363288 223038
rect 363236 222974 363288 222980
rect 362592 221876 362644 221882
rect 362592 221818 362644 221824
rect 362500 221740 362552 221746
rect 362500 221682 362552 221688
rect 361672 220108 361724 220114
rect 361672 220050 361724 220056
rect 361684 217410 361712 220050
rect 362512 217410 362540 221682
rect 363248 217410 363276 222974
rect 364168 220114 364196 231662
rect 364444 230382 364472 231676
rect 365010 231662 365392 231690
rect 364432 230376 364484 230382
rect 364432 230318 364484 230324
rect 365364 229094 365392 231662
rect 365548 230466 365576 231676
rect 366114 231662 366588 231690
rect 366666 231662 366864 231690
rect 365548 230438 365852 230466
rect 365628 230376 365680 230382
rect 365628 230318 365680 230324
rect 365364 229066 365484 229094
rect 365456 225622 365484 229066
rect 365260 225616 365312 225622
rect 365260 225558 365312 225564
rect 365444 225616 365496 225622
rect 365444 225558 365496 225564
rect 364340 221604 364392 221610
rect 364340 221546 364392 221552
rect 364156 220108 364208 220114
rect 364156 220050 364208 220056
rect 364352 217410 364380 221546
rect 365272 220794 365300 225558
rect 365640 221610 365668 230318
rect 365824 229906 365852 230438
rect 365812 229900 365864 229906
rect 365812 229842 365864 229848
rect 366560 229094 366588 231662
rect 366468 229066 366588 229094
rect 365812 227044 365864 227050
rect 365812 226986 365864 226992
rect 365628 221604 365680 221610
rect 365628 221546 365680 221552
rect 365260 220788 365312 220794
rect 365260 220730 365312 220736
rect 365168 220244 365220 220250
rect 365168 220186 365220 220192
rect 365180 217410 365208 220186
rect 365824 217410 365852 226986
rect 366468 220386 366496 229066
rect 366836 227050 366864 231662
rect 367204 227322 367232 231676
rect 367756 229294 367784 231676
rect 368124 231662 368322 231690
rect 367744 229288 367796 229294
rect 367744 229230 367796 229236
rect 367192 227316 367244 227322
rect 367192 227258 367244 227264
rect 366824 227044 366876 227050
rect 366824 226986 366876 226992
rect 367376 222896 367428 222902
rect 367376 222838 367428 222844
rect 366640 220788 366692 220794
rect 366640 220730 366692 220736
rect 366456 220380 366508 220386
rect 366456 220322 366508 220328
rect 366652 217410 366680 220730
rect 367388 217410 367416 222838
rect 368124 220250 368152 231662
rect 368388 230036 368440 230042
rect 368388 229978 368440 229984
rect 368400 224534 368428 229978
rect 368388 224528 368440 224534
rect 368388 224470 368440 224476
rect 368480 224392 368532 224398
rect 368480 224334 368532 224340
rect 368112 220244 368164 220250
rect 368112 220186 368164 220192
rect 368492 217410 368520 224334
rect 368860 223446 368888 231676
rect 369412 230246 369440 231676
rect 369400 230240 369452 230246
rect 369400 230182 369452 230188
rect 369584 229764 369636 229770
rect 369584 229706 369636 229712
rect 369596 223582 369624 229706
rect 369964 228546 369992 231676
rect 369952 228540 370004 228546
rect 369952 228482 370004 228488
rect 370516 224942 370544 231676
rect 370504 224936 370556 224942
rect 370504 224878 370556 224884
rect 369584 223576 369636 223582
rect 369584 223518 369636 223524
rect 368848 223440 368900 223446
rect 368848 223382 368900 223388
rect 369860 223168 369912 223174
rect 369860 223110 369912 223116
rect 369032 223032 369084 223038
rect 369032 222974 369084 222980
rect 369044 217410 369072 222974
rect 369872 217410 369900 223110
rect 371068 222902 371096 231676
rect 371620 230382 371648 231676
rect 371608 230376 371660 230382
rect 371608 230318 371660 230324
rect 371884 230240 371936 230246
rect 371884 230182 371936 230188
rect 371516 227180 371568 227186
rect 371516 227122 371568 227128
rect 371056 222896 371108 222902
rect 371056 222838 371108 222844
rect 370780 221468 370832 221474
rect 370780 221410 370832 221416
rect 370792 217410 370820 221410
rect 371528 217410 371556 227122
rect 371896 221746 371924 230182
rect 372172 227458 372200 231676
rect 372724 230042 372752 231676
rect 372712 230036 372764 230042
rect 372712 229978 372764 229984
rect 373276 228410 373304 231676
rect 373632 230376 373684 230382
rect 373632 230318 373684 230324
rect 373080 228404 373132 228410
rect 373080 228346 373132 228352
rect 373264 228404 373316 228410
rect 373264 228346 373316 228352
rect 372160 227452 372212 227458
rect 372160 227394 372212 227400
rect 372712 224256 372764 224262
rect 372712 224198 372764 224204
rect 371884 221740 371936 221746
rect 371884 221682 371936 221688
rect 372724 217410 372752 224198
rect 373092 219434 373120 228346
rect 373644 223038 373672 230318
rect 373828 229158 373856 231676
rect 373816 229152 373868 229158
rect 373816 229094 373868 229100
rect 374184 228676 374236 228682
rect 374184 228618 374236 228624
rect 374000 223576 374052 223582
rect 374000 223518 374052 223524
rect 373632 223032 373684 223038
rect 373632 222974 373684 222980
rect 373092 219406 373212 219434
rect 373184 217410 373212 219406
rect 374012 217870 374040 223518
rect 374000 217864 374052 217870
rect 374000 217806 374052 217812
rect 374196 217410 374224 228618
rect 374380 223174 374408 231676
rect 374932 230178 374960 231676
rect 375498 231662 375880 231690
rect 376050 231662 376432 231690
rect 374920 230172 374972 230178
rect 374920 230114 374972 230120
rect 374644 229152 374696 229158
rect 374644 229094 374696 229100
rect 374368 223168 374420 223174
rect 374368 223110 374420 223116
rect 374656 221474 374684 229094
rect 375656 228812 375708 228818
rect 375656 228754 375708 228760
rect 374644 221468 374696 221474
rect 374644 221410 374696 221416
rect 374920 217864 374972 217870
rect 374920 217806 374972 217812
rect 374932 217410 374960 217806
rect 375668 217410 375696 228754
rect 375852 224670 375880 231662
rect 376116 224936 376168 224942
rect 376116 224878 376168 224884
rect 375840 224664 375892 224670
rect 375840 224606 375892 224612
rect 376128 220522 376156 224878
rect 376404 224398 376432 231662
rect 376588 230382 376616 231676
rect 376576 230376 376628 230382
rect 376576 230318 376628 230324
rect 377140 229770 377168 231676
rect 377128 229764 377180 229770
rect 377128 229706 377180 229712
rect 377692 228682 377720 231676
rect 378244 230382 378272 231676
rect 377864 230376 377916 230382
rect 377864 230318 377916 230324
rect 378232 230376 378284 230382
rect 378232 230318 378284 230324
rect 377680 228676 377732 228682
rect 377680 228618 377732 228624
rect 376760 224528 376812 224534
rect 376760 224470 376812 224476
rect 376392 224392 376444 224398
rect 376392 224334 376444 224340
rect 376116 220516 376168 220522
rect 376116 220458 376168 220464
rect 376772 217410 376800 224470
rect 377876 223310 377904 230318
rect 378048 229900 378100 229906
rect 378048 229842 378100 229848
rect 378060 225010 378088 229842
rect 378796 229430 378824 231676
rect 379152 230376 379204 230382
rect 379152 230318 379204 230324
rect 378784 229424 378836 229430
rect 378784 229366 378836 229372
rect 378968 225752 379020 225758
rect 378968 225694 379020 225700
rect 378048 225004 378100 225010
rect 378048 224946 378100 224952
rect 377864 223304 377916 223310
rect 377864 223246 377916 223252
rect 377404 221876 377456 221882
rect 377404 221818 377456 221824
rect 377416 217410 377444 221818
rect 378232 220108 378284 220114
rect 378232 220050 378284 220056
rect 378244 217410 378272 220050
rect 378980 217410 379008 225694
rect 379164 221882 379192 230318
rect 379348 224618 379376 231676
rect 379900 226166 379928 231676
rect 379888 226160 379940 226166
rect 379888 226102 379940 226108
rect 379796 225004 379848 225010
rect 379796 224946 379848 224952
rect 379348 224590 379560 224618
rect 379336 223440 379388 223446
rect 379336 223382 379388 223388
rect 379348 223174 379376 223382
rect 379336 223168 379388 223174
rect 379336 223110 379388 223116
rect 379152 221876 379204 221882
rect 379152 221818 379204 221824
rect 379532 220114 379560 224590
rect 379520 220108 379572 220114
rect 379520 220050 379572 220056
rect 379808 217410 379836 224946
rect 380452 224262 380480 231676
rect 381004 230314 381032 231676
rect 381570 231662 381952 231690
rect 380992 230308 381044 230314
rect 380992 230250 381044 230256
rect 381176 230172 381228 230178
rect 381176 230114 381228 230120
rect 381188 226030 381216 230114
rect 381176 226024 381228 226030
rect 381176 225966 381228 225972
rect 380440 224256 380492 224262
rect 380440 224198 380492 224204
rect 381924 222154 381952 231662
rect 382108 227186 382136 231676
rect 382280 230036 382332 230042
rect 382280 229978 382332 229984
rect 382292 228818 382320 229978
rect 382464 229084 382516 229090
rect 382464 229026 382516 229032
rect 382280 228812 382332 228818
rect 382280 228754 382332 228760
rect 382096 227180 382148 227186
rect 382096 227122 382148 227128
rect 381912 222148 381964 222154
rect 381912 222090 381964 222096
rect 380900 221604 380952 221610
rect 380900 221546 380952 221552
rect 380912 217410 380940 221546
rect 381544 220380 381596 220386
rect 381544 220322 381596 220328
rect 381556 217410 381584 220322
rect 382476 217870 382504 229026
rect 382660 225894 382688 231676
rect 383212 230110 383240 231676
rect 383778 231662 384160 231690
rect 383200 230104 383252 230110
rect 383200 230046 383252 230052
rect 383936 229424 383988 229430
rect 383936 229366 383988 229372
rect 383948 227594 383976 229366
rect 383936 227588 383988 227594
rect 383936 227530 383988 227536
rect 383936 227044 383988 227050
rect 383936 226986 383988 226992
rect 382648 225888 382700 225894
rect 382648 225830 382700 225836
rect 382648 225616 382700 225622
rect 382648 225558 382700 225564
rect 382464 217864 382516 217870
rect 382464 217806 382516 217812
rect 382660 217410 382688 225558
rect 383200 217864 383252 217870
rect 383200 217806 383252 217812
rect 383212 217410 383240 217806
rect 383948 217410 383976 226986
rect 384132 224534 384160 231662
rect 384316 229090 384344 231676
rect 384868 229498 384896 231676
rect 385434 231662 385816 231690
rect 384856 229492 384908 229498
rect 384856 229434 384908 229440
rect 384304 229084 384356 229090
rect 384304 229026 384356 229032
rect 385592 227316 385644 227322
rect 385592 227258 385644 227264
rect 384120 224528 384172 224534
rect 384120 224470 384172 224476
rect 385040 220244 385092 220250
rect 385040 220186 385092 220192
rect 385052 217410 385080 220186
rect 385604 217410 385632 227258
rect 385788 223174 385816 231662
rect 385972 229362 386000 231676
rect 386538 231662 386920 231690
rect 387090 231662 387564 231690
rect 385960 229356 386012 229362
rect 385960 229298 386012 229304
rect 386604 228540 386656 228546
rect 386604 228482 386656 228488
rect 385776 223168 385828 223174
rect 385776 223110 385828 223116
rect 386616 217410 386644 228482
rect 386892 225758 386920 231662
rect 386880 225752 386932 225758
rect 386880 225694 386932 225700
rect 387248 223576 387300 223582
rect 387248 223518 387300 223524
rect 387260 217410 387288 223518
rect 387536 221610 387564 231662
rect 387628 229650 387656 231676
rect 388180 230450 388208 231676
rect 388168 230444 388220 230450
rect 388168 230386 388220 230392
rect 387628 229634 387748 229650
rect 387628 229628 387760 229634
rect 387628 229622 387708 229628
rect 387708 229570 387760 229576
rect 388444 229492 388496 229498
rect 388444 229434 388496 229440
rect 388456 225570 388484 229434
rect 388732 227050 388760 231676
rect 389088 230308 389140 230314
rect 389088 230250 389140 230256
rect 388720 227044 388772 227050
rect 388720 226986 388772 226992
rect 388456 225542 388668 225570
rect 388444 222148 388496 222154
rect 388444 222090 388496 222096
rect 387524 221604 387576 221610
rect 387524 221546 387576 221552
rect 388168 220516 388220 220522
rect 388168 220458 388220 220464
rect 388180 217410 388208 220458
rect 388456 220386 388484 222090
rect 388640 222018 388668 225542
rect 389100 222494 389128 230250
rect 389284 229906 389312 231676
rect 389272 229900 389324 229906
rect 389272 229842 389324 229848
rect 389836 229226 389864 231676
rect 390388 230110 390416 231676
rect 390744 230444 390796 230450
rect 390744 230386 390796 230392
rect 390008 230104 390060 230110
rect 390008 230046 390060 230052
rect 390376 230104 390428 230110
rect 390376 230046 390428 230052
rect 389824 229220 389876 229226
rect 389824 229162 389876 229168
rect 389732 227452 389784 227458
rect 389732 227394 389784 227400
rect 389088 222488 389140 222494
rect 389088 222430 389140 222436
rect 388628 222012 388680 222018
rect 388628 221954 388680 221960
rect 389180 221740 389232 221746
rect 389180 221682 389232 221688
rect 388444 220380 388496 220386
rect 388444 220322 388496 220328
rect 389192 217410 389220 221682
rect 389744 217410 389772 227394
rect 390020 222630 390048 230046
rect 390756 229974 390784 230386
rect 390744 229968 390796 229974
rect 390744 229910 390796 229916
rect 390468 229900 390520 229906
rect 390468 229842 390520 229848
rect 390008 222624 390060 222630
rect 390008 222566 390060 222572
rect 390480 221746 390508 229842
rect 390940 228954 390968 231676
rect 391492 230382 391520 231676
rect 391480 230376 391532 230382
rect 391480 230318 391532 230324
rect 391756 229628 391808 229634
rect 391756 229570 391808 229576
rect 390928 228948 390980 228954
rect 390928 228890 390980 228896
rect 390744 228812 390796 228818
rect 390744 228754 390796 228760
rect 390468 221740 390520 221746
rect 390468 221682 390520 221688
rect 390756 217870 390784 228754
rect 390928 222896 390980 222902
rect 390928 222838 390980 222844
rect 390744 217864 390796 217870
rect 390744 217806 390796 217812
rect 390940 217410 390968 222838
rect 391768 222766 391796 229570
rect 392044 229362 392072 231676
rect 392610 231662 393084 231690
rect 392584 230376 392636 230382
rect 392584 230318 392636 230324
rect 392216 229832 392268 229838
rect 392216 229774 392268 229780
rect 392228 229498 392256 229774
rect 392216 229492 392268 229498
rect 392216 229434 392268 229440
rect 392032 229356 392084 229362
rect 392032 229298 392084 229304
rect 392216 223032 392268 223038
rect 392216 222974 392268 222980
rect 391756 222760 391808 222766
rect 391756 222702 391808 222708
rect 391480 217864 391532 217870
rect 391480 217806 391532 217812
rect 391492 217410 391520 217806
rect 392228 217410 392256 222974
rect 392596 221338 392624 230318
rect 392860 229220 392912 229226
rect 392860 229162 392912 229168
rect 392872 223582 392900 229162
rect 392860 223576 392912 223582
rect 392860 223518 392912 223524
rect 392584 221332 392636 221338
rect 392584 221274 392636 221280
rect 393056 220658 393084 231662
rect 393148 229094 393176 231676
rect 393148 229066 393268 229094
rect 393240 228546 393268 229066
rect 393228 228540 393280 228546
rect 393228 228482 393280 228488
rect 393320 228404 393372 228410
rect 393320 228346 393372 228352
rect 393044 220652 393096 220658
rect 393044 220594 393096 220600
rect 393332 217870 393360 228346
rect 393700 225622 393728 231676
rect 394252 230246 394280 231676
rect 394818 231662 395200 231690
rect 394056 230240 394108 230246
rect 394056 230182 394108 230188
rect 394240 230240 394292 230246
rect 394240 230182 394292 230188
rect 394068 229566 394096 230182
rect 395172 229906 395200 231662
rect 395160 229900 395212 229906
rect 395160 229842 395212 229848
rect 394700 229832 394752 229838
rect 394700 229774 394752 229780
rect 394056 229560 394108 229566
rect 394056 229502 394108 229508
rect 394056 229356 394108 229362
rect 394056 229298 394108 229304
rect 393688 225616 393740 225622
rect 393688 225558 393740 225564
rect 393504 223440 393556 223446
rect 393504 223382 393556 223388
rect 393320 217864 393372 217870
rect 393320 217806 393372 217812
rect 393516 217410 393544 223382
rect 394068 223038 394096 229298
rect 394712 224806 394740 229774
rect 395160 229696 395212 229702
rect 395160 229638 395212 229644
rect 394884 226024 394936 226030
rect 394884 225966 394936 225972
rect 394700 224800 394752 224806
rect 394700 224742 394752 224748
rect 394056 223032 394108 223038
rect 394056 222974 394108 222980
rect 393964 217864 394016 217870
rect 393964 217806 394016 217812
rect 344296 217382 344632 217410
rect 345400 217382 345460 217410
rect 345952 217382 346288 217410
rect 346688 217382 347116 217410
rect 347884 217382 347944 217410
rect 348344 217382 348772 217410
rect 349264 217382 349600 217410
rect 350000 217382 350428 217410
rect 350920 217382 351256 217410
rect 351932 217382 352084 217410
rect 352484 217382 352912 217410
rect 353496 217382 353740 217410
rect 354232 217382 354568 217410
rect 355060 217382 355396 217410
rect 356164 217382 356224 217410
rect 356716 217382 357052 217410
rect 357452 217382 357880 217410
rect 358372 217382 358708 217410
rect 359108 217382 359536 217410
rect 360212 217382 360364 217410
rect 360764 217382 361192 217410
rect 361684 217382 362020 217410
rect 362512 217382 362848 217410
rect 363248 217382 363676 217410
rect 364352 217382 364504 217410
rect 365180 217382 365332 217410
rect 365824 217382 366160 217410
rect 366652 217382 366988 217410
rect 367388 217382 367816 217410
rect 368492 217382 368644 217410
rect 369044 217382 369472 217410
rect 369872 217382 370300 217410
rect 370792 217382 371128 217410
rect 371528 217382 371956 217410
rect 372724 217382 372784 217410
rect 373184 217382 373612 217410
rect 374196 217382 374440 217410
rect 374932 217382 375268 217410
rect 375668 217382 376096 217410
rect 376772 217382 376924 217410
rect 377416 217382 377752 217410
rect 378244 217382 378580 217410
rect 378980 217382 379408 217410
rect 379808 217382 380236 217410
rect 380912 217382 381064 217410
rect 381556 217382 381892 217410
rect 382660 217382 382720 217410
rect 383212 217382 383548 217410
rect 383948 217382 384376 217410
rect 385052 217382 385204 217410
rect 385604 217382 386032 217410
rect 386616 217382 386860 217410
rect 387260 217382 387688 217410
rect 388180 217382 388516 217410
rect 389192 217382 389344 217410
rect 389744 217382 390172 217410
rect 390940 217382 391000 217410
rect 391492 217382 391828 217410
rect 392228 217382 392656 217410
rect 393484 217382 393544 217410
rect 393976 217410 394004 217806
rect 394896 217410 394924 225966
rect 395172 220794 395200 229638
rect 395356 227458 395384 231676
rect 395908 230382 395936 231676
rect 395896 230376 395948 230382
rect 395896 230318 395948 230324
rect 396460 229770 396488 231676
rect 397026 231662 397408 231690
rect 396724 230376 396776 230382
rect 396724 230318 396776 230324
rect 396448 229764 396500 229770
rect 396448 229706 396500 229712
rect 395344 227452 395396 227458
rect 395344 227394 395396 227400
rect 396356 223304 396408 223310
rect 396356 223246 396408 223252
rect 395620 221468 395672 221474
rect 395620 221410 395672 221416
rect 395160 220788 395212 220794
rect 395160 220730 395212 220736
rect 395632 217410 395660 221410
rect 396368 217410 396396 223246
rect 396736 221202 396764 230318
rect 397184 230240 397236 230246
rect 397184 230182 397236 230188
rect 397196 223310 397224 230182
rect 397184 223304 397236 223310
rect 397184 223246 397236 223252
rect 396724 221196 396776 221202
rect 396724 221138 396776 221144
rect 397380 220522 397408 231662
rect 397564 228410 397592 231676
rect 398130 231662 398604 231690
rect 397920 230036 397972 230042
rect 397920 229978 397972 229984
rect 397552 228404 397604 228410
rect 397552 228346 397604 228352
rect 397932 224670 397960 229978
rect 397552 224664 397604 224670
rect 397552 224606 397604 224612
rect 397920 224664 397972 224670
rect 397920 224606 397972 224612
rect 397368 220516 397420 220522
rect 397368 220458 397420 220464
rect 397564 217410 397592 224606
rect 398576 221474 398604 231662
rect 398668 230194 398696 231676
rect 398668 230178 398788 230194
rect 398668 230172 398800 230178
rect 398668 230166 398748 230172
rect 398748 230114 398800 230120
rect 399220 230042 399248 231676
rect 399208 230036 399260 230042
rect 399208 229978 399260 229984
rect 399484 229560 399536 229566
rect 399484 229502 399536 229508
rect 398840 227588 398892 227594
rect 398840 227530 398892 227536
rect 398564 221468 398616 221474
rect 398564 221410 398616 221416
rect 398104 220788 398156 220794
rect 398104 220730 398156 220736
rect 398116 217410 398144 220730
rect 398852 217870 398880 227530
rect 399024 224392 399076 224398
rect 399024 224334 399076 224340
rect 398840 217864 398892 217870
rect 398840 217806 398892 217812
rect 399036 217410 399064 224334
rect 399496 224126 399524 229502
rect 399772 226914 399800 231676
rect 400338 231662 400720 231690
rect 400496 228676 400548 228682
rect 400496 228618 400548 228624
rect 399760 226908 399812 226914
rect 399760 226850 399812 226856
rect 399484 224120 399536 224126
rect 399484 224062 399536 224068
rect 399760 217864 399812 217870
rect 399760 217806 399812 217812
rect 399772 217410 399800 217806
rect 400508 217410 400536 228618
rect 400692 226030 400720 231662
rect 400876 229906 400904 231676
rect 400864 229900 400916 229906
rect 400864 229842 400916 229848
rect 400680 226024 400732 226030
rect 400680 225966 400732 225972
rect 401428 220250 401456 231676
rect 401692 229764 401744 229770
rect 401692 229706 401744 229712
rect 401704 223446 401732 229706
rect 401980 228818 402008 231676
rect 402546 231662 402744 231690
rect 401968 228812 402020 228818
rect 401968 228754 402020 228760
rect 401692 223440 401744 223446
rect 401692 223382 401744 223388
rect 402716 222154 402744 231662
rect 403084 229498 403112 231676
rect 403256 230444 403308 230450
rect 403256 230386 403308 230392
rect 403072 229492 403124 229498
rect 403072 229434 403124 229440
rect 402980 226160 403032 226166
rect 402980 226102 403032 226108
rect 402704 222148 402756 222154
rect 402704 222090 402756 222096
rect 402244 221876 402296 221882
rect 402244 221818 402296 221824
rect 401416 220244 401468 220250
rect 401416 220186 401468 220192
rect 401600 220108 401652 220114
rect 401600 220050 401652 220056
rect 401612 217410 401640 220050
rect 402256 217410 402284 221818
rect 402992 217870 403020 226102
rect 403268 223990 403296 230386
rect 403636 230382 403664 231676
rect 403624 230376 403676 230382
rect 403624 230318 403676 230324
rect 404188 228682 404216 231676
rect 404740 229634 404768 231676
rect 405004 230376 405056 230382
rect 405004 230318 405056 230324
rect 404728 229628 404780 229634
rect 404728 229570 404780 229576
rect 404176 228676 404228 228682
rect 404176 228618 404228 228624
rect 403256 223984 403308 223990
rect 403256 223926 403308 223932
rect 403164 222488 403216 222494
rect 403164 222430 403216 222436
rect 402980 217864 403032 217870
rect 402980 217806 403032 217812
rect 403176 217410 403204 222430
rect 405016 220386 405044 230318
rect 405292 222902 405320 231676
rect 405844 229770 405872 231676
rect 406396 230382 406424 231676
rect 406384 230376 406436 230382
rect 406384 230318 406436 230324
rect 406660 230036 406712 230042
rect 406660 229978 406712 229984
rect 405832 229764 405884 229770
rect 405832 229706 405884 229712
rect 406672 224262 406700 229978
rect 405740 224256 405792 224262
rect 405740 224198 405792 224204
rect 406660 224256 406712 224262
rect 406660 224198 406712 224204
rect 405280 222896 405332 222902
rect 405280 222838 405332 222844
rect 404728 220380 404780 220386
rect 404728 220322 404780 220328
rect 405004 220380 405056 220386
rect 405004 220322 405056 220328
rect 403900 217864 403952 217870
rect 403900 217806 403952 217812
rect 403912 217410 403940 217806
rect 404740 217410 404768 220322
rect 405752 217410 405780 224198
rect 406948 222630 406976 231676
rect 407304 227180 407356 227186
rect 407304 227122 407356 227128
rect 406292 222624 406344 222630
rect 406292 222566 406344 222572
rect 406936 222624 406988 222630
rect 406936 222566 406988 222572
rect 406304 217410 406332 222566
rect 407316 217410 407344 227122
rect 407500 225214 407528 231676
rect 408052 229094 408080 231676
rect 408408 230376 408460 230382
rect 408408 230318 408460 230324
rect 408052 229066 408172 229094
rect 407488 225208 407540 225214
rect 407488 225150 407540 225156
rect 407948 224528 408000 224534
rect 407948 224470 408000 224476
rect 407960 217410 407988 224470
rect 408144 220114 408172 229066
rect 408420 227730 408448 230318
rect 408408 227724 408460 227730
rect 408408 227666 408460 227672
rect 408604 226166 408632 231676
rect 409170 231662 409644 231690
rect 408776 230444 408828 230450
rect 408776 230386 408828 230392
rect 408788 229634 408816 230386
rect 408776 229628 408828 229634
rect 408776 229570 408828 229576
rect 408592 226160 408644 226166
rect 408592 226102 408644 226108
rect 408776 225888 408828 225894
rect 408776 225830 408828 225836
rect 408132 220108 408184 220114
rect 408132 220050 408184 220056
rect 408788 217410 408816 225830
rect 409616 221882 409644 231662
rect 409708 230058 409736 231676
rect 409708 230042 409828 230058
rect 409708 230036 409840 230042
rect 409708 230030 409788 230036
rect 409788 229978 409840 229984
rect 409788 229764 409840 229770
rect 409788 229706 409840 229712
rect 409800 224942 409828 229706
rect 410260 229226 410288 231676
rect 410248 229220 410300 229226
rect 410248 229162 410300 229168
rect 410432 229084 410484 229090
rect 410432 229026 410484 229032
rect 409788 224936 409840 224942
rect 409788 224878 409840 224884
rect 409972 223168 410024 223174
rect 409972 223110 410024 223116
rect 409604 221876 409656 221882
rect 409604 221818 409656 221824
rect 409984 217410 410012 223110
rect 410444 217410 410472 229026
rect 410812 225486 410840 231676
rect 411378 231662 411760 231690
rect 410800 225480 410852 225486
rect 410800 225422 410852 225428
rect 411260 224800 411312 224806
rect 411260 224742 411312 224748
rect 411272 217410 411300 224742
rect 411732 222494 411760 231662
rect 411916 223174 411944 231676
rect 412468 224806 412496 231676
rect 412732 229220 412784 229226
rect 412732 229162 412784 229168
rect 412456 224800 412508 224806
rect 412456 224742 412508 224748
rect 412744 223854 412772 229162
rect 413020 226302 413048 231676
rect 413192 230172 413244 230178
rect 413192 230114 413244 230120
rect 413008 226296 413060 226302
rect 413008 226238 413060 226244
rect 412732 223848 412784 223854
rect 412732 223790 412784 223796
rect 411904 223168 411956 223174
rect 411904 223110 411956 223116
rect 413204 222766 413232 230114
rect 413572 229362 413600 231676
rect 414124 230314 414152 231676
rect 414112 230308 414164 230314
rect 414112 230250 414164 230256
rect 413560 229356 413612 229362
rect 413560 229298 413612 229304
rect 414676 229094 414704 231676
rect 414676 229066 414796 229094
rect 414020 225752 414072 225758
rect 414020 225694 414072 225700
rect 412916 222760 412968 222766
rect 412916 222702 412968 222708
rect 413192 222760 413244 222766
rect 413192 222702 413244 222708
rect 411720 222488 411772 222494
rect 411720 222430 411772 222436
rect 412180 222012 412232 222018
rect 412180 221954 412232 221960
rect 412192 217410 412220 221954
rect 412928 217410 412956 222702
rect 414032 217410 414060 225694
rect 414768 224670 414796 229066
rect 415228 227594 415256 231676
rect 415216 227588 415268 227594
rect 415216 227530 415268 227536
rect 415780 227322 415808 231676
rect 416044 230444 416096 230450
rect 416044 230386 416096 230392
rect 415768 227316 415820 227322
rect 415768 227258 415820 227264
rect 414572 224664 414624 224670
rect 414572 224606 414624 224612
rect 414756 224664 414808 224670
rect 414756 224606 414808 224612
rect 414584 217410 414612 224606
rect 415584 221604 415636 221610
rect 415584 221546 415636 221552
rect 415596 217410 415624 221546
rect 416056 221066 416084 230386
rect 416332 223718 416360 231676
rect 416884 229634 416912 231676
rect 417240 229900 417292 229906
rect 417240 229842 417292 229848
rect 416872 229628 416924 229634
rect 416872 229570 416924 229576
rect 417252 229498 417280 229842
rect 417240 229492 417292 229498
rect 417240 229434 417292 229440
rect 417056 227044 417108 227050
rect 417056 226986 417108 226992
rect 416320 223712 416372 223718
rect 416320 223654 416372 223660
rect 416228 223576 416280 223582
rect 416228 223518 416280 223524
rect 416044 221060 416096 221066
rect 416044 221002 416096 221008
rect 416240 217410 416268 223518
rect 417068 217410 417096 226986
rect 417436 225350 417464 231676
rect 417804 231662 418002 231690
rect 417424 225344 417476 225350
rect 417424 225286 417476 225292
rect 417804 222018 417832 231662
rect 418540 229226 418568 231676
rect 419092 229498 419120 231676
rect 419080 229492 419132 229498
rect 419080 229434 419132 229440
rect 418804 229356 418856 229362
rect 418804 229298 418856 229304
rect 418528 229220 418580 229226
rect 418528 229162 418580 229168
rect 418816 229094 418844 229298
rect 418816 229066 419028 229094
rect 418160 224120 418212 224126
rect 418160 224062 418212 224068
rect 417792 222012 417844 222018
rect 417792 221954 417844 221960
rect 418172 217410 418200 224062
rect 418804 221740 418856 221746
rect 418804 221682 418856 221688
rect 418816 217410 418844 221682
rect 419000 220930 419028 229066
rect 419644 229022 419672 231676
rect 419632 229016 419684 229022
rect 419632 228958 419684 228964
rect 419448 228948 419500 228954
rect 419448 228890 419500 228896
rect 419460 228834 419488 228890
rect 419460 228806 419580 228834
rect 418988 220924 419040 220930
rect 418988 220866 419040 220872
rect 419552 217870 419580 228806
rect 420196 227186 420224 231676
rect 420748 230178 420776 231676
rect 421300 230450 421328 231676
rect 421288 230444 421340 230450
rect 421288 230386 421340 230392
rect 420736 230172 420788 230178
rect 420736 230114 420788 230120
rect 420920 229764 420972 229770
rect 420920 229706 420972 229712
rect 420184 227180 420236 227186
rect 420184 227122 420236 227128
rect 419724 223032 419776 223038
rect 419724 222974 419776 222980
rect 419540 217864 419592 217870
rect 419540 217806 419592 217812
rect 419736 217410 419764 222974
rect 420932 222358 420960 229706
rect 421852 229634 421880 231676
rect 422404 230450 422432 231676
rect 422970 231662 423352 231690
rect 422208 230444 422260 230450
rect 422208 230386 422260 230392
rect 422392 230444 422444 230450
rect 422392 230386 422444 230392
rect 421840 229628 421892 229634
rect 421840 229570 421892 229576
rect 421104 225208 421156 225214
rect 421104 225150 421156 225156
rect 420920 222352 420972 222358
rect 420920 222294 420972 222300
rect 421116 219706 421144 225150
rect 422220 221746 422248 230386
rect 422944 229288 422996 229294
rect 422944 229230 422996 229236
rect 422956 229094 422984 229230
rect 423324 229094 423352 231662
rect 423508 229094 423536 231676
rect 422956 229066 423260 229094
rect 423324 229066 423444 229094
rect 423508 229066 423720 229094
rect 423036 225616 423088 225622
rect 423036 225558 423088 225564
rect 422852 223304 422904 223310
rect 422852 223246 422904 223252
rect 422208 221740 422260 221746
rect 422208 221682 422260 221688
rect 422300 221332 422352 221338
rect 422300 221274 422352 221280
rect 421288 220652 421340 220658
rect 421288 220594 421340 220600
rect 421104 219700 421156 219706
rect 421104 219642 421156 219648
rect 420460 217864 420512 217870
rect 420460 217806 420512 217812
rect 420472 217410 420500 217806
rect 421300 217410 421328 220594
rect 422312 217410 422340 221274
rect 422864 217410 422892 223246
rect 423048 220794 423076 225558
rect 423232 221338 423260 229066
rect 423416 224534 423444 229066
rect 423404 224528 423456 224534
rect 423404 224470 423456 224476
rect 423692 224398 423720 229066
rect 424060 228954 424088 231676
rect 424232 229900 424284 229906
rect 424232 229842 424284 229848
rect 424048 228948 424100 228954
rect 424048 228890 424100 228896
rect 423956 228540 424008 228546
rect 423956 228482 424008 228488
rect 423680 224392 423732 224398
rect 423680 224334 423732 224340
rect 423772 222624 423824 222630
rect 423772 222566 423824 222572
rect 423220 221332 423272 221338
rect 423220 221274 423272 221280
rect 423036 220788 423088 220794
rect 423036 220730 423088 220736
rect 423784 219570 423812 222566
rect 423772 219564 423824 219570
rect 423772 219506 423824 219512
rect 423968 219434 423996 228482
rect 424244 223582 424272 229842
rect 424612 229226 424640 231676
rect 424600 229220 424652 229226
rect 424600 229162 424652 229168
rect 425164 226030 425192 231676
rect 425730 231662 426112 231690
rect 425520 229764 425572 229770
rect 425520 229706 425572 229712
rect 425152 226024 425204 226030
rect 425152 225966 425204 225972
rect 425532 223990 425560 229706
rect 425796 225888 425848 225894
rect 425796 225830 425848 225836
rect 424692 223984 424744 223990
rect 424692 223926 424744 223932
rect 425520 223984 425572 223990
rect 425520 223926 425572 223932
rect 424232 223576 424284 223582
rect 424232 223518 424284 223524
rect 423876 219406 423996 219434
rect 423876 217410 423904 219406
rect 424704 217410 424732 223926
rect 425428 220788 425480 220794
rect 425428 220730 425480 220736
rect 425440 217410 425468 220730
rect 425808 220658 425836 225830
rect 426084 223038 426112 231662
rect 426268 227050 426296 231676
rect 426820 229362 426848 231676
rect 427372 229906 427400 231676
rect 427728 230308 427780 230314
rect 427728 230250 427780 230256
rect 427544 230036 427596 230042
rect 427544 229978 427596 229984
rect 427360 229900 427412 229906
rect 427360 229842 427412 229848
rect 426808 229356 426860 229362
rect 426808 229298 426860 229304
rect 426440 227452 426492 227458
rect 426440 227394 426492 227400
rect 426256 227044 426308 227050
rect 426256 226986 426308 226992
rect 426072 223032 426124 223038
rect 426072 222974 426124 222980
rect 425796 220652 425848 220658
rect 425796 220594 425848 220600
rect 426452 217870 426480 227394
rect 426624 223440 426676 223446
rect 426624 223382 426676 223388
rect 426440 217864 426492 217870
rect 426440 217806 426492 217812
rect 426636 217410 426664 223382
rect 427556 223310 427584 229978
rect 427740 226778 427768 230250
rect 427728 226772 427780 226778
rect 427728 226714 427780 226720
rect 427924 225894 427952 231676
rect 428476 228274 428504 231676
rect 429028 229770 429056 231676
rect 429580 230314 429608 231676
rect 430146 231662 430436 231690
rect 429568 230308 429620 230314
rect 429568 230250 429620 230256
rect 429016 229764 429068 229770
rect 429016 229706 429068 229712
rect 430028 229764 430080 229770
rect 430028 229706 430080 229712
rect 430212 229764 430264 229770
rect 430212 229706 430264 229712
rect 430040 229498 430068 229706
rect 429844 229492 429896 229498
rect 429844 229434 429896 229440
rect 430028 229492 430080 229498
rect 430028 229434 430080 229440
rect 428464 228268 428516 228274
rect 428464 228210 428516 228216
rect 427912 225888 427964 225894
rect 427912 225830 427964 225836
rect 429856 224126 429884 229434
rect 430224 229226 430252 229706
rect 430212 229220 430264 229226
rect 430212 229162 430264 229168
rect 429844 224120 429896 224126
rect 429844 224062 429896 224068
rect 429200 223712 429252 223718
rect 429200 223654 429252 223660
rect 427544 223304 427596 223310
rect 427544 223246 427596 223252
rect 428096 222488 428148 222494
rect 428096 222430 428148 222436
rect 427912 220516 427964 220522
rect 427912 220458 427964 220464
rect 427084 217864 427136 217870
rect 427084 217806 427136 217812
rect 393976 217382 394312 217410
rect 394896 217382 395140 217410
rect 395632 217382 395968 217410
rect 396368 217382 396796 217410
rect 397564 217382 397624 217410
rect 398116 217382 398452 217410
rect 399036 217382 399280 217410
rect 399772 217382 400108 217410
rect 400508 217382 400936 217410
rect 401612 217382 401764 217410
rect 402256 217382 402592 217410
rect 403176 217382 403420 217410
rect 403912 217382 404248 217410
rect 404740 217382 405076 217410
rect 405752 217382 405904 217410
rect 406304 217382 406732 217410
rect 407316 217382 407560 217410
rect 407960 217382 408388 217410
rect 408788 217382 409216 217410
rect 409984 217382 410044 217410
rect 410444 217382 410872 217410
rect 411272 217382 411700 217410
rect 412192 217382 412528 217410
rect 412928 217382 413356 217410
rect 414032 217382 414184 217410
rect 414584 217382 415012 217410
rect 415596 217382 415840 217410
rect 416240 217382 416668 217410
rect 417068 217382 417496 217410
rect 418172 217382 418324 217410
rect 418816 217382 419152 217410
rect 419736 217382 419980 217410
rect 420472 217382 420808 217410
rect 421300 217382 421636 217410
rect 422312 217382 422464 217410
rect 422864 217382 423292 217410
rect 423876 217382 424120 217410
rect 424704 217382 424948 217410
rect 425440 217382 425776 217410
rect 426604 217382 426664 217410
rect 427096 217410 427124 217806
rect 427924 217410 427952 220458
rect 428108 219978 428136 222430
rect 428740 221196 428792 221202
rect 428740 221138 428792 221144
rect 428096 219972 428148 219978
rect 428096 219914 428148 219920
rect 428752 217410 428780 221138
rect 429212 220794 429240 223654
rect 429476 222760 429528 222766
rect 429476 222702 429528 222708
rect 429200 220788 429252 220794
rect 429200 220730 429252 220736
rect 429488 217410 429516 222702
rect 430408 219434 430436 231662
rect 430684 229226 430712 231676
rect 431250 231662 431724 231690
rect 431696 229378 431724 231662
rect 431788 230058 431816 231676
rect 432340 230314 432368 231676
rect 432144 230308 432196 230314
rect 432144 230250 432196 230256
rect 432328 230308 432380 230314
rect 432328 230250 432380 230256
rect 431788 230042 431908 230058
rect 431788 230036 431920 230042
rect 431788 230030 431868 230036
rect 431868 229978 431920 229984
rect 431696 229350 431816 229378
rect 430672 229220 430724 229226
rect 430672 229162 430724 229168
rect 431592 229220 431644 229226
rect 431592 229162 431644 229168
rect 430580 228404 430632 228410
rect 430580 228346 430632 228352
rect 430396 219428 430448 219434
rect 430396 219370 430448 219376
rect 430592 217410 430620 228346
rect 431132 224256 431184 224262
rect 431132 224198 431184 224204
rect 431144 217410 431172 224198
rect 431604 219298 431632 229162
rect 431592 219292 431644 219298
rect 431592 219234 431644 219240
rect 431788 219162 431816 229350
rect 432156 227458 432184 230250
rect 432892 229906 432920 231676
rect 432604 229900 432656 229906
rect 432604 229842 432656 229848
rect 432880 229900 432932 229906
rect 432880 229842 432932 229848
rect 432420 229492 432472 229498
rect 432420 229434 432472 229440
rect 432432 229226 432460 229434
rect 432420 229220 432472 229226
rect 432420 229162 432472 229168
rect 432616 228546 432644 229842
rect 433444 229226 433472 231676
rect 433616 229764 433668 229770
rect 433616 229706 433668 229712
rect 433800 229764 433852 229770
rect 433800 229706 433852 229712
rect 433432 229220 433484 229226
rect 433432 229162 433484 229168
rect 432604 228540 432656 228546
rect 432604 228482 432656 228488
rect 433628 228410 433656 229706
rect 433812 229362 433840 229706
rect 433800 229356 433852 229362
rect 433800 229298 433852 229304
rect 433616 228404 433668 228410
rect 433616 228346 433668 228352
rect 432144 227452 432196 227458
rect 432144 227394 432196 227400
rect 433616 226908 433668 226914
rect 433616 226850 433668 226856
rect 432788 222352 432840 222358
rect 432788 222294 432840 222300
rect 432052 221468 432104 221474
rect 432052 221410 432104 221416
rect 431776 219156 431828 219162
rect 431776 219098 431828 219104
rect 432064 217410 432092 221410
rect 432800 217410 432828 222294
rect 433628 217410 433656 226850
rect 433996 225622 434024 231676
rect 434548 229362 434576 231676
rect 434536 229356 434588 229362
rect 434536 229298 434588 229304
rect 435100 229226 435128 231676
rect 434352 229220 434404 229226
rect 434352 229162 434404 229168
rect 435088 229220 435140 229226
rect 435088 229162 435140 229168
rect 433984 225616 434036 225622
rect 433984 225558 434036 225564
rect 434364 219026 434392 229162
rect 434720 228812 434772 228818
rect 434720 228754 434772 228760
rect 434732 220522 434760 228754
rect 435652 224262 435680 231676
rect 436218 231662 436600 231690
rect 436192 229764 436244 229770
rect 436192 229706 436244 229712
rect 436008 229220 436060 229226
rect 436008 229162 436060 229168
rect 435640 224256 435692 224262
rect 435640 224198 435692 224204
rect 436020 221474 436048 229162
rect 436204 226914 436232 229706
rect 436192 226908 436244 226914
rect 436192 226850 436244 226856
rect 436192 223576 436244 223582
rect 436192 223518 436244 223524
rect 436008 221468 436060 221474
rect 436008 221410 436060 221416
rect 435548 220652 435600 220658
rect 435548 220594 435600 220600
rect 434720 220516 434772 220522
rect 434720 220458 434772 220464
rect 434812 220244 434864 220250
rect 434812 220186 434864 220192
rect 434352 219020 434404 219026
rect 434352 218962 434404 218968
rect 434824 217410 434852 220186
rect 435560 217410 435588 220594
rect 436204 217410 436232 223518
rect 436572 223446 436600 231662
rect 436756 229226 436784 231676
rect 436744 229220 436796 229226
rect 436744 229162 436796 229168
rect 436744 225344 436796 225350
rect 436744 225286 436796 225292
rect 436560 223440 436612 223446
rect 436560 223382 436612 223388
rect 436756 219706 436784 225286
rect 437308 221241 437336 231676
rect 437874 231662 438256 231690
rect 438032 230580 438084 230586
rect 438032 230522 438084 230528
rect 437848 230308 437900 230314
rect 437848 230250 437900 230256
rect 437860 229906 437888 230250
rect 438044 229906 438072 230522
rect 437848 229900 437900 229906
rect 437848 229842 437900 229848
rect 438032 229900 438084 229906
rect 438032 229842 438084 229848
rect 438032 229764 438084 229770
rect 438032 229706 438084 229712
rect 438044 229362 438072 229706
rect 438032 229356 438084 229362
rect 438032 229298 438084 229304
rect 438228 225758 438256 231662
rect 438216 225752 438268 225758
rect 438216 225694 438268 225700
rect 437480 225480 437532 225486
rect 437480 225422 437532 225428
rect 437294 221232 437350 221241
rect 437294 221167 437350 221176
rect 437020 220516 437072 220522
rect 437020 220458 437072 220464
rect 436744 219700 436796 219706
rect 436744 219642 436796 219648
rect 437032 217410 437060 220458
rect 437492 220250 437520 225422
rect 438412 222426 438440 231676
rect 438964 229634 438992 231676
rect 439530 231662 439912 231690
rect 438584 229628 438636 229634
rect 438584 229570 438636 229576
rect 438952 229628 439004 229634
rect 438952 229570 439004 229576
rect 438596 229362 438624 229570
rect 438584 229356 438636 229362
rect 438584 229298 438636 229304
rect 439596 229356 439648 229362
rect 439596 229298 439648 229304
rect 439412 222896 439464 222902
rect 439412 222838 439464 222844
rect 438400 222420 438452 222426
rect 438400 222362 438452 222368
rect 438860 222148 438912 222154
rect 438860 222090 438912 222096
rect 437848 220380 437900 220386
rect 437848 220322 437900 220328
rect 437480 220244 437532 220250
rect 437480 220186 437532 220192
rect 437860 217410 437888 220322
rect 438872 217410 438900 222090
rect 439424 217410 439452 222838
rect 439608 221202 439636 229298
rect 439884 222902 439912 231662
rect 440068 225214 440096 231676
rect 440620 229362 440648 231676
rect 441172 229634 441200 231676
rect 441738 231662 442120 231690
rect 442290 231662 442672 231690
rect 441896 229900 441948 229906
rect 441896 229842 441948 229848
rect 441160 229628 441212 229634
rect 441160 229570 441212 229576
rect 440792 229492 440844 229498
rect 440792 229434 440844 229440
rect 440608 229356 440660 229362
rect 440608 229298 440660 229304
rect 440424 228676 440476 228682
rect 440424 228618 440476 228624
rect 440056 225208 440108 225214
rect 440056 225150 440108 225156
rect 439872 222896 439924 222902
rect 439872 222838 439924 222844
rect 439596 221196 439648 221202
rect 439596 221138 439648 221144
rect 440436 217410 440464 228618
rect 440804 228138 440832 229434
rect 441436 229356 441488 229362
rect 441436 229298 441488 229304
rect 440792 228132 440844 228138
rect 440792 228074 440844 228080
rect 441068 224936 441120 224942
rect 441068 224878 441120 224884
rect 441080 217410 441108 224878
rect 441448 220386 441476 229298
rect 441908 228682 441936 229842
rect 441896 228676 441948 228682
rect 441896 228618 441948 228624
rect 442092 222766 442120 231662
rect 442264 230444 442316 230450
rect 442264 230386 442316 230392
rect 442276 229906 442304 230386
rect 442264 229900 442316 229906
rect 442264 229842 442316 229848
rect 442264 229084 442316 229090
rect 442264 229026 442316 229032
rect 442276 228818 442304 229026
rect 442264 228812 442316 228818
rect 442264 228754 442316 228760
rect 442644 225350 442672 231662
rect 442632 225344 442684 225350
rect 442632 225286 442684 225292
rect 442828 224942 442856 231676
rect 443394 231662 443776 231690
rect 443552 227724 443604 227730
rect 443552 227666 443604 227672
rect 442816 224936 442868 224942
rect 442816 224878 442868 224884
rect 442080 222760 442132 222766
rect 442080 222702 442132 222708
rect 442908 222420 442960 222426
rect 442908 222362 442960 222368
rect 441988 221060 442040 221066
rect 441988 221002 442040 221008
rect 441436 220380 441488 220386
rect 441436 220322 441488 220328
rect 442000 217410 442028 221002
rect 442920 220153 442948 222362
rect 442906 220144 442962 220153
rect 442906 220079 442962 220088
rect 443000 219836 443052 219842
rect 443000 219778 443052 219784
rect 443012 217410 443040 219778
rect 443564 217410 443592 227666
rect 443748 223582 443776 231662
rect 443932 230450 443960 231676
rect 443920 230444 443972 230450
rect 443920 230386 443972 230392
rect 444484 229362 444512 231676
rect 444852 231662 445050 231690
rect 445496 231662 445602 231690
rect 444472 229356 444524 229362
rect 444472 229298 444524 229304
rect 443736 223576 443788 223582
rect 443736 223518 443788 223524
rect 444196 223576 444248 223582
rect 444196 223518 444248 223524
rect 444208 223174 444236 223518
rect 444012 223168 444064 223174
rect 444012 223110 444064 223116
rect 444196 223168 444248 223174
rect 444196 223110 444248 223116
rect 444024 220658 444052 223110
rect 444852 222358 444880 231662
rect 445300 224528 445352 224534
rect 445300 224470 445352 224476
rect 444840 222352 444892 222358
rect 444840 222294 444892 222300
rect 444012 220652 444064 220658
rect 444012 220594 444064 220600
rect 445312 220522 445340 224470
rect 445300 220516 445352 220522
rect 445300 220458 445352 220464
rect 444564 220108 444616 220114
rect 444564 220050 444616 220056
rect 444576 217410 444604 220050
rect 445300 219564 445352 219570
rect 445300 219506 445352 219512
rect 445312 217410 445340 219506
rect 445496 218754 445524 231662
rect 445944 230444 445996 230450
rect 445944 230386 445996 230392
rect 445668 229356 445720 229362
rect 445668 229298 445720 229304
rect 445680 221610 445708 229298
rect 445956 225078 445984 230386
rect 445944 225072 445996 225078
rect 445944 225014 445996 225020
rect 446140 224534 446168 231676
rect 446706 231662 446904 231690
rect 446128 224528 446180 224534
rect 446128 224470 446180 224476
rect 446036 223304 446088 223310
rect 446036 223246 446088 223252
rect 445668 221604 445720 221610
rect 445668 221546 445720 221552
rect 445668 220516 445720 220522
rect 445668 220458 445720 220464
rect 445680 219570 445708 220458
rect 445668 219564 445720 219570
rect 445668 219506 445720 219512
rect 445484 218748 445536 218754
rect 445484 218690 445536 218696
rect 446048 217410 446076 223246
rect 446876 222154 446904 231662
rect 447244 230450 447272 231676
rect 447232 230444 447284 230450
rect 447232 230386 447284 230392
rect 447796 229094 447824 231676
rect 448060 230444 448112 230450
rect 448060 230386 448112 230392
rect 447796 229066 447916 229094
rect 447048 226160 447100 226166
rect 447048 226102 447100 226108
rect 446864 222148 446916 222154
rect 446864 222090 446916 222096
rect 447060 219434 447088 226102
rect 447692 223848 447744 223854
rect 447692 223790 447744 223796
rect 447060 219406 447180 219434
rect 447152 217410 447180 219406
rect 447704 217410 447732 223790
rect 447888 223310 447916 229066
rect 447876 223304 447928 223310
rect 447876 223246 447928 223252
rect 448072 218890 448100 230386
rect 448348 222630 448376 231676
rect 448900 225486 448928 231676
rect 449466 231662 449848 231690
rect 449820 229094 449848 231662
rect 449728 229066 449848 229094
rect 450004 229094 450032 231676
rect 450004 229066 450124 229094
rect 449072 226296 449124 226302
rect 449072 226238 449124 226244
rect 448888 225480 448940 225486
rect 448888 225422 448940 225428
rect 448336 222624 448388 222630
rect 448336 222566 448388 222572
rect 448612 221876 448664 221882
rect 448612 221818 448664 221824
rect 448060 218884 448112 218890
rect 448060 218826 448112 218832
rect 448624 217410 448652 221818
rect 449084 219570 449112 226238
rect 449728 220658 449756 229066
rect 449900 223440 449952 223446
rect 449900 223382 449952 223388
rect 449440 220652 449492 220658
rect 449440 220594 449492 220600
rect 449716 220652 449768 220658
rect 449716 220594 449768 220600
rect 449072 219564 449124 219570
rect 449072 219506 449124 219512
rect 449452 217410 449480 220594
rect 449912 220425 449940 223382
rect 450096 222494 450124 229066
rect 450556 226506 450584 231676
rect 450924 231662 451122 231690
rect 450544 226500 450596 226506
rect 450544 226442 450596 226448
rect 450084 222488 450136 222494
rect 450084 222430 450136 222436
rect 449898 220416 449954 220425
rect 449898 220351 449954 220360
rect 450924 220250 450952 231662
rect 451464 230172 451516 230178
rect 451464 230114 451516 230120
rect 451280 229084 451332 229090
rect 451280 229026 451332 229032
rect 451292 228818 451320 229026
rect 451280 228812 451332 228818
rect 451280 228754 451332 228760
rect 451476 224806 451504 230114
rect 451660 228818 451688 231676
rect 451648 228812 451700 228818
rect 451648 228754 451700 228760
rect 451280 224800 451332 224806
rect 451280 224742 451332 224748
rect 451464 224800 451516 224806
rect 451464 224742 451516 224748
rect 450268 220244 450320 220250
rect 450268 220186 450320 220192
rect 450912 220244 450964 220250
rect 450912 220186 450964 220192
rect 450280 217410 450308 220186
rect 451292 217410 451320 224742
rect 452212 223446 452240 231676
rect 452568 227588 452620 227594
rect 452568 227530 452620 227536
rect 452200 223440 452252 223446
rect 452200 223382 452252 223388
rect 452580 220658 452608 227530
rect 452764 226778 452792 231676
rect 453316 230450 453344 231676
rect 453684 231662 453882 231690
rect 454434 231662 454816 231690
rect 453304 230444 453356 230450
rect 453304 230386 453356 230392
rect 453684 229094 453712 231662
rect 454500 230444 454552 230450
rect 454500 230386 454552 230392
rect 453408 229066 453712 229094
rect 453948 229084 454000 229090
rect 452752 226772 452804 226778
rect 452752 226714 452804 226720
rect 452752 226636 452804 226642
rect 452752 226578 452804 226584
rect 452568 220652 452620 220658
rect 452568 220594 452620 220600
rect 451924 219972 451976 219978
rect 451924 219914 451976 219920
rect 451936 217410 451964 219914
rect 452764 217410 452792 226578
rect 427096 217382 427432 217410
rect 427924 217382 428260 217410
rect 428752 217382 429088 217410
rect 429488 217382 429916 217410
rect 430592 217382 430744 217410
rect 431144 217382 431572 217410
rect 432064 217382 432400 217410
rect 432800 217382 433228 217410
rect 433628 217382 434056 217410
rect 434824 217382 434884 217410
rect 435560 217382 435712 217410
rect 436204 217382 436540 217410
rect 437032 217382 437368 217410
rect 437860 217382 438196 217410
rect 438872 217382 439024 217410
rect 439424 217382 439852 217410
rect 440436 217382 440680 217410
rect 441080 217382 441508 217410
rect 442000 217382 442336 217410
rect 443012 217382 443164 217410
rect 443564 217382 443992 217410
rect 444576 217382 444820 217410
rect 445312 217382 445648 217410
rect 446048 217382 446476 217410
rect 447152 217382 447304 217410
rect 447704 217382 448132 217410
rect 448624 217382 448960 217410
rect 449452 217382 449788 217410
rect 450280 217382 450616 217410
rect 451292 217382 451444 217410
rect 451936 217382 452272 217410
rect 452764 217382 453100 217410
rect 185216 217252 185268 217258
rect 185216 217194 185268 217200
rect 178040 217116 178092 217122
rect 178040 217058 178092 217064
rect 453408 216986 453436 229066
rect 453948 229026 454000 229032
rect 453960 220114 453988 229026
rect 454512 228002 454540 230386
rect 454500 227996 454552 228002
rect 454500 227938 454552 227944
rect 454316 224664 454368 224670
rect 454316 224606 454368 224612
rect 453948 220108 454000 220114
rect 453948 220050 454000 220056
rect 453580 219564 453632 219570
rect 453580 219506 453632 219512
rect 453592 217410 453620 219506
rect 454328 217410 454356 224606
rect 454788 223854 454816 231662
rect 454972 230178 455000 231676
rect 455538 231662 455920 231690
rect 454960 230172 455012 230178
rect 454960 230114 455012 230120
rect 455696 228268 455748 228274
rect 455696 228210 455748 228216
rect 455708 227866 455736 228210
rect 455696 227860 455748 227866
rect 455696 227802 455748 227808
rect 454776 223848 454828 223854
rect 454776 223790 454828 223796
rect 455892 223310 455920 231662
rect 456076 226642 456104 231676
rect 456628 230450 456656 231676
rect 457194 231662 457576 231690
rect 457746 231662 458036 231690
rect 456616 230444 456668 230450
rect 456616 230386 456668 230392
rect 457076 228948 457128 228954
rect 457076 228890 457128 228896
rect 456248 228812 456300 228818
rect 456248 228754 456300 228760
rect 456260 228138 456288 228754
rect 456248 228132 456300 228138
rect 456248 228074 456300 228080
rect 456064 226636 456116 226642
rect 456064 226578 456116 226584
rect 457088 224954 457116 228890
rect 457088 224926 457208 224954
rect 455696 223304 455748 223310
rect 455696 223246 455748 223252
rect 455880 223304 455932 223310
rect 455880 223246 455932 223252
rect 455420 220924 455472 220930
rect 455420 220866 455472 220872
rect 455432 217410 455460 220866
rect 455708 219978 455736 223246
rect 456064 220788 456116 220794
rect 456064 220730 456116 220736
rect 455696 219972 455748 219978
rect 455696 219914 455748 219920
rect 456076 217410 456104 220730
rect 457180 220658 457208 224926
rect 456984 220652 457036 220658
rect 456984 220594 457036 220600
rect 457168 220652 457220 220658
rect 457168 220594 457220 220600
rect 456996 217410 457024 220594
rect 453592 217382 453928 217410
rect 454328 217382 454756 217410
rect 455432 217382 455584 217410
rect 456076 217382 456412 217410
rect 456996 217382 457240 217410
rect 174360 216980 174412 216986
rect 174360 216922 174412 216928
rect 453396 216980 453448 216986
rect 453396 216922 453448 216928
rect 457548 216850 457576 231662
rect 458008 229094 458036 231662
rect 458008 229066 458128 229094
rect 457720 223984 457772 223990
rect 457720 223926 457772 223932
rect 457732 217410 457760 223926
rect 458100 222057 458128 229066
rect 458284 228954 458312 231676
rect 458836 229090 458864 231676
rect 458824 229084 458876 229090
rect 458824 229026 458876 229032
rect 458272 228948 458324 228954
rect 458272 228890 458324 228896
rect 458456 227316 458508 227322
rect 458456 227258 458508 227264
rect 458086 222048 458142 222057
rect 458086 221983 458142 221992
rect 458468 217410 458496 227258
rect 459388 225321 459416 231676
rect 459560 230172 459612 230178
rect 459560 230114 459612 230120
rect 459572 227866 459600 230114
rect 459560 227860 459612 227866
rect 459560 227802 459612 227808
rect 459744 227724 459796 227730
rect 459744 227666 459796 227672
rect 459374 225312 459430 225321
rect 459374 225247 459430 225256
rect 459560 221332 459612 221338
rect 459560 221274 459612 221280
rect 459572 217410 459600 221274
rect 459756 219570 459784 227666
rect 459940 221066 459968 231676
rect 460492 224670 460520 231676
rect 461044 227730 461072 231676
rect 461228 231662 461610 231690
rect 461032 227724 461084 227730
rect 461032 227666 461084 227672
rect 460480 224664 460532 224670
rect 460480 224606 460532 224612
rect 461032 224120 461084 224126
rect 461032 224062 461084 224068
rect 459928 221060 459980 221066
rect 459928 221002 459980 221008
rect 460204 219836 460256 219842
rect 460204 219778 460256 219784
rect 459744 219564 459796 219570
rect 459744 219506 459796 219512
rect 460216 217410 460244 219778
rect 461044 217410 461072 224062
rect 461228 220862 461256 231662
rect 461584 224528 461636 224534
rect 461584 224470 461636 224476
rect 461596 224126 461624 224470
rect 461584 224120 461636 224126
rect 461584 224062 461636 224068
rect 462148 223990 462176 231676
rect 462700 229094 462728 231676
rect 463252 230178 463280 231676
rect 463818 231662 464200 231690
rect 463240 230172 463292 230178
rect 463240 230114 463292 230120
rect 462700 229066 462820 229094
rect 462136 223984 462188 223990
rect 462136 223926 462188 223932
rect 462792 222873 462820 229066
rect 463884 228404 463936 228410
rect 463884 228346 463936 228352
rect 463896 228290 463924 228346
rect 463344 228274 463924 228290
rect 463332 228268 463924 228274
rect 463384 228262 463924 228268
rect 463332 228210 463384 228216
rect 462964 224800 463016 224806
rect 462964 224742 463016 224748
rect 462778 222864 462834 222873
rect 462778 222799 462834 222808
rect 461860 222012 461912 222018
rect 461860 221954 461912 221960
rect 461216 220856 461268 220862
rect 461216 220798 461268 220804
rect 461872 217410 461900 221954
rect 462976 217410 463004 224742
rect 464172 223038 464200 231662
rect 464356 224942 464384 231676
rect 464908 228818 464936 231676
rect 464896 228812 464948 228818
rect 464896 228754 464948 228760
rect 465264 227316 465316 227322
rect 465264 227258 465316 227264
rect 464988 227180 465040 227186
rect 464988 227122 465040 227128
rect 465000 226914 465028 227122
rect 464988 226908 465040 226914
rect 464988 226850 465040 226856
rect 464344 224936 464396 224942
rect 464344 224878 464396 224884
rect 465080 224800 465132 224806
rect 465080 224742 465132 224748
rect 463884 223032 463936 223038
rect 463884 222974 463936 222980
rect 464160 223032 464212 223038
rect 464160 222974 464212 222980
rect 463700 220108 463752 220114
rect 463700 220050 463752 220056
rect 463712 217410 463740 220050
rect 463896 219842 463924 222974
rect 464344 221740 464396 221746
rect 464344 221682 464396 221688
rect 463884 219836 463936 219842
rect 463884 219778 463936 219784
rect 464356 217410 464384 221682
rect 465092 220114 465120 224742
rect 465080 220108 465132 220114
rect 465080 220050 465132 220056
rect 465276 217410 465304 227258
rect 465460 224534 465488 231676
rect 465816 230444 465868 230450
rect 465816 230386 465868 230392
rect 465828 229094 465856 230386
rect 466012 229226 466040 231676
rect 466564 230450 466592 231676
rect 466552 230444 466604 230450
rect 466552 230386 466604 230392
rect 466000 229220 466052 229226
rect 466000 229162 466052 229168
rect 465828 229066 465948 229094
rect 465724 226908 465776 226914
rect 465724 226850 465776 226856
rect 465736 226642 465764 226850
rect 465920 226642 465948 229066
rect 465724 226636 465776 226642
rect 465724 226578 465776 226584
rect 465908 226636 465960 226642
rect 465908 226578 465960 226584
rect 467116 224806 467144 231676
rect 467576 231662 467682 231690
rect 467576 226137 467604 231662
rect 467748 230444 467800 230450
rect 467748 230386 467800 230392
rect 467562 226128 467618 226137
rect 467562 226063 467618 226072
rect 467104 224800 467156 224806
rect 467104 224742 467156 224748
rect 465448 224528 465500 224534
rect 465448 224470 465500 224476
rect 466460 224120 466512 224126
rect 466460 224062 466512 224068
rect 466472 219706 466500 224062
rect 467760 221202 467788 230386
rect 468220 227594 468248 231676
rect 468392 228676 468444 228682
rect 468392 228618 468444 228624
rect 468208 227588 468260 227594
rect 468208 227530 468260 227536
rect 467932 224392 467984 224398
rect 467932 224334 467984 224340
rect 466828 221196 466880 221202
rect 466828 221138 466880 221144
rect 467748 221196 467800 221202
rect 467748 221138 467800 221144
rect 466000 219700 466052 219706
rect 466000 219642 466052 219648
rect 466460 219700 466512 219706
rect 466460 219642 466512 219648
rect 466012 217410 466040 219642
rect 466840 217410 466868 221138
rect 467944 217410 467972 224334
rect 468404 217410 468432 228618
rect 468772 224126 468800 231676
rect 469324 226302 469352 231676
rect 469890 231662 470364 231690
rect 470336 229094 470364 231662
rect 470244 229066 470364 229094
rect 469312 226296 469364 226302
rect 469312 226238 469364 226244
rect 469312 226024 469364 226030
rect 469312 225966 469364 225972
rect 468760 224120 468812 224126
rect 468760 224062 468812 224068
rect 469324 217410 469352 225966
rect 470244 221338 470272 229066
rect 470428 224398 470456 231676
rect 470994 231662 471468 231690
rect 471546 231662 471928 231690
rect 472098 231662 472480 231690
rect 470416 224392 470468 224398
rect 470416 224334 470468 224340
rect 470232 221332 470284 221338
rect 470232 221274 470284 221280
rect 470140 220652 470192 220658
rect 470140 220594 470192 220600
rect 470152 217410 470180 220594
rect 471440 219842 471468 231662
rect 471900 228682 471928 231662
rect 471888 228676 471940 228682
rect 471888 228618 471940 228624
rect 471980 228268 472032 228274
rect 471980 228210 472032 228216
rect 471796 224936 471848 224942
rect 471796 224878 471848 224884
rect 471808 220522 471836 224878
rect 471796 220516 471848 220522
rect 471796 220458 471848 220464
rect 470968 219836 471020 219842
rect 470968 219778 471020 219784
rect 471428 219836 471480 219842
rect 471428 219778 471480 219784
rect 470980 217410 471008 219778
rect 471992 217410 472020 228210
rect 472256 224936 472308 224942
rect 472256 224878 472308 224884
rect 472268 224534 472296 224878
rect 472256 224528 472308 224534
rect 472256 224470 472308 224476
rect 472452 223718 472480 231662
rect 472636 230586 472664 231676
rect 472624 230580 472676 230586
rect 472624 230522 472676 230528
rect 472808 228540 472860 228546
rect 472808 228482 472860 228488
rect 472624 224392 472676 224398
rect 472624 224334 472676 224340
rect 472636 224126 472664 224334
rect 472624 224120 472676 224126
rect 472624 224062 472676 224068
rect 472440 223712 472492 223718
rect 472440 223654 472492 223660
rect 472820 219434 472848 228482
rect 473188 222018 473216 231676
rect 473740 228546 473768 231676
rect 474306 231662 474688 231690
rect 474660 230722 474688 231662
rect 474648 230716 474700 230722
rect 474648 230658 474700 230664
rect 474844 229226 474872 231676
rect 474648 229220 474700 229226
rect 474648 229162 474700 229168
rect 474832 229220 474884 229226
rect 474832 229162 474884 229168
rect 473728 228540 473780 228546
rect 473728 228482 473780 228488
rect 474660 228274 474688 229162
rect 474924 228404 474976 228410
rect 474924 228346 474976 228352
rect 474648 228268 474700 228274
rect 474648 228210 474700 228216
rect 473544 227044 473596 227050
rect 473544 226986 473596 226992
rect 473176 222012 473228 222018
rect 473176 221954 473228 221960
rect 472544 219406 472848 219434
rect 472544 217410 472572 219406
rect 473556 217410 473584 226986
rect 474188 225888 474240 225894
rect 474188 225830 474240 225836
rect 474200 217410 474228 225830
rect 474464 219836 474516 219842
rect 474464 219778 474516 219784
rect 474476 219609 474504 219778
rect 474462 219600 474518 219609
rect 474462 219535 474518 219544
rect 474936 219434 474964 228346
rect 475396 227322 475424 231676
rect 475384 227316 475436 227322
rect 475384 227258 475436 227264
rect 475108 226024 475160 226030
rect 475108 225966 475160 225972
rect 475120 225622 475148 225966
rect 475108 225616 475160 225622
rect 475108 225558 475160 225564
rect 475384 224528 475436 224534
rect 475384 224470 475436 224476
rect 475568 224528 475620 224534
rect 475568 224470 475620 224476
rect 475396 224126 475424 224470
rect 475384 224120 475436 224126
rect 475384 224062 475436 224068
rect 475580 223718 475608 224470
rect 475568 223712 475620 223718
rect 475568 223654 475620 223660
rect 475948 221746 475976 231676
rect 476500 230450 476528 231676
rect 476488 230444 476540 230450
rect 476488 230386 476540 230392
rect 476212 227452 476264 227458
rect 476212 227394 476264 227400
rect 476224 224954 476252 227394
rect 476224 224926 476344 224954
rect 475936 221740 475988 221746
rect 475936 221682 475988 221688
rect 475384 221604 475436 221610
rect 475384 221546 475436 221552
rect 475396 220522 475424 221546
rect 475200 220516 475252 220522
rect 475200 220458 475252 220464
rect 475384 220516 475436 220522
rect 475384 220458 475436 220464
rect 475212 220266 475240 220458
rect 475212 220238 475792 220266
rect 475764 220114 475792 220238
rect 475568 220108 475620 220114
rect 475568 220050 475620 220056
rect 475752 220108 475804 220114
rect 475752 220050 475804 220056
rect 475580 219706 475608 220050
rect 475568 219700 475620 219706
rect 475568 219642 475620 219648
rect 474936 219406 475056 219434
rect 475028 217410 475056 219406
rect 475936 219428 475988 219434
rect 475936 219370 475988 219376
rect 475752 219292 475804 219298
rect 475752 219234 475804 219240
rect 475764 217530 475792 219234
rect 475948 217666 475976 219370
rect 476316 219178 476344 224926
rect 477052 223718 477080 231676
rect 477408 230444 477460 230450
rect 477408 230386 477460 230392
rect 477224 229220 477276 229226
rect 477224 229162 477276 229168
rect 477236 227458 477264 229162
rect 477224 227452 477276 227458
rect 477224 227394 477276 227400
rect 477040 223712 477092 223718
rect 477040 223654 477092 223660
rect 477420 221882 477448 230386
rect 477604 228410 477632 231676
rect 477880 231662 478170 231690
rect 477592 228404 477644 228410
rect 477592 228346 477644 228352
rect 477408 221876 477460 221882
rect 477408 221818 477460 221824
rect 477880 221610 477908 231662
rect 478052 230716 478104 230722
rect 478052 230658 478104 230664
rect 478064 230450 478092 230658
rect 478052 230444 478104 230450
rect 478052 230386 478104 230392
rect 478328 227180 478380 227186
rect 478328 227122 478380 227128
rect 477868 221604 477920 221610
rect 477868 221546 477920 221552
rect 476578 219600 476634 219609
rect 476578 219535 476580 219544
rect 476632 219535 476634 219544
rect 476580 219506 476632 219512
rect 476764 219428 476816 219434
rect 476764 219370 476816 219376
rect 476074 219156 476126 219162
rect 476316 219150 476620 219178
rect 476074 219098 476126 219104
rect 476086 219042 476114 219098
rect 476086 219014 476436 219042
rect 476408 218754 476436 219014
rect 476396 218748 476448 218754
rect 476396 218690 476448 218696
rect 475936 217660 475988 217666
rect 475936 217602 475988 217608
rect 475752 217524 475804 217530
rect 475752 217466 475804 217472
rect 476592 217410 476620 219150
rect 457732 217382 458068 217410
rect 458468 217382 458896 217410
rect 459572 217382 459724 217410
rect 460216 217382 460552 217410
rect 461044 217382 461380 217410
rect 461872 217382 462208 217410
rect 462976 217382 463036 217410
rect 463712 217382 463864 217410
rect 464356 217382 464692 217410
rect 465276 217382 465520 217410
rect 466012 217382 466348 217410
rect 466840 217382 467176 217410
rect 467944 217382 468004 217410
rect 468404 217382 468832 217410
rect 469324 217382 469660 217410
rect 470152 217382 470488 217410
rect 470980 217382 471316 217410
rect 471992 217382 472144 217410
rect 472544 217382 472972 217410
rect 473556 217382 473800 217410
rect 474200 217382 474628 217410
rect 475028 217382 475456 217410
rect 476284 217382 476620 217410
rect 476776 217410 476804 219370
rect 477914 217660 477966 217666
rect 477914 217602 477966 217608
rect 476776 217382 477112 217410
rect 477926 217396 477954 217602
rect 478340 217410 478368 227122
rect 478708 226166 478736 231676
rect 479260 229226 479288 231676
rect 479248 229220 479300 229226
rect 479248 229162 479300 229168
rect 479812 227186 479840 231676
rect 480076 230444 480128 230450
rect 480076 230386 480128 230392
rect 480088 229094 480116 230386
rect 479996 229066 480116 229094
rect 479800 227180 479852 227186
rect 479800 227122 479852 227128
rect 478696 226160 478748 226166
rect 478696 226102 478748 226108
rect 479996 224369 480024 229066
rect 480364 225622 480392 231676
rect 480916 230382 480944 231676
rect 481100 231662 481482 231690
rect 480904 230376 480956 230382
rect 480904 230318 480956 230324
rect 480536 230308 480588 230314
rect 480536 230250 480588 230256
rect 480548 227050 480576 230250
rect 480536 227044 480588 227050
rect 480536 226986 480588 226992
rect 480352 225616 480404 225622
rect 480352 225558 480404 225564
rect 481100 224641 481128 231662
rect 481272 230716 481324 230722
rect 481272 230658 481324 230664
rect 481086 224632 481142 224641
rect 481086 224567 481142 224576
rect 479982 224360 480038 224369
rect 479982 224295 480038 224304
rect 481086 224360 481142 224369
rect 481086 224295 481142 224304
rect 481100 224126 481128 224295
rect 480904 224120 480956 224126
rect 480904 224062 480956 224068
rect 481088 224120 481140 224126
rect 481088 224062 481140 224068
rect 480916 223718 480944 224062
rect 480904 223712 480956 223718
rect 480904 223654 480956 223660
rect 480352 220652 480404 220658
rect 480352 220594 480404 220600
rect 480364 219609 480392 220594
rect 481088 220516 481140 220522
rect 481088 220458 481140 220464
rect 481100 220402 481128 220458
rect 480548 220374 481128 220402
rect 480548 220114 480576 220374
rect 481284 220114 481312 230658
rect 481824 230036 481876 230042
rect 481824 229978 481876 229984
rect 481836 224954 481864 229978
rect 482020 225894 482048 231676
rect 482572 230178 482600 231676
rect 483138 231662 483520 231690
rect 483690 231662 484072 231690
rect 483296 230376 483348 230382
rect 483294 230344 483296 230353
rect 483348 230344 483350 230353
rect 483294 230279 483350 230288
rect 482560 230172 482612 230178
rect 482560 230114 482612 230120
rect 483296 230036 483348 230042
rect 483296 229978 483348 229984
rect 483308 229537 483336 229978
rect 483294 229528 483350 229537
rect 483294 229463 483350 229472
rect 483492 229094 483520 231662
rect 483756 230308 483808 230314
rect 483756 230250 483808 230256
rect 483400 229066 483520 229094
rect 482008 225888 482060 225894
rect 482008 225830 482060 225836
rect 481836 224926 482508 224954
rect 481454 224632 481510 224641
rect 481454 224567 481510 224576
rect 481468 221241 481496 224567
rect 481454 221232 481510 221241
rect 481454 221167 481510 221176
rect 480536 220108 480588 220114
rect 480536 220050 480588 220056
rect 480720 220108 480772 220114
rect 480720 220050 480772 220056
rect 481272 220108 481324 220114
rect 481272 220050 481324 220056
rect 481456 220108 481508 220114
rect 481456 220050 481508 220056
rect 480350 219600 480406 219609
rect 480350 219535 480406 219544
rect 479892 219428 479944 219434
rect 479892 219370 479944 219376
rect 479904 217410 479932 219370
rect 480732 217410 480760 220050
rect 481468 219570 481496 220050
rect 481456 219564 481508 219570
rect 481456 219506 481508 219512
rect 481732 218748 481784 218754
rect 481732 218690 481784 218696
rect 481226 217524 481278 217530
rect 481226 217466 481278 217472
rect 478340 217382 478768 217410
rect 479596 217382 479932 217410
rect 480424 217382 480760 217410
rect 481238 217396 481266 217466
rect 481744 217410 481772 218690
rect 482480 217410 482508 224926
rect 483400 223145 483428 229066
rect 483572 226024 483624 226030
rect 483572 225966 483624 225972
rect 483386 223136 483442 223145
rect 483386 223071 483442 223080
rect 483584 219298 483612 225966
rect 483572 219292 483624 219298
rect 483572 219234 483624 219240
rect 483768 217410 483796 230250
rect 484044 226030 484072 231662
rect 484228 230042 484256 231676
rect 484780 230625 484808 231676
rect 484766 230616 484822 230625
rect 484766 230551 484822 230560
rect 484216 230036 484268 230042
rect 484216 229978 484268 229984
rect 484860 229900 484912 229906
rect 484860 229842 484912 229848
rect 484676 227044 484728 227050
rect 484676 226986 484728 226992
rect 484032 226024 484084 226030
rect 484032 225966 484084 225972
rect 484688 219162 484716 226986
rect 484676 219156 484728 219162
rect 484676 219098 484728 219104
rect 484872 217410 484900 229842
rect 485332 227050 485360 231676
rect 485884 229906 485912 231676
rect 485872 229900 485924 229906
rect 485872 229842 485924 229848
rect 486436 227769 486464 231676
rect 486422 227760 486478 227769
rect 486422 227695 486478 227704
rect 485320 227044 485372 227050
rect 485320 226986 485372 226992
rect 486988 225622 487016 231676
rect 487540 229770 487568 231676
rect 488092 230314 488120 231676
rect 507504 230722 507532 237895
rect 510724 233918 510752 240615
rect 511092 238754 511120 247959
rect 513300 246362 513328 249766
rect 513288 246356 513340 246362
rect 513288 246298 513340 246304
rect 511814 245576 511870 245585
rect 511870 245534 512040 245562
rect 511814 245511 511870 245520
rect 511262 243128 511318 243137
rect 511262 243063 511318 243072
rect 511276 242350 511304 243063
rect 511264 242344 511316 242350
rect 511264 242286 511316 242292
rect 512012 242214 512040 245534
rect 512000 242208 512052 242214
rect 512000 242150 512052 242156
rect 511092 238726 511304 238754
rect 511276 238066 511304 238726
rect 514036 238202 514064 259966
rect 519544 256760 519596 256766
rect 519544 256702 519596 256708
rect 519556 240786 519584 256702
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 519544 240780 519596 240786
rect 519544 240722 519596 240728
rect 514024 238196 514076 238202
rect 514024 238138 514076 238144
rect 511264 238060 511316 238066
rect 511264 238002 511316 238008
rect 510894 235784 510950 235793
rect 510894 235719 510950 235728
rect 510908 234054 510936 235719
rect 510896 234048 510948 234054
rect 510896 233990 510948 233996
rect 510712 233912 510764 233918
rect 510712 233854 510764 233860
rect 510618 233336 510674 233345
rect 510618 233271 510674 233280
rect 507492 230716 507544 230722
rect 507492 230658 507544 230664
rect 491390 230616 491446 230625
rect 491390 230551 491446 230560
rect 488446 230344 488502 230353
rect 488080 230308 488132 230314
rect 488446 230279 488502 230288
rect 488080 230250 488132 230256
rect 488460 230178 488488 230279
rect 488448 230172 488500 230178
rect 488448 230114 488500 230120
rect 487344 229764 487396 229770
rect 487344 229706 487396 229712
rect 487528 229764 487580 229770
rect 487528 229706 487580 229712
rect 487356 229094 487384 229706
rect 490380 229628 490432 229634
rect 490380 229570 490432 229576
rect 490564 229628 490616 229634
rect 490564 229570 490616 229576
rect 489182 229528 489238 229537
rect 489182 229463 489238 229472
rect 488908 229356 488960 229362
rect 488908 229298 488960 229304
rect 487356 229066 487568 229094
rect 486792 225616 486844 225622
rect 486792 225558 486844 225564
rect 486976 225616 487028 225622
rect 486976 225558 487028 225564
rect 486804 225049 486832 225558
rect 486790 225040 486846 225049
rect 486790 224975 486846 224984
rect 485226 224496 485282 224505
rect 485226 224431 485282 224440
rect 485240 224262 485268 224431
rect 485228 224256 485280 224262
rect 485228 224198 485280 224204
rect 485780 224120 485832 224126
rect 485608 224068 485780 224074
rect 485608 224062 485832 224068
rect 485608 224046 485820 224062
rect 485228 223576 485280 223582
rect 485228 223518 485280 223524
rect 485240 223394 485268 223518
rect 485608 223394 485636 224046
rect 485872 223576 485924 223582
rect 485872 223518 485924 223524
rect 485240 223366 485636 223394
rect 485884 223258 485912 223518
rect 485746 223230 485912 223258
rect 485746 223174 485774 223230
rect 485734 223168 485786 223174
rect 485872 223168 485924 223174
rect 485734 223110 485786 223116
rect 485870 223136 485872 223145
rect 485924 223136 485926 223145
rect 485870 223071 485926 223080
rect 485872 222896 485924 222902
rect 485872 222838 485924 222844
rect 485884 221626 485912 222838
rect 486424 222760 486476 222766
rect 486424 222702 486476 222708
rect 485884 221598 486188 221626
rect 485734 221468 485786 221474
rect 485734 221410 485786 221416
rect 485872 221468 485924 221474
rect 485872 221410 485924 221416
rect 485746 221082 485774 221410
rect 485884 221241 485912 221410
rect 485870 221232 485926 221241
rect 485870 221167 485926 221176
rect 485746 221054 485912 221082
rect 485884 220697 485912 221054
rect 485870 220688 485926 220697
rect 485870 220623 485926 220632
rect 485870 219600 485926 219609
rect 485870 219535 485872 219544
rect 485924 219535 485926 219544
rect 485872 219506 485924 219512
rect 485780 219292 485832 219298
rect 485780 219234 485832 219240
rect 485044 219156 485096 219162
rect 485044 219098 485096 219104
rect 481744 217382 482080 217410
rect 482480 217382 482908 217410
rect 483736 217382 483796 217410
rect 484564 217382 484900 217410
rect 485056 217410 485084 219098
rect 485056 217382 485544 217410
rect 171140 216844 171192 216850
rect 171140 216786 171192 216792
rect 457536 216844 457588 216850
rect 457536 216786 457588 216792
rect 484872 216753 484900 217382
rect 484858 216744 484914 216753
rect 85468 216708 85632 216714
rect 85468 216702 85580 216708
rect 85580 216650 85632 216656
rect 168656 216708 168708 216714
rect 484858 216679 484914 216688
rect 168656 216650 168708 216656
rect 485516 216442 485544 217382
rect 485792 217025 485820 219234
rect 486160 219094 486188 221598
rect 486436 219230 486464 222702
rect 486424 219224 486476 219230
rect 486424 219166 486476 219172
rect 486148 219088 486200 219094
rect 486148 219030 486200 219036
rect 485964 219020 486016 219026
rect 485964 218962 486016 218968
rect 485976 217410 486004 218962
rect 487540 217410 487568 229066
rect 488920 222834 488948 229298
rect 489196 229094 489224 229463
rect 490392 229362 490420 229570
rect 490380 229356 490432 229362
rect 490380 229298 490432 229304
rect 489196 229066 489316 229094
rect 489090 224496 489146 224505
rect 489090 224431 489146 224440
rect 488908 222828 488960 222834
rect 488908 222770 488960 222776
rect 488538 220688 488594 220697
rect 488538 220623 488594 220632
rect 488552 217938 488580 220623
rect 488540 217932 488592 217938
rect 488540 217874 488592 217880
rect 488552 217410 488580 217874
rect 489104 217410 489132 224431
rect 489288 223145 489316 229066
rect 489918 226672 489974 226681
rect 489918 226607 489974 226616
rect 489932 226522 489960 226607
rect 489886 226506 489960 226522
rect 489874 226500 489960 226506
rect 489926 226494 489960 226500
rect 489874 226442 489926 226448
rect 489550 226400 489606 226409
rect 489550 226335 489606 226344
rect 490010 226400 490066 226409
rect 490010 226335 490066 226344
rect 489564 226030 489592 226335
rect 489552 226024 489604 226030
rect 489552 225966 489604 225972
rect 489736 226024 489788 226030
rect 489736 225966 489788 225972
rect 489748 225049 489776 225966
rect 490024 225758 490052 226335
rect 489874 225752 489926 225758
rect 489874 225694 489926 225700
rect 490012 225752 490064 225758
rect 490012 225694 490064 225700
rect 489886 225570 489914 225694
rect 489886 225542 490052 225570
rect 490024 225350 490052 225542
rect 489874 225344 489926 225350
rect 489874 225286 489926 225292
rect 490012 225344 490064 225350
rect 490012 225286 490064 225292
rect 489886 225162 489914 225286
rect 489886 225134 489960 225162
rect 489932 225049 489960 225134
rect 489734 225040 489790 225049
rect 489734 224975 489790 224984
rect 489918 225040 489974 225049
rect 489918 224975 489974 224984
rect 490576 224954 490604 229570
rect 490930 226672 490986 226681
rect 490930 226607 490986 226616
rect 490944 226506 490972 226607
rect 490932 226500 490984 226506
rect 490932 226442 490984 226448
rect 490116 224926 490604 224954
rect 489274 223136 489330 223145
rect 489274 223071 489330 223080
rect 490116 219434 490144 224926
rect 490838 223408 490894 223417
rect 490838 223343 490894 223352
rect 490852 222850 490880 223343
rect 491404 223038 491432 230551
rect 510632 229634 510660 233271
rect 544384 230512 544436 230518
rect 544384 230454 544436 230460
rect 542452 230308 542504 230314
rect 542452 230250 542504 230256
rect 542084 230172 542136 230178
rect 542084 230114 542136 230120
rect 510620 229628 510672 229634
rect 510620 229570 510672 229576
rect 494704 229492 494756 229498
rect 494704 229434 494756 229440
rect 494716 229094 494744 229434
rect 497464 229356 497516 229362
rect 497464 229298 497516 229304
rect 494716 229066 495112 229094
rect 491574 227760 491630 227769
rect 491574 227695 491630 227704
rect 491392 223032 491444 223038
rect 491392 222974 491444 222980
rect 491588 222902 491616 227695
rect 492588 225344 492640 225350
rect 492588 225286 492640 225292
rect 492772 225344 492824 225350
rect 492772 225286 492824 225292
rect 491576 222896 491628 222902
rect 490852 222834 490972 222850
rect 491576 222838 491628 222844
rect 490852 222828 490984 222834
rect 490852 222822 490932 222828
rect 490932 222770 490984 222776
rect 490286 220416 490342 220425
rect 490286 220351 490342 220360
rect 490104 219428 490156 219434
rect 490104 219370 490156 219376
rect 490300 218113 490328 220351
rect 490286 218104 490342 218113
rect 490286 218039 490342 218048
rect 490300 217410 490328 218039
rect 490944 217410 490972 222770
rect 491666 220960 491722 220969
rect 491666 220895 491722 220904
rect 491680 218074 491708 220895
rect 492600 219450 492628 225286
rect 492784 225049 492812 225286
rect 492770 225040 492826 225049
rect 492770 224975 492826 224984
rect 493322 220144 493378 220153
rect 493322 220079 493378 220088
rect 492600 219422 492720 219450
rect 491668 218068 491720 218074
rect 491668 218010 491720 218016
rect 491680 217410 491708 218010
rect 492692 217410 492720 219422
rect 493336 217841 493364 220079
rect 494060 219088 494112 219094
rect 494060 219030 494112 219036
rect 494072 218346 494100 219030
rect 495084 218385 495112 229066
rect 495532 226500 495584 226506
rect 495532 226442 495584 226448
rect 495254 223136 495310 223145
rect 495254 223071 495310 223080
rect 495268 221626 495296 223071
rect 495268 221598 495434 221626
rect 495406 221474 495434 221598
rect 495256 221468 495308 221474
rect 495256 221410 495308 221416
rect 495394 221468 495446 221474
rect 495394 221410 495446 221416
rect 495268 221241 495296 221410
rect 495254 221232 495310 221241
rect 495254 221167 495310 221176
rect 495254 220552 495310 220561
rect 495254 220487 495310 220496
rect 495268 220386 495296 220487
rect 495256 220380 495308 220386
rect 495256 220322 495308 220328
rect 495394 220380 495446 220386
rect 495394 220322 495446 220328
rect 495406 220266 495434 220322
rect 495268 220238 495434 220266
rect 495268 219570 495296 220238
rect 495544 219706 495572 226442
rect 495716 225208 495768 225214
rect 495716 225150 495768 225156
rect 495532 219700 495584 219706
rect 495532 219642 495584 219648
rect 495256 219564 495308 219570
rect 495256 219506 495308 219512
rect 494794 218376 494850 218385
rect 494060 218340 494112 218346
rect 494794 218311 494850 218320
rect 495070 218376 495126 218385
rect 495070 218311 495126 218320
rect 495256 218340 495308 218346
rect 494060 218282 494112 218288
rect 493322 217832 493378 217841
rect 493322 217767 493378 217776
rect 493336 217410 493364 217767
rect 494808 217410 494836 218311
rect 495256 218282 495308 218288
rect 485976 217382 486220 217410
rect 487540 217396 487876 217410
rect 487540 217382 487890 217396
rect 488552 217382 488704 217410
rect 489104 217382 489532 217410
rect 490300 217382 490360 217410
rect 490944 217382 491188 217410
rect 491680 217382 492016 217410
rect 492692 217382 492844 217410
rect 493336 217382 493672 217410
rect 494500 217382 494836 217410
rect 495268 217410 495296 218282
rect 495728 217410 495756 225150
rect 496818 220552 496874 220561
rect 496818 220487 496874 220496
rect 496832 219366 496860 220487
rect 496820 219360 496872 219366
rect 496820 219302 496872 219308
rect 496832 217410 496860 219302
rect 497476 218657 497504 229298
rect 522580 229220 522632 229226
rect 522580 229162 522632 229168
rect 513196 228132 513248 228138
rect 513196 228074 513248 228080
rect 509516 225480 509568 225486
rect 509516 225422 509568 225428
rect 499028 225344 499080 225350
rect 499028 225286 499080 225292
rect 498292 219224 498344 219230
rect 498292 219166 498344 219172
rect 497462 218648 497518 218657
rect 497462 218583 497518 218592
rect 497476 217410 497504 218583
rect 498304 218482 498332 219166
rect 498292 218476 498344 218482
rect 498292 218418 498344 218424
rect 498304 217410 498332 218418
rect 499040 217410 499068 225286
rect 501512 225072 501564 225078
rect 501512 225014 501564 225020
rect 499578 224632 499634 224641
rect 499578 224567 499634 224576
rect 499592 224482 499620 224567
rect 499500 224454 499620 224482
rect 499302 224360 499358 224369
rect 499302 224295 499358 224304
rect 499316 223718 499344 224295
rect 499500 224262 499528 224454
rect 499670 224360 499726 224369
rect 499670 224295 499726 224304
rect 499488 224256 499540 224262
rect 499488 224198 499540 224204
rect 499684 224194 499712 224295
rect 499672 224188 499724 224194
rect 499672 224130 499724 224136
rect 499488 224120 499540 224126
rect 499488 224062 499540 224068
rect 499500 223836 499528 224062
rect 499948 223848 500000 223854
rect 499500 223808 499948 223836
rect 499948 223790 500000 223796
rect 499304 223712 499356 223718
rect 499304 223654 499356 223660
rect 499534 223644 499586 223650
rect 499534 223586 499586 223592
rect 499304 223576 499356 223582
rect 499304 223518 499356 223524
rect 499316 223145 499344 223518
rect 499546 223417 499574 223586
rect 499532 223408 499588 223417
rect 499532 223343 499588 223352
rect 499302 223136 499358 223145
rect 499302 223071 499358 223080
rect 499670 223136 499726 223145
rect 499670 223071 499726 223080
rect 499684 222630 499712 223071
rect 499868 222686 501092 222714
rect 499488 222624 499540 222630
rect 499488 222566 499540 222572
rect 499672 222624 499724 222630
rect 499672 222566 499724 222572
rect 499500 222442 499528 222566
rect 499868 222442 499896 222686
rect 501064 222630 501092 222686
rect 500868 222624 500920 222630
rect 500868 222566 500920 222572
rect 501052 222624 501104 222630
rect 501052 222566 501104 222572
rect 499500 222414 499896 222442
rect 499592 222278 499988 222306
rect 499592 222154 499620 222278
rect 499580 222148 499632 222154
rect 499580 222090 499632 222096
rect 499764 222148 499816 222154
rect 499764 222090 499816 222096
rect 499776 221241 499804 222090
rect 499960 221241 499988 222278
rect 499762 221232 499818 221241
rect 499762 221167 499818 221176
rect 499946 221232 500002 221241
rect 499946 221167 500002 221176
rect 499948 219564 500000 219570
rect 499948 219506 500000 219512
rect 495268 217382 495328 217410
rect 495728 217382 496156 217410
rect 496832 217382 496984 217410
rect 497476 217382 497812 217410
rect 498304 217382 498640 217410
rect 499040 217382 499468 217410
rect 487862 217274 487890 217382
rect 488170 217288 488226 217297
rect 487862 217260 488170 217274
rect 487876 217246 488170 217260
rect 488170 217223 488226 217232
rect 485778 217016 485834 217025
rect 485778 216951 485834 216960
rect 486882 217016 486938 217025
rect 486938 216974 487048 217002
rect 486882 216951 486938 216960
rect 499960 216458 499988 219506
rect 500880 219434 500908 222566
rect 500880 219406 501092 219434
rect 501064 219162 501092 219406
rect 501052 219156 501104 219162
rect 501052 219098 501104 219104
rect 501064 217410 501092 219098
rect 501524 217410 501552 225014
rect 505190 224632 505246 224641
rect 505190 224567 505246 224576
rect 505204 224262 505232 224567
rect 505192 224256 505244 224262
rect 505192 224198 505244 224204
rect 504916 224188 504968 224194
rect 504916 224130 504968 224136
rect 504732 223712 504784 223718
rect 504732 223654 504784 223660
rect 504744 223417 504772 223654
rect 504928 223530 504956 224130
rect 504928 223514 505416 223530
rect 504928 223508 505428 223514
rect 504928 223502 505376 223508
rect 505376 223450 505428 223456
rect 505192 223440 505244 223446
rect 504730 223408 504786 223417
rect 505192 223382 505244 223388
rect 504730 223343 504786 223352
rect 505204 222630 505232 223382
rect 503444 222624 503496 222630
rect 503444 222566 503496 222572
rect 505192 222624 505244 222630
rect 505192 222566 505244 222572
rect 503456 222358 503484 222566
rect 505008 222488 505060 222494
rect 505192 222488 505244 222494
rect 505060 222448 505192 222476
rect 505008 222430 505060 222436
rect 505192 222430 505244 222436
rect 503168 222352 503220 222358
rect 503168 222294 503220 222300
rect 503444 222352 503496 222358
rect 503444 222294 503496 222300
rect 508504 222352 508556 222358
rect 508504 222294 508556 222300
rect 502340 220652 502392 220658
rect 502340 220594 502392 220600
rect 502352 220017 502380 220594
rect 502338 220008 502394 220017
rect 502338 219943 502394 219952
rect 502352 217410 502380 219943
rect 503180 219026 503208 222294
rect 504730 221232 504786 221241
rect 504730 221167 504786 221176
rect 504364 220652 504416 220658
rect 504364 220594 504416 220600
rect 504376 220386 504404 220594
rect 504364 220380 504416 220386
rect 504364 220322 504416 220328
rect 504548 220380 504600 220386
rect 504548 220322 504600 220328
rect 504560 219706 504588 220322
rect 504744 219706 504772 221167
rect 506032 220782 506612 220810
rect 506032 220658 506060 220782
rect 506020 220652 506072 220658
rect 506020 220594 506072 220600
rect 506204 220652 506256 220658
rect 506204 220594 506256 220600
rect 505098 219872 505154 219881
rect 505098 219807 505100 219816
rect 505152 219807 505154 219816
rect 505100 219778 505152 219784
rect 504548 219700 504600 219706
rect 504548 219642 504600 219648
rect 504732 219700 504784 219706
rect 504732 219642 504784 219648
rect 503168 219020 503220 219026
rect 503168 218962 503220 218968
rect 503628 219020 503680 219026
rect 503628 218962 503680 218968
rect 503640 217410 503668 218962
rect 504364 218748 504416 218754
rect 504364 218690 504416 218696
rect 504178 217832 504234 217841
rect 504178 217767 504234 217776
rect 501064 217382 501124 217410
rect 501524 217382 501952 217410
rect 502352 217382 502780 217410
rect 503608 217382 503668 217410
rect 504192 217297 504220 217767
rect 504376 217410 504404 218690
rect 505112 217410 505140 219778
rect 506216 219638 506244 220594
rect 506584 219842 506612 220782
rect 507768 219972 507820 219978
rect 507768 219914 507820 219920
rect 506572 219836 506624 219842
rect 506572 219778 506624 219784
rect 506204 219632 506256 219638
rect 506204 219574 506256 219580
rect 506216 217410 506244 219574
rect 507780 219473 507808 219914
rect 507766 219464 507822 219473
rect 507766 219399 507822 219408
rect 506572 218884 506624 218890
rect 506572 218826 506624 218832
rect 504376 217382 504436 217410
rect 505112 217382 505264 217410
rect 506092 217382 506244 217410
rect 506584 217410 506612 218826
rect 507780 217410 507808 219399
rect 508516 218618 508544 222294
rect 508504 218612 508556 218618
rect 508504 218554 508556 218560
rect 506584 217382 506920 217410
rect 507748 217382 507808 217410
rect 508516 217410 508544 218554
rect 509528 217410 509556 225422
rect 509884 224120 509936 224126
rect 509884 224062 509936 224068
rect 509896 223854 509924 224062
rect 509884 223848 509936 223854
rect 509884 223790 509936 223796
rect 510068 223848 510120 223854
rect 510068 223790 510120 223796
rect 510080 223417 510108 223790
rect 510066 223408 510122 223417
rect 510066 223343 510122 223352
rect 510712 222488 510764 222494
rect 510712 222430 510764 222436
rect 509976 219836 510028 219842
rect 509976 219778 510028 219784
rect 508516 217382 508576 217410
rect 509404 217382 509556 217410
rect 509988 217410 510016 219778
rect 510724 218210 510752 222430
rect 511540 220380 511592 220386
rect 511540 220322 511592 220328
rect 510712 218204 510764 218210
rect 510712 218146 510764 218152
rect 510724 217410 510752 218146
rect 511552 217410 511580 220322
rect 511998 220280 512054 220289
rect 511998 220215 512000 220224
rect 512052 220215 512054 220224
rect 512642 220280 512698 220289
rect 512642 220215 512698 220224
rect 512000 220186 512052 220192
rect 512656 217410 512684 220215
rect 509988 217382 510384 217410
rect 510724 217382 511060 217410
rect 511552 217382 511888 217410
rect 512656 217382 512716 217410
rect 504178 217288 504234 217297
rect 504178 217223 504234 217232
rect 510356 217122 510384 217382
rect 510344 217116 510396 217122
rect 510344 217058 510396 217064
rect 513208 216458 513236 228074
rect 514760 227996 514812 228002
rect 514760 227938 514812 227944
rect 513380 226772 513432 226778
rect 513380 226714 513432 226720
rect 513392 220386 513420 226714
rect 514576 223848 514628 223854
rect 514576 223790 514628 223796
rect 514588 223417 514616 223790
rect 514574 223408 514630 223417
rect 514574 223343 514630 223352
rect 514024 222624 514076 222630
rect 514024 222566 514076 222572
rect 513380 220380 513432 220386
rect 513380 220322 513432 220328
rect 514036 217410 514064 222566
rect 514772 217666 514800 227938
rect 518072 227860 518124 227866
rect 518072 227802 518124 227808
rect 516784 223848 516836 223854
rect 516784 223790 516836 223796
rect 516796 223514 516824 223790
rect 516784 223508 516836 223514
rect 516784 223450 516836 223456
rect 517426 223408 517482 223417
rect 517426 223343 517482 223352
rect 515588 220380 515640 220386
rect 515588 220322 515640 220328
rect 515600 219298 515628 220322
rect 517440 219450 517468 223343
rect 517440 219422 517652 219450
rect 515588 219292 515640 219298
rect 515588 219234 515640 219240
rect 514760 217660 514812 217666
rect 514760 217602 514812 217608
rect 515600 217410 515628 219234
rect 516002 217660 516054 217666
rect 516002 217602 516054 217608
rect 514036 217382 514372 217410
rect 515200 217382 515628 217410
rect 516014 217410 516042 217602
rect 517624 217410 517652 219422
rect 518084 217410 518112 227802
rect 519176 226908 519228 226914
rect 519176 226850 519228 226856
rect 518992 223304 519044 223310
rect 518992 223246 519044 223252
rect 519004 217410 519032 223246
rect 519188 217666 519216 226850
rect 520556 226636 520608 226642
rect 520556 226578 520608 226584
rect 519544 223304 519596 223310
rect 519544 223246 519596 223252
rect 519556 222766 519584 223246
rect 519544 222760 519596 222766
rect 519544 222702 519596 222708
rect 519728 222284 519780 222290
rect 519728 222226 519780 222232
rect 519544 222148 519596 222154
rect 519544 222090 519596 222096
rect 519556 221474 519584 222090
rect 519740 221474 519768 222226
rect 519544 221468 519596 221474
rect 519544 221410 519596 221416
rect 519728 221468 519780 221474
rect 519728 221410 519780 221416
rect 519176 217660 519228 217666
rect 519176 217602 519228 217608
rect 520142 217660 520194 217666
rect 520142 217602 520194 217608
rect 516014 217396 516364 217410
rect 516028 217382 516364 217396
rect 517624 217382 517684 217410
rect 518084 217382 518848 217410
rect 519004 217382 519340 217410
rect 516140 216708 516192 216714
rect 516140 216650 516192 216656
rect 513838 216472 513894 216481
rect 499960 216442 500632 216458
rect 485504 216436 485556 216442
rect 499960 216436 500644 216442
rect 499960 216430 500592 216436
rect 485504 216378 485556 216384
rect 513208 216430 513838 216458
rect 516152 216442 516180 216650
rect 516336 216442 516364 217382
rect 516520 216986 516856 217002
rect 516508 216980 516856 216986
rect 516560 216974 516856 216980
rect 516508 216922 516560 216928
rect 518624 216708 518676 216714
rect 518624 216650 518676 216656
rect 518636 216442 518664 216650
rect 518820 216442 518848 217382
rect 520154 216730 520182 217602
rect 520568 217410 520596 226578
rect 522592 223446 522620 229162
rect 524052 229084 524104 229090
rect 524052 229026 524104 229032
rect 523132 228948 523184 228954
rect 523132 228890 523184 228896
rect 522580 223440 522632 223446
rect 522580 223382 522632 223388
rect 523144 222426 523172 228890
rect 523132 222420 523184 222426
rect 523132 222362 523184 222368
rect 523684 222420 523736 222426
rect 523684 222362 523736 222368
rect 521658 222048 521714 222057
rect 521658 221983 521714 221992
rect 521672 219774 521700 221983
rect 521660 219768 521712 219774
rect 521660 219710 521712 219716
rect 522580 219768 522632 219774
rect 522580 219710 522632 219716
rect 522592 217410 522620 219710
rect 523696 217410 523724 222362
rect 520568 217382 521240 217410
rect 522592 217382 522652 217410
rect 523480 217382 523724 217410
rect 524064 217410 524092 229026
rect 532700 228812 532752 228818
rect 532700 228754 532752 228760
rect 527824 227724 527876 227730
rect 527824 227666 527876 227672
rect 525062 225312 525118 225321
rect 525062 225247 525118 225256
rect 524236 224664 524288 224670
rect 524234 224632 524236 224641
rect 524374 224664 524426 224670
rect 524288 224632 524290 224641
rect 524374 224606 524426 224612
rect 524234 224567 524290 224576
rect 524386 224482 524414 224606
rect 524248 224454 524414 224482
rect 524248 223854 524276 224454
rect 524236 223848 524288 223854
rect 524236 223790 524288 223796
rect 524374 223848 524426 223854
rect 524374 223790 524426 223796
rect 524386 223666 524414 223790
rect 524248 223638 524414 223666
rect 524248 223417 524276 223638
rect 524234 223408 524290 223417
rect 524234 223343 524290 223352
rect 525076 220017 525104 225247
rect 526350 224632 526406 224641
rect 526350 224567 526406 224576
rect 526168 221060 526220 221066
rect 526168 221002 526220 221008
rect 525062 220008 525118 220017
rect 525062 219943 525118 219952
rect 525076 217410 525104 219943
rect 526180 217410 526208 221002
rect 524064 217382 524308 217410
rect 525076 217382 525136 217410
rect 525964 217382 526208 217410
rect 526364 217410 526392 224567
rect 527836 219638 527864 227666
rect 528836 223984 528888 223990
rect 528836 223926 528888 223932
rect 528376 220856 528428 220862
rect 528376 220798 528428 220804
rect 527824 219632 527876 219638
rect 527824 219574 527876 219580
rect 527836 217410 527864 219574
rect 526364 217382 526792 217410
rect 527620 217382 527864 217410
rect 528388 217410 528416 220798
rect 528560 220652 528612 220658
rect 528560 220594 528612 220600
rect 528572 218754 528600 220594
rect 528560 218748 528612 218754
rect 528560 218690 528612 218696
rect 528848 217410 528876 223926
rect 531320 223304 531372 223310
rect 531320 223246 531372 223252
rect 530398 222864 530454 222873
rect 530398 222799 530454 222808
rect 530412 219910 530440 222799
rect 530768 222148 530820 222154
rect 530768 222090 530820 222096
rect 530400 219904 530452 219910
rect 530400 219846 530452 219852
rect 530412 217410 530440 219846
rect 528388 217382 528448 217410
rect 528848 217382 529276 217410
rect 530104 217382 530440 217410
rect 520154 216716 520320 216730
rect 520168 216714 520320 216716
rect 520168 216708 520332 216714
rect 520168 216702 520280 216708
rect 520280 216650 520332 216656
rect 520646 216472 520702 216481
rect 513838 216407 513894 216416
rect 516140 216436 516192 216442
rect 500592 216378 500644 216384
rect 516140 216378 516192 216384
rect 516324 216436 516376 216442
rect 516324 216378 516376 216384
rect 518624 216436 518676 216442
rect 518624 216378 518676 216384
rect 518808 216436 518860 216442
rect 521212 216442 521240 217382
rect 526444 217116 526496 217122
rect 526444 217058 526496 217064
rect 521672 216850 521824 216866
rect 521660 216844 521824 216850
rect 521712 216838 521824 216844
rect 525432 216844 525484 216850
rect 521660 216786 521712 216792
rect 525432 216786 525484 216792
rect 525444 216578 525472 216786
rect 525432 216572 525484 216578
rect 525432 216514 525484 216520
rect 526074 216472 526130 216481
rect 520646 216407 520648 216416
rect 518808 216378 518860 216384
rect 520700 216407 520702 216416
rect 521200 216436 521252 216442
rect 520648 216378 520700 216384
rect 526456 216442 526484 217058
rect 530780 217002 530808 222090
rect 531332 217410 531360 223246
rect 532516 220380 532568 220386
rect 532516 220322 532568 220328
rect 532528 217410 532556 220322
rect 531332 217382 531760 217410
rect 532528 217382 532588 217410
rect 531240 217246 531452 217274
rect 531240 217122 531268 217246
rect 531228 217116 531280 217122
rect 531228 217058 531280 217064
rect 530780 216986 531268 217002
rect 530780 216980 531280 216986
rect 530780 216974 531228 216980
rect 531228 216922 531280 216928
rect 531424 216578 531452 217246
rect 531872 216844 531924 216850
rect 531872 216786 531924 216792
rect 531412 216572 531464 216578
rect 531412 216514 531464 216520
rect 531226 216472 531282 216481
rect 526074 216407 526076 216416
rect 521200 216378 521252 216384
rect 526128 216407 526130 216416
rect 526444 216436 526496 216442
rect 526076 216378 526128 216384
rect 531884 216442 531912 216786
rect 532712 216578 532740 228754
rect 540336 228540 540388 228546
rect 540336 228482 540388 228488
rect 540348 228274 540376 228482
rect 534724 228268 534776 228274
rect 534724 228210 534776 228216
rect 540336 228268 540388 228274
rect 540336 228210 540388 228216
rect 534172 224936 534224 224942
rect 534172 224878 534224 224884
rect 533344 224664 533396 224670
rect 533344 224606 533396 224612
rect 533356 224398 533384 224606
rect 533160 224392 533212 224398
rect 533160 224334 533212 224340
rect 533344 224392 533396 224398
rect 533344 224334 533396 224340
rect 533172 223990 533200 224334
rect 533160 223984 533212 223990
rect 533160 223926 533212 223932
rect 533526 220008 533582 220017
rect 533080 219966 533526 219994
rect 533080 219745 533108 219966
rect 533526 219943 533582 219952
rect 533066 219736 533122 219745
rect 533066 219671 533122 219680
rect 534184 217410 534212 224878
rect 534736 220522 534764 228210
rect 538220 227588 538272 227594
rect 538220 227530 538272 227536
rect 537482 226128 537538 226137
rect 537482 226063 537538 226072
rect 536380 224800 536432 224806
rect 536380 224742 536432 224748
rect 535552 221196 535604 221202
rect 535552 221138 535604 221144
rect 534724 220516 534776 220522
rect 534724 220458 534776 220464
rect 534736 217410 534764 220458
rect 535368 219496 535420 219502
rect 535368 219438 535420 219444
rect 535380 218929 535408 219438
rect 535366 218920 535422 218929
rect 535366 218855 535422 218864
rect 535564 217410 535592 221138
rect 536392 217410 536420 224742
rect 537496 219502 537524 226063
rect 537484 219496 537536 219502
rect 537484 219438 537536 219444
rect 537496 217410 537524 219438
rect 537668 217660 537720 217666
rect 537668 217602 537720 217608
rect 534184 217382 534244 217410
rect 534736 217382 535072 217410
rect 535564 217382 536236 217410
rect 536392 217382 536728 217410
rect 537496 217382 537556 217410
rect 536208 217122 536236 217382
rect 536196 217116 536248 217122
rect 536196 217058 536248 217064
rect 533416 216578 533752 216594
rect 532700 216572 532752 216578
rect 533416 216572 533764 216578
rect 533416 216566 533712 216572
rect 532700 216514 532752 216520
rect 533712 216514 533764 216520
rect 537390 216472 537446 216481
rect 531226 216407 531228 216416
rect 526444 216378 526496 216384
rect 531280 216407 531282 216416
rect 531872 216436 531924 216442
rect 531228 216378 531280 216384
rect 537680 216442 537708 217602
rect 538232 217274 538260 227530
rect 540336 226296 540388 226302
rect 540336 226238 540388 226244
rect 538864 223984 538916 223990
rect 538864 223926 538916 223932
rect 538680 217524 538732 217530
rect 538680 217466 538732 217472
rect 538232 217258 538384 217274
rect 538220 217252 538384 217258
rect 538272 217246 538384 217252
rect 538220 217194 538272 217200
rect 538036 216844 538088 216850
rect 538036 216786 538088 216792
rect 538048 216442 538076 216786
rect 538692 216442 538720 217466
rect 538876 217410 538904 223926
rect 540348 220250 540376 226238
rect 542096 224398 542124 230114
rect 542464 228682 542492 230250
rect 542452 228676 542504 228682
rect 542452 228618 542504 228624
rect 542820 228540 542872 228546
rect 542820 228482 542872 228488
rect 542832 224954 542860 228482
rect 544396 224954 544424 230454
rect 549904 230036 549956 230042
rect 549904 229978 549956 229984
rect 546500 228268 546552 228274
rect 546500 228210 546552 228216
rect 542832 224926 542952 224954
rect 544396 224926 544608 224954
rect 541348 224392 541400 224398
rect 541348 224334 541400 224340
rect 542084 224392 542136 224398
rect 542084 224334 542136 224340
rect 540520 221332 540572 221338
rect 540520 221274 540572 221280
rect 540336 220244 540388 220250
rect 540336 220186 540388 220192
rect 539600 218884 539652 218890
rect 539600 218826 539652 218832
rect 538876 217382 539212 217410
rect 539612 216578 539640 218826
rect 540348 217410 540376 220186
rect 540040 217382 540376 217410
rect 540532 217410 540560 221274
rect 541162 217560 541218 217569
rect 541162 217495 541218 217504
rect 540532 217396 540868 217410
rect 540532 217382 540882 217396
rect 540854 216866 540882 217382
rect 540854 216852 541020 216866
rect 540868 216850 541020 216852
rect 539784 216844 539836 216850
rect 540868 216844 541032 216850
rect 540868 216838 540980 216844
rect 539784 216786 539836 216792
rect 540980 216786 541032 216792
rect 539796 216578 539824 216786
rect 539600 216572 539652 216578
rect 539600 216514 539652 216520
rect 539784 216572 539836 216578
rect 539784 216514 539836 216520
rect 541176 216442 541204 217495
rect 541360 217410 541388 224334
rect 542544 220516 542596 220522
rect 542544 220458 542596 220464
rect 542360 220108 542412 220114
rect 542360 220050 542412 220056
rect 541716 217796 541768 217802
rect 541716 217738 541768 217744
rect 541728 217530 541756 217738
rect 542082 217662 542138 217671
rect 541912 217620 542082 217648
rect 541716 217524 541768 217530
rect 541716 217466 541768 217472
rect 541360 217382 541696 217410
rect 541912 216560 541940 217620
rect 542082 217597 542138 217606
rect 542176 217524 542228 217530
rect 542176 217466 542228 217472
rect 542188 216578 542216 217466
rect 542372 217410 542400 220050
rect 542556 220046 542584 220458
rect 542544 220040 542596 220046
rect 542544 219982 542596 219988
rect 542542 219192 542598 219201
rect 542542 219127 542598 219136
rect 542556 217682 542584 219127
rect 542728 217796 542780 217802
rect 542728 217738 542780 217744
rect 542556 217654 542676 217682
rect 542496 217560 542552 217569
rect 542496 217495 542552 217504
rect 542510 217410 542538 217495
rect 542372 217396 542538 217410
rect 542372 217382 542524 217396
rect 542648 216730 542676 217654
rect 542740 217274 542768 217738
rect 542924 217410 542952 224926
rect 543924 224528 543976 224534
rect 543924 224470 543976 224476
rect 543462 219192 543518 219201
rect 543462 219127 543518 219136
rect 543096 217796 543148 217802
rect 543096 217738 543148 217744
rect 543108 217530 543136 217738
rect 543096 217524 543148 217530
rect 543096 217466 543148 217472
rect 543326 217524 543378 217530
rect 543326 217466 543378 217472
rect 543338 217410 543366 217466
rect 542924 217396 543366 217410
rect 542924 217382 543352 217396
rect 542740 217246 543044 217274
rect 542648 216702 542768 216730
rect 542176 216572 542228 216578
rect 541912 216532 542032 216560
rect 542004 216442 542032 216532
rect 542176 216514 542228 216520
rect 542740 216510 542768 216702
rect 542728 216504 542780 216510
rect 542728 216446 542780 216452
rect 543016 216442 543044 217246
rect 543476 216442 543504 219127
rect 543646 217560 543702 217569
rect 543646 217495 543702 217504
rect 543660 216442 543688 217495
rect 543936 217410 543964 224470
rect 544580 220522 544608 224926
rect 545764 222012 545816 222018
rect 545764 221954 545816 221960
rect 545776 220833 545804 221954
rect 545762 220824 545818 220833
rect 545762 220759 545818 220768
rect 544568 220516 544620 220522
rect 544568 220458 544620 220464
rect 544382 219192 544438 219201
rect 544382 219127 544438 219136
rect 544396 217802 544424 219127
rect 544384 217796 544436 217802
rect 544384 217738 544436 217744
rect 544580 217410 544608 220458
rect 545580 217660 545632 217666
rect 545580 217602 545632 217608
rect 543936 217382 544180 217410
rect 544580 217382 545008 217410
rect 545592 217394 545620 217602
rect 545776 217410 545804 220759
rect 546132 218884 546184 218890
rect 546132 218826 546184 218832
rect 546316 218884 546368 218890
rect 546316 218826 546368 218832
rect 546144 217569 546172 218826
rect 546328 217802 546356 218826
rect 546316 217796 546368 217802
rect 546316 217738 546368 217744
rect 546130 217560 546186 217569
rect 546130 217495 546186 217504
rect 546512 217410 546540 228210
rect 547972 227452 548024 227458
rect 547972 227394 548024 227400
rect 547420 224256 547472 224262
rect 547420 224198 547472 224204
rect 547432 222358 547460 224198
rect 547420 222352 547472 222358
rect 547420 222294 547472 222300
rect 547432 217410 547460 222294
rect 547984 219434 548012 227394
rect 548708 227316 548760 227322
rect 548708 227258 548760 227264
rect 548340 220652 548392 220658
rect 548340 220594 548392 220600
rect 548154 220552 548210 220561
rect 548154 220487 548156 220496
rect 548208 220487 548210 220496
rect 548156 220458 548208 220464
rect 548352 219502 548380 220594
rect 548524 220516 548576 220522
rect 548524 220458 548576 220464
rect 548536 220046 548564 220458
rect 548524 220040 548576 220046
rect 548524 219982 548576 219988
rect 548340 219496 548392 219502
rect 548340 219438 548392 219444
rect 547984 219406 548196 219434
rect 547970 217560 548026 217569
rect 547970 217495 548026 217504
rect 545580 217388 545632 217394
rect 545776 217382 545836 217410
rect 546512 217382 546664 217410
rect 547432 217382 547492 217410
rect 545580 217330 545632 217336
rect 547984 216578 548012 217495
rect 548168 217410 548196 219406
rect 548524 218884 548576 218890
rect 548524 218826 548576 218832
rect 548536 217802 548564 218826
rect 548524 217796 548576 217802
rect 548524 217738 548576 217744
rect 548720 217410 548748 227258
rect 549916 222018 549944 229978
rect 558184 229900 558236 229906
rect 558184 229842 558236 229848
rect 552296 228404 552348 228410
rect 552296 228346 552348 228352
rect 551284 224120 551336 224126
rect 551284 224062 551336 224068
rect 549904 222012 549956 222018
rect 549904 221954 549956 221960
rect 550640 221876 550692 221882
rect 550640 221818 550692 221824
rect 549996 221740 550048 221746
rect 549996 221682 550048 221688
rect 549350 220824 549406 220833
rect 549350 220759 549406 220768
rect 548890 220552 548946 220561
rect 548890 220487 548946 220496
rect 548904 220046 548932 220487
rect 548892 220040 548944 220046
rect 548892 219982 548944 219988
rect 549364 219434 549392 220759
rect 550008 219502 550036 221682
rect 549996 219496 550048 219502
rect 549996 219438 550048 219444
rect 549364 219406 549484 219434
rect 548168 217394 548564 217410
rect 548168 217388 548576 217394
rect 548168 217382 548524 217388
rect 548720 217382 549148 217410
rect 548524 217330 548576 217336
rect 547972 216572 548024 216578
rect 547972 216514 548024 216520
rect 549456 216481 549484 219406
rect 550008 217410 550036 219438
rect 550652 217841 550680 221818
rect 551296 218054 551324 224062
rect 552308 218890 552336 228346
rect 554780 227180 554832 227186
rect 554780 227122 554832 227128
rect 553676 226160 553728 226166
rect 553676 226102 553728 226108
rect 553308 221332 553360 221338
rect 553308 221274 553360 221280
rect 552662 219192 552718 219201
rect 552662 219127 552718 219136
rect 552296 218884 552348 218890
rect 552296 218826 552348 218832
rect 550928 218026 551324 218054
rect 550638 217832 550694 217841
rect 550638 217767 550694 217776
rect 549976 217382 550036 217410
rect 550652 217410 550680 217767
rect 550652 217382 550804 217410
rect 545670 216472 545726 216481
rect 537390 216407 537392 216416
rect 531872 216378 531924 216384
rect 537444 216407 537446 216416
rect 537668 216436 537720 216442
rect 537392 216378 537444 216384
rect 537668 216378 537720 216384
rect 538036 216436 538088 216442
rect 538036 216378 538088 216384
rect 538680 216436 538732 216442
rect 538680 216378 538732 216384
rect 541164 216436 541216 216442
rect 541164 216378 541216 216384
rect 541992 216436 542044 216442
rect 541992 216378 542044 216384
rect 543004 216436 543056 216442
rect 543004 216378 543056 216384
rect 543464 216436 543516 216442
rect 543464 216378 543516 216384
rect 543648 216436 543700 216442
rect 543648 216378 543700 216384
rect 545120 216436 545172 216442
rect 545488 216436 545540 216442
rect 545172 216396 545488 216424
rect 545120 216378 545172 216384
rect 545670 216407 545672 216416
rect 545488 216378 545540 216384
rect 545724 216407 545726 216416
rect 546774 216472 546830 216481
rect 546774 216407 546776 216416
rect 545672 216378 545724 216384
rect 546828 216407 546830 216416
rect 549442 216472 549498 216481
rect 550928 216458 550956 218026
rect 552308 217410 552336 218826
rect 552308 217382 552460 217410
rect 550928 216430 551632 216458
rect 552676 216442 552704 219127
rect 553320 217410 553348 221274
rect 553490 219192 553546 219201
rect 553490 219127 553546 219136
rect 553504 217802 553532 219127
rect 553492 217796 553544 217802
rect 553492 217738 553544 217744
rect 553288 217382 553348 217410
rect 553688 217410 553716 226102
rect 554792 222630 554820 227122
rect 556160 226024 556212 226030
rect 556160 225966 556212 225972
rect 554964 223440 555016 223446
rect 554964 223382 555016 223388
rect 554780 222624 554832 222630
rect 554780 222566 554832 222572
rect 554976 220561 555004 223382
rect 555424 222624 555476 222630
rect 555424 222566 555476 222572
rect 555436 222494 555464 222566
rect 555424 222488 555476 222494
rect 555424 222430 555476 222436
rect 554962 220552 555018 220561
rect 554962 220487 555018 220496
rect 554976 217410 555004 220487
rect 553688 217382 554116 217410
rect 554944 217382 555004 217410
rect 555436 217410 555464 222430
rect 556172 217410 556200 225966
rect 557356 224392 557408 224398
rect 557356 224334 557408 224340
rect 557368 222630 557396 224334
rect 557356 222624 557408 222630
rect 557356 222566 557408 222572
rect 556986 219192 557042 219201
rect 556986 219127 557042 219136
rect 556802 217832 556858 217841
rect 556802 217767 556804 217776
rect 556856 217767 556858 217776
rect 556804 217738 556856 217744
rect 555436 217382 555772 217410
rect 556172 217382 556600 217410
rect 557000 216481 557028 219127
rect 557368 217410 557396 222566
rect 558196 221882 558224 229842
rect 559472 228676 559524 228682
rect 559472 228618 559524 228624
rect 558920 225888 558972 225894
rect 558920 225830 558972 225836
rect 558184 221876 558236 221882
rect 558184 221818 558236 221824
rect 558368 221332 558420 221338
rect 558368 221274 558420 221280
rect 558380 221218 558408 221274
rect 558012 221202 558408 221218
rect 558000 221196 558408 221202
rect 558052 221190 558408 221196
rect 558000 221138 558052 221144
rect 558380 217410 558408 221190
rect 557368 217382 557428 217410
rect 558256 217382 558408 217410
rect 558932 217410 558960 225830
rect 559484 217410 559512 228618
rect 561220 225752 561272 225758
rect 561220 225694 561272 225700
rect 560392 223168 560444 223174
rect 560392 223110 560444 223116
rect 560114 217832 560170 217841
rect 560114 217767 560170 217776
rect 560128 217410 560156 217767
rect 558932 217382 559084 217410
rect 559484 217382 560156 217410
rect 560404 217410 560432 223110
rect 560576 222012 560628 222018
rect 560576 221954 560628 221960
rect 560588 220833 560616 221954
rect 560574 220824 560630 220833
rect 560574 220759 560630 220768
rect 561034 217832 561090 217841
rect 561034 217767 561090 217776
rect 561048 217410 561076 217767
rect 560404 217382 561076 217410
rect 561232 217410 561260 225694
rect 562336 224262 562364 252554
rect 567200 240780 567252 240786
rect 567200 240722 567252 240728
rect 565084 229764 565136 229770
rect 565084 229706 565136 229712
rect 563888 227044 563940 227050
rect 563888 226986 563940 226992
rect 562324 224256 562376 224262
rect 562324 224198 562376 224204
rect 563612 223032 563664 223038
rect 563612 222974 563664 222980
rect 563624 222194 563652 222974
rect 563624 222166 563744 222194
rect 562322 221096 562378 221105
rect 562322 221031 562378 221040
rect 562138 220824 562194 220833
rect 562138 220759 562194 220768
rect 562152 217410 562180 220759
rect 562336 219910 562364 221031
rect 562508 220652 562560 220658
rect 562508 220594 562560 220600
rect 562966 220654 563022 220663
rect 562520 219910 562548 220594
rect 562966 220589 563022 220598
rect 562324 219904 562376 219910
rect 562324 219846 562376 219852
rect 562508 219904 562560 219910
rect 562508 219846 562560 219852
rect 562876 219904 562928 219910
rect 562876 219846 562928 219852
rect 563060 219904 563112 219910
rect 563060 219846 563112 219852
rect 562888 219450 562916 219846
rect 563072 219638 563100 219846
rect 563060 219632 563112 219638
rect 563060 219574 563112 219580
rect 562888 219422 563284 219450
rect 563256 219298 563284 219422
rect 563060 219292 563112 219298
rect 563060 219234 563112 219240
rect 563244 219292 563296 219298
rect 563244 219234 563296 219240
rect 562506 219192 562562 219201
rect 563072 219178 563100 219234
rect 563426 219192 563482 219201
rect 563072 219150 563426 219178
rect 562506 219127 562562 219136
rect 563426 219127 563482 219136
rect 561232 217382 561568 217410
rect 562152 217382 562396 217410
rect 562520 216578 562548 219127
rect 563026 218198 563468 218226
rect 563026 218074 563054 218198
rect 563014 218068 563066 218074
rect 563014 218010 563066 218016
rect 563152 218068 563204 218074
rect 563152 218010 563204 218016
rect 563164 217841 563192 218010
rect 563440 217841 563468 218198
rect 563716 217841 563744 222166
rect 563900 218054 563928 226986
rect 564716 221876 564768 221882
rect 564716 221818 564768 221824
rect 564728 221610 564756 221818
rect 565096 221746 565124 229706
rect 567212 229094 567240 240722
rect 567212 229066 568160 229094
rect 566096 225616 566148 225622
rect 566096 225558 566148 225564
rect 565728 222896 565780 222902
rect 565728 222838 565780 222844
rect 565740 222630 565768 222838
rect 565728 222624 565780 222630
rect 565728 222566 565780 222572
rect 565740 222194 565768 222566
rect 565648 222166 565768 222194
rect 565084 221740 565136 221746
rect 565084 221682 565136 221688
rect 564716 221604 564768 221610
rect 564716 221546 564768 221552
rect 564070 221096 564126 221105
rect 564070 221031 564126 221040
rect 564084 219366 564112 221031
rect 564072 219360 564124 219366
rect 564072 219302 564124 219308
rect 563808 218026 563928 218054
rect 563808 217954 563836 218026
rect 563808 217926 563928 217954
rect 563150 217832 563206 217841
rect 563150 217767 563206 217776
rect 563426 217832 563482 217841
rect 563426 217767 563482 217776
rect 563702 217832 563758 217841
rect 563702 217767 563758 217776
rect 563716 217410 563744 217767
rect 563224 217382 563744 217410
rect 563900 217410 563928 217926
rect 564728 217410 564756 221546
rect 565648 217410 565676 222166
rect 566108 217410 566136 225558
rect 568132 224954 568160 229066
rect 568132 224926 568436 224954
rect 567384 221740 567436 221746
rect 567384 221682 567436 221688
rect 567396 217410 567424 221682
rect 567936 219904 567988 219910
rect 567936 219846 567988 219852
rect 568408 219858 568436 224926
rect 568592 221474 568620 261462
rect 571340 249076 571392 249082
rect 571340 249018 571392 249024
rect 569960 246356 570012 246362
rect 569960 246298 570012 246304
rect 568764 238196 568816 238202
rect 568764 238138 568816 238144
rect 568580 221468 568632 221474
rect 568580 221410 568632 221416
rect 567948 219756 567976 219846
rect 568408 219830 568528 219858
rect 568304 219768 568356 219774
rect 567948 219728 568304 219756
rect 568304 219710 568356 219716
rect 568500 217410 568528 219830
rect 563900 217382 564052 217410
rect 564728 217382 564880 217410
rect 565648 217382 565708 217410
rect 566108 217382 566536 217410
rect 567364 217382 567424 217410
rect 568192 217382 568528 217410
rect 568776 217410 568804 238138
rect 569972 229094 570000 246298
rect 571352 229094 571380 249018
rect 628564 242344 628616 242350
rect 628564 242286 628616 242292
rect 577504 234048 577556 234054
rect 577504 233990 577556 233996
rect 569972 229066 570644 229094
rect 571352 229066 572024 229094
rect 569500 221468 569552 221474
rect 569500 221410 569552 221416
rect 569512 217410 569540 221410
rect 570420 217660 570472 217666
rect 570420 217602 570472 217608
rect 568776 217382 569020 217410
rect 569512 217382 569848 217410
rect 570432 217122 570460 217602
rect 570616 217410 570644 229066
rect 571340 224256 571392 224262
rect 571340 224198 571392 224204
rect 571352 217410 571380 224198
rect 571996 222194 572024 229066
rect 571628 222166 572024 222194
rect 571628 218192 571656 222166
rect 572272 220918 572668 220946
rect 572272 220425 572300 220918
rect 572640 220833 572668 220918
rect 572442 220824 572498 220833
rect 572442 220759 572498 220768
rect 572626 220824 572682 220833
rect 572626 220759 572682 220768
rect 575110 220824 575166 220833
rect 575110 220759 575166 220768
rect 572456 220674 572484 220759
rect 572456 220646 572714 220674
rect 572534 220552 572590 220561
rect 572686 220522 572714 220646
rect 572534 220487 572536 220496
rect 572588 220487 572590 220496
rect 572674 220516 572726 220522
rect 572536 220458 572588 220464
rect 572674 220458 572726 220464
rect 572258 220416 572314 220425
rect 572258 220351 572314 220360
rect 572442 220280 572498 220289
rect 572442 220215 572498 220224
rect 572456 219745 572484 220215
rect 574928 219904 574980 219910
rect 574928 219846 574980 219852
rect 572442 219736 572498 219745
rect 572442 219671 572498 219680
rect 572168 219496 572220 219502
rect 572168 219438 572220 219444
rect 572180 219201 572208 219438
rect 572996 219292 573048 219298
rect 572996 219234 573048 219240
rect 572166 219192 572222 219201
rect 572166 219127 572222 219136
rect 571812 218470 572484 218498
rect 571812 218346 571840 218470
rect 572456 218346 572484 218470
rect 571800 218340 571852 218346
rect 571800 218282 571852 218288
rect 572444 218340 572496 218346
rect 572444 218282 572496 218288
rect 571628 218164 571748 218192
rect 571720 218054 571748 218164
rect 573008 218054 573036 219234
rect 573730 219192 573786 219201
rect 573730 219127 573786 219136
rect 571720 218026 571932 218054
rect 571904 217410 571932 218026
rect 572640 218026 573036 218054
rect 573364 218068 573416 218074
rect 572640 217841 572668 218026
rect 573364 218010 573416 218016
rect 572626 217832 572682 217841
rect 572626 217767 572682 217776
rect 573376 217666 573404 218010
rect 573364 217660 573416 217666
rect 573364 217602 573416 217608
rect 570616 217382 570676 217410
rect 571352 217382 571504 217410
rect 571904 217382 572332 217410
rect 567844 217116 567896 217122
rect 567844 217058 567896 217064
rect 570420 217116 570472 217122
rect 570420 217058 570472 217064
rect 566188 216708 566240 216714
rect 566188 216650 566240 216656
rect 562508 216572 562560 216578
rect 562508 216514 562560 216520
rect 553950 216472 554006 216481
rect 552664 216436 552716 216442
rect 549442 216407 549498 216416
rect 546776 216378 546828 216384
rect 553950 216407 553952 216416
rect 552664 216378 552716 216384
rect 554004 216407 554006 216416
rect 556986 216472 557042 216481
rect 566200 216442 566228 216650
rect 567856 216442 567884 217058
rect 573744 216986 573772 219127
rect 574650 218376 574706 218385
rect 574650 218311 574706 218320
rect 574468 218068 574520 218074
rect 574664 218054 574692 218311
rect 574940 218054 574968 219846
rect 574664 218026 574876 218054
rect 574940 218026 575060 218054
rect 574468 218010 574520 218016
rect 574480 217841 574508 218010
rect 574466 217832 574522 217841
rect 574466 217767 574522 217776
rect 574466 217560 574522 217569
rect 574466 217495 574522 217504
rect 573548 216980 573600 216986
rect 573548 216922 573600 216928
rect 573732 216980 573784 216986
rect 573732 216922 573784 216928
rect 573560 216866 573588 216922
rect 573560 216838 574324 216866
rect 556986 216407 557042 216416
rect 566188 216436 566240 216442
rect 553952 216378 554004 216384
rect 566188 216378 566240 216384
rect 567844 216436 567896 216442
rect 567844 216378 567896 216384
rect 573732 216436 573784 216442
rect 573732 216378 573784 216384
rect 573744 216050 573772 216378
rect 574008 216368 574060 216374
rect 574008 216310 574060 216316
rect 574020 216209 574048 216310
rect 574006 216200 574062 216209
rect 574006 216135 574062 216144
rect 573744 216022 574140 216050
rect 573916 215620 573968 215626
rect 573916 215562 573968 215568
rect 573732 215348 573784 215354
rect 573732 215290 573784 215296
rect 573744 214606 573772 215290
rect 573928 214742 573956 215562
rect 573916 214736 573968 214742
rect 573916 214678 573968 214684
rect 573732 214600 573784 214606
rect 573732 214542 573784 214548
rect 574112 213518 574140 216022
rect 574296 215778 574324 216838
rect 574480 216209 574508 217495
rect 574466 216200 574522 216209
rect 574466 216135 574522 216144
rect 574558 215928 574614 215937
rect 574558 215863 574614 215872
rect 574296 215750 574508 215778
rect 574480 213654 574508 215750
rect 574572 214418 574600 215863
rect 574848 215642 574876 218026
rect 574756 215614 574876 215642
rect 574756 214742 574784 215614
rect 575032 214826 575060 218026
rect 574940 214798 575060 214826
rect 574940 214742 574968 214798
rect 574744 214736 574796 214742
rect 574744 214678 574796 214684
rect 574928 214736 574980 214742
rect 574928 214678 574980 214684
rect 574836 214464 574888 214470
rect 574572 214390 574692 214418
rect 574836 214406 574888 214412
rect 574664 213790 574692 214390
rect 574652 213784 574704 213790
rect 574652 213726 574704 213732
rect 574468 213648 574520 213654
rect 574468 213590 574520 213596
rect 574100 213512 574152 213518
rect 574100 213454 574152 213460
rect 574848 213246 574876 214406
rect 575124 214334 575152 220759
rect 575846 220552 575902 220561
rect 575846 220487 575902 220496
rect 575296 219904 575348 219910
rect 575296 219846 575348 219852
rect 575308 219502 575336 219846
rect 575860 219774 575888 220487
rect 576030 220280 576086 220289
rect 576030 220215 576086 220224
rect 575664 219768 575716 219774
rect 575664 219710 575716 219716
rect 575848 219768 575900 219774
rect 575848 219710 575900 219716
rect 575296 219496 575348 219502
rect 575296 219438 575348 219444
rect 575296 216980 575348 216986
rect 575296 216922 575348 216928
rect 575308 214470 575336 216922
rect 575478 216200 575534 216209
rect 575478 216135 575534 216144
rect 575296 214464 575348 214470
rect 575296 214406 575348 214412
rect 575112 214328 575164 214334
rect 575112 214270 575164 214276
rect 575492 213382 575520 216135
rect 575676 214878 575704 219710
rect 576044 219434 576072 220215
rect 575860 219406 576072 219434
rect 575664 214872 575716 214878
rect 575664 214814 575716 214820
rect 575860 214606 575888 219406
rect 576766 216472 576822 216481
rect 576766 216407 576822 216416
rect 576780 216102 576808 216407
rect 576584 216096 576636 216102
rect 576584 216038 576636 216044
rect 576768 216096 576820 216102
rect 576768 216038 576820 216044
rect 576596 215914 576624 216038
rect 576596 215886 576854 215914
rect 576582 215792 576638 215801
rect 576826 215762 576854 215886
rect 576582 215727 576638 215736
rect 576814 215756 576866 215762
rect 576030 215384 576086 215393
rect 576596 215354 576624 215727
rect 576814 215698 576866 215704
rect 576030 215319 576086 215328
rect 576584 215348 576636 215354
rect 576044 215014 576072 215319
rect 576584 215290 576636 215296
rect 576032 215008 576084 215014
rect 576032 214950 576084 214956
rect 575848 214600 575900 214606
rect 575848 214542 575900 214548
rect 575480 213376 575532 213382
rect 575480 213318 575532 213324
rect 574836 213240 574888 213246
rect 574836 213182 574888 213188
rect 51724 211200 51776 211206
rect 51724 211142 51776 211148
rect 50344 204604 50396 204610
rect 50344 204546 50396 204552
rect 48964 204332 49016 204338
rect 48964 204274 49016 204280
rect 47582 203280 47638 203289
rect 47582 203215 47638 203224
rect 44548 191820 44600 191826
rect 44548 191762 44600 191768
rect 44364 191684 44416 191690
rect 44364 191626 44416 191632
rect 42432 183524 42484 183530
rect 42432 183466 42484 183472
rect 44180 183524 44232 183530
rect 44180 183466 44232 183472
rect 41786 183424 41842 183433
rect 41786 183359 41842 183368
rect 41800 183124 41828 183359
rect 42444 182491 42472 183466
rect 42182 182463 42472 182491
rect 577516 97986 577544 233990
rect 617708 223848 617760 223854
rect 617708 223790 617760 223796
rect 611360 222624 611412 222630
rect 611360 222566 611412 222572
rect 608600 222488 608652 222494
rect 608600 222430 608652 222436
rect 601700 222216 601752 222222
rect 601700 222158 601752 222164
rect 596732 221740 596784 221746
rect 596732 221682 596784 221688
rect 596744 220862 596772 221682
rect 597100 221332 597152 221338
rect 597100 221274 597152 221280
rect 597112 221066 597140 221274
rect 597100 221060 597152 221066
rect 597100 221002 597152 221008
rect 596732 220856 596784 220862
rect 596732 220798 596784 220804
rect 591304 220720 591356 220726
rect 590948 220668 591304 220674
rect 590948 220662 591356 220668
rect 590948 220646 591344 220662
rect 596272 220652 596324 220658
rect 590948 220522 590976 220646
rect 596272 220594 596324 220600
rect 590936 220516 590988 220522
rect 590936 220458 590988 220464
rect 596284 219162 596312 220594
rect 601516 220040 601568 220046
rect 601516 219982 601568 219988
rect 597560 219768 597612 219774
rect 597560 219710 597612 219716
rect 596088 219156 596140 219162
rect 596088 219098 596140 219104
rect 596272 219156 596324 219162
rect 596272 219098 596324 219104
rect 587900 219020 587952 219026
rect 587900 218962 587952 218968
rect 591304 219020 591356 219026
rect 591304 218962 591356 218968
rect 587532 218476 587584 218482
rect 587532 218418 587584 218424
rect 580356 218340 580408 218346
rect 580356 218282 580408 218288
rect 581644 218340 581696 218346
rect 581644 218282 581696 218288
rect 578698 216064 578754 216073
rect 578698 215999 578754 216008
rect 578514 212800 578570 212809
rect 578514 212735 578570 212744
rect 578528 211342 578556 212735
rect 578516 211336 578568 211342
rect 578516 211278 578568 211284
rect 578712 208350 578740 215999
rect 579250 214296 579306 214305
rect 579250 214231 579306 214240
rect 579264 212022 579292 214231
rect 580368 213926 580396 218282
rect 581656 218074 581684 218282
rect 587544 218074 587572 218418
rect 587912 218346 587940 218962
rect 591316 218482 591344 218962
rect 596100 218906 596128 219098
rect 596100 218878 596220 218906
rect 591304 218476 591356 218482
rect 591304 218418 591356 218424
rect 587900 218340 587952 218346
rect 587900 218282 587952 218288
rect 596192 218074 596220 218878
rect 597572 218754 597600 219710
rect 597376 218748 597428 218754
rect 597376 218690 597428 218696
rect 597560 218748 597612 218754
rect 597560 218690 597612 218696
rect 597388 218482 597416 218690
rect 598480 218612 598532 218618
rect 598480 218554 598532 218560
rect 597376 218476 597428 218482
rect 597376 218418 597428 218424
rect 597928 218476 597980 218482
rect 597928 218418 597980 218424
rect 597560 218340 597612 218346
rect 597560 218282 597612 218288
rect 581644 218068 581696 218074
rect 581644 218010 581696 218016
rect 587532 218068 587584 218074
rect 587532 218010 587584 218016
rect 595352 218068 595404 218074
rect 595352 218010 595404 218016
rect 596180 218068 596232 218074
rect 596180 218010 596232 218016
rect 596824 218068 596876 218074
rect 596824 218010 596876 218016
rect 594800 217932 594852 217938
rect 594800 217874 594852 217880
rect 586702 215520 586758 215529
rect 586474 215484 586526 215490
rect 586702 215455 586704 215464
rect 586474 215426 586526 215432
rect 586756 215455 586758 215464
rect 586704 215426 586756 215432
rect 586486 215370 586514 215426
rect 586486 215342 586652 215370
rect 586624 215257 586652 215342
rect 586610 215248 586666 215257
rect 586610 215183 586666 215192
rect 594062 215248 594118 215257
rect 594062 215183 594118 215192
rect 581644 215144 581696 215150
rect 581644 215086 581696 215092
rect 581460 215008 581512 215014
rect 581460 214950 581512 214956
rect 581472 214742 581500 214950
rect 581460 214736 581512 214742
rect 581460 214678 581512 214684
rect 581656 214334 581684 215086
rect 581644 214328 581696 214334
rect 581644 214270 581696 214276
rect 580356 213920 580408 213926
rect 580356 213862 580408 213868
rect 579252 212016 579304 212022
rect 579252 211958 579304 211964
rect 581920 212016 581972 212022
rect 581920 211958 581972 211964
rect 578884 211200 578936 211206
rect 578882 211168 578884 211177
rect 580908 211200 580960 211206
rect 578936 211168 578938 211177
rect 580908 211142 580960 211148
rect 578882 211103 578938 211112
rect 579252 209840 579304 209846
rect 579250 209808 579252 209817
rect 579304 209808 579306 209817
rect 579250 209743 579306 209752
rect 578700 208344 578752 208350
rect 578422 208312 578478 208321
rect 578700 208286 578752 208292
rect 578422 208247 578478 208256
rect 578436 208078 578464 208247
rect 578424 208072 578476 208078
rect 578424 208014 578476 208020
rect 580632 208072 580684 208078
rect 580632 208014 580684 208020
rect 578698 206816 578754 206825
rect 578698 206751 578754 206760
rect 578712 205698 578740 206751
rect 578700 205692 578752 205698
rect 578700 205634 578752 205640
rect 579066 205320 579122 205329
rect 579066 205255 579068 205264
rect 579120 205255 579122 205264
rect 579068 205226 579120 205232
rect 578698 203824 578754 203833
rect 578698 203759 578754 203768
rect 578712 202910 578740 203759
rect 578700 202904 578752 202910
rect 578700 202846 578752 202852
rect 578238 202328 578294 202337
rect 578238 202263 578294 202272
rect 578252 201686 578280 202263
rect 578240 201680 578292 201686
rect 578240 201622 578292 201628
rect 578514 200832 578570 200841
rect 578514 200767 578570 200776
rect 578528 200462 578556 200767
rect 578516 200456 578568 200462
rect 578516 200398 578568 200404
rect 580644 200054 580672 208014
rect 580920 204202 580948 211142
rect 581644 209840 581696 209846
rect 581644 209782 581696 209788
rect 580908 204196 580960 204202
rect 580908 204138 580960 204144
rect 581656 202774 581684 209782
rect 581932 206990 581960 211958
rect 583300 211336 583352 211342
rect 583300 211278 583352 211284
rect 581920 206984 581972 206990
rect 581920 206926 581972 206932
rect 581828 205692 581880 205698
rect 581828 205634 581880 205640
rect 581644 202768 581696 202774
rect 581644 202710 581696 202716
rect 580908 201680 580960 201686
rect 580908 201622 580960 201628
rect 580632 200048 580684 200054
rect 580632 199990 580684 199996
rect 578882 199336 578938 199345
rect 578882 199271 578938 199280
rect 578896 198762 578924 199271
rect 578884 198756 578936 198762
rect 578884 198698 578936 198704
rect 578330 197840 578386 197849
rect 578330 197775 578386 197784
rect 578344 197470 578372 197775
rect 578332 197464 578384 197470
rect 578332 197406 578384 197412
rect 580264 197464 580316 197470
rect 580264 197406 580316 197412
rect 579250 196344 579306 196353
rect 579250 196279 579306 196288
rect 579264 196178 579292 196279
rect 579252 196172 579304 196178
rect 579252 196114 579304 196120
rect 578882 194848 578938 194857
rect 578882 194783 578938 194792
rect 578514 193488 578570 193497
rect 578514 193423 578516 193432
rect 578568 193423 578570 193432
rect 578516 193394 578568 193400
rect 578238 190360 578294 190369
rect 578238 190295 578294 190304
rect 578252 189106 578280 190295
rect 578240 189100 578292 189106
rect 578240 189042 578292 189048
rect 578514 187368 578570 187377
rect 578514 187303 578570 187312
rect 578528 187202 578556 187303
rect 578516 187196 578568 187202
rect 578516 187138 578568 187144
rect 578896 186250 578924 194783
rect 579528 191888 579580 191894
rect 579526 191856 579528 191865
rect 579580 191856 579582 191865
rect 579526 191791 579582 191800
rect 579250 188864 579306 188873
rect 579250 188799 579252 188808
rect 579304 188799 579306 188808
rect 579252 188770 579304 188776
rect 580276 187610 580304 197406
rect 580920 194546 580948 201622
rect 581840 200802 581868 205634
rect 583312 205630 583340 211278
rect 594076 210202 594104 215183
rect 594812 210202 594840 217874
rect 595364 213790 595392 218010
rect 596270 215928 596326 215937
rect 596270 215863 596326 215872
rect 595810 215792 595866 215801
rect 595866 215750 596128 215778
rect 596284 215762 596312 215863
rect 595810 215727 595866 215736
rect 596100 215744 596128 215750
rect 596272 215756 596324 215762
rect 596100 215716 596174 215744
rect 595994 215656 596050 215665
rect 595994 215591 596050 215600
rect 596008 215490 596036 215591
rect 596146 215506 596174 215716
rect 596272 215698 596324 215704
rect 596456 215756 596508 215762
rect 596456 215698 596508 215704
rect 596468 215506 596496 215698
rect 596638 215656 596694 215665
rect 596638 215591 596640 215600
rect 596692 215591 596694 215600
rect 596640 215562 596692 215568
rect 595996 215484 596048 215490
rect 596146 215478 596496 215506
rect 595996 215426 596048 215432
rect 595720 213920 595772 213926
rect 595720 213862 595772 213868
rect 596364 213920 596416 213926
rect 596364 213862 596416 213868
rect 595168 213784 595220 213790
rect 595168 213726 595220 213732
rect 595352 213784 595404 213790
rect 595352 213726 595404 213732
rect 595180 210202 595208 213726
rect 595732 210202 595760 213862
rect 596376 210202 596404 213862
rect 596836 210202 596864 218010
rect 597572 210202 597600 218282
rect 597940 210202 597968 218418
rect 598492 210202 598520 218554
rect 599032 218204 599084 218210
rect 599032 218146 599084 218152
rect 599044 210202 599072 218146
rect 600780 216504 600832 216510
rect 600780 216446 600832 216452
rect 600964 216504 601016 216510
rect 600964 216446 601016 216452
rect 600792 216102 600820 216446
rect 600976 216238 601004 216446
rect 600964 216232 601016 216238
rect 600964 216174 601016 216180
rect 600780 216096 600832 216102
rect 600780 216038 600832 216044
rect 601528 215966 601556 219982
rect 601240 215960 601292 215966
rect 600502 215928 600558 215937
rect 599584 215892 599636 215898
rect 601240 215902 601292 215908
rect 601516 215960 601568 215966
rect 601516 215902 601568 215908
rect 600502 215863 600558 215872
rect 599584 215834 599636 215840
rect 599596 210202 599624 215834
rect 600516 215490 600544 215863
rect 600688 215756 600740 215762
rect 600688 215698 600740 215704
rect 600320 215484 600372 215490
rect 600320 215426 600372 215432
rect 600504 215484 600556 215490
rect 600504 215426 600556 215432
rect 600332 210202 600360 215426
rect 600700 210202 600728 215698
rect 601252 210202 601280 215902
rect 601712 210202 601740 222158
rect 603448 221740 603500 221746
rect 603448 221682 603500 221688
rect 602252 220924 602304 220930
rect 602252 220866 602304 220872
rect 602068 217252 602120 217258
rect 602068 217194 602120 217200
rect 602080 213790 602108 217194
rect 602068 213784 602120 213790
rect 602068 213726 602120 213732
rect 602264 210202 602292 220866
rect 602896 220516 602948 220522
rect 602896 220458 602948 220464
rect 602908 216102 602936 220458
rect 603080 216844 603132 216850
rect 603080 216786 603132 216792
rect 602896 216096 602948 216102
rect 602896 216038 602948 216044
rect 603092 213926 603120 216786
rect 603080 213920 603132 213926
rect 603080 213862 603132 213868
rect 603460 210202 603488 221682
rect 607220 220380 607272 220386
rect 607220 220322 607272 220328
rect 605288 217524 605340 217530
rect 605288 217466 605340 217472
rect 604000 215484 604052 215490
rect 604000 215426 604052 215432
rect 603632 213648 603684 213654
rect 603632 213590 603684 213596
rect 594076 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599596 210174 599932 210202
rect 600332 210174 600484 210202
rect 600700 210174 601036 210202
rect 601252 210174 601588 210202
rect 601712 210174 602140 210202
rect 602264 210174 602692 210202
rect 603244 210174 603488 210202
rect 603644 210202 603672 213590
rect 604012 210202 604040 215426
rect 605300 213790 605328 217466
rect 607232 217326 607260 220322
rect 607864 217796 607916 217802
rect 607864 217738 607916 217744
rect 607404 217456 607456 217462
rect 607404 217398 607456 217404
rect 607220 217320 607272 217326
rect 607220 217262 607272 217268
rect 606760 216504 606812 216510
rect 606760 216446 606812 216452
rect 605932 213920 605984 213926
rect 605932 213862 605984 213868
rect 605104 213784 605156 213790
rect 605104 213726 605156 213732
rect 605288 213784 605340 213790
rect 605288 213726 605340 213732
rect 604552 213512 604604 213518
rect 604552 213454 604604 213460
rect 604564 210202 604592 213454
rect 605116 210202 605144 213726
rect 605944 210202 605972 213862
rect 606208 213784 606260 213790
rect 606208 213726 606260 213732
rect 606220 210202 606248 213726
rect 606772 210202 606800 216446
rect 607416 210202 607444 217398
rect 607876 210202 607904 217738
rect 603644 210174 603796 210202
rect 604012 210174 604348 210202
rect 604564 210174 604900 210202
rect 605116 210174 605452 210202
rect 605944 210174 606004 210202
rect 606220 210174 606556 210202
rect 606772 210174 607108 210202
rect 607416 210174 607660 210202
rect 607876 210174 608212 210202
rect 608612 210118 608640 222430
rect 608968 221196 609020 221202
rect 608968 221138 609020 221144
rect 608784 221060 608836 221066
rect 608784 221002 608836 221008
rect 608796 214470 608824 221002
rect 608784 214464 608836 214470
rect 608784 214406 608836 214412
rect 608980 210202 609008 221138
rect 610348 219904 610400 219910
rect 610348 219846 610400 219852
rect 609244 219292 609296 219298
rect 609244 219234 609296 219240
rect 609256 213926 609284 219234
rect 609888 217660 609940 217666
rect 609888 217602 609940 217608
rect 609520 214464 609572 214470
rect 609520 214406 609572 214412
rect 609244 213920 609296 213926
rect 609244 213862 609296 213868
rect 608764 210174 609008 210202
rect 609532 210202 609560 214406
rect 609900 212650 609928 217602
rect 610360 217462 610388 219846
rect 610348 217456 610400 217462
rect 610348 217398 610400 217404
rect 610624 213920 610676 213926
rect 610624 213862 610676 213868
rect 609900 212622 610112 212650
rect 610084 210202 610112 212622
rect 610636 210202 610664 213862
rect 611372 210202 611400 222566
rect 614026 220008 614082 220017
rect 614026 219943 614082 219952
rect 613382 218920 613438 218929
rect 613382 218855 613438 218864
rect 612278 218104 612334 218113
rect 612278 218039 612334 218048
rect 611726 217016 611782 217025
rect 611726 216951 611782 216960
rect 611740 210202 611768 216951
rect 612292 210202 612320 218039
rect 612830 217288 612886 217297
rect 612830 217223 612886 217232
rect 612844 210202 612872 217223
rect 613396 210202 613424 218855
rect 614040 216850 614068 219943
rect 614946 219736 615002 219745
rect 614946 219671 615002 219680
rect 614028 216844 614080 216850
rect 614028 216786 614080 216792
rect 614488 216844 614540 216850
rect 614488 216786 614540 216792
rect 614120 215620 614172 215626
rect 614120 215562 614172 215568
rect 614132 210202 614160 215562
rect 614500 210202 614528 216786
rect 614960 210202 614988 219671
rect 615498 219464 615554 219473
rect 615498 219399 615554 219408
rect 615512 210202 615540 219399
rect 617248 219020 617300 219026
rect 617248 218962 617300 218968
rect 616144 217116 616196 217122
rect 616144 217058 616196 217064
rect 616156 210202 616184 217058
rect 616696 216232 616748 216238
rect 616696 216174 616748 216180
rect 616708 213042 616736 216174
rect 616880 215144 616932 215150
rect 616880 215086 616932 215092
rect 616696 213036 616748 213042
rect 616696 212978 616748 212984
rect 616892 210202 616920 215086
rect 617260 210202 617288 218962
rect 617720 210202 617748 223790
rect 626540 222624 626592 222630
rect 626540 222566 626592 222572
rect 623964 222352 624016 222358
rect 623964 222294 624016 222300
rect 620284 221468 620336 221474
rect 620284 221410 620336 221416
rect 620296 221202 620324 221410
rect 620284 221196 620336 221202
rect 620284 221138 620336 221144
rect 622676 220244 622728 220250
rect 622676 220186 622728 220192
rect 621664 218748 621716 218754
rect 621664 218690 621716 218696
rect 620560 217456 620612 217462
rect 620560 217398 620612 217404
rect 618352 216708 618404 216714
rect 618352 216650 618404 216656
rect 618364 210202 618392 216650
rect 618904 215008 618956 215014
rect 618904 214950 618956 214956
rect 618916 210202 618944 214950
rect 620008 214872 620060 214878
rect 620008 214814 620060 214820
rect 619640 214736 619692 214742
rect 619640 214678 619692 214684
rect 619652 210202 619680 214678
rect 620020 210202 620048 214814
rect 620572 210202 620600 217398
rect 621112 217320 621164 217326
rect 621112 217262 621164 217268
rect 621124 210202 621152 217262
rect 621676 210202 621704 218690
rect 622400 214600 622452 214606
rect 622400 214542 622452 214548
rect 622412 210202 622440 214542
rect 622688 210202 622716 220186
rect 623780 215960 623832 215966
rect 623780 215902 623832 215908
rect 623320 213036 623372 213042
rect 623320 212978 623372 212984
rect 623332 210202 623360 212978
rect 623792 210202 623820 215902
rect 623976 210338 624004 222294
rect 624148 219496 624200 219502
rect 624148 219438 624200 219444
rect 624160 213926 624188 219438
rect 625528 218884 625580 218890
rect 625528 218826 625580 218832
rect 624148 213920 624200 213926
rect 624148 213862 624200 213868
rect 625252 213920 625304 213926
rect 625252 213862 625304 213868
rect 623976 210310 624372 210338
rect 624344 210202 624372 210310
rect 625264 210202 625292 213862
rect 625540 210202 625568 218826
rect 626080 216096 626132 216102
rect 626080 216038 626132 216044
rect 626092 210202 626120 216038
rect 626552 210202 626580 222566
rect 628196 221332 628248 221338
rect 628196 221274 628248 221280
rect 628012 221196 628064 221202
rect 628012 221138 628064 221144
rect 628024 219162 628052 221138
rect 627828 219156 627880 219162
rect 627828 219098 627880 219104
rect 628012 219156 628064 219162
rect 628012 219098 628064 219104
rect 627840 219042 627868 219098
rect 627840 219014 627960 219042
rect 627184 216368 627236 216374
rect 627184 216310 627236 216316
rect 627196 210202 627224 216310
rect 627932 210202 627960 219014
rect 628208 210202 628236 221274
rect 628576 213926 628604 242286
rect 633440 242208 633492 242214
rect 633440 242150 633492 242156
rect 632704 238060 632756 238066
rect 632704 238002 632756 238008
rect 629944 233912 629996 233918
rect 629944 233854 629996 233860
rect 629956 229094 629984 233854
rect 629956 229066 630076 229094
rect 629852 223644 629904 223650
rect 629852 223586 629904 223592
rect 628840 219156 628892 219162
rect 628840 219098 628892 219104
rect 628564 213920 628616 213926
rect 628564 213862 628616 213868
rect 628852 210202 628880 219098
rect 629392 213376 629444 213382
rect 629392 213318 629444 213324
rect 629404 210202 629432 213318
rect 629864 210202 629892 223586
rect 630048 212702 630076 229066
rect 631046 218648 631102 218657
rect 631046 218583 631102 218592
rect 630680 213240 630732 213246
rect 630680 213182 630732 213188
rect 630036 212696 630088 212702
rect 630036 212638 630088 212644
rect 630692 210202 630720 213182
rect 631060 210202 631088 218583
rect 631598 216744 631654 216753
rect 631598 216679 631654 216688
rect 631612 210202 631640 216679
rect 632716 212838 632744 238002
rect 632704 212832 632756 212838
rect 632704 212774 632756 212780
rect 632704 212696 632756 212702
rect 632704 212638 632756 212644
rect 632716 210202 632744 212638
rect 633452 210202 633480 242150
rect 641812 230988 641864 230994
rect 641812 230930 641864 230936
rect 633808 213920 633860 213926
rect 633808 213862 633860 213868
rect 639972 213920 640024 213926
rect 639972 213862 640024 213868
rect 633820 210202 633848 213862
rect 638868 213784 638920 213790
rect 638868 213726 638920 213732
rect 638316 213648 638368 213654
rect 638316 213590 638368 213596
rect 636660 213512 636712 213518
rect 636660 213454 636712 213460
rect 635556 213376 635608 213382
rect 635556 213318 635608 213324
rect 634360 212832 634412 212838
rect 634360 212774 634412 212780
rect 634372 210202 634400 212774
rect 635568 210202 635596 213318
rect 636672 210202 636700 213454
rect 637212 213240 637264 213246
rect 637212 213182 637264 213188
rect 637224 210202 637252 213182
rect 638328 210202 638356 213590
rect 638880 210202 638908 213726
rect 639984 210202 640012 213862
rect 640248 213104 640300 213110
rect 640248 213046 640300 213052
rect 640260 210202 640288 213046
rect 641628 212968 641680 212974
rect 641628 212910 641680 212916
rect 641640 210202 641668 212910
rect 609532 210174 609868 210202
rect 610084 210174 610420 210202
rect 610636 210174 610972 210202
rect 611372 210174 611524 210202
rect 611740 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 614960 210174 615388 210202
rect 615512 210174 615940 210202
rect 616156 210174 616492 210202
rect 616892 210174 617044 210202
rect 617260 210174 617596 210202
rect 617720 210174 618148 210202
rect 618364 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620020 210174 620356 210202
rect 620572 210174 620908 210202
rect 621124 210174 621460 210202
rect 621676 210174 622012 210202
rect 622412 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623792 210174 624220 210202
rect 624344 210174 624772 210202
rect 625264 210174 625324 210202
rect 625540 210174 625876 210202
rect 626092 210174 626428 210202
rect 626552 210174 626980 210202
rect 627196 210174 627532 210202
rect 627932 210174 628084 210202
rect 628208 210174 628636 210202
rect 628852 210174 629188 210202
rect 629404 210174 629740 210202
rect 629864 210174 630292 210202
rect 630692 210174 630844 210202
rect 631060 210174 631396 210202
rect 631612 210174 631948 210202
rect 632716 210174 633052 210202
rect 633452 210174 633604 210202
rect 633820 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210174 635596 210202
rect 636364 210174 636700 210202
rect 636916 210174 637252 210202
rect 638020 210174 638356 210202
rect 638572 210174 638908 210202
rect 639676 210174 640012 210202
rect 640228 210174 640288 210202
rect 641332 210174 641668 210202
rect 641824 210202 641852 230930
rect 642008 229094 642036 278015
rect 642744 271153 642772 277780
rect 643744 274712 643796 274718
rect 643744 274654 643796 274660
rect 642730 271144 642786 271153
rect 642730 271079 642786 271088
rect 643756 265674 643784 274654
rect 643940 273970 643968 277780
rect 643928 273964 643980 273970
rect 643928 273906 643980 273912
rect 643744 265668 643796 265674
rect 643744 265610 643796 265616
rect 643100 231668 643152 231674
rect 643100 231610 643152 231616
rect 642008 229066 642588 229094
rect 642560 210202 642588 229066
rect 643112 210202 643140 231610
rect 644480 231260 644532 231266
rect 644480 231202 644532 231208
rect 644492 229094 644520 231202
rect 644492 229066 644612 229094
rect 644584 212534 644612 229066
rect 644492 212506 644612 212534
rect 644492 211070 644520 212506
rect 644480 211064 644532 211070
rect 644480 211006 644532 211012
rect 644676 210746 644704 278394
rect 645136 274718 645164 277780
rect 645872 277766 646346 277794
rect 647252 277766 647542 277794
rect 645124 274712 645176 274718
rect 645124 274654 645176 274660
rect 645872 268530 645900 277766
rect 647252 269822 647280 277766
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 648632 276842 648660 277366
rect 648540 276814 648660 276842
rect 648540 276570 648568 276814
rect 648710 276720 648766 276729
rect 648710 276655 648766 276664
rect 648540 276542 648660 276570
rect 648632 275346 648660 276542
rect 648540 275330 648660 275346
rect 648528 275324 648660 275330
rect 648580 275318 648660 275324
rect 648528 275266 648580 275272
rect 647240 269816 647292 269822
rect 647240 269758 647292 269764
rect 645860 268524 645912 268530
rect 645860 268466 645912 268472
rect 646044 231804 646096 231810
rect 646044 231746 646096 231752
rect 645860 231396 645912 231402
rect 645860 231338 645912 231344
rect 644848 211064 644900 211070
rect 644848 211006 644900 211012
rect 644584 210718 644704 210746
rect 644584 210202 644612 210718
rect 644860 210202 644888 211006
rect 645872 210202 645900 231338
rect 646056 229094 646084 231746
rect 648724 229094 648752 276655
rect 648908 229094 648936 990082
rect 646056 229066 646452 229094
rect 648724 229066 648844 229094
rect 648908 229066 649028 229094
rect 646424 210202 646452 229066
rect 647330 228848 647386 228857
rect 647330 228783 647386 228792
rect 647344 215294 647372 228783
rect 648066 227216 648122 227225
rect 648066 227151 648122 227160
rect 647344 215266 647556 215294
rect 647528 210202 647556 215266
rect 648080 210202 648108 227151
rect 648816 215294 648844 229066
rect 649000 215294 649028 229066
rect 648816 215266 648936 215294
rect 649000 215266 649120 215294
rect 648908 210338 648936 215266
rect 649092 213382 649120 215266
rect 650012 213790 650040 993006
rect 651380 992928 651432 992934
rect 651380 992870 651432 992876
rect 650736 991500 650788 991506
rect 650736 991442 650788 991448
rect 650184 988780 650236 988786
rect 650184 988722 650236 988728
rect 650000 213784 650052 213790
rect 650000 213726 650052 213732
rect 650196 213518 650224 988722
rect 650368 984632 650420 984638
rect 650368 984574 650420 984580
rect 650184 213512 650236 213518
rect 650184 213454 650236 213460
rect 649080 213376 649132 213382
rect 649080 213318 649132 213324
rect 650380 212974 650408 984574
rect 650552 231532 650604 231538
rect 650552 231474 650604 231480
rect 650368 212968 650420 212974
rect 650368 212910 650420 212916
rect 648908 210310 649212 210338
rect 649184 210202 649212 210310
rect 650564 210202 650592 231474
rect 650748 213246 650776 991442
rect 650920 987420 650972 987426
rect 650920 987362 650972 987368
rect 650736 213240 650788 213246
rect 650736 213182 650788 213188
rect 650932 213110 650960 987362
rect 651102 227488 651158 227497
rect 651102 227423 651158 227432
rect 650920 213104 650972 213110
rect 650920 213046 650972 213052
rect 641824 210174 641884 210202
rect 642560 210174 642988 210202
rect 643112 210174 643540 210202
rect 644584 210174 644644 210202
rect 644860 210174 645196 210202
rect 645872 210174 646300 210202
rect 646424 210174 646852 210202
rect 647528 210174 647956 210202
rect 648080 210174 648508 210202
rect 649184 210174 649612 210202
rect 650164 210174 650592 210202
rect 651116 210202 651144 227423
rect 651392 213926 651420 992870
rect 651748 991636 651800 991642
rect 651748 991578 651800 991584
rect 651562 975896 651618 975905
rect 651562 975831 651618 975840
rect 651576 975730 651604 975831
rect 651564 975724 651616 975730
rect 651564 975666 651616 975672
rect 651562 962568 651618 962577
rect 651562 962503 651618 962512
rect 651576 961926 651604 962503
rect 651564 961920 651616 961926
rect 651564 961862 651616 961868
rect 651562 949376 651618 949385
rect 651562 949311 651618 949320
rect 651576 948122 651604 949311
rect 651564 948116 651616 948122
rect 651564 948058 651616 948064
rect 651564 937032 651616 937038
rect 651564 936974 651616 936980
rect 651576 936193 651604 936974
rect 651562 936184 651618 936193
rect 651562 936119 651618 936128
rect 651562 922720 651618 922729
rect 651562 922655 651618 922664
rect 651576 921874 651604 922655
rect 651564 921868 651616 921874
rect 651564 921810 651616 921816
rect 651562 909528 651618 909537
rect 651562 909463 651564 909472
rect 651616 909463 651618 909472
rect 651564 909434 651616 909440
rect 651562 896200 651618 896209
rect 651562 896135 651618 896144
rect 651576 895694 651604 896135
rect 651564 895688 651616 895694
rect 651564 895630 651616 895636
rect 651562 869680 651618 869689
rect 651562 869615 651618 869624
rect 651576 869446 651604 869615
rect 651564 869440 651616 869446
rect 651564 869382 651616 869388
rect 651562 856352 651618 856361
rect 651562 856287 651618 856296
rect 651576 855642 651604 856287
rect 651564 855636 651616 855642
rect 651564 855578 651616 855584
rect 651562 843024 651618 843033
rect 651562 842959 651618 842968
rect 651576 841838 651604 842959
rect 651564 841832 651616 841838
rect 651564 841774 651616 841780
rect 651562 829832 651618 829841
rect 651562 829767 651618 829776
rect 651576 829462 651604 829767
rect 651564 829456 651616 829462
rect 651564 829398 651616 829404
rect 651562 816504 651618 816513
rect 651562 816439 651618 816448
rect 651576 815658 651604 816439
rect 651564 815652 651616 815658
rect 651564 815594 651616 815600
rect 651562 803312 651618 803321
rect 651562 803247 651564 803256
rect 651616 803247 651618 803256
rect 651564 803218 651616 803224
rect 651562 789984 651618 789993
rect 651562 789919 651618 789928
rect 651576 789410 651604 789919
rect 651564 789404 651616 789410
rect 651564 789346 651616 789352
rect 651562 776656 651618 776665
rect 651562 776591 651618 776600
rect 651576 775606 651604 776591
rect 651564 775600 651616 775606
rect 651564 775542 651616 775548
rect 651562 763328 651618 763337
rect 651562 763263 651564 763272
rect 651616 763263 651618 763272
rect 651564 763234 651616 763240
rect 651562 750136 651618 750145
rect 651562 750071 651618 750080
rect 651576 749426 651604 750071
rect 651564 749420 651616 749426
rect 651564 749362 651616 749368
rect 651562 736808 651618 736817
rect 651562 736743 651618 736752
rect 651576 735622 651604 736743
rect 651564 735616 651616 735622
rect 651564 735558 651616 735564
rect 651562 723480 651618 723489
rect 651562 723415 651618 723424
rect 651576 723178 651604 723415
rect 651564 723172 651616 723178
rect 651564 723114 651616 723120
rect 651562 710288 651618 710297
rect 651562 710223 651618 710232
rect 651576 709374 651604 710223
rect 651564 709368 651616 709374
rect 651564 709310 651616 709316
rect 651564 696992 651616 696998
rect 651562 696960 651564 696969
rect 651616 696960 651618 696969
rect 651562 696895 651618 696904
rect 651562 683632 651618 683641
rect 651562 683567 651618 683576
rect 651576 683194 651604 683567
rect 651564 683188 651616 683194
rect 651564 683130 651616 683136
rect 651562 670440 651618 670449
rect 651562 670375 651618 670384
rect 651576 669390 651604 670375
rect 651564 669384 651616 669390
rect 651564 669326 651616 669332
rect 651562 657112 651618 657121
rect 651562 657047 651618 657056
rect 651576 656946 651604 657047
rect 651564 656940 651616 656946
rect 651564 656882 651616 656888
rect 651562 643784 651618 643793
rect 651562 643719 651618 643728
rect 651576 643142 651604 643719
rect 651564 643136 651616 643142
rect 651564 643078 651616 643084
rect 651562 630592 651618 630601
rect 651562 630527 651618 630536
rect 651576 629338 651604 630527
rect 651564 629332 651616 629338
rect 651564 629274 651616 629280
rect 651562 617264 651618 617273
rect 651562 617199 651618 617208
rect 651576 616894 651604 617199
rect 651564 616888 651616 616894
rect 651564 616830 651616 616836
rect 651562 590744 651618 590753
rect 651562 590679 651564 590688
rect 651616 590679 651618 590688
rect 651564 590650 651616 590656
rect 651562 577416 651618 577425
rect 651562 577351 651618 577360
rect 651576 576910 651604 577351
rect 651564 576904 651616 576910
rect 651564 576846 651616 576852
rect 651562 550896 651618 550905
rect 651562 550831 651618 550840
rect 651576 550662 651604 550831
rect 651564 550656 651616 550662
rect 651564 550598 651616 550604
rect 651562 537568 651618 537577
rect 651562 537503 651618 537512
rect 651576 536858 651604 537503
rect 651564 536852 651616 536858
rect 651564 536794 651616 536800
rect 651562 524240 651618 524249
rect 651562 524175 651618 524184
rect 651576 523054 651604 524175
rect 651564 523048 651616 523054
rect 651564 522990 651616 522996
rect 651562 511048 651618 511057
rect 651562 510983 651618 510992
rect 651576 510678 651604 510983
rect 651564 510672 651616 510678
rect 651564 510614 651616 510620
rect 651562 497720 651618 497729
rect 651562 497655 651618 497664
rect 651576 496874 651604 497655
rect 651564 496868 651616 496874
rect 651564 496810 651616 496816
rect 651562 484528 651618 484537
rect 651562 484463 651564 484472
rect 651616 484463 651618 484472
rect 651564 484434 651616 484440
rect 651562 471200 651618 471209
rect 651562 471135 651618 471144
rect 651576 470626 651604 471135
rect 651564 470620 651616 470626
rect 651564 470562 651616 470568
rect 651562 457872 651618 457881
rect 651562 457807 651618 457816
rect 651576 456822 651604 457807
rect 651564 456816 651616 456822
rect 651564 456758 651616 456764
rect 651562 444544 651618 444553
rect 651562 444479 651564 444488
rect 651616 444479 651618 444488
rect 651564 444450 651616 444456
rect 651562 431352 651618 431361
rect 651562 431287 651618 431296
rect 651576 430642 651604 431287
rect 651564 430636 651616 430642
rect 651564 430578 651616 430584
rect 651562 418024 651618 418033
rect 651562 417959 651618 417968
rect 651576 416838 651604 417959
rect 651564 416832 651616 416838
rect 651564 416774 651616 416780
rect 651562 404696 651618 404705
rect 651562 404631 651618 404640
rect 651576 404394 651604 404631
rect 651564 404388 651616 404394
rect 651564 404330 651616 404336
rect 651562 391504 651618 391513
rect 651562 391439 651618 391448
rect 651576 390590 651604 391439
rect 651564 390584 651616 390590
rect 651564 390526 651616 390532
rect 651564 378208 651616 378214
rect 651562 378176 651564 378185
rect 651616 378176 651618 378185
rect 651562 378111 651618 378120
rect 651562 364848 651618 364857
rect 651562 364783 651618 364792
rect 651576 364410 651604 364783
rect 651564 364404 651616 364410
rect 651564 364346 651616 364352
rect 651562 325000 651618 325009
rect 651562 324935 651618 324944
rect 651576 324358 651604 324935
rect 651564 324352 651616 324358
rect 651564 324294 651616 324300
rect 651562 311808 651618 311817
rect 651562 311743 651618 311752
rect 651576 310554 651604 311743
rect 651564 310548 651616 310554
rect 651564 310490 651616 310496
rect 651562 285288 651618 285297
rect 651562 285223 651618 285232
rect 651576 284374 651604 285223
rect 651564 284368 651616 284374
rect 651564 284310 651616 284316
rect 651562 228304 651618 228313
rect 651562 228239 651618 228248
rect 651380 213920 651432 213926
rect 651380 213862 651432 213868
rect 651576 210202 651604 228239
rect 651760 213654 651788 991578
rect 658924 985992 658976 985998
rect 658924 985934 658976 985940
rect 658936 937242 658964 985934
rect 660304 984904 660356 984910
rect 660304 984846 660356 984852
rect 660316 937378 660344 984846
rect 661684 975724 661736 975730
rect 661684 975666 661736 975672
rect 660488 957772 660540 957778
rect 660488 957714 660540 957720
rect 660304 937372 660356 937378
rect 660304 937314 660356 937320
rect 658924 937236 658976 937242
rect 658924 937178 658976 937184
rect 660500 937038 660528 957714
rect 661696 938466 661724 975666
rect 663064 961920 663116 961926
rect 663064 961862 663116 961868
rect 663076 941866 663104 961862
rect 663064 941860 663116 941866
rect 663064 941802 663116 941808
rect 661684 938460 661736 938466
rect 661684 938402 661736 938408
rect 660488 937032 660540 937038
rect 660488 936974 660540 936980
rect 661684 921868 661736 921874
rect 661684 921810 661736 921816
rect 652390 882872 652446 882881
rect 652390 882807 652446 882816
rect 652404 881890 652432 882807
rect 652392 881884 652444 881890
rect 652392 881826 652444 881832
rect 658924 869440 658976 869446
rect 658924 869382 658976 869388
rect 658936 715018 658964 869382
rect 659108 841832 659160 841838
rect 659108 841774 659160 841780
rect 659120 715154 659148 841774
rect 660304 829456 660356 829462
rect 660304 829398 660356 829404
rect 660316 779006 660344 829398
rect 660304 779000 660356 779006
rect 660304 778942 660356 778948
rect 660488 775600 660540 775606
rect 660488 775542 660540 775548
rect 660304 763224 660356 763230
rect 660304 763166 660356 763172
rect 659292 723172 659344 723178
rect 659292 723114 659344 723120
rect 659108 715148 659160 715154
rect 659108 715090 659160 715096
rect 658924 715012 658976 715018
rect 658924 714954 658976 714960
rect 658924 709368 658976 709374
rect 658924 709310 658976 709316
rect 652574 603936 652630 603945
rect 652574 603871 652630 603880
rect 652588 603158 652616 603871
rect 652576 603152 652628 603158
rect 652576 603094 652628 603100
rect 658936 579834 658964 709310
rect 659304 689314 659332 723114
rect 659292 689308 659344 689314
rect 659292 689250 659344 689256
rect 659108 683188 659160 683194
rect 659108 683130 659160 683136
rect 658924 579828 658976 579834
rect 658924 579770 658976 579776
rect 659120 579698 659148 683130
rect 660316 625190 660344 763166
rect 660500 734874 660528 775542
rect 661696 760578 661724 921810
rect 664444 909492 664496 909498
rect 664444 909434 664496 909440
rect 663064 895688 663116 895694
rect 663064 895630 663116 895636
rect 661868 815652 661920 815658
rect 661868 815594 661920 815600
rect 661684 760572 661736 760578
rect 661684 760514 661736 760520
rect 660488 734868 660540 734874
rect 660488 734810 660540 734816
rect 661880 670750 661908 815594
rect 662052 789404 662104 789410
rect 662052 789346 662104 789352
rect 661868 670744 661920 670750
rect 661868 670686 661920 670692
rect 662064 669390 662092 789346
rect 663076 760442 663104 895630
rect 663248 803276 663300 803282
rect 663248 803218 663300 803224
rect 663064 760436 663116 760442
rect 663064 760378 663116 760384
rect 663064 735616 663116 735622
rect 663064 735558 663116 735564
rect 661868 669384 661920 669390
rect 661868 669326 661920 669332
rect 662052 669384 662104 669390
rect 662052 669326 662104 669332
rect 661684 656940 661736 656946
rect 661684 656882 661736 656888
rect 660304 625184 660356 625190
rect 660304 625126 660356 625132
rect 660488 616888 660540 616894
rect 660488 616830 660540 616836
rect 660304 603152 660356 603158
rect 660304 603094 660356 603100
rect 659108 579692 659160 579698
rect 659108 579634 659160 579640
rect 659292 576904 659344 576910
rect 659292 576846 659344 576852
rect 652390 564088 652446 564097
rect 652390 564023 652446 564032
rect 652404 563106 652432 564023
rect 652392 563100 652444 563106
rect 652392 563042 652444 563048
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 658936 554062 658964 563042
rect 658924 554056 658976 554062
rect 658924 553998 658976 554004
rect 658924 550656 658976 550662
rect 658924 550598 658976 550604
rect 658936 403034 658964 550598
rect 659108 496868 659160 496874
rect 659108 496810 659160 496816
rect 658924 403028 658976 403034
rect 658924 402970 658976 402976
rect 659120 357746 659148 496810
rect 659304 491366 659332 576846
rect 660316 491502 660344 603094
rect 660500 599622 660528 616830
rect 660488 599616 660540 599622
rect 660488 599558 660540 599564
rect 661696 535498 661724 656882
rect 661880 643754 661908 669326
rect 661868 643748 661920 643754
rect 661868 643690 661920 643696
rect 661868 629332 661920 629338
rect 661868 629274 661920 629280
rect 661684 535492 661736 535498
rect 661684 535434 661736 535440
rect 661880 534274 661908 629274
rect 663076 625462 663104 735558
rect 663260 670886 663288 803218
rect 664456 760918 664484 909434
rect 664444 760912 664496 760918
rect 664444 760854 664496 760860
rect 664444 749420 664496 749426
rect 664444 749362 664496 749368
rect 663248 670880 663300 670886
rect 663248 670822 663300 670828
rect 663248 643136 663300 643142
rect 663248 643078 663300 643084
rect 663064 625456 663116 625462
rect 663064 625398 663116 625404
rect 663064 536852 663116 536858
rect 663064 536794 663116 536800
rect 661868 534268 661920 534274
rect 661868 534210 661920 534216
rect 661684 523048 661736 523054
rect 661684 522990 661736 522996
rect 660488 510672 660540 510678
rect 660488 510614 660540 510620
rect 660304 491496 660356 491502
rect 660304 491438 660356 491444
rect 659292 491360 659344 491366
rect 659292 491302 659344 491308
rect 660304 430636 660356 430642
rect 660304 430578 660356 430584
rect 659292 404388 659344 404394
rect 659292 404330 659344 404336
rect 659108 357740 659160 357746
rect 659108 357682 659160 357688
rect 652022 351656 652078 351665
rect 652022 351591 652078 351600
rect 651748 213648 651800 213654
rect 651748 213590 651800 213596
rect 652036 210458 652064 351591
rect 652206 338328 652262 338337
rect 652206 338263 652262 338272
rect 652220 338162 652248 338263
rect 652208 338156 652260 338162
rect 652208 338098 652260 338104
rect 652206 298480 652262 298489
rect 652206 298415 652262 298424
rect 652024 210452 652076 210458
rect 652024 210394 652076 210400
rect 651116 210174 651268 210202
rect 651576 210174 651820 210202
rect 608600 210112 608652 210118
rect 608600 210054 608652 210060
rect 608968 210112 609020 210118
rect 609020 210060 609316 210066
rect 608968 210054 609316 210060
rect 608980 210038 609316 210054
rect 591304 209840 591356 209846
rect 591304 209782 591356 209788
rect 632152 209840 632204 209846
rect 632204 209788 632500 209794
rect 632152 209782 632500 209788
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208185 589504 208286
rect 589462 208176 589518 208185
rect 589462 208111 589518 208120
rect 589464 206984 589516 206990
rect 589464 206926 589516 206932
rect 589476 206553 589504 206926
rect 589462 206544 589518 206553
rect 589462 206479 589518 206488
rect 583300 205624 583352 205630
rect 583300 205566 583352 205572
rect 589464 205624 589516 205630
rect 589464 205566 589516 205572
rect 584404 205284 584456 205290
rect 584404 205226 584456 205232
rect 583208 202904 583260 202910
rect 583208 202846 583260 202852
rect 581828 200796 581880 200802
rect 581828 200738 581880 200744
rect 581736 200456 581788 200462
rect 581736 200398 581788 200404
rect 581748 196654 581776 200398
rect 583024 198756 583076 198762
rect 583024 198698 583076 198704
rect 581736 196648 581788 196654
rect 581736 196590 581788 196596
rect 581644 196172 581696 196178
rect 581644 196114 581696 196120
rect 580908 194540 580960 194546
rect 580908 194482 580960 194488
rect 581656 188970 581684 196114
rect 583036 190466 583064 198698
rect 583220 195974 583248 202846
rect 584416 197334 584444 205226
rect 589476 204921 589504 205566
rect 589462 204912 589518 204921
rect 589462 204847 589518 204856
rect 589464 204196 589516 204202
rect 589464 204138 589516 204144
rect 589476 203289 589504 204138
rect 589462 203280 589518 203289
rect 589462 203215 589518 203224
rect 589372 202768 589424 202774
rect 589372 202710 589424 202716
rect 589384 201657 589412 202710
rect 589370 201648 589426 201657
rect 589370 201583 589426 201592
rect 590384 200796 590436 200802
rect 590384 200738 590436 200744
rect 589464 200048 589516 200054
rect 589462 200016 589464 200025
rect 589516 200016 589518 200025
rect 589462 199951 589518 199960
rect 590396 198393 590424 200738
rect 590382 198384 590438 198393
rect 590382 198319 590438 198328
rect 584404 197328 584456 197334
rect 584404 197270 584456 197276
rect 589464 197328 589516 197334
rect 589464 197270 589516 197276
rect 589476 196761 589504 197270
rect 589462 196752 589518 196761
rect 589462 196687 589518 196696
rect 589648 196648 589700 196654
rect 589648 196590 589700 196596
rect 583208 195968 583260 195974
rect 583208 195910 583260 195916
rect 589464 195968 589516 195974
rect 589464 195910 589516 195916
rect 589476 195129 589504 195910
rect 589462 195120 589518 195129
rect 589462 195055 589518 195064
rect 589464 194540 589516 194546
rect 589464 194482 589516 194488
rect 589476 193497 589504 194482
rect 589462 193488 589518 193497
rect 583760 193452 583812 193458
rect 589462 193423 589518 193432
rect 583760 193394 583812 193400
rect 583772 191146 583800 193394
rect 588544 191888 588596 191894
rect 588544 191830 588596 191836
rect 583760 191140 583812 191146
rect 583760 191082 583812 191088
rect 583024 190460 583076 190466
rect 583024 190402 583076 190408
rect 585968 189100 586020 189106
rect 585968 189042 586020 189048
rect 581644 188964 581696 188970
rect 581644 188906 581696 188912
rect 581828 188828 581880 188834
rect 581828 188770 581880 188776
rect 580264 187604 580316 187610
rect 580264 187546 580316 187552
rect 578884 186244 578936 186250
rect 578884 186186 578936 186192
rect 578330 185872 578386 185881
rect 578330 185807 578386 185816
rect 578344 185298 578372 185807
rect 578332 185292 578384 185298
rect 578332 185234 578384 185240
rect 580448 185292 580500 185298
rect 580448 185234 580500 185240
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579540 183598 579568 184311
rect 579528 183592 579580 183598
rect 579528 183534 579580 183540
rect 578882 182880 578938 182889
rect 578882 182815 578938 182824
rect 578896 182238 578924 182815
rect 578884 182232 578936 182238
rect 578884 182174 578936 182180
rect 578514 181384 578570 181393
rect 578514 181319 578516 181328
rect 578568 181319 578570 181328
rect 578516 181290 578568 181296
rect 578974 179888 579030 179897
rect 578974 179823 579030 179832
rect 578988 179722 579016 179823
rect 578976 179716 579028 179722
rect 578976 179658 579028 179664
rect 578606 178392 578662 178401
rect 578606 178327 578608 178336
rect 578660 178327 578662 178336
rect 580264 178356 580316 178362
rect 578608 178298 578660 178304
rect 580264 178298 580316 178304
rect 579526 176896 579582 176905
rect 579526 176831 579528 176840
rect 579580 176831 579582 176840
rect 579528 176802 579580 176808
rect 579434 175536 579490 175545
rect 579490 175494 579660 175522
rect 579434 175471 579490 175480
rect 579632 174554 579660 175494
rect 579620 174548 579672 174554
rect 579620 174490 579672 174496
rect 578330 173904 578386 173913
rect 578330 173839 578386 173848
rect 578344 172582 578372 173839
rect 578332 172576 578384 172582
rect 578332 172518 578384 172524
rect 579066 172408 579122 172417
rect 579066 172343 579122 172352
rect 579080 171698 579108 172343
rect 579068 171692 579120 171698
rect 579068 171634 579120 171640
rect 579526 170912 579582 170921
rect 579526 170847 579582 170856
rect 579540 169794 579568 170847
rect 579528 169788 579580 169794
rect 579528 169730 579580 169736
rect 578238 169416 578294 169425
rect 578238 169351 578294 169360
rect 578252 168434 578280 169351
rect 578240 168428 578292 168434
rect 578240 168370 578292 168376
rect 580276 168298 580304 178298
rect 580460 176594 580488 185234
rect 581644 181348 581696 181354
rect 581644 181290 581696 181296
rect 580448 176588 580500 176594
rect 580448 176530 580500 176536
rect 581656 171018 581684 181290
rect 581840 179314 581868 188770
rect 584588 187196 584640 187202
rect 584588 187138 584640 187144
rect 583024 182232 583076 182238
rect 583024 182174 583076 182180
rect 581828 179308 581880 179314
rect 581828 179250 581880 179256
rect 583036 172446 583064 182174
rect 584600 178022 584628 187138
rect 585980 180810 586008 189042
rect 587164 183592 587216 183598
rect 587164 183534 587216 183540
rect 585968 180804 586020 180810
rect 585968 180746 586020 180752
rect 585784 179716 585836 179722
rect 585784 179658 585836 179664
rect 584588 178016 584640 178022
rect 584588 177958 584640 177964
rect 584404 176860 584456 176866
rect 584404 176802 584456 176808
rect 583208 172576 583260 172582
rect 583208 172518 583260 172524
rect 583024 172440 583076 172446
rect 583024 172382 583076 172388
rect 581828 171692 581880 171698
rect 581828 171634 581880 171640
rect 581644 171012 581696 171018
rect 581644 170954 581696 170960
rect 580448 168428 580500 168434
rect 580448 168370 580500 168376
rect 580264 168292 580316 168298
rect 580264 168234 580316 168240
rect 579434 167920 579490 167929
rect 579490 167878 579660 167906
rect 579434 167855 579490 167864
rect 579066 166424 579122 166433
rect 579066 166359 579122 166368
rect 579080 165646 579108 166359
rect 579632 166326 579660 167878
rect 579620 166320 579672 166326
rect 579620 166262 579672 166268
rect 579068 165640 579120 165646
rect 579068 165582 579120 165588
rect 579526 164384 579582 164393
rect 579526 164319 579528 164328
rect 579580 164319 579582 164328
rect 579528 164290 579580 164296
rect 578698 163432 578754 163441
rect 578698 163367 578754 163376
rect 578712 162926 578740 163367
rect 578700 162920 578752 162926
rect 578700 162862 578752 162868
rect 578882 161936 578938 161945
rect 578882 161871 578938 161880
rect 578514 160440 578570 160449
rect 578514 160375 578570 160384
rect 578528 160274 578556 160375
rect 578516 160268 578568 160274
rect 578516 160210 578568 160216
rect 578698 152960 578754 152969
rect 578698 152895 578754 152904
rect 578712 152318 578740 152895
rect 578700 152312 578752 152318
rect 578700 152254 578752 152260
rect 578896 150346 578924 161871
rect 580264 160268 580316 160274
rect 580264 160210 580316 160216
rect 579526 158944 579582 158953
rect 579526 158879 579582 158888
rect 579540 158778 579568 158879
rect 579528 158772 579580 158778
rect 579528 158714 579580 158720
rect 579434 157448 579490 157457
rect 579490 157406 579660 157434
rect 579434 157383 579490 157392
rect 579632 156670 579660 157406
rect 579620 156664 579672 156670
rect 579620 156606 579672 156612
rect 579250 155952 579306 155961
rect 579250 155887 579306 155896
rect 579264 154630 579292 155887
rect 579252 154624 579304 154630
rect 579252 154566 579304 154572
rect 579250 154456 579306 154465
rect 579250 154391 579306 154400
rect 579264 153338 579292 154391
rect 579252 153332 579304 153338
rect 579252 153274 579304 153280
rect 579158 151464 579214 151473
rect 579158 151399 579214 151408
rect 579172 150482 579200 151399
rect 579160 150476 579212 150482
rect 579160 150418 579212 150424
rect 578884 150340 578936 150346
rect 578884 150282 578936 150288
rect 578882 149968 578938 149977
rect 578882 149903 578938 149912
rect 578896 149122 578924 149903
rect 578884 149116 578936 149122
rect 578884 149058 578936 149064
rect 579526 148472 579582 148481
rect 579526 148407 579582 148416
rect 579540 147694 579568 148407
rect 579528 147688 579580 147694
rect 579528 147630 579580 147636
rect 579252 147552 579304 147558
rect 579252 147494 579304 147500
rect 579264 146985 579292 147494
rect 580276 147422 580304 160210
rect 580460 158642 580488 168370
rect 581644 162920 581696 162926
rect 581644 162862 581696 162868
rect 580448 158636 580500 158642
rect 580448 158578 580500 158584
rect 581656 151706 581684 162862
rect 581840 161430 581868 171634
rect 583024 164348 583076 164354
rect 583024 164290 583076 164296
rect 581828 161424 581880 161430
rect 581828 161366 581880 161372
rect 583036 153134 583064 164290
rect 583220 162858 583248 172518
rect 584416 165510 584444 176802
rect 585796 169658 585824 179658
rect 587176 173874 587204 183534
rect 588556 182073 588584 191830
rect 589660 191729 589688 196590
rect 589646 191720 589702 191729
rect 589646 191655 589702 191664
rect 590384 191140 590436 191146
rect 590384 191082 590436 191088
rect 589464 190460 589516 190466
rect 589464 190402 589516 190408
rect 589476 190233 589504 190402
rect 589462 190224 589518 190233
rect 589462 190159 589518 190168
rect 589464 188964 589516 188970
rect 589464 188906 589516 188912
rect 589476 188601 589504 188906
rect 589462 188592 589518 188601
rect 589462 188527 589518 188536
rect 589372 187604 589424 187610
rect 589372 187546 589424 187552
rect 589384 186969 589412 187546
rect 589370 186960 589426 186969
rect 589370 186895 589426 186904
rect 589464 186244 589516 186250
rect 589464 186186 589516 186192
rect 589476 185337 589504 186186
rect 589462 185328 589518 185337
rect 589462 185263 589518 185272
rect 590396 183569 590424 191082
rect 590382 183560 590438 183569
rect 590382 183495 590438 183504
rect 588542 182064 588598 182073
rect 588542 181999 588598 182008
rect 589464 180804 589516 180810
rect 589464 180746 589516 180752
rect 589476 180441 589504 180746
rect 589462 180432 589518 180441
rect 589462 180367 589518 180376
rect 589556 179308 589608 179314
rect 589556 179250 589608 179256
rect 589568 178809 589596 179250
rect 589554 178800 589610 178809
rect 589554 178735 589610 178744
rect 589464 178016 589516 178022
rect 589464 177958 589516 177964
rect 589476 177177 589504 177958
rect 589462 177168 589518 177177
rect 589462 177103 589518 177112
rect 589464 176588 589516 176594
rect 589464 176530 589516 176536
rect 589476 175545 589504 176530
rect 589462 175536 589518 175545
rect 589462 175471 589518 175480
rect 589924 174548 589976 174554
rect 589924 174490 589976 174496
rect 589278 173904 589334 173913
rect 587164 173868 587216 173874
rect 589278 173839 589280 173848
rect 587164 173810 587216 173816
rect 589332 173839 589334 173848
rect 589280 173810 589332 173816
rect 589372 172440 589424 172446
rect 589372 172382 589424 172388
rect 589384 172281 589412 172382
rect 589370 172272 589426 172281
rect 589370 172207 589426 172216
rect 589464 171012 589516 171018
rect 589464 170954 589516 170960
rect 589476 170649 589504 170954
rect 589462 170640 589518 170649
rect 589462 170575 589518 170584
rect 588728 169788 588780 169794
rect 588728 169730 588780 169736
rect 585784 169652 585836 169658
rect 585784 169594 585836 169600
rect 584588 165640 584640 165646
rect 584588 165582 584640 165588
rect 584404 165504 584456 165510
rect 584404 165446 584456 165452
rect 583208 162852 583260 162858
rect 583208 162794 583260 162800
rect 584600 154494 584628 165582
rect 588740 159225 588768 169730
rect 589464 169652 589516 169658
rect 589464 169594 589516 169600
rect 589476 169017 589504 169594
rect 589462 169008 589518 169017
rect 589462 168943 589518 168952
rect 589464 168292 589516 168298
rect 589464 168234 589516 168240
rect 589476 167385 589504 168234
rect 589462 167376 589518 167385
rect 589462 167311 589518 167320
rect 589462 165608 589518 165617
rect 589462 165543 589464 165552
rect 589516 165543 589518 165552
rect 589464 165514 589516 165520
rect 589936 164121 589964 174490
rect 590384 166320 590436 166326
rect 590384 166262 590436 166268
rect 589922 164112 589978 164121
rect 589922 164047 589978 164056
rect 589464 162852 589516 162858
rect 589464 162794 589516 162800
rect 589476 162489 589504 162794
rect 589462 162480 589518 162489
rect 589462 162415 589518 162424
rect 589464 161424 589516 161430
rect 589464 161366 589516 161372
rect 589476 160857 589504 161366
rect 589462 160848 589518 160857
rect 589462 160783 589518 160792
rect 588726 159216 588782 159225
rect 588726 159151 588782 159160
rect 588544 158772 588596 158778
rect 588544 158714 588596 158720
rect 587348 154624 587400 154630
rect 587348 154566 587400 154572
rect 584588 154488 584640 154494
rect 584588 154430 584640 154436
rect 585784 153332 585836 153338
rect 585784 153274 585836 153280
rect 583024 153128 583076 153134
rect 583024 153070 583076 153076
rect 584404 152312 584456 152318
rect 584404 152254 584456 152260
rect 581644 151700 581696 151706
rect 581644 151642 581696 151648
rect 583208 150476 583260 150482
rect 583208 150418 583260 150424
rect 581644 149116 581696 149122
rect 581644 149058 581696 149064
rect 580264 147416 580316 147422
rect 580264 147358 580316 147364
rect 579250 146976 579306 146985
rect 579250 146911 579306 146920
rect 579434 145480 579490 145489
rect 579490 145438 579660 145466
rect 579434 145415 579490 145424
rect 579632 144226 579660 145438
rect 579620 144220 579672 144226
rect 579620 144162 579672 144168
rect 578514 143984 578570 143993
rect 578514 143919 578570 143928
rect 578528 143682 578556 143919
rect 578516 143676 578568 143682
rect 578516 143618 578568 143624
rect 580264 143676 580316 143682
rect 580264 143618 580316 143624
rect 579526 142488 579582 142497
rect 579526 142423 579582 142432
rect 579540 142186 579568 142423
rect 579528 142180 579580 142186
rect 579528 142122 579580 142128
rect 578882 140992 578938 141001
rect 578882 140927 578938 140936
rect 578238 135008 578294 135017
rect 578238 134943 578294 134952
rect 578252 134570 578280 134943
rect 578240 134564 578292 134570
rect 578240 134506 578292 134512
rect 578514 133512 578570 133521
rect 578514 133447 578570 133456
rect 578528 132938 578556 133447
rect 578516 132932 578568 132938
rect 578516 132874 578568 132880
rect 578422 132016 578478 132025
rect 578422 131951 578478 131960
rect 578436 130422 578464 131951
rect 578606 130520 578662 130529
rect 578606 130455 578662 130464
rect 578424 130416 578476 130422
rect 578424 130358 578476 130364
rect 578620 129946 578648 130455
rect 578608 129940 578660 129946
rect 578608 129882 578660 129888
rect 578896 128382 578924 140927
rect 579526 139496 579582 139505
rect 579526 139431 579528 139440
rect 579580 139431 579582 139440
rect 579528 139402 579580 139408
rect 579250 138000 579306 138009
rect 579250 137935 579252 137944
rect 579304 137935 579306 137944
rect 579252 137906 579304 137912
rect 579066 136504 579122 136513
rect 579066 136439 579122 136448
rect 579080 135386 579108 136439
rect 579068 135380 579120 135386
rect 579068 135322 579120 135328
rect 580276 132394 580304 143618
rect 581656 136542 581684 149058
rect 583220 137970 583248 150418
rect 584416 140758 584444 152254
rect 585796 142050 585824 153274
rect 587360 143546 587388 154566
rect 588556 146169 588584 158714
rect 589464 158636 589516 158642
rect 589464 158578 589516 158584
rect 589476 157593 589504 158578
rect 589462 157584 589518 157593
rect 589462 157519 589518 157528
rect 589924 156664 589976 156670
rect 589924 156606 589976 156612
rect 589372 154488 589424 154494
rect 589372 154430 589424 154436
rect 589384 154329 589412 154430
rect 589370 154320 589426 154329
rect 589370 154255 589426 154264
rect 589464 153128 589516 153134
rect 589464 153070 589516 153076
rect 589476 152697 589504 153070
rect 589462 152688 589518 152697
rect 589462 152623 589518 152632
rect 589464 151700 589516 151706
rect 589464 151642 589516 151648
rect 589476 151065 589504 151642
rect 589462 151056 589518 151065
rect 589462 150991 589518 151000
rect 589464 150340 589516 150346
rect 589464 150282 589516 150288
rect 589476 149433 589504 150282
rect 589462 149424 589518 149433
rect 589462 149359 589518 149368
rect 588728 147688 588780 147694
rect 588728 147630 588780 147636
rect 589462 147656 589518 147665
rect 588542 146160 588598 146169
rect 588542 146095 588598 146104
rect 587348 143540 587400 143546
rect 587348 143482 587400 143488
rect 587164 142180 587216 142186
rect 587164 142122 587216 142128
rect 585784 142044 585836 142050
rect 585784 141986 585836 141992
rect 584404 140752 584456 140758
rect 584404 140694 584456 140700
rect 584588 139460 584640 139466
rect 584588 139402 584640 139408
rect 583024 137964 583076 137970
rect 583024 137906 583076 137912
rect 583208 137964 583260 137970
rect 583208 137906 583260 137912
rect 581644 136536 581696 136542
rect 581644 136478 581696 136484
rect 581092 135380 581144 135386
rect 581092 135322 581144 135328
rect 581104 133210 581132 135322
rect 581092 133204 581144 133210
rect 581092 133146 581144 133152
rect 581644 132932 581696 132938
rect 581644 132874 581696 132880
rect 580264 132388 580316 132394
rect 580264 132330 580316 132336
rect 580448 129940 580500 129946
rect 580448 129882 580500 129888
rect 579434 129024 579490 129033
rect 579434 128959 579490 128968
rect 578884 128376 578936 128382
rect 578884 128318 578936 128324
rect 578330 127528 578386 127537
rect 578330 127463 578386 127472
rect 578344 127022 578372 127463
rect 578332 127016 578384 127022
rect 578332 126958 578384 126964
rect 579448 126274 579476 128959
rect 580264 127016 580316 127022
rect 580264 126958 580316 126964
rect 579436 126268 579488 126274
rect 579436 126210 579488 126216
rect 578514 126032 578570 126041
rect 578514 125967 578570 125976
rect 578528 125866 578556 125967
rect 578516 125860 578568 125866
rect 578516 125802 578568 125808
rect 578882 124536 578938 124545
rect 578882 124471 578938 124480
rect 578896 124234 578924 124471
rect 578884 124228 578936 124234
rect 578884 124170 578936 124176
rect 578882 123040 578938 123049
rect 578882 122975 578938 122984
rect 578330 117056 578386 117065
rect 578330 116991 578332 117000
rect 578384 116991 578386 117000
rect 578332 116962 578384 116968
rect 578896 109002 578924 122975
rect 579526 121544 579582 121553
rect 579526 121479 579528 121488
rect 579580 121479 579582 121488
rect 579528 121450 579580 121456
rect 580276 120766 580304 126958
rect 580264 120760 580316 120766
rect 580264 120702 580316 120708
rect 579250 120048 579306 120057
rect 579250 119983 579306 119992
rect 579264 118726 579292 119983
rect 579252 118720 579304 118726
rect 579252 118662 579304 118668
rect 579066 118552 579122 118561
rect 579066 118487 579122 118496
rect 579080 117366 579108 118487
rect 579068 117360 579120 117366
rect 579068 117302 579120 117308
rect 580460 117230 580488 129882
rect 581656 120086 581684 132874
rect 583036 124098 583064 137906
rect 584600 129742 584628 139402
rect 585968 134564 586020 134570
rect 585968 134506 586020 134512
rect 584588 129736 584640 129742
rect 584588 129678 584640 129684
rect 584404 125860 584456 125866
rect 584404 125802 584456 125808
rect 583024 124092 583076 124098
rect 583024 124034 583076 124040
rect 583024 121508 583076 121514
rect 583024 121450 583076 121456
rect 581644 120080 581696 120086
rect 581644 120022 581696 120028
rect 581644 117360 581696 117366
rect 581644 117302 581696 117308
rect 580448 117224 580500 117230
rect 580448 117166 580500 117172
rect 580264 117020 580316 117026
rect 580264 116962 580316 116968
rect 578884 108996 578936 109002
rect 578884 108938 578936 108944
rect 580276 102134 580304 116962
rect 581656 104854 581684 117302
rect 583036 107642 583064 121450
rect 584416 111790 584444 125802
rect 585980 124914 586008 134506
rect 587176 126954 587204 142122
rect 588740 134745 588768 147630
rect 589462 147591 589518 147600
rect 589476 147422 589504 147591
rect 589464 147416 589516 147422
rect 589464 147358 589516 147364
rect 589936 144537 589964 156606
rect 590396 155961 590424 166262
rect 590382 155952 590438 155961
rect 590382 155887 590438 155896
rect 591316 147558 591344 209782
rect 632164 209766 632500 209782
rect 652220 209574 652248 298415
rect 658280 278180 658332 278186
rect 658280 278122 658332 278128
rect 656898 276992 656954 277001
rect 656898 276927 656954 276936
rect 655520 276684 655572 276690
rect 655520 276626 655572 276632
rect 652760 231124 652812 231130
rect 652760 231066 652812 231072
rect 652772 210202 652800 231066
rect 654138 230072 654194 230081
rect 654138 230007 654194 230016
rect 653034 228576 653090 228585
rect 653034 228511 653090 228520
rect 653048 210202 653076 228511
rect 654152 210202 654180 230007
rect 654322 229800 654378 229809
rect 654322 229735 654378 229744
rect 654336 229094 654364 229735
rect 654336 229066 654732 229094
rect 654704 210202 654732 229066
rect 655532 214606 655560 276626
rect 655704 264240 655756 264246
rect 655704 264182 655756 264188
rect 655716 229094 655744 264182
rect 656912 229094 656940 276927
rect 655716 229066 655836 229094
rect 656912 229066 657492 229094
rect 655520 214600 655572 214606
rect 655520 214542 655572 214548
rect 655808 210202 655836 229066
rect 656440 214600 656492 214606
rect 656440 214542 656492 214548
rect 656452 210202 656480 214542
rect 657464 210202 657492 229066
rect 658292 210202 658320 278122
rect 659304 268054 659332 404330
rect 659660 278044 659712 278050
rect 659660 277986 659712 277992
rect 659292 268048 659344 268054
rect 659292 267990 659344 267996
rect 658462 265568 658518 265577
rect 658462 265503 658518 265512
rect 658476 229094 658504 265503
rect 658476 229066 659148 229094
rect 659120 210202 659148 229066
rect 659672 214606 659700 277986
rect 660316 267918 660344 430578
rect 660500 357474 660528 510614
rect 660672 444440 660724 444446
rect 660672 444382 660724 444388
rect 660488 357468 660540 357474
rect 660488 357410 660540 357416
rect 660684 312050 660712 444382
rect 661696 403170 661724 522990
rect 661868 470620 661920 470626
rect 661868 470562 661920 470568
rect 661684 403164 661736 403170
rect 661684 403106 661736 403112
rect 661684 390584 661736 390590
rect 661684 390526 661736 390532
rect 660672 312044 660724 312050
rect 660672 311986 660724 311992
rect 661040 278316 661092 278322
rect 661040 278258 661092 278264
rect 660304 267912 660356 267918
rect 660304 267854 660356 267860
rect 659842 226944 659898 226953
rect 659842 226879 659898 226888
rect 659660 214600 659712 214606
rect 659660 214542 659712 214548
rect 659856 210202 659884 226879
rect 660304 214600 660356 214606
rect 660304 214542 660356 214548
rect 660316 210202 660344 214542
rect 661052 210202 661080 278258
rect 661316 230852 661368 230858
rect 661316 230794 661368 230800
rect 661328 214606 661356 230794
rect 661498 225856 661554 225865
rect 661498 225791 661554 225800
rect 661316 214600 661368 214606
rect 661316 214542 661368 214548
rect 661512 210202 661540 225791
rect 661696 222630 661724 390526
rect 661880 313342 661908 470562
rect 663076 403306 663104 536794
rect 663260 535634 663288 643078
rect 664456 625734 664484 749362
rect 664628 696992 664680 696998
rect 664628 696934 664680 696940
rect 664444 625728 664496 625734
rect 664444 625670 664496 625676
rect 663524 608660 663576 608666
rect 663524 608602 663576 608608
rect 663248 535628 663300 535634
rect 663248 535570 663300 535576
rect 663536 531486 663564 608602
rect 664444 590708 664496 590714
rect 664444 590650 664496 590656
rect 663708 564460 663760 564466
rect 663708 564402 663760 564408
rect 663524 531480 663576 531486
rect 663524 531422 663576 531428
rect 663720 485858 663748 564402
rect 664456 491638 664484 590650
rect 664640 581058 664668 696934
rect 664996 654152 665048 654158
rect 664996 654094 665048 654100
rect 664628 581052 664680 581058
rect 664628 580994 664680 581000
rect 665008 574122 665036 654094
rect 664996 574116 665048 574122
rect 664996 574058 665048 574064
rect 664996 564596 665048 564602
rect 664996 564538 665048 564544
rect 664444 491632 664496 491638
rect 664444 491574 664496 491580
rect 663708 485852 663760 485858
rect 663708 485794 663760 485800
rect 665008 484430 665036 564538
rect 664812 484424 664864 484430
rect 664812 484366 664864 484372
rect 664996 484424 665048 484430
rect 664996 484366 665048 484372
rect 663248 456816 663300 456822
rect 663248 456758 663300 456764
rect 663064 403300 663116 403306
rect 663064 403242 663116 403248
rect 663064 378208 663116 378214
rect 663064 378150 663116 378156
rect 661868 313336 661920 313342
rect 661868 313278 661920 313284
rect 662418 225584 662474 225593
rect 662418 225519 662474 225528
rect 661684 222624 661736 222630
rect 661684 222566 661736 222572
rect 661960 214600 662012 214606
rect 661960 214542 662012 214548
rect 661972 210202 662000 214542
rect 662432 210202 662460 225519
rect 662878 222592 662934 222601
rect 662878 222527 662934 222536
rect 662892 219434 662920 222527
rect 663076 222494 663104 378150
rect 663260 313478 663288 456758
rect 664444 416832 664496 416838
rect 664444 416774 664496 416780
rect 663248 313472 663300 313478
rect 663248 313414 663300 313420
rect 664260 311908 664312 311914
rect 664260 311850 664312 311856
rect 664272 266558 664300 311850
rect 664456 268190 664484 416774
rect 664628 364404 664680 364410
rect 664628 364346 664680 364352
rect 664444 268184 664496 268190
rect 664444 268126 664496 268132
rect 664260 266552 664312 266558
rect 664260 266494 664312 266500
rect 664444 266416 664496 266422
rect 664444 266358 664496 266364
rect 664260 264988 664312 264994
rect 664260 264930 664312 264936
rect 663064 222488 663116 222494
rect 663064 222430 663116 222436
rect 663798 221504 663854 221513
rect 663798 221439 663854 221448
rect 662892 219406 663012 219434
rect 662984 210202 663012 219406
rect 663812 210202 663840 221439
rect 664272 221134 664300 264930
rect 664456 222222 664484 266358
rect 664640 222358 664668 364346
rect 664824 357610 664852 484366
rect 664812 357604 664864 357610
rect 664812 357546 664864 357552
rect 664996 309188 665048 309194
rect 664996 309130 665048 309136
rect 664812 284368 664864 284374
rect 664812 284310 664864 284316
rect 664628 222352 664680 222358
rect 664628 222294 664680 222300
rect 664444 222216 664496 222222
rect 664444 222158 664496 222164
rect 664260 221128 664312 221134
rect 664260 221070 664312 221076
rect 664168 215348 664220 215354
rect 664168 215290 664220 215296
rect 664180 210202 664208 215290
rect 664824 211138 664852 284310
rect 665008 265130 665036 309130
rect 665192 273737 665220 993142
rect 665456 990276 665508 990282
rect 665456 990218 665508 990224
rect 665468 287054 665496 990218
rect 665640 984768 665692 984774
rect 665640 984710 665692 984716
rect 665652 287054 665680 984710
rect 666376 742484 666428 742490
rect 666376 742426 666428 742432
rect 666100 692912 666152 692918
rect 666100 692854 666152 692860
rect 665916 641776 665968 641782
rect 665916 641718 665968 641724
rect 665928 570042 665956 641718
rect 666112 619682 666140 692854
rect 666388 665242 666416 742426
rect 666376 665236 666428 665242
rect 666376 665178 666428 665184
rect 666284 641912 666336 641918
rect 666284 641854 666336 641860
rect 666100 619676 666152 619682
rect 666100 619618 666152 619624
rect 666100 596216 666152 596222
rect 666100 596158 666152 596164
rect 665916 570036 665968 570042
rect 665916 569978 665968 569984
rect 666112 528630 666140 596158
rect 666296 574258 666324 641854
rect 666284 574252 666336 574258
rect 666284 574194 666336 574200
rect 666376 557592 666428 557598
rect 666376 557534 666428 557540
rect 666100 528624 666152 528630
rect 666100 528566 666152 528572
rect 666388 485994 666416 557534
rect 666376 485988 666428 485994
rect 666376 485930 666428 485936
rect 666376 310752 666428 310758
rect 666376 310694 666428 310700
rect 665468 287026 665588 287054
rect 665652 287026 665772 287054
rect 665178 273728 665234 273737
rect 665178 273663 665234 273672
rect 665560 273465 665588 287026
rect 665744 273737 665772 287026
rect 665730 273728 665786 273737
rect 665730 273663 665786 273672
rect 665546 273456 665602 273465
rect 665546 273391 665602 273400
rect 666388 266694 666416 310694
rect 666376 266688 666428 266694
rect 666376 266630 666428 266636
rect 666008 265260 666060 265266
rect 666008 265202 666060 265208
rect 664996 265124 665048 265130
rect 664996 265066 665048 265072
rect 665088 263628 665140 263634
rect 665088 263570 665140 263576
rect 665100 219638 665128 263570
rect 666020 219774 666048 265202
rect 666376 259616 666428 259622
rect 666376 259558 666428 259564
rect 666192 259480 666244 259486
rect 666192 259422 666244 259428
rect 666204 242894 666232 259422
rect 666192 242888 666244 242894
rect 666192 242830 666244 242836
rect 666388 237386 666416 259558
rect 666376 237380 666428 237386
rect 666376 237322 666428 237328
rect 666008 219768 666060 219774
rect 666008 219710 666060 219716
rect 665088 219632 665140 219638
rect 665088 219574 665140 219580
rect 664812 211132 664864 211138
rect 664812 211074 664864 211080
rect 652772 210174 652924 210202
rect 653048 210174 653476 210202
rect 654152 210174 654580 210202
rect 654704 210174 655132 210202
rect 655808 210174 656236 210202
rect 656452 210174 656788 210202
rect 657464 210174 657892 210202
rect 658292 210174 658444 210202
rect 659120 210174 659548 210202
rect 659856 210174 660100 210202
rect 660316 210174 660652 210202
rect 661052 210174 661204 210202
rect 661512 210174 661756 210202
rect 661972 210174 662308 210202
rect 662432 210174 662860 210202
rect 662984 210174 663412 210202
rect 663812 210174 663964 210202
rect 664180 210174 664516 210202
rect 652208 209568 652260 209574
rect 652208 209510 652260 209516
rect 666572 184249 666600 994230
rect 666928 993336 666980 993342
rect 666928 993278 666980 993284
rect 666744 990412 666796 990418
rect 666744 990354 666796 990360
rect 666756 245721 666784 990354
rect 666742 245712 666798 245721
rect 666742 245647 666798 245656
rect 666742 245440 666798 245449
rect 666940 245426 666968 993278
rect 667124 972914 667152 994366
rect 668032 991772 668084 991778
rect 668032 991714 668084 991720
rect 666798 245398 666968 245426
rect 667032 972886 667152 972914
rect 666742 245375 666798 245384
rect 666742 223952 666798 223961
rect 666742 223887 666798 223896
rect 666558 184240 666614 184249
rect 666558 184175 666614 184184
rect 591304 147552 591356 147558
rect 591304 147494 591356 147500
rect 589922 144528 589978 144537
rect 589922 144463 589978 144472
rect 590384 144220 590436 144226
rect 590384 144162 590436 144168
rect 590016 143540 590068 143546
rect 590016 143482 590068 143488
rect 590028 142905 590056 143482
rect 590014 142896 590070 142905
rect 590014 142831 590070 142840
rect 589464 142044 589516 142050
rect 589464 141986 589516 141992
rect 589476 141273 589504 141986
rect 589462 141264 589518 141273
rect 589462 141199 589518 141208
rect 589464 140752 589516 140758
rect 589464 140694 589516 140700
rect 589476 139641 589504 140694
rect 589462 139632 589518 139641
rect 589462 139567 589518 139576
rect 589462 138000 589518 138009
rect 589462 137935 589464 137944
rect 589516 137935 589518 137944
rect 589464 137906 589516 137912
rect 589372 136536 589424 136542
rect 589372 136478 589424 136484
rect 589384 136377 589412 136478
rect 589370 136368 589426 136377
rect 589370 136303 589426 136312
rect 588726 134736 588782 134745
rect 588726 134671 588782 134680
rect 589924 133204 589976 133210
rect 589924 133146 589976 133152
rect 589464 132388 589516 132394
rect 589464 132330 589516 132336
rect 589476 131481 589504 132330
rect 589462 131472 589518 131481
rect 589462 131407 589518 131416
rect 588544 130416 588596 130422
rect 588544 130358 588596 130364
rect 587164 126948 587216 126954
rect 587164 126890 587216 126896
rect 587348 126268 587400 126274
rect 587348 126210 587400 126216
rect 585968 124908 586020 124914
rect 585968 124850 586020 124856
rect 585784 124228 585836 124234
rect 585784 124170 585836 124176
rect 585796 114510 585824 124170
rect 587164 118720 587216 118726
rect 587164 118662 587216 118668
rect 585784 114504 585836 114510
rect 585784 114446 585836 114452
rect 584404 111784 584456 111790
rect 584404 111726 584456 111732
rect 583024 107636 583076 107642
rect 583024 107578 583076 107584
rect 587176 106282 587204 118662
rect 587360 115938 587388 126210
rect 588556 118425 588584 130358
rect 589464 129736 589516 129742
rect 589462 129704 589464 129713
rect 589516 129704 589518 129713
rect 589462 129639 589518 129648
rect 589464 128240 589516 128246
rect 589462 128208 589464 128217
rect 589516 128208 589518 128217
rect 589462 128143 589518 128152
rect 589740 126948 589792 126954
rect 589740 126890 589792 126896
rect 589752 126585 589780 126890
rect 589738 126576 589794 126585
rect 589738 126511 589794 126520
rect 589936 124953 589964 133146
rect 590396 133113 590424 144162
rect 590382 133104 590438 133113
rect 590382 133039 590438 133048
rect 589922 124944 589978 124953
rect 589922 124879 589978 124888
rect 590384 124908 590436 124914
rect 590384 124850 590436 124856
rect 589464 124092 589516 124098
rect 589464 124034 589516 124040
rect 589476 123321 589504 124034
rect 589462 123312 589518 123321
rect 589462 123247 589518 123256
rect 590396 121689 590424 124850
rect 590382 121680 590438 121689
rect 590382 121615 590438 121624
rect 589924 120760 589976 120766
rect 589924 120702 589976 120708
rect 589464 120080 589516 120086
rect 589462 120048 589464 120057
rect 589516 120048 589518 120057
rect 589462 119983 589518 119992
rect 588542 118416 588598 118425
rect 588542 118351 588598 118360
rect 589464 117224 589516 117230
rect 589464 117166 589516 117172
rect 589476 116793 589504 117166
rect 589462 116784 589518 116793
rect 589462 116719 589518 116728
rect 587348 115932 587400 115938
rect 587348 115874 587400 115880
rect 589280 115932 589332 115938
rect 589280 115874 589332 115880
rect 589292 115161 589320 115874
rect 589278 115152 589334 115161
rect 589278 115087 589334 115096
rect 589464 114504 589516 114510
rect 589464 114446 589516 114452
rect 589476 113529 589504 114446
rect 589462 113520 589518 113529
rect 589462 113455 589518 113464
rect 589464 111784 589516 111790
rect 589462 111752 589464 111761
rect 589516 111752 589518 111761
rect 589462 111687 589518 111696
rect 589936 110265 589964 120702
rect 589922 110256 589978 110265
rect 589922 110191 589978 110200
rect 666756 109381 666784 223887
rect 667032 187649 667060 972886
rect 667664 732828 667716 732834
rect 667664 732770 667716 732776
rect 667676 665378 667704 732770
rect 667846 684992 667902 685001
rect 667846 684927 667902 684936
rect 667664 665372 667716 665378
rect 667664 665314 667716 665320
rect 667860 615913 667888 684927
rect 667846 615904 667902 615913
rect 667846 615839 667902 615848
rect 667848 603152 667900 603158
rect 667848 603094 667900 603100
rect 667860 530126 667888 603094
rect 667848 530120 667900 530126
rect 667848 530062 667900 530068
rect 667848 353660 667900 353666
rect 667848 353602 667900 353608
rect 667388 338156 667440 338162
rect 667388 338098 667440 338104
rect 667204 310548 667256 310554
rect 667204 310490 667256 310496
rect 667018 187640 667074 187649
rect 667018 187575 667074 187584
rect 667216 132938 667244 310490
rect 667400 178294 667428 338098
rect 667860 325514 667888 353602
rect 667848 325508 667900 325514
rect 667848 325450 667900 325456
rect 668044 245721 668072 991714
rect 672724 990548 672776 990554
rect 672724 990490 672776 990496
rect 668216 988916 668268 988922
rect 668216 988858 668268 988864
rect 668030 245712 668086 245721
rect 668030 245647 668086 245656
rect 667848 220856 667900 220862
rect 667848 220798 667900 220804
rect 667572 211132 667624 211138
rect 667572 211074 667624 211080
rect 667388 178288 667440 178294
rect 667388 178230 667440 178236
rect 667204 132932 667256 132938
rect 667204 132874 667256 132880
rect 667584 132802 667612 211074
rect 667860 175438 667888 220798
rect 668228 197441 668256 988858
rect 669964 987692 670016 987698
rect 669964 987634 670016 987640
rect 668400 987556 668452 987562
rect 668400 987498 668452 987504
rect 668412 245857 668440 987498
rect 669976 935950 670004 987634
rect 671344 948116 671396 948122
rect 671344 948058 671396 948064
rect 671356 938602 671384 948058
rect 672736 938738 672764 990490
rect 675404 966521 675432 966723
rect 675390 966512 675446 966521
rect 675390 966447 675446 966456
rect 673368 966204 673420 966210
rect 673368 966146 673420 966152
rect 675116 966204 675168 966210
rect 675116 966146 675168 966152
rect 672998 959168 673054 959177
rect 672998 959103 673054 959112
rect 672724 938732 672776 938738
rect 672724 938674 672776 938680
rect 671344 938596 671396 938602
rect 671344 938538 671396 938544
rect 671528 937576 671580 937582
rect 671528 937518 671580 937524
rect 671160 937100 671212 937106
rect 671160 937042 671212 937048
rect 669964 935944 670016 935950
rect 669964 935886 670016 935892
rect 669780 928804 669832 928810
rect 669780 928746 669832 928752
rect 669596 879096 669648 879102
rect 669596 879038 669648 879044
rect 669228 866720 669280 866726
rect 669228 866662 669280 866668
rect 668768 782536 668820 782542
rect 668768 782478 668820 782484
rect 668582 773800 668638 773809
rect 668582 773735 668638 773744
rect 668596 709782 668624 773735
rect 668584 709776 668636 709782
rect 668584 709718 668636 709724
rect 668780 709374 668808 782478
rect 669240 753001 669268 866662
rect 669608 754662 669636 879038
rect 669596 754656 669648 754662
rect 669596 754598 669648 754604
rect 669226 752992 669282 753001
rect 669226 752927 669282 752936
rect 669596 750100 669648 750106
rect 669596 750042 669648 750048
rect 669228 743708 669280 743714
rect 669228 743650 669280 743656
rect 669042 730144 669098 730153
rect 669042 730079 669098 730088
rect 668768 709368 668820 709374
rect 668768 709310 668820 709316
rect 668768 699712 668820 699718
rect 668768 699654 668820 699660
rect 668780 618322 668808 699654
rect 669056 663513 669084 730079
rect 669240 663814 669268 743650
rect 669412 685908 669464 685914
rect 669412 685850 669464 685856
rect 669228 663808 669280 663814
rect 669228 663750 669280 663756
rect 669042 663504 669098 663513
rect 669042 663439 669098 663448
rect 668952 649120 669004 649126
rect 668952 649062 669004 649068
rect 668768 618316 668820 618322
rect 668768 618258 668820 618264
rect 668584 616820 668636 616826
rect 668584 616762 668636 616768
rect 668398 245848 668454 245857
rect 668398 245783 668454 245792
rect 668400 222760 668452 222766
rect 668400 222702 668452 222708
rect 668412 222494 668440 222702
rect 668400 222488 668452 222494
rect 668400 222430 668452 222436
rect 668398 222320 668454 222329
rect 668398 222255 668454 222264
rect 668214 197432 668270 197441
rect 668032 197396 668084 197402
rect 668214 197367 668270 197376
rect 668032 197338 668084 197344
rect 667848 175432 667900 175438
rect 667848 175374 667900 175380
rect 668044 163169 668072 197338
rect 668216 184884 668268 184890
rect 668216 184826 668268 184832
rect 668030 163160 668086 163169
rect 668030 163095 668086 163104
rect 668032 138032 668084 138038
rect 668032 137974 668084 137980
rect 667572 132796 667624 132802
rect 667572 132738 667624 132744
rect 668044 124001 668072 137974
rect 668228 135425 668256 184826
rect 668214 135416 668270 135425
rect 668214 135351 668270 135360
rect 668412 131238 668440 222255
rect 668596 182753 668624 616762
rect 668768 595264 668820 595270
rect 668768 595206 668820 595212
rect 668780 589286 668808 595206
rect 668768 589280 668820 589286
rect 668964 589274 668992 649062
rect 669228 647760 669280 647766
rect 669228 647702 669280 647708
rect 668964 589246 669176 589274
rect 668768 589222 668820 589228
rect 669148 579986 669176 589246
rect 669056 579958 669176 579986
rect 669056 579816 669084 579958
rect 668964 579788 669084 579816
rect 668964 576854 668992 579788
rect 668872 576826 668992 576854
rect 668872 572762 668900 576826
rect 668860 572756 668912 572762
rect 668860 572698 668912 572704
rect 669240 572121 669268 647702
rect 669424 619886 669452 685850
rect 669412 619880 669464 619886
rect 669412 619822 669464 619828
rect 669412 589280 669464 589286
rect 669412 589222 669464 589228
rect 669226 572112 669282 572121
rect 669226 572047 669282 572056
rect 669424 569954 669452 589222
rect 669056 569926 669452 569954
rect 668766 563952 668822 563961
rect 668766 563887 668822 563896
rect 668582 182744 668638 182753
rect 668582 182679 668638 182688
rect 668584 178016 668636 178022
rect 668584 177958 668636 177964
rect 668596 177857 668624 177958
rect 668582 177848 668638 177857
rect 668582 177783 668638 177792
rect 668780 158273 668808 563887
rect 669056 529990 669084 569926
rect 669044 529984 669096 529990
rect 669044 529926 669096 529932
rect 669320 403436 669372 403442
rect 669320 403378 669372 403384
rect 669332 402966 669360 403378
rect 669320 402960 669372 402966
rect 669320 402902 669372 402908
rect 668952 268048 669004 268054
rect 668952 267990 669004 267996
rect 668964 267782 668992 267990
rect 668952 267776 669004 267782
rect 668952 267718 669004 267724
rect 669320 265600 669372 265606
rect 669320 265542 669372 265548
rect 669332 264926 669360 265542
rect 669320 264920 669372 264926
rect 669320 264862 669372 264868
rect 669228 259752 669280 259758
rect 669228 259694 669280 259700
rect 669240 241738 669268 259694
rect 669412 245200 669464 245206
rect 669412 245142 669464 245148
rect 669424 242894 669452 245142
rect 669412 242888 669464 242894
rect 669412 242830 669464 242836
rect 669228 241732 669280 241738
rect 669228 241674 669280 241680
rect 668950 223680 669006 223689
rect 668950 223615 669006 223624
rect 668766 158264 668822 158273
rect 668766 158199 668822 158208
rect 668766 148472 668822 148481
rect 668766 148407 668822 148416
rect 668780 148238 668808 148407
rect 668768 148232 668820 148238
rect 668768 148174 668820 148180
rect 668768 146260 668820 146266
rect 668768 146202 668820 146208
rect 668780 145217 668808 146202
rect 668766 145208 668822 145217
rect 668766 145143 668822 145152
rect 668768 144220 668820 144226
rect 668768 144162 668820 144168
rect 668780 143585 668808 144162
rect 668766 143576 668822 143585
rect 668766 143511 668822 143520
rect 668768 140752 668820 140758
rect 668768 140694 668820 140700
rect 668780 140321 668808 140694
rect 668766 140312 668822 140321
rect 668766 140247 668822 140256
rect 668768 139392 668820 139398
rect 668768 139334 668820 139340
rect 668780 138689 668808 139334
rect 668766 138680 668822 138689
rect 668766 138615 668822 138624
rect 668584 137352 668636 137358
rect 668584 137294 668636 137300
rect 668400 131232 668452 131238
rect 668400 131174 668452 131180
rect 668308 131096 668360 131102
rect 668308 131038 668360 131044
rect 668320 130529 668348 131038
rect 668306 130520 668362 130529
rect 668306 130455 668362 130464
rect 668596 129946 668624 137294
rect 668768 131232 668820 131238
rect 668768 131174 668820 131180
rect 668584 129940 668636 129946
rect 668584 129882 668636 129888
rect 668216 129260 668268 129266
rect 668216 129202 668268 129208
rect 668228 125633 668256 129202
rect 668214 125624 668270 125633
rect 668214 125559 668270 125568
rect 668030 123992 668086 124001
rect 668030 123927 668086 123936
rect 668308 112872 668360 112878
rect 668308 112814 668360 112820
rect 668320 112577 668348 112814
rect 668306 112568 668362 112577
rect 668306 112503 668362 112512
rect 666742 109372 666798 109381
rect 666742 109307 666798 109316
rect 589464 108996 589516 109002
rect 589464 108938 589516 108944
rect 589476 108633 589504 108938
rect 589462 108624 589518 108633
rect 589462 108559 589518 108568
rect 589372 107636 589424 107642
rect 589372 107578 589424 107584
rect 589384 107001 589412 107578
rect 589370 106992 589426 107001
rect 589370 106927 589426 106936
rect 587164 106276 587216 106282
rect 587164 106218 587216 106224
rect 589280 106276 589332 106282
rect 589280 106218 589332 106224
rect 589292 105369 589320 106218
rect 589278 105360 589334 105369
rect 589278 105295 589334 105304
rect 581644 104848 581696 104854
rect 581644 104790 581696 104796
rect 589372 104848 589424 104854
rect 589372 104790 589424 104796
rect 589384 103737 589412 104790
rect 589370 103728 589426 103737
rect 589370 103663 589426 103672
rect 668596 102785 668624 129882
rect 668780 106049 668808 131174
rect 668964 128382 668992 223615
rect 669134 221776 669190 221785
rect 669134 221711 669190 221720
rect 669148 137358 669176 221711
rect 669318 209944 669374 209953
rect 669318 209879 669374 209888
rect 669332 209794 669360 209879
rect 669240 209766 669360 209794
rect 669240 190346 669268 209766
rect 669412 209092 669464 209098
rect 669412 209034 669464 209040
rect 669240 190330 669314 190346
rect 669240 190324 669326 190330
rect 669240 190318 669274 190324
rect 669274 190266 669326 190272
rect 669136 137352 669188 137358
rect 669136 137294 669188 137300
rect 669228 133816 669280 133822
rect 669226 133784 669228 133793
rect 669280 133784 669282 133793
rect 669226 133719 669282 133728
rect 669424 133414 669452 209034
rect 669608 208321 669636 750042
rect 669792 616826 669820 928746
rect 670608 927444 670660 927450
rect 670608 927386 670660 927392
rect 670422 872264 670478 872273
rect 670422 872199 670478 872208
rect 670240 789404 670292 789410
rect 670240 789346 670292 789352
rect 670054 775024 670110 775033
rect 670054 774959 670110 774968
rect 670068 710705 670096 774959
rect 670054 710696 670110 710705
rect 670054 710631 670110 710640
rect 670252 709646 670280 789346
rect 670436 752729 670464 872199
rect 670422 752720 670478 752729
rect 670422 752655 670478 752664
rect 670424 728680 670476 728686
rect 670424 728622 670476 728628
rect 670240 709640 670292 709646
rect 670240 709582 670292 709588
rect 669964 705084 670016 705090
rect 669964 705026 670016 705032
rect 669780 616820 669832 616826
rect 669780 616762 669832 616768
rect 669780 349308 669832 349314
rect 669780 349250 669832 349256
rect 669792 332654 669820 349250
rect 669780 332648 669832 332654
rect 669780 332590 669832 332596
rect 669780 256624 669832 256630
rect 669780 256566 669832 256572
rect 669594 208312 669650 208321
rect 669594 208247 669650 208256
rect 669596 208140 669648 208146
rect 669596 208082 669648 208088
rect 669608 205634 669636 208082
rect 669608 205606 669728 205634
rect 669700 135254 669728 205606
rect 669608 135226 669728 135254
rect 669412 133408 669464 133414
rect 669412 133350 669464 133356
rect 669228 129668 669280 129674
rect 669228 129610 669280 129616
rect 669240 128897 669268 129610
rect 669608 129146 669636 135226
rect 669792 129266 669820 256566
rect 669976 169697 670004 705026
rect 670436 664902 670464 728622
rect 670424 664896 670476 664902
rect 670424 664838 670476 664844
rect 670240 644496 670292 644502
rect 670240 644438 670292 644444
rect 670252 611354 670280 644438
rect 670424 641776 670476 641782
rect 670424 641718 670476 641724
rect 670436 641306 670464 641718
rect 670424 641300 670476 641306
rect 670424 641242 670476 641248
rect 670424 616140 670476 616146
rect 670424 616082 670476 616088
rect 670436 611354 670464 616082
rect 670160 611326 670280 611354
rect 670344 611326 670464 611354
rect 670160 607209 670188 611326
rect 670146 607200 670202 607209
rect 670344 607170 670372 611326
rect 670146 607135 670202 607144
rect 670332 607164 670384 607170
rect 670332 607106 670384 607112
rect 670330 606928 670386 606937
rect 670148 606892 670200 606898
rect 670330 606863 670386 606872
rect 670148 606834 670200 606840
rect 670160 606778 670188 606834
rect 670344 606778 670372 606863
rect 670068 606750 670188 606778
rect 670252 606750 670372 606778
rect 670068 205634 670096 606750
rect 670252 572898 670280 606750
rect 670424 601724 670476 601730
rect 670424 601666 670476 601672
rect 670240 572892 670292 572898
rect 670240 572834 670292 572840
rect 670238 548448 670294 548457
rect 670238 548383 670294 548392
rect 670252 485654 670280 548383
rect 670436 526862 670464 601666
rect 670424 526856 670476 526862
rect 670424 526798 670476 526804
rect 670240 485648 670292 485654
rect 670240 485590 670292 485596
rect 670424 396092 670476 396098
rect 670424 396034 670476 396040
rect 670436 379506 670464 396034
rect 670424 379500 670476 379506
rect 670424 379442 670476 379448
rect 670424 352572 670476 352578
rect 670424 352514 670476 352520
rect 670238 342272 670294 342281
rect 670238 342207 670294 342216
rect 670252 325650 670280 342207
rect 670436 333946 670464 352514
rect 670424 333940 670476 333946
rect 670424 333882 670476 333888
rect 670240 325644 670292 325650
rect 670240 325586 670292 325592
rect 670424 310412 670476 310418
rect 670424 310354 670476 310360
rect 670240 302252 670292 302258
rect 670240 302194 670292 302200
rect 670252 205634 670280 302194
rect 670436 265878 670464 310354
rect 670424 265872 670476 265878
rect 670424 265814 670476 265820
rect 670424 259276 670476 259282
rect 670424 259218 670476 259224
rect 670436 242894 670464 259218
rect 670424 242888 670476 242894
rect 670424 242830 670476 242836
rect 670424 216708 670476 216714
rect 670424 216650 670476 216656
rect 670436 215294 670464 216650
rect 670436 215266 670556 215294
rect 670528 205634 670556 215266
rect 670620 212786 670648 927386
rect 670976 866856 671028 866862
rect 670976 866798 671028 866804
rect 670792 788044 670844 788050
rect 670792 787986 670844 787992
rect 670804 785234 670832 787986
rect 670804 785206 670924 785234
rect 670896 756254 670924 785206
rect 670804 756226 670924 756254
rect 670804 746594 670832 756226
rect 670988 753438 671016 866798
rect 671172 759558 671200 937042
rect 671344 881884 671396 881890
rect 671344 881826 671396 881832
rect 671356 869038 671384 881826
rect 671344 869032 671396 869038
rect 671344 868974 671396 868980
rect 671344 855636 671396 855642
rect 671344 855578 671396 855584
rect 671160 759552 671212 759558
rect 671160 759494 671212 759500
rect 671160 759076 671212 759082
rect 671160 759018 671212 759024
rect 670976 753432 671028 753438
rect 670976 753374 671028 753380
rect 670804 746566 671016 746594
rect 670792 735004 670844 735010
rect 670792 734946 670844 734952
rect 670804 662046 670832 734946
rect 670988 711278 671016 746566
rect 671172 714542 671200 759018
rect 671356 716582 671384 855578
rect 671540 760306 671568 937518
rect 672080 935808 672132 935814
rect 672080 935750 672132 935756
rect 671802 868048 671858 868057
rect 671802 867983 671858 867992
rect 671528 760300 671580 760306
rect 671528 760242 671580 760248
rect 671528 759892 671580 759898
rect 671528 759834 671580 759840
rect 671344 716576 671396 716582
rect 671344 716518 671396 716524
rect 671540 715358 671568 759834
rect 671816 751806 671844 867983
rect 672092 758742 672120 935750
rect 672448 935672 672500 935678
rect 672448 935614 672500 935620
rect 672264 782672 672316 782678
rect 672264 782614 672316 782620
rect 672080 758736 672132 758742
rect 672080 758678 672132 758684
rect 672080 757444 672132 757450
rect 672080 757386 672132 757392
rect 671804 751800 671856 751806
rect 671804 751742 671856 751748
rect 671896 742824 671948 742830
rect 671896 742766 671948 742772
rect 671710 733680 671766 733689
rect 671710 733615 671766 733624
rect 671528 715352 671580 715358
rect 671528 715294 671580 715300
rect 671528 714876 671580 714882
rect 671528 714818 671580 714824
rect 671160 714536 671212 714542
rect 671160 714478 671212 714484
rect 671160 713244 671212 713250
rect 671160 713186 671212 713192
rect 670976 711272 671028 711278
rect 670976 711214 671028 711220
rect 671172 698294 671200 713186
rect 671344 712428 671396 712434
rect 671344 712370 671396 712376
rect 671356 707954 671384 712370
rect 671356 707926 671476 707954
rect 671080 698266 671200 698294
rect 671080 668574 671108 698266
rect 671252 687472 671304 687478
rect 671252 687414 671304 687420
rect 671068 668568 671120 668574
rect 671068 668510 671120 668516
rect 671068 668432 671120 668438
rect 671068 668374 671120 668380
rect 670792 662040 670844 662046
rect 670792 661982 670844 661988
rect 670792 661156 670844 661162
rect 670792 661098 670844 661104
rect 670804 229094 670832 661098
rect 671080 660090 671108 668374
rect 671080 660062 671200 660090
rect 670976 660000 671028 660006
rect 670976 659942 671028 659948
rect 670988 229094 671016 659942
rect 671172 624374 671200 660062
rect 671264 649994 671292 687414
rect 671448 678974 671476 707926
rect 671356 678946 671476 678974
rect 671356 669474 671384 678946
rect 671540 669662 671568 714818
rect 671724 673454 671752 733615
rect 671724 673426 671844 673454
rect 671528 669656 671580 669662
rect 671528 669598 671580 669604
rect 671620 669520 671672 669526
rect 671356 669446 671476 669474
rect 671620 669462 671672 669468
rect 671448 667758 671476 669446
rect 671436 667752 671488 667758
rect 671436 667694 671488 667700
rect 671632 659654 671660 669462
rect 671816 661638 671844 673426
rect 671908 669314 671936 742766
rect 672092 712910 672120 757386
rect 672276 753494 672304 782614
rect 672460 757926 672488 935614
rect 673012 933366 673040 959103
rect 673184 956412 673236 956418
rect 673184 956354 673236 956360
rect 673000 933360 673052 933366
rect 673000 933302 673052 933308
rect 673196 930170 673224 956354
rect 673380 933026 673408 966146
rect 675128 966090 675156 966146
rect 675128 966062 675418 966090
rect 675772 965161 675800 965435
rect 675758 965152 675814 965161
rect 675758 965087 675814 965096
rect 675220 963581 675418 963609
rect 675220 963393 675248 963581
rect 675206 963384 675262 963393
rect 675206 963319 675262 963328
rect 675312 963070 675432 963098
rect 675312 963030 675340 963070
rect 674668 963002 675340 963030
rect 675404 963016 675432 963070
rect 674288 961920 674340 961926
rect 674288 961862 674340 961868
rect 674102 952232 674158 952241
rect 674102 952167 674158 952176
rect 674116 933473 674144 952167
rect 674102 933464 674158 933473
rect 674102 933399 674158 933408
rect 673368 933020 673420 933026
rect 673368 932962 673420 932968
rect 674300 932249 674328 961862
rect 674472 957908 674524 957914
rect 674472 957850 674524 957856
rect 674286 932240 674342 932249
rect 674286 932175 674342 932184
rect 674484 931433 674512 957850
rect 674668 932657 674696 963002
rect 675128 962390 675418 962418
rect 675128 961926 675156 962390
rect 675758 962024 675814 962033
rect 675758 961959 675814 961968
rect 675116 961920 675168 961926
rect 675116 961862 675168 961868
rect 675772 961755 675800 961959
rect 674930 959440 674986 959449
rect 674930 959375 674986 959384
rect 674944 951538 674972 959375
rect 675128 959262 675418 959290
rect 675128 959177 675156 959262
rect 675114 959168 675170 959177
rect 675114 959103 675170 959112
rect 675772 958361 675800 958732
rect 675758 958352 675814 958361
rect 675758 958287 675814 958296
rect 675312 958174 675432 958202
rect 675312 958066 675340 958174
rect 675128 958038 675340 958066
rect 675404 958052 675432 958174
rect 675128 957914 675156 958038
rect 675116 957908 675168 957914
rect 675116 957850 675168 957856
rect 675128 957426 675418 957454
rect 675128 956418 675156 957426
rect 675300 957364 675352 957370
rect 675300 957306 675352 957312
rect 675116 956412 675168 956418
rect 675116 956354 675168 956360
rect 675312 955482 675340 957306
rect 675758 956448 675814 956457
rect 675758 956383 675814 956392
rect 675772 956216 675800 956383
rect 675312 955454 675524 955482
rect 675496 955060 675524 955454
rect 675220 954366 675418 954394
rect 674944 951510 675156 951538
rect 674930 948968 674986 948977
rect 674930 948903 674986 948912
rect 674944 941905 674972 948903
rect 675128 946694 675156 951510
rect 675220 948784 675248 954366
rect 675404 953442 675432 953768
rect 675312 953414 675432 953442
rect 675312 949454 675340 953414
rect 675496 952241 675524 952544
rect 675482 952232 675538 952241
rect 675482 952167 675538 952176
rect 677506 951552 677562 951561
rect 677506 951487 677562 951496
rect 675852 949476 675904 949482
rect 675312 949426 675852 949454
rect 675852 949418 675904 949424
rect 675852 948796 675904 948802
rect 675220 948756 675852 948784
rect 675852 948738 675904 948744
rect 675128 946666 675248 946694
rect 674930 941896 674986 941905
rect 675220 941848 675248 946666
rect 675850 941896 675906 941905
rect 674930 941831 674986 941840
rect 675128 941820 675248 941848
rect 675484 941860 675536 941866
rect 674930 939584 674986 939593
rect 674930 939519 674986 939528
rect 674944 938466 674972 939519
rect 674932 938460 674984 938466
rect 674932 938402 674984 938408
rect 674930 937952 674986 937961
rect 674930 937887 674986 937896
rect 674944 937242 674972 937887
rect 674932 937236 674984 937242
rect 674932 937178 674984 937184
rect 675128 934153 675156 941820
rect 675850 941831 675906 941840
rect 675484 941802 675536 941808
rect 675496 940001 675524 941802
rect 675482 939992 675538 940001
rect 675482 939927 675538 939936
rect 675298 939176 675354 939185
rect 675298 939111 675354 939120
rect 675312 938602 675340 939111
rect 675482 938768 675538 938777
rect 675482 938703 675484 938712
rect 675536 938703 675538 938712
rect 675484 938674 675536 938680
rect 675300 938596 675352 938602
rect 675300 938538 675352 938544
rect 675482 938360 675538 938369
rect 675482 938295 675538 938304
rect 675496 937582 675524 938295
rect 675484 937576 675536 937582
rect 675298 937544 675354 937553
rect 675484 937518 675536 937524
rect 675298 937479 675354 937488
rect 675312 937106 675340 937479
rect 675484 937372 675536 937378
rect 675484 937314 675536 937320
rect 675496 937145 675524 937314
rect 675482 937136 675538 937145
rect 675300 937100 675352 937106
rect 675482 937071 675538 937080
rect 675300 937042 675352 937048
rect 675666 936728 675722 936737
rect 675666 936663 675722 936672
rect 675482 936320 675538 936329
rect 675482 936255 675538 936264
rect 675496 935950 675524 936255
rect 675484 935944 675536 935950
rect 675298 935912 675354 935921
rect 675484 935886 675536 935892
rect 675298 935847 675354 935856
rect 675312 935678 675340 935847
rect 675484 935808 675536 935814
rect 675680 935762 675708 936663
rect 675536 935756 675708 935762
rect 675484 935750 675708 935756
rect 675496 935734 675708 935750
rect 675300 935672 675352 935678
rect 675300 935614 675352 935620
rect 675864 934697 675892 941831
rect 675850 934688 675906 934697
rect 675850 934623 675906 934632
rect 675114 934144 675170 934153
rect 675114 934079 675170 934088
rect 675482 933872 675538 933881
rect 675482 933807 675538 933816
rect 675496 933366 675524 933807
rect 675484 933360 675536 933366
rect 675484 933302 675536 933308
rect 675482 933056 675538 933065
rect 675482 932991 675484 933000
rect 675536 932991 675538 933000
rect 675484 932962 675536 932968
rect 674654 932648 674710 932657
rect 674654 932583 674710 932592
rect 674470 931424 674526 931433
rect 674470 931359 674526 931368
rect 677520 931161 677548 951487
rect 683302 950056 683358 950065
rect 683302 949991 683358 950000
rect 678244 949476 678296 949482
rect 678244 949418 678296 949424
rect 677506 931152 677562 931161
rect 677506 931087 677562 931096
rect 675482 930200 675538 930209
rect 673184 930164 673236 930170
rect 675482 930135 675484 930144
rect 673184 930106 673236 930112
rect 675536 930135 675538 930144
rect 675484 930106 675536 930112
rect 678256 930102 678284 949418
rect 682384 948796 682436 948802
rect 682384 948738 682436 948744
rect 682396 935241 682424 948738
rect 683316 935649 683344 949991
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 683302 935640 683358 935649
rect 683302 935575 683358 935584
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 678244 930096 678296 930102
rect 678244 930038 678296 930044
rect 683120 930096 683172 930102
rect 683120 930038 683172 930044
rect 675482 929792 675538 929801
rect 675482 929727 675538 929736
rect 675496 928810 675524 929727
rect 683132 929529 683160 930038
rect 683118 929520 683174 929529
rect 683118 929455 683174 929464
rect 675484 928804 675536 928810
rect 675484 928746 675536 928752
rect 675482 928568 675538 928577
rect 675482 928503 675538 928512
rect 675496 927450 675524 928503
rect 675484 927444 675536 927450
rect 675484 927386 675536 927392
rect 675300 879096 675352 879102
rect 675300 879038 675352 879044
rect 675312 877146 675340 879038
rect 675772 877169 675800 877540
rect 675758 877160 675814 877169
rect 675312 877118 675432 877146
rect 675404 876860 675432 877118
rect 675758 877095 675814 877104
rect 675298 876480 675354 876489
rect 675298 876415 675354 876424
rect 675312 876262 675340 876415
rect 675312 876234 675418 876262
rect 675404 874041 675432 874412
rect 675390 874032 675446 874041
rect 675390 873967 675446 873976
rect 675404 873633 675432 873868
rect 672630 873624 672686 873633
rect 672630 873559 672686 873568
rect 675390 873624 675446 873633
rect 675390 873559 675446 873568
rect 672448 757920 672500 757926
rect 672448 757862 672500 757868
rect 672644 754254 672672 873559
rect 674024 873174 675418 873202
rect 673000 869440 673052 869446
rect 673000 869382 673052 869388
rect 672816 778388 672868 778394
rect 672816 778330 672868 778336
rect 672632 754248 672684 754254
rect 672632 754190 672684 754196
rect 672276 753466 672580 753494
rect 672354 751360 672410 751369
rect 672354 751295 672410 751304
rect 672368 746450 672396 751295
rect 672184 746422 672396 746450
rect 672184 727274 672212 746422
rect 672552 746178 672580 753466
rect 672276 746150 672580 746178
rect 672276 736934 672304 746150
rect 672276 736906 672396 736934
rect 672184 727246 672304 727274
rect 672080 712904 672132 712910
rect 672080 712846 672132 712852
rect 672276 712722 672304 727246
rect 672184 712694 672304 712722
rect 671908 669286 672028 669314
rect 672000 666126 672028 669286
rect 671988 666120 672040 666126
rect 671988 666062 672040 666068
rect 671804 661632 671856 661638
rect 671804 661574 671856 661580
rect 671540 659626 671660 659654
rect 671264 649966 671384 649994
rect 671160 624368 671212 624374
rect 671160 624310 671212 624316
rect 671356 618186 671384 649966
rect 671540 624986 671568 659626
rect 671896 651432 671948 651438
rect 671896 651374 671948 651380
rect 671710 643512 671766 643521
rect 671710 643447 671766 643456
rect 671528 624980 671580 624986
rect 671528 624922 671580 624928
rect 671528 623076 671580 623082
rect 671528 623018 671580 623024
rect 671344 618180 671396 618186
rect 671344 618122 671396 618128
rect 671344 577312 671396 577318
rect 671344 577254 671396 577260
rect 671160 576904 671212 576910
rect 671160 576846 671212 576852
rect 671356 576854 671384 577254
rect 671540 577046 671568 623018
rect 671528 577040 671580 577046
rect 671528 576982 671580 576988
rect 671172 532574 671200 576846
rect 671356 576826 671568 576854
rect 671344 569628 671396 569634
rect 671344 569570 671396 569576
rect 671160 532568 671212 532574
rect 671160 532510 671212 532516
rect 671160 397316 671212 397322
rect 671160 397258 671212 397264
rect 671172 377777 671200 397258
rect 671158 377768 671214 377777
rect 671158 377703 671214 377712
rect 671160 348492 671212 348498
rect 671160 348434 671212 348440
rect 670804 229066 670924 229094
rect 670988 229066 671108 229094
rect 670620 212758 670740 212786
rect 670712 212514 670740 212758
rect 670620 212486 670740 212514
rect 670620 209658 670648 212486
rect 670896 210497 670924 229066
rect 671080 212673 671108 229066
rect 671172 215294 671200 348434
rect 671172 215266 671292 215294
rect 671066 212664 671122 212673
rect 671066 212599 671122 212608
rect 670882 210488 670938 210497
rect 670882 210423 670938 210432
rect 670976 210316 671028 210322
rect 670976 210258 671028 210264
rect 670790 209672 670846 209681
rect 670620 209630 670790 209658
rect 670790 209607 670846 209616
rect 670068 205606 670188 205634
rect 670252 205606 670372 205634
rect 670528 205606 670648 205634
rect 670160 197402 670188 205606
rect 670148 197396 670200 197402
rect 670148 197338 670200 197344
rect 670344 195974 670372 205606
rect 670252 195946 670372 195974
rect 669962 169688 670018 169697
rect 669962 169623 670018 169632
rect 669964 166864 670016 166870
rect 669964 166806 670016 166812
rect 669780 129260 669832 129266
rect 669780 129202 669832 129208
rect 669608 129118 669728 129146
rect 669226 128888 669282 128897
rect 669226 128823 669282 128832
rect 668952 128376 669004 128382
rect 668952 128318 669004 128324
rect 668964 113174 668992 128318
rect 669700 120737 669728 129118
rect 669686 120728 669742 120737
rect 669686 120663 669742 120672
rect 669228 120080 669280 120086
rect 669228 120022 669280 120028
rect 669240 119105 669268 120022
rect 669226 119096 669282 119105
rect 669226 119031 669282 119040
rect 669976 117473 670004 166806
rect 670252 131102 670280 195946
rect 670620 193633 670648 205606
rect 670606 193624 670662 193633
rect 670606 193559 670662 193568
rect 670988 178158 671016 210258
rect 671264 195974 671292 215266
rect 671172 195946 671292 195974
rect 670976 178152 671028 178158
rect 670976 178094 671028 178100
rect 670424 171148 670476 171154
rect 670424 171090 670476 171096
rect 670436 154970 670464 171090
rect 670608 169108 670660 169114
rect 670608 169050 670660 169056
rect 670424 154964 670476 154970
rect 670424 154906 670476 154912
rect 670620 150414 670648 169050
rect 671172 162602 671200 195946
rect 671356 166994 671384 569570
rect 671540 533390 671568 576826
rect 671724 571266 671752 643447
rect 671908 621014 671936 651374
rect 672184 625161 672212 712694
rect 672368 707606 672396 736906
rect 672538 734224 672594 734233
rect 672538 734159 672594 734168
rect 672356 707600 672408 707606
rect 672356 707542 672408 707548
rect 672356 668092 672408 668098
rect 672356 668034 672408 668040
rect 672170 625152 672226 625161
rect 672170 625087 672226 625096
rect 672368 623558 672396 668034
rect 672552 662862 672580 734159
rect 672828 706790 672856 778330
rect 673012 752214 673040 869382
rect 673368 862912 673420 862918
rect 673368 862854 673420 862860
rect 673184 758260 673236 758266
rect 673184 758202 673236 758208
rect 673000 752208 673052 752214
rect 673000 752150 673052 752156
rect 673000 714060 673052 714066
rect 673000 714002 673052 714008
rect 672816 706784 672868 706790
rect 672816 706726 672868 706732
rect 672816 690056 672868 690062
rect 672816 689998 672868 690004
rect 672828 688786 672856 689998
rect 672828 688758 672948 688786
rect 672722 688664 672778 688673
rect 672722 688599 672778 688608
rect 672540 662856 672592 662862
rect 672540 662798 672592 662804
rect 672538 645416 672594 645425
rect 672538 645351 672594 645360
rect 672356 623552 672408 623558
rect 672356 623494 672408 623500
rect 672080 622260 672132 622266
rect 672080 622202 672132 622208
rect 672092 622146 672120 622202
rect 671816 620986 671936 621014
rect 672000 622118 672120 622146
rect 671816 576854 671844 620986
rect 672000 577182 672028 622118
rect 672172 614916 672224 614922
rect 672172 614858 672224 614864
rect 671988 577176 672040 577182
rect 671988 577118 672040 577124
rect 671816 576826 671936 576854
rect 671908 575550 671936 576826
rect 671896 575544 671948 575550
rect 671896 575486 671948 575492
rect 671712 571260 671764 571266
rect 671712 571202 671764 571208
rect 671804 554804 671856 554810
rect 671804 554746 671856 554752
rect 671528 533384 671580 533390
rect 671528 533326 671580 533332
rect 671816 482798 671844 554746
rect 671986 553480 672042 553489
rect 671986 553415 672042 553424
rect 671804 482792 671856 482798
rect 671804 482734 671856 482740
rect 672000 482390 672028 553415
rect 671988 482384 672040 482390
rect 671988 482326 672040 482332
rect 671528 480684 671580 480690
rect 671528 480626 671580 480632
rect 671540 470594 671568 480626
rect 670804 162574 671200 162602
rect 671264 166966 671384 166994
rect 671448 470566 671568 470594
rect 670804 154574 670832 162574
rect 671264 155145 671292 166966
rect 671250 155136 671306 155145
rect 671250 155071 671306 155080
rect 670804 154546 671200 154574
rect 670608 150408 670660 150414
rect 670608 150350 670660 150356
rect 671172 139398 671200 154546
rect 671448 146266 671476 470566
rect 671620 392420 671672 392426
rect 671620 392362 671672 392368
rect 671436 146260 671488 146266
rect 671436 146202 671488 146208
rect 671632 140758 671660 392362
rect 671804 353388 671856 353394
rect 671804 353330 671856 353336
rect 671816 338094 671844 353330
rect 671804 338088 671856 338094
rect 671804 338030 671856 338036
rect 671804 261316 671856 261322
rect 671804 261258 671856 261264
rect 671816 247081 671844 261258
rect 671802 247072 671858 247081
rect 671802 247007 671858 247016
rect 671988 216844 672040 216850
rect 671988 216786 672040 216792
rect 671804 213716 671856 213722
rect 671804 213658 671856 213664
rect 671816 201278 671844 213658
rect 671804 201272 671856 201278
rect 671804 201214 671856 201220
rect 672000 198694 672028 216786
rect 672184 215294 672212 614858
rect 672354 586256 672410 586265
rect 672354 586191 672410 586200
rect 672368 393281 672396 586191
rect 672552 574394 672580 645351
rect 672736 616622 672764 688599
rect 672920 678974 672948 688758
rect 672828 678946 672948 678974
rect 672828 649994 672856 678946
rect 673012 669798 673040 714002
rect 673196 713726 673224 758202
rect 673380 755070 673408 862854
rect 673644 779816 673696 779822
rect 673644 779758 673696 779764
rect 673368 755064 673420 755070
rect 673368 755006 673420 755012
rect 673458 732728 673514 732737
rect 673458 732663 673514 732672
rect 673184 713720 673236 713726
rect 673184 713662 673236 713668
rect 673000 669792 673052 669798
rect 673000 669734 673052 669740
rect 673276 667276 673328 667282
rect 673276 667218 673328 667224
rect 673288 659654 673316 667218
rect 673472 663270 673500 732663
rect 673656 707198 673684 779758
rect 673828 779136 673880 779142
rect 673828 779078 673880 779084
rect 673840 708014 673868 779078
rect 674024 756294 674052 873174
rect 675404 872273 675432 872576
rect 675390 872264 675446 872273
rect 675390 872199 675446 872208
rect 675680 869689 675708 870060
rect 675666 869680 675722 869689
rect 675666 869615 675722 869624
rect 674838 869544 674894 869553
rect 674838 869479 674894 869488
rect 675128 869502 675418 869530
rect 674656 868080 674708 868086
rect 674656 868022 674708 868028
rect 674472 864680 674524 864686
rect 674472 864622 674524 864628
rect 674288 784168 674340 784174
rect 674288 784110 674340 784116
rect 674300 777186 674328 784110
rect 674300 777158 674420 777186
rect 674196 777028 674248 777034
rect 674196 776970 674248 776976
rect 674012 756288 674064 756294
rect 674012 756230 674064 756236
rect 674012 738676 674064 738682
rect 674012 738618 674064 738624
rect 673828 708008 673880 708014
rect 673828 707950 673880 707956
rect 673644 707192 673696 707198
rect 673644 707134 673696 707140
rect 673644 694204 673696 694210
rect 673644 694146 673696 694152
rect 673460 663264 673512 663270
rect 673460 663206 673512 663212
rect 673288 659626 673408 659654
rect 672828 649966 673224 649994
rect 673196 627914 673224 649966
rect 673380 640334 673408 659626
rect 673656 640626 673684 694146
rect 673828 693388 673880 693394
rect 673828 693330 673880 693336
rect 673840 640626 673868 693330
rect 674024 683097 674052 738618
rect 674208 727569 674236 776970
rect 674392 756254 674420 777158
rect 674484 772290 674512 864622
rect 674668 772449 674696 868022
rect 674852 856994 674880 869479
rect 675128 869446 675156 869502
rect 675116 869440 675168 869446
rect 675116 869382 675168 869388
rect 675024 869032 675076 869038
rect 674944 868980 675024 868986
rect 674944 868974 675076 868980
rect 674944 868958 675064 868974
rect 674944 866538 674972 868958
rect 675128 868861 675418 868889
rect 675128 868086 675156 868861
rect 675116 868080 675168 868086
rect 675496 868057 675524 868224
rect 675116 868022 675168 868028
rect 675482 868048 675538 868057
rect 675482 867983 675538 867992
rect 675128 867021 675418 867049
rect 675128 866862 675156 867021
rect 675116 866856 675168 866862
rect 675116 866798 675168 866804
rect 674944 866510 675340 866538
rect 675024 866448 675076 866454
rect 675024 866390 675076 866396
rect 675036 864566 675064 866390
rect 675312 865858 675340 866510
rect 675312 865830 675418 865858
rect 675312 865181 675418 865209
rect 675312 864686 675340 865181
rect 675300 864680 675352 864686
rect 675300 864622 675352 864628
rect 675036 864538 675418 864566
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675128 863314 675340 863342
rect 675404 863328 675432 863382
rect 675128 862918 675156 863314
rect 675116 862912 675168 862918
rect 675116 862854 675168 862860
rect 674852 856966 675340 856994
rect 675312 799034 675340 856966
rect 674852 799006 675340 799034
rect 674852 775946 674880 799006
rect 675116 789404 675168 789410
rect 674944 789352 675116 789374
rect 674944 789346 675168 789352
rect 674944 787693 674972 789346
rect 675128 788310 675418 788338
rect 675128 788050 675156 788310
rect 675116 788044 675168 788050
rect 675116 787986 675168 787992
rect 674944 787665 675418 787693
rect 674944 787018 675418 787046
rect 674944 776030 674972 787018
rect 675128 785182 675418 785210
rect 675128 784174 675156 785182
rect 675312 784638 675418 784666
rect 675312 784281 675340 784638
rect 675298 784272 675354 784281
rect 675298 784207 675354 784216
rect 675116 784168 675168 784174
rect 675116 784110 675168 784116
rect 675312 784094 675432 784122
rect 675114 784000 675170 784009
rect 675312 783986 675340 784094
rect 675170 783958 675340 783986
rect 675404 783972 675432 784094
rect 675114 783935 675170 783944
rect 675128 783346 675418 783374
rect 675128 782678 675156 783346
rect 675116 782672 675168 782678
rect 675116 782614 675168 782620
rect 675300 782536 675352 782542
rect 675300 782478 675352 782484
rect 675312 781402 675340 782478
rect 675312 781374 675432 781402
rect 675404 780844 675432 781374
rect 675312 780422 675432 780450
rect 675312 780314 675340 780422
rect 675128 780286 675340 780314
rect 675404 780300 675432 780422
rect 675128 779822 675156 780286
rect 675116 779816 675168 779822
rect 675116 779758 675168 779764
rect 675128 779674 675418 779702
rect 675128 779142 675156 779674
rect 675116 779136 675168 779142
rect 675116 779078 675168 779084
rect 675312 779062 675432 779090
rect 675116 779000 675168 779006
rect 675116 778942 675168 778948
rect 675128 776642 675156 778942
rect 675312 778394 675340 779062
rect 675404 779008 675432 779062
rect 675300 778388 675352 778394
rect 675300 778330 675352 778336
rect 675404 777322 675432 777852
rect 675312 777294 675432 777322
rect 675312 777034 675340 777294
rect 675300 777028 675352 777034
rect 675300 776970 675352 776976
rect 675128 776614 675418 776642
rect 674944 776002 675064 776030
rect 674840 775940 674892 775946
rect 674840 775882 674892 775888
rect 675036 775810 675064 776002
rect 675208 775940 675260 775946
rect 675208 775882 675260 775888
rect 675024 775804 675076 775810
rect 675024 775746 675076 775752
rect 675220 775690 675248 775882
rect 675128 775662 675248 775690
rect 674840 775600 674892 775606
rect 674840 775542 674892 775548
rect 674852 772970 674880 775542
rect 674852 772942 674972 772970
rect 674654 772440 674710 772449
rect 674654 772375 674710 772384
rect 674484 772262 674696 772290
rect 674668 772177 674696 772262
rect 674654 772168 674710 772177
rect 674654 772103 674710 772112
rect 674944 766601 674972 772942
rect 675128 770681 675156 775662
rect 675404 775554 675432 776016
rect 675312 775526 675432 775554
rect 675312 772814 675340 775526
rect 675496 775033 675524 775336
rect 675482 775024 675538 775033
rect 675482 774959 675538 774968
rect 675496 773809 675524 774180
rect 675482 773800 675538 773809
rect 675482 773735 675538 773744
rect 675312 772786 675432 772814
rect 675114 770672 675170 770681
rect 675114 770607 675170 770616
rect 674930 766592 674986 766601
rect 674930 766527 674986 766536
rect 675404 766426 675432 772786
rect 679622 772712 679678 772721
rect 679622 772647 679678 772656
rect 676034 772440 676090 772449
rect 676034 772375 676090 772384
rect 676048 772274 676076 772375
rect 676036 772268 676088 772274
rect 676036 772210 676088 772216
rect 675850 772168 675906 772177
rect 675850 772103 675852 772112
rect 675904 772103 675906 772112
rect 675852 772074 675904 772080
rect 675850 770672 675906 770681
rect 675850 770607 675906 770616
rect 674932 766420 674984 766426
rect 674932 766362 674984 766368
rect 675392 766420 675444 766426
rect 675392 766362 675444 766368
rect 674300 756226 674420 756254
rect 674300 746594 674328 756226
rect 674944 752457 674972 766362
rect 675482 761560 675538 761569
rect 675482 761495 675538 761504
rect 675298 761152 675354 761161
rect 675298 761087 675354 761096
rect 675312 760578 675340 761087
rect 675496 760918 675524 761495
rect 675484 760912 675536 760918
rect 675484 760854 675536 760860
rect 675482 760744 675538 760753
rect 675482 760679 675538 760688
rect 675300 760572 675352 760578
rect 675300 760514 675352 760520
rect 675496 760442 675524 760679
rect 675484 760436 675536 760442
rect 675484 760378 675536 760384
rect 675298 760336 675354 760345
rect 675298 760271 675300 760280
rect 675352 760271 675354 760280
rect 675300 760242 675352 760248
rect 675482 759928 675538 759937
rect 675482 759863 675484 759872
rect 675536 759863 675538 759872
rect 675484 759834 675536 759840
rect 675484 759552 675536 759558
rect 675482 759520 675484 759529
rect 675536 759520 675538 759529
rect 675482 759455 675538 759464
rect 675482 759112 675538 759121
rect 675482 759047 675484 759056
rect 675536 759047 675538 759056
rect 675484 759018 675536 759024
rect 675484 758736 675536 758742
rect 675482 758704 675484 758713
rect 675536 758704 675538 758713
rect 675482 758639 675538 758648
rect 675482 758296 675538 758305
rect 675482 758231 675484 758240
rect 675536 758231 675538 758240
rect 675484 758202 675536 758208
rect 675484 757920 675536 757926
rect 675482 757888 675484 757897
rect 675536 757888 675538 757897
rect 675482 757823 675538 757832
rect 675482 757480 675538 757489
rect 675482 757415 675484 757424
rect 675536 757415 675538 757424
rect 675484 757386 675536 757392
rect 675116 756288 675168 756294
rect 675116 756230 675168 756236
rect 675128 753817 675156 756230
rect 675864 755857 675892 770607
rect 679636 756265 679664 772647
rect 683304 772268 683356 772274
rect 683304 772210 683356 772216
rect 682382 768768 682438 768777
rect 682382 768703 682438 768712
rect 679622 756256 679678 756265
rect 679622 756191 679678 756200
rect 675850 755848 675906 755857
rect 675850 755783 675906 755792
rect 682396 755449 682424 768703
rect 682382 755440 682438 755449
rect 682382 755375 682438 755384
rect 675484 755064 675536 755070
rect 675482 755032 675484 755041
rect 675536 755032 675538 755041
rect 675482 754967 675538 754976
rect 675484 754656 675536 754662
rect 675482 754624 675484 754633
rect 675536 754624 675538 754633
rect 675482 754559 675538 754568
rect 675484 754248 675536 754254
rect 675482 754216 675484 754225
rect 675536 754216 675538 754225
rect 675482 754151 675538 754160
rect 675114 753808 675170 753817
rect 675114 753743 675170 753752
rect 675484 753432 675536 753438
rect 675482 753400 675484 753409
rect 675536 753400 675538 753409
rect 675482 753335 675538 753344
rect 683316 753001 683344 772210
rect 684132 772132 684184 772138
rect 684132 772074 684184 772080
rect 684144 756673 684172 772074
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 684130 756664 684186 756673
rect 684130 756599 684186 756608
rect 675850 752992 675906 753001
rect 675850 752927 675906 752936
rect 683302 752992 683358 753001
rect 683302 752927 683358 752936
rect 674930 752448 674986 752457
rect 674930 752383 674986 752392
rect 675484 752208 675536 752214
rect 675482 752176 675484 752185
rect 675536 752176 675538 752185
rect 675482 752111 675538 752120
rect 675484 751800 675536 751806
rect 675482 751768 675484 751777
rect 675536 751768 675538 751777
rect 675482 751703 675538 751712
rect 675864 750990 675892 752927
rect 675852 750984 675904 750990
rect 675852 750926 675904 750932
rect 683120 750984 683172 750990
rect 683120 750926 683172 750932
rect 683132 750757 683160 750926
rect 683118 750748 683174 750757
rect 683118 750683 683174 750692
rect 675482 750136 675538 750145
rect 675482 750071 675484 750080
rect 675536 750071 675538 750080
rect 675484 750042 675536 750048
rect 674300 746566 674696 746594
rect 674472 739764 674524 739770
rect 674472 739706 674524 739712
rect 674194 727560 674250 727569
rect 674194 727495 674250 727504
rect 674196 687948 674248 687954
rect 674196 687890 674248 687896
rect 674010 683088 674066 683097
rect 674010 683023 674066 683032
rect 674208 649994 674236 687890
rect 674484 664057 674512 739706
rect 674668 728113 674696 746566
rect 675116 743708 675168 743714
rect 675116 743650 675168 743656
rect 675128 742710 675156 743650
rect 675312 743294 675418 743322
rect 675312 742830 675340 743294
rect 675300 742824 675352 742830
rect 675300 742766 675352 742772
rect 675128 742682 675340 742710
rect 675312 742642 675340 742682
rect 675404 742642 675432 742696
rect 675312 742614 675432 742642
rect 675300 742484 675352 742490
rect 675300 742426 675352 742432
rect 674840 741668 674892 741674
rect 674840 741610 674892 741616
rect 674654 728104 674710 728113
rect 674654 728039 674710 728048
rect 674852 721585 674880 741610
rect 675312 740194 675340 742426
rect 675496 741674 675524 742016
rect 675484 741668 675536 741674
rect 675484 741610 675536 741616
rect 675312 740166 675418 740194
rect 675116 739764 675168 739770
rect 675116 739706 675168 739712
rect 675128 739650 675156 739706
rect 675128 739622 675418 739650
rect 675404 738682 675432 739024
rect 675392 738676 675444 738682
rect 675392 738618 675444 738624
rect 675128 738330 675418 738358
rect 675128 738177 675156 738330
rect 675114 738168 675170 738177
rect 675114 738103 675170 738112
rect 675128 735882 675340 735910
rect 675128 733009 675156 735882
rect 675312 735842 675340 735882
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 675312 735305 675418 735333
rect 675312 735010 675340 735305
rect 675300 735004 675352 735010
rect 675300 734946 675352 734952
rect 675300 734868 675352 734874
rect 675300 734810 675352 734816
rect 675114 733000 675170 733009
rect 675114 732935 675170 732944
rect 675116 732828 675168 732834
rect 675116 732770 675168 732776
rect 675128 731014 675156 732770
rect 675312 732034 675340 734810
rect 675496 734233 675524 734672
rect 675482 734224 675538 734233
rect 675482 734159 675538 734168
rect 675496 733689 675524 734031
rect 675482 733680 675538 733689
rect 675482 733615 675538 733624
rect 675496 732737 675524 732836
rect 675482 732728 675538 732737
rect 675482 732663 675538 732672
rect 675312 732006 675432 732034
rect 675404 731612 675432 732006
rect 675128 730986 675418 731014
rect 675128 730337 675418 730365
rect 675128 730153 675156 730337
rect 675114 730144 675170 730153
rect 675114 730079 675170 730088
rect 675128 729150 675418 729178
rect 675128 728686 675156 729150
rect 675116 728680 675168 728686
rect 675116 728622 675168 728628
rect 675850 728104 675906 728113
rect 675850 728039 675906 728048
rect 677506 728104 677562 728113
rect 677506 728039 677562 728048
rect 675864 726850 675892 728039
rect 676034 727560 676090 727569
rect 676034 727495 676090 727504
rect 675852 726844 675904 726850
rect 675852 726786 675904 726792
rect 676048 726578 676076 727495
rect 676036 726572 676088 726578
rect 676036 726514 676088 726520
rect 674838 721576 674894 721585
rect 674838 721511 674894 721520
rect 675484 716576 675536 716582
rect 675482 716544 675484 716553
rect 675536 716544 675538 716553
rect 675482 716479 675538 716488
rect 675298 716136 675354 716145
rect 675298 716071 675354 716080
rect 675116 715352 675168 715358
rect 675114 715320 675116 715329
rect 675168 715320 675170 715329
rect 675114 715255 675170 715264
rect 675312 715018 675340 716071
rect 675482 715728 675538 715737
rect 675482 715663 675538 715672
rect 675496 715154 675524 715663
rect 675484 715148 675536 715154
rect 675484 715090 675536 715096
rect 675300 715012 675352 715018
rect 675300 714954 675352 714960
rect 675482 714912 675538 714921
rect 675482 714847 675484 714856
rect 675536 714847 675538 714856
rect 675484 714818 675536 714824
rect 675484 714536 675536 714542
rect 675482 714504 675484 714513
rect 675536 714504 675538 714513
rect 675482 714439 675538 714448
rect 675482 714096 675538 714105
rect 675482 714031 675484 714040
rect 675536 714031 675538 714040
rect 675484 714002 675536 714008
rect 675484 713720 675536 713726
rect 675482 713688 675484 713697
rect 675536 713688 675538 713697
rect 675482 713623 675538 713632
rect 676770 713488 676826 713497
rect 676770 713423 676826 713432
rect 675482 713280 675538 713289
rect 675482 713215 675484 713224
rect 675536 713215 675538 713224
rect 675484 713186 675536 713192
rect 675484 712904 675536 712910
rect 675482 712872 675484 712881
rect 675536 712872 675538 712881
rect 675482 712807 675538 712816
rect 675482 712464 675538 712473
rect 675482 712399 675484 712408
rect 675536 712399 675538 712408
rect 675484 712370 675536 712376
rect 676220 712088 676272 712094
rect 676034 712056 676090 712065
rect 676090 712036 676220 712042
rect 676090 712030 676272 712036
rect 676090 712014 676260 712030
rect 676034 711991 676090 712000
rect 676784 711890 676812 713423
rect 677520 712094 677548 728039
rect 683394 727832 683450 727841
rect 683394 727767 683450 727776
rect 683212 726572 683264 726578
rect 683212 726514 683264 726520
rect 677508 712088 677560 712094
rect 677508 712030 677560 712036
rect 676036 711884 676088 711890
rect 676036 711826 676088 711832
rect 676772 711884 676824 711890
rect 676772 711826 676824 711832
rect 676048 711657 676076 711826
rect 676034 711648 676090 711657
rect 676034 711583 676090 711592
rect 675484 711272 675536 711278
rect 675482 711240 675484 711249
rect 675536 711240 675538 711249
rect 675482 711175 675538 711184
rect 675850 710696 675906 710705
rect 675850 710631 675906 710640
rect 675298 710424 675354 710433
rect 675298 710359 675354 710368
rect 675312 709374 675340 710359
rect 675482 710016 675538 710025
rect 675482 709951 675538 709960
rect 675496 709782 675524 709951
rect 675484 709776 675536 709782
rect 675484 709718 675536 709724
rect 675484 709640 675536 709646
rect 675482 709608 675484 709617
rect 675536 709608 675538 709617
rect 675482 709543 675538 709552
rect 675300 709368 675352 709374
rect 675300 709310 675352 709316
rect 675484 708008 675536 708014
rect 675482 707976 675484 707985
rect 675536 707976 675538 707985
rect 675482 707911 675538 707920
rect 675484 707600 675536 707606
rect 675482 707568 675484 707577
rect 675536 707568 675538 707577
rect 675482 707503 675538 707512
rect 675484 707192 675536 707198
rect 675482 707160 675484 707169
rect 675536 707160 675538 707169
rect 675482 707095 675538 707104
rect 675484 706784 675536 706790
rect 675482 706752 675484 706761
rect 675536 706752 675538 706761
rect 675482 706687 675538 706696
rect 675864 705226 675892 710631
rect 683224 708393 683252 726514
rect 683408 709209 683436 727767
rect 684224 726844 684276 726850
rect 684224 726786 684276 726792
rect 684236 710841 684264 726786
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 684222 710832 684278 710841
rect 684222 710767 684278 710776
rect 683394 709200 683450 709209
rect 683394 709135 683450 709144
rect 683210 708384 683266 708393
rect 683210 708319 683266 708328
rect 683118 705528 683174 705537
rect 683118 705463 683174 705472
rect 683132 705226 683160 705463
rect 675852 705220 675904 705226
rect 675852 705162 675904 705168
rect 683120 705220 683172 705226
rect 683120 705162 683172 705168
rect 675482 705120 675538 705129
rect 675482 705055 675484 705064
rect 675536 705055 675538 705064
rect 675484 705026 675536 705032
rect 675116 699712 675168 699718
rect 675116 699654 675168 699660
rect 675128 697694 675156 699654
rect 675390 698592 675446 698601
rect 675390 698527 675446 698536
rect 675404 698323 675432 698527
rect 675128 697666 675418 697694
rect 675404 696833 675432 697035
rect 675390 696824 675446 696833
rect 675390 696759 675446 696768
rect 675128 695181 675418 695209
rect 675128 694210 675156 695181
rect 675680 694385 675708 694620
rect 675666 694376 675722 694385
rect 675666 694311 675722 694320
rect 675116 694204 675168 694210
rect 675116 694146 675168 694152
rect 675128 693994 675418 694022
rect 675128 693394 675156 693994
rect 675116 693388 675168 693394
rect 675116 693330 675168 693336
rect 675496 693138 675524 693328
rect 675404 693110 675524 693138
rect 675404 693054 675432 693110
rect 674656 693048 674708 693054
rect 674656 692990 674708 692996
rect 675392 693048 675444 693054
rect 675392 692990 675444 692996
rect 674470 664048 674526 664057
rect 674470 663983 674526 663992
rect 674208 649966 674328 649994
rect 674102 644328 674158 644337
rect 674102 644263 674158 644272
rect 674116 642649 674144 644263
rect 674116 642621 674236 642649
rect 673644 640620 673696 640626
rect 673644 640562 673696 640568
rect 673828 640620 673880 640626
rect 673828 640562 673880 640568
rect 674010 640520 674066 640529
rect 673104 627886 673224 627914
rect 673288 640306 673408 640334
rect 673472 640478 674010 640506
rect 672908 624708 672960 624714
rect 672908 624650 672960 624656
rect 672724 616616 672776 616622
rect 672724 616558 672776 616564
rect 672920 611354 672948 624650
rect 673104 622724 673132 627886
rect 673288 622826 673316 640306
rect 673472 622946 673500 640478
rect 674010 640455 674066 640464
rect 673644 640348 673696 640354
rect 673644 640290 673696 640296
rect 673828 640348 673880 640354
rect 674208 640334 674236 642621
rect 673828 640290 673880 640296
rect 674116 640306 674236 640334
rect 673656 637129 673684 640290
rect 673642 637120 673698 637129
rect 673642 637055 673698 637064
rect 673460 622940 673512 622946
rect 673460 622882 673512 622888
rect 673288 622798 673684 622826
rect 673656 622742 673684 622798
rect 673460 622736 673512 622742
rect 673104 622696 673316 622724
rect 673092 619132 673144 619138
rect 673092 619074 673144 619080
rect 673104 611354 673132 619074
rect 673288 617030 673316 622696
rect 673460 622678 673512 622684
rect 673644 622736 673696 622742
rect 673644 622678 673696 622684
rect 673276 617024 673328 617030
rect 673276 616966 673328 616972
rect 672920 611326 673040 611354
rect 673104 611326 673316 611354
rect 672722 598496 672778 598505
rect 672722 598431 672778 598440
rect 672540 574388 672592 574394
rect 672540 574330 672592 574336
rect 672540 532772 672592 532778
rect 672540 532714 672592 532720
rect 672552 488714 672580 532714
rect 672736 526454 672764 598431
rect 673012 580038 673040 611326
rect 673000 580032 673052 580038
rect 673000 579974 673052 579980
rect 673288 578542 673316 611326
rect 673472 592929 673500 622678
rect 673840 618633 673868 640290
rect 673826 618624 673882 618633
rect 673826 618559 673882 618568
rect 673644 603492 673696 603498
rect 673644 603434 673696 603440
rect 673458 592920 673514 592929
rect 673458 592855 673514 592864
rect 673276 578536 673328 578542
rect 673276 578478 673328 578484
rect 673092 578400 673144 578406
rect 673092 578342 673144 578348
rect 672908 578264 672960 578270
rect 672908 578206 672960 578212
rect 672920 534410 672948 578206
rect 673104 534614 673132 578342
rect 673460 577652 673512 577658
rect 673460 577594 673512 577600
rect 673472 577130 673500 577594
rect 673380 577102 673500 577130
rect 673380 577046 673408 577102
rect 673368 577040 673420 577046
rect 673368 576982 673420 576988
rect 673276 557728 673328 557734
rect 673276 557670 673328 557676
rect 673092 534608 673144 534614
rect 673092 534550 673144 534556
rect 672908 534404 672960 534410
rect 672908 534346 672960 534352
rect 673000 534132 673052 534138
rect 673000 534074 673052 534080
rect 672724 526448 672776 526454
rect 672724 526390 672776 526396
rect 673012 490074 673040 534074
rect 673000 490068 673052 490074
rect 673000 490010 673052 490016
rect 672540 488708 672592 488714
rect 672540 488650 672592 488656
rect 673288 483206 673316 557670
rect 673460 554192 673512 554198
rect 673460 554134 673512 554140
rect 673472 483614 673500 554134
rect 673656 528494 673684 603434
rect 673918 599176 673974 599185
rect 673918 599111 673974 599120
rect 673932 597530 673960 599111
rect 674116 598934 674144 640306
rect 674300 617817 674328 649966
rect 674470 644736 674526 644745
rect 674470 644671 674526 644680
rect 674286 617808 674342 617817
rect 674286 617743 674342 617752
rect 674288 604376 674340 604382
rect 674288 604318 674340 604324
rect 674116 598906 674236 598934
rect 673932 597502 674052 597530
rect 673826 597408 673882 597417
rect 673826 597343 673882 597352
rect 673644 528488 673696 528494
rect 673644 528430 673696 528436
rect 673840 528086 673868 597343
rect 673828 528080 673880 528086
rect 673828 528022 673880 528028
rect 674024 527649 674052 597502
rect 674208 591297 674236 598906
rect 674300 592090 674328 604318
rect 674484 592249 674512 644671
rect 674668 640334 674696 692990
rect 675116 692912 675168 692918
rect 675116 692854 675168 692860
rect 675128 690894 675156 692854
rect 675128 690866 675418 690894
rect 675128 690322 675340 690350
rect 675128 690062 675156 690322
rect 675312 690282 675340 690322
rect 675404 690282 675432 690336
rect 675312 690254 675432 690282
rect 675116 690056 675168 690062
rect 675116 689998 675168 690004
rect 675312 689710 675432 689738
rect 674932 689308 674984 689314
rect 674932 689250 674984 689256
rect 674944 686678 674972 689250
rect 675312 687954 675340 689710
rect 675404 689656 675432 689710
rect 675496 688673 675524 689044
rect 675482 688664 675538 688673
rect 675482 688599 675538 688608
rect 675300 687948 675352 687954
rect 675300 687890 675352 687896
rect 675128 687806 675418 687834
rect 675128 687478 675156 687806
rect 675116 687472 675168 687478
rect 675116 687414 675168 687420
rect 674944 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675128 685970 675418 685998
rect 675128 685794 675156 685970
rect 674852 685766 675156 685794
rect 674852 678974 674880 685766
rect 675300 685568 675352 685574
rect 675300 685510 675352 685516
rect 675022 685264 675078 685273
rect 675022 685199 675078 685208
rect 675036 679130 675064 685199
rect 675312 684162 675340 685510
rect 675496 685001 675524 685372
rect 675482 684992 675538 685001
rect 675482 684927 675538 684936
rect 675312 684134 675418 684162
rect 675850 683088 675906 683097
rect 675850 683023 675906 683032
rect 675864 682446 675892 683023
rect 675852 682440 675904 682446
rect 675852 682382 675904 682388
rect 683396 682440 683448 682446
rect 683396 682382 683448 682388
rect 675036 679102 675156 679130
rect 674852 678946 675064 678974
rect 674840 669792 674892 669798
rect 674840 669734 674892 669740
rect 674852 669361 674880 669734
rect 674838 669352 674894 669361
rect 674838 669287 674894 669296
rect 674838 649224 674894 649233
rect 674838 649159 674840 649168
rect 674892 649159 674894 649168
rect 674840 649130 674892 649136
rect 674840 644496 674892 644502
rect 674840 644438 674892 644444
rect 674852 643113 674880 644438
rect 674838 643104 674894 643113
rect 674838 643039 674894 643048
rect 674840 641912 674892 641918
rect 674840 641854 674892 641860
rect 674576 640306 674696 640334
rect 674576 630674 674604 640306
rect 674852 639441 674880 641854
rect 674838 639432 674894 639441
rect 674838 639367 674894 639376
rect 675036 637401 675064 678946
rect 675128 640334 675156 679102
rect 678242 678328 678298 678337
rect 678242 678263 678298 678272
rect 675298 671392 675354 671401
rect 675298 671327 675354 671336
rect 675312 670886 675340 671327
rect 675482 670984 675538 670993
rect 675482 670919 675538 670928
rect 675300 670880 675352 670886
rect 675300 670822 675352 670828
rect 675496 670750 675524 670919
rect 675484 670744 675536 670750
rect 675484 670686 675536 670692
rect 675666 670576 675722 670585
rect 675666 670511 675722 670520
rect 675298 670168 675354 670177
rect 675298 670103 675354 670112
rect 675312 669662 675340 670103
rect 675482 669760 675538 669769
rect 675482 669695 675538 669704
rect 675300 669656 675352 669662
rect 675300 669598 675352 669604
rect 675496 669526 675524 669695
rect 675484 669520 675536 669526
rect 675484 669462 675536 669468
rect 675484 669384 675536 669390
rect 675680 669338 675708 670511
rect 675536 669332 675708 669338
rect 675484 669326 675708 669332
rect 675496 669310 675708 669326
rect 675298 668944 675354 668953
rect 675298 668879 675354 668888
rect 675312 668438 675340 668879
rect 675484 668568 675536 668574
rect 675482 668536 675484 668545
rect 675536 668536 675538 668545
rect 675482 668471 675538 668480
rect 675300 668432 675352 668438
rect 675300 668374 675352 668380
rect 675482 668128 675538 668137
rect 675482 668063 675484 668072
rect 675536 668063 675538 668072
rect 675484 668034 675536 668040
rect 675484 667752 675536 667758
rect 675482 667720 675484 667729
rect 675536 667720 675538 667729
rect 675482 667655 675538 667664
rect 675482 667312 675538 667321
rect 675482 667247 675484 667256
rect 675536 667247 675538 667256
rect 675484 667218 675536 667224
rect 678256 667049 678284 678263
rect 683210 674112 683266 674121
rect 683210 674047 683266 674056
rect 678242 667040 678298 667049
rect 678242 666975 678298 666984
rect 675298 666496 675354 666505
rect 675298 666431 675354 666440
rect 675312 665378 675340 666431
rect 675484 666120 675536 666126
rect 675482 666088 675484 666097
rect 675536 666088 675538 666097
rect 675482 666023 675538 666032
rect 675482 665680 675538 665689
rect 675482 665615 675538 665624
rect 675300 665372 675352 665378
rect 675300 665314 675352 665320
rect 675496 665242 675524 665615
rect 675484 665236 675536 665242
rect 675484 665178 675536 665184
rect 675484 664896 675536 664902
rect 675482 664864 675484 664873
rect 675536 664864 675538 664873
rect 675482 664799 675538 664808
rect 675482 664456 675538 664465
rect 675482 664391 675538 664400
rect 675496 663814 675524 664391
rect 675484 663808 675536 663814
rect 675484 663750 675536 663756
rect 675850 663504 675906 663513
rect 675850 663439 675906 663448
rect 675484 663264 675536 663270
rect 675482 663232 675484 663241
rect 675536 663232 675538 663241
rect 675482 663167 675538 663176
rect 675484 662856 675536 662862
rect 675482 662824 675484 662833
rect 675536 662824 675538 662833
rect 675482 662759 675538 662768
rect 675484 662040 675536 662046
rect 675482 662008 675484 662017
rect 675536 662008 675538 662017
rect 675482 661943 675538 661952
rect 675484 661632 675536 661638
rect 675482 661600 675484 661609
rect 675536 661600 675538 661609
rect 675482 661535 675538 661544
rect 675482 661192 675538 661201
rect 675482 661127 675484 661136
rect 675536 661127 675538 661136
rect 675484 661098 675536 661104
rect 675484 660000 675536 660006
rect 675482 659968 675484 659977
rect 675536 659968 675538 659977
rect 675482 659903 675538 659912
rect 675864 659870 675892 663439
rect 683224 662561 683252 674047
rect 683408 663785 683436 682382
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683394 663776 683450 663785
rect 683394 663711 683450 663720
rect 683210 662552 683266 662561
rect 683210 662487 683266 662496
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 683132 659870 683160 660039
rect 675852 659864 675904 659870
rect 675852 659806 675904 659812
rect 683120 659864 683172 659870
rect 683120 659806 683172 659812
rect 675300 654152 675352 654158
rect 675300 654094 675352 654100
rect 675312 653018 675340 654094
rect 675312 652990 675432 653018
rect 675404 652460 675432 652990
rect 675588 652905 675616 653140
rect 675574 652896 675630 652905
rect 675574 652831 675630 652840
rect 675312 651834 675418 651862
rect 675312 651438 675340 651834
rect 675300 651432 675352 651438
rect 675300 651374 675352 651380
rect 675220 649998 675340 650026
rect 675220 647234 675248 649998
rect 675312 649994 675340 649998
rect 675404 649994 675432 650012
rect 675312 649966 675432 649994
rect 675496 649233 675524 649468
rect 675482 649224 675538 649233
rect 675482 649159 675538 649168
rect 675588 648689 675616 648788
rect 675574 648680 675630 648689
rect 675574 648615 675630 648624
rect 675404 647766 675432 648176
rect 675392 647760 675444 647766
rect 675392 647702 675444 647708
rect 675220 647206 675340 647234
rect 675312 645833 675340 647206
rect 675298 645824 675354 645833
rect 675298 645759 675354 645768
rect 675496 645425 675524 645660
rect 675482 645416 675538 645425
rect 675482 645351 675538 645360
rect 675404 644745 675432 645116
rect 675390 644736 675446 644745
rect 675390 644671 675446 644680
rect 675404 644337 675432 644475
rect 675390 644328 675446 644337
rect 675390 644263 675446 644272
rect 675300 643680 675352 643686
rect 675300 643622 675352 643628
rect 675312 641458 675340 643622
rect 675496 643521 675524 643824
rect 675482 643512 675538 643521
rect 675482 643447 675538 643456
rect 675482 643104 675538 643113
rect 675482 643039 675538 643048
rect 675496 642635 675524 643039
rect 675312 641430 675418 641458
rect 675300 641300 675352 641306
rect 675300 641242 675352 641248
rect 675128 640306 675248 640334
rect 675220 638217 675248 640306
rect 675312 640166 675340 641242
rect 675496 640529 675524 640795
rect 675482 640520 675538 640529
rect 675482 640455 675538 640464
rect 675312 640138 675418 640166
rect 675390 639432 675446 639441
rect 675390 639367 675446 639376
rect 675404 638928 675432 639367
rect 675206 638208 675262 638217
rect 675206 638143 675262 638152
rect 675758 638208 675814 638217
rect 675758 638143 675814 638152
rect 675298 637800 675354 637809
rect 675298 637735 675354 637744
rect 675312 637574 675340 637735
rect 675574 637664 675630 637673
rect 675574 637599 675630 637608
rect 675220 637546 675340 637574
rect 675022 637392 675078 637401
rect 675022 637327 675078 637336
rect 675220 633706 675248 637546
rect 675220 633678 675340 633706
rect 674576 630646 674696 630674
rect 674668 617409 674696 630646
rect 675114 625968 675170 625977
rect 675114 625903 675170 625912
rect 675128 625190 675156 625903
rect 675116 625184 675168 625190
rect 675116 625126 675168 625132
rect 674838 623928 674894 623937
rect 674838 623863 674894 623872
rect 674852 619138 674880 623863
rect 675312 621014 675340 633678
rect 675588 631417 675616 637599
rect 675772 637574 675800 638143
rect 675772 637546 675892 637574
rect 675864 633622 675892 637546
rect 676036 637560 676088 637566
rect 676036 637502 676088 637508
rect 682384 637560 682436 637566
rect 682384 637502 682436 637508
rect 676048 637401 676076 637502
rect 676034 637392 676090 637401
rect 676034 637327 676090 637336
rect 676034 637120 676090 637129
rect 676034 637055 676090 637064
rect 676048 636886 676076 637055
rect 676036 636880 676088 636886
rect 676036 636822 676088 636828
rect 675852 633616 675904 633622
rect 675852 633558 675904 633564
rect 675574 631408 675630 631417
rect 675574 631343 675630 631352
rect 675482 626376 675538 626385
rect 675482 626311 675538 626320
rect 675496 625734 675524 626311
rect 675484 625728 675536 625734
rect 675484 625670 675536 625676
rect 675482 625560 675538 625569
rect 675482 625495 675538 625504
rect 675496 625326 675524 625495
rect 675484 625320 675536 625326
rect 675484 625262 675536 625268
rect 675482 625152 675538 625161
rect 675482 625087 675538 625096
rect 675496 624986 675524 625087
rect 675484 624980 675536 624986
rect 675484 624922 675536 624928
rect 675482 624744 675538 624753
rect 675482 624679 675484 624688
rect 675536 624679 675538 624688
rect 675484 624650 675536 624656
rect 675484 624368 675536 624374
rect 675482 624336 675484 624345
rect 675536 624336 675538 624345
rect 675482 624271 675538 624280
rect 675484 623552 675536 623558
rect 675482 623520 675484 623529
rect 675536 623520 675538 623529
rect 675482 623455 675538 623464
rect 675482 623112 675538 623121
rect 675482 623047 675484 623056
rect 675536 623047 675538 623056
rect 675484 623018 675536 623024
rect 675484 622736 675536 622742
rect 675482 622704 675484 622713
rect 675536 622704 675538 622713
rect 675482 622639 675538 622648
rect 675482 622296 675538 622305
rect 675482 622231 675484 622240
rect 675536 622231 675538 622240
rect 675484 622202 675536 622208
rect 682396 621625 682424 637502
rect 683304 636880 683356 636886
rect 683304 636822 683356 636828
rect 682568 633616 682620 633622
rect 682568 633558 682620 633564
rect 682580 622033 682608 633558
rect 682566 622024 682622 622033
rect 682566 621959 682622 621968
rect 682382 621616 682438 621625
rect 682382 621551 682438 621560
rect 675220 620986 675340 621014
rect 675024 619880 675076 619886
rect 675022 619848 675024 619857
rect 675076 619848 675078 619857
rect 675022 619783 675078 619792
rect 674840 619132 674892 619138
rect 674840 619074 674892 619080
rect 674654 617400 674710 617409
rect 674654 617335 674710 617344
rect 675220 611354 675248 620986
rect 683316 620809 683344 636822
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683302 620800 683358 620809
rect 683302 620735 683358 620744
rect 675482 620256 675538 620265
rect 675482 620191 675538 620200
rect 675496 619682 675524 620191
rect 675484 619676 675536 619682
rect 675484 619618 675536 619624
rect 675482 619440 675538 619449
rect 675482 619375 675538 619384
rect 675496 618322 675524 619375
rect 675484 618316 675536 618322
rect 675484 618258 675536 618264
rect 675666 618216 675722 618225
rect 675496 618186 675666 618202
rect 675484 618180 675666 618186
rect 675536 618174 675666 618180
rect 675666 618151 675722 618160
rect 675484 618122 675536 618128
rect 675484 617024 675536 617030
rect 675482 616992 675484 617001
rect 675536 616992 675538 617001
rect 675482 616927 675538 616936
rect 675484 616616 675536 616622
rect 675482 616584 675484 616593
rect 675536 616584 675538 616593
rect 675482 616519 675538 616528
rect 675482 616176 675538 616185
rect 675482 616111 675484 616120
rect 675536 616111 675538 616120
rect 675484 616082 675536 616088
rect 675850 615904 675906 615913
rect 675850 615839 675906 615848
rect 675864 615670 675892 615839
rect 675852 615664 675904 615670
rect 675852 615606 675904 615612
rect 683120 615664 683172 615670
rect 683120 615606 683172 615612
rect 683132 615505 683160 615606
rect 683118 615496 683174 615505
rect 683118 615431 683174 615440
rect 675482 614952 675538 614961
rect 675482 614887 675484 614896
rect 675536 614887 675538 614896
rect 675484 614858 675536 614864
rect 675036 611326 675248 611354
rect 674840 603152 674892 603158
rect 674840 603094 674892 603100
rect 674852 601225 674880 603094
rect 674838 601216 674894 601225
rect 674838 601151 674894 601160
rect 675036 601066 675064 611326
rect 675208 608864 675260 608870
rect 675208 608806 675260 608812
rect 675220 606846 675248 608806
rect 675404 607889 675432 608124
rect 675390 607880 675446 607889
rect 675390 607815 675446 607824
rect 675772 607345 675800 607479
rect 675758 607336 675814 607345
rect 675758 607271 675814 607280
rect 675220 606818 675418 606846
rect 674944 601038 675064 601066
rect 675128 604982 675418 605010
rect 674944 597689 674972 601038
rect 674930 597680 674986 597689
rect 674930 597615 674986 597624
rect 675128 597530 675156 604982
rect 675312 604438 675418 604466
rect 675312 604382 675340 604438
rect 675300 604376 675352 604382
rect 675300 604318 675352 604324
rect 675496 603514 675524 603772
rect 675404 603498 675524 603514
rect 675392 603492 675524 603498
rect 675444 603486 675524 603492
rect 675392 603434 675444 603440
rect 675312 603146 675418 603174
rect 675312 602993 675340 603146
rect 675298 602984 675354 602993
rect 675298 602919 675354 602928
rect 675300 601724 675352 601730
rect 675220 601672 675300 601694
rect 675220 601666 675352 601672
rect 675220 600522 675248 601666
rect 675390 601216 675446 601225
rect 675390 601151 675446 601160
rect 675404 600644 675432 601151
rect 675220 600494 675432 600522
rect 675404 600100 675432 600494
rect 675300 599616 675352 599622
rect 675300 599558 675352 599564
rect 675036 597502 675156 597530
rect 674748 596216 674800 596222
rect 674800 596164 674880 596170
rect 674748 596158 674880 596164
rect 674760 596142 674880 596158
rect 674852 595082 674880 596142
rect 674760 595066 674880 595082
rect 674748 595060 674880 595066
rect 674800 595054 674880 595060
rect 674748 595002 674800 595008
rect 675036 594946 675064 597502
rect 675312 596442 675340 599558
rect 675496 599185 675524 599488
rect 675482 599176 675538 599185
rect 675482 599111 675538 599120
rect 675496 598505 675524 598808
rect 675482 598496 675538 598505
rect 675482 598431 675538 598440
rect 675496 597417 675524 597652
rect 675482 597408 675538 597417
rect 675482 597343 675538 597352
rect 675312 596414 675418 596442
rect 675404 595490 675432 595816
rect 675312 595462 675432 595490
rect 675312 595270 675340 595462
rect 675300 595264 675352 595270
rect 675300 595206 675352 595212
rect 675300 595060 675352 595066
rect 675300 595002 675352 595008
rect 675036 594918 675248 594946
rect 675022 594552 675078 594561
rect 675022 594487 675078 594496
rect 674470 592240 674526 592249
rect 674470 592175 674526 592184
rect 674300 592062 674604 592090
rect 674194 591288 674250 591297
rect 674194 591223 674250 591232
rect 674576 582374 674604 592062
rect 675036 589274 675064 594487
rect 675220 589274 675248 594918
rect 675312 593858 675340 595002
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675404 593858 675432 593980
rect 675312 593830 675432 593858
rect 675850 592920 675906 592929
rect 675850 592855 675906 592864
rect 675864 592686 675892 592855
rect 675852 592680 675904 592686
rect 675852 592622 675904 592628
rect 683304 592680 683356 592686
rect 683304 592622 683356 592628
rect 675852 592544 675904 592550
rect 675850 592512 675852 592521
rect 678244 592544 678296 592550
rect 675904 592512 675906 592521
rect 678244 592486 678296 592492
rect 675850 592447 675906 592456
rect 675850 592240 675906 592249
rect 675850 592175 675906 592184
rect 675864 591462 675892 592175
rect 675852 591456 675904 591462
rect 675852 591398 675904 591404
rect 675852 591320 675904 591326
rect 675850 591288 675852 591297
rect 675904 591288 675906 591297
rect 675850 591223 675906 591232
rect 675036 589246 675156 589274
rect 675220 589246 675340 589274
rect 674208 582346 674604 582374
rect 674208 547369 674236 582346
rect 674930 580680 674986 580689
rect 674930 580615 674986 580624
rect 674944 579834 674972 580615
rect 674932 579828 674984 579834
rect 674932 579770 674984 579776
rect 674930 579456 674986 579465
rect 674930 579391 674986 579400
rect 674944 578270 674972 579391
rect 674932 578264 674984 578270
rect 674932 578206 674984 578212
rect 674656 558272 674708 558278
rect 674656 558214 674708 558220
rect 674472 549772 674524 549778
rect 674472 549714 674524 549720
rect 674194 547360 674250 547369
rect 674194 547295 674250 547304
rect 674484 545494 674512 549714
rect 674472 545488 674524 545494
rect 674472 545430 674524 545436
rect 674470 535120 674526 535129
rect 674470 535055 674526 535064
rect 674484 534274 674512 535055
rect 674472 534268 674524 534274
rect 674472 534210 674524 534216
rect 674286 533624 674342 533633
rect 674286 533559 674342 533568
rect 674010 527640 674066 527649
rect 674010 527575 674066 527584
rect 673736 525836 673788 525842
rect 673736 525778 673788 525784
rect 673460 483608 673512 483614
rect 673460 483550 673512 483556
rect 673276 483200 673328 483206
rect 673276 483142 673328 483148
rect 672630 474872 672686 474881
rect 672630 474807 672686 474816
rect 672644 394346 672672 474807
rect 672816 400580 672868 400586
rect 672816 400522 672868 400528
rect 672828 398834 672856 400522
rect 673184 399764 673236 399770
rect 673184 399706 673236 399712
rect 672736 398806 672856 398834
rect 672736 396074 672764 398806
rect 672736 396046 672948 396074
rect 672644 394318 672764 394346
rect 672540 394188 672592 394194
rect 672540 394130 672592 394136
rect 672354 393272 672410 393281
rect 672354 393207 672410 393216
rect 672552 364334 672580 394130
rect 672736 391218 672764 394318
rect 672920 394194 672948 396046
rect 672908 394188 672960 394194
rect 672908 394130 672960 394136
rect 673000 394052 673052 394058
rect 673000 393994 673052 394000
rect 672460 364306 672580 364334
rect 672644 391190 672764 391218
rect 672460 355910 672488 364306
rect 672448 355904 672500 355910
rect 672448 355846 672500 355852
rect 672448 355428 672500 355434
rect 672448 355370 672500 355376
rect 672460 350534 672488 355370
rect 672460 350506 672580 350534
rect 672356 347268 672408 347274
rect 672356 347210 672408 347216
rect 672368 340874 672396 347210
rect 672368 340846 672488 340874
rect 672460 273254 672488 340846
rect 672552 316554 672580 350506
rect 672644 317414 672672 391190
rect 672814 389328 672870 389337
rect 672814 389263 672870 389272
rect 672828 372570 672856 389263
rect 673012 376650 673040 393994
rect 673000 376644 673052 376650
rect 673000 376586 673052 376592
rect 672816 372564 672868 372570
rect 672816 372506 672868 372512
rect 673196 355094 673224 399706
rect 673368 394460 673420 394466
rect 673368 394402 673420 394408
rect 673380 377874 673408 394402
rect 673368 377868 673420 377874
rect 673368 377810 673420 377816
rect 673184 355088 673236 355094
rect 673184 355030 673236 355036
rect 673184 354612 673236 354618
rect 673184 354554 673236 354560
rect 673000 348900 673052 348906
rect 673000 348842 673052 348848
rect 673012 331770 673040 348842
rect 673000 331764 673052 331770
rect 673000 331706 673052 331712
rect 672644 317386 673040 317414
rect 672552 316526 672764 316554
rect 672736 310865 672764 316526
rect 672722 310856 672778 310865
rect 672722 310791 672778 310800
rect 673012 307754 673040 317386
rect 673196 310078 673224 354554
rect 673368 350124 673420 350130
rect 673368 350066 673420 350072
rect 673380 336054 673408 350066
rect 673552 349716 673604 349722
rect 673552 349658 673604 349664
rect 673368 336048 673420 336054
rect 673368 335990 673420 335996
rect 673564 335918 673592 349658
rect 673552 335912 673604 335918
rect 673552 335854 673604 335860
rect 673552 324352 673604 324358
rect 673552 324294 673604 324300
rect 673184 310072 673236 310078
rect 673184 310014 673236 310020
rect 672644 307726 673040 307754
rect 672460 273226 672580 273254
rect 672356 258460 672408 258466
rect 672356 258402 672408 258408
rect 672092 215266 672212 215294
rect 672092 205634 672120 215266
rect 672368 213466 672396 258402
rect 672552 234614 672580 273226
rect 672460 234586 672580 234614
rect 672460 215294 672488 234586
rect 672644 217433 672672 307726
rect 673276 305516 673328 305522
rect 673276 305458 673328 305464
rect 673092 303884 673144 303890
rect 673092 303826 673144 303832
rect 672816 303476 672868 303482
rect 672816 303418 672868 303424
rect 672630 217424 672686 217433
rect 672630 217359 672686 217368
rect 672460 215266 672580 215294
rect 672368 213438 672488 213466
rect 672264 213308 672316 213314
rect 672264 213250 672316 213256
rect 672092 205606 672212 205634
rect 671988 198688 672040 198694
rect 671988 198630 672040 198636
rect 672184 176654 672212 205606
rect 672092 176626 672212 176654
rect 671804 169516 671856 169522
rect 671804 169458 671856 169464
rect 671816 167090 671844 169458
rect 672092 168337 672120 176626
rect 672078 168328 672134 168337
rect 672078 168263 672134 168272
rect 671986 168056 672042 168065
rect 671986 167991 672042 168000
rect 671724 167062 671844 167090
rect 671724 164098 671752 167062
rect 671724 164070 671844 164098
rect 671816 162110 671844 164070
rect 671804 162104 671856 162110
rect 671804 162046 671856 162052
rect 672000 159338 672028 167991
rect 671816 159310 672028 159338
rect 671620 140752 671672 140758
rect 671620 140694 671672 140700
rect 671160 139392 671212 139398
rect 671160 139334 671212 139340
rect 670240 131096 670292 131102
rect 670240 131038 670292 131044
rect 671344 130892 671396 130898
rect 671344 130834 671396 130840
rect 670148 122460 670200 122466
rect 670148 122402 670200 122408
rect 669962 117464 670018 117473
rect 669962 117399 670018 117408
rect 669228 115864 669280 115870
rect 669226 115832 669228 115841
rect 669280 115832 669282 115841
rect 669226 115767 669282 115776
rect 669226 114200 669282 114209
rect 669226 114135 669228 114144
rect 669280 114135 669282 114144
rect 669228 114106 669280 114112
rect 668872 113146 668992 113174
rect 668872 110786 668900 113146
rect 670160 112878 670188 122402
rect 670148 112872 670200 112878
rect 670148 112814 670200 112820
rect 669044 111784 669096 111790
rect 669044 111726 669096 111732
rect 669056 110945 669084 111726
rect 669042 110936 669098 110945
rect 669042 110871 669098 110880
rect 668872 110758 668992 110786
rect 668766 106040 668822 106049
rect 668766 105975 668822 105984
rect 668964 104417 668992 110758
rect 671356 109002 671384 130834
rect 671528 121440 671580 121446
rect 671528 121382 671580 121388
rect 671540 111790 671568 121382
rect 671816 120086 671844 159310
rect 672276 142154 672304 213250
rect 672460 195974 672488 213438
rect 672184 142126 672304 142154
rect 672368 195946 672488 195974
rect 672184 138038 672212 142126
rect 672172 138032 672224 138038
rect 672172 137974 672224 137980
rect 672368 129674 672396 195946
rect 672552 184890 672580 215266
rect 672828 212534 672856 303418
rect 673104 286521 673132 303826
rect 673090 286512 673146 286521
rect 673090 286447 673146 286456
rect 673288 285569 673316 305458
rect 673274 285560 673330 285569
rect 673274 285495 673330 285504
rect 673090 278760 673146 278769
rect 673090 278695 673146 278704
rect 673104 214577 673132 278695
rect 673276 262948 673328 262954
rect 673276 262890 673328 262896
rect 673288 247761 673316 262890
rect 673274 247752 673330 247761
rect 673274 247687 673330 247696
rect 673276 220992 673328 220998
rect 673276 220934 673328 220940
rect 673090 214568 673146 214577
rect 673090 214503 673146 214512
rect 673092 214124 673144 214130
rect 673092 214066 673144 214072
rect 672736 212506 672856 212534
rect 672736 205634 672764 212506
rect 672736 205606 672856 205634
rect 672540 184884 672592 184890
rect 672540 184826 672592 184832
rect 672538 183560 672594 183569
rect 672538 183495 672594 183504
rect 672552 178022 672580 183495
rect 672540 178016 672592 178022
rect 672540 177958 672592 177964
rect 672632 167068 672684 167074
rect 672632 167010 672684 167016
rect 672356 129668 672408 129674
rect 672356 129610 672408 129616
rect 671804 120080 671856 120086
rect 671804 120022 671856 120028
rect 672644 115870 672672 167010
rect 672828 133822 672856 205606
rect 673104 197810 673132 214066
rect 673288 200841 673316 220934
rect 673274 200832 673330 200841
rect 673274 200767 673330 200776
rect 673092 197804 673144 197810
rect 673092 197746 673144 197752
rect 673564 177750 673592 324294
rect 673748 215393 673776 525778
rect 674300 490113 674328 533559
rect 674470 531992 674526 532001
rect 674470 531927 674526 531936
rect 674286 490104 674342 490113
rect 674286 490039 674342 490048
rect 674484 488481 674512 531927
rect 674470 488472 674526 488481
rect 674470 488407 674526 488416
rect 674668 484401 674696 558214
rect 675128 557534 675156 589246
rect 675312 586265 675340 589246
rect 675298 586256 675354 586265
rect 675298 586191 675354 586200
rect 675482 581088 675538 581097
rect 675482 581023 675484 581032
rect 675536 581023 675538 581032
rect 675484 580994 675536 581000
rect 675298 580272 675354 580281
rect 675298 580207 675354 580216
rect 675312 579698 675340 580207
rect 675484 580032 675536 580038
rect 675484 579974 675536 579980
rect 675496 579873 675524 579974
rect 675482 579864 675538 579873
rect 675482 579799 675538 579808
rect 675300 579692 675352 579698
rect 675300 579634 675352 579640
rect 675298 579048 675354 579057
rect 675298 578983 675354 578992
rect 675312 578542 675340 578983
rect 675482 578640 675538 578649
rect 675482 578575 675538 578584
rect 675300 578536 675352 578542
rect 675300 578478 675352 578484
rect 675496 578406 675524 578575
rect 675484 578400 675536 578406
rect 675484 578342 675536 578348
rect 675482 578232 675538 578241
rect 675482 578167 675538 578176
rect 675298 577824 675354 577833
rect 675298 577759 675354 577768
rect 675312 577318 675340 577759
rect 675496 577658 675524 578167
rect 675484 577652 675536 577658
rect 675484 577594 675536 577600
rect 675482 577416 675538 577425
rect 675482 577351 675538 577360
rect 675300 577312 675352 577318
rect 675300 577254 675352 577260
rect 675496 577182 675524 577351
rect 675484 577176 675536 577182
rect 675484 577118 675536 577124
rect 675482 577008 675538 577017
rect 675482 576943 675484 576952
rect 675536 576943 675538 576952
rect 675484 576914 675536 576920
rect 675482 576600 675538 576609
rect 675482 576535 675538 576544
rect 675496 575550 675524 576535
rect 678256 575657 678284 592486
rect 682382 589248 682438 589257
rect 682382 589183 682438 589192
rect 682396 576065 682424 589183
rect 683316 576473 683344 592622
rect 683488 591456 683540 591462
rect 683488 591398 683540 591404
rect 683302 576464 683358 576473
rect 683302 576399 683358 576408
rect 682382 576056 682438 576065
rect 682382 575991 682438 576000
rect 678242 575648 678298 575657
rect 678242 575583 678298 575592
rect 675484 575544 675536 575550
rect 675484 575486 675536 575492
rect 675482 574968 675538 574977
rect 675482 574903 675538 574912
rect 675298 574560 675354 574569
rect 675298 574495 675354 574504
rect 675312 574258 675340 574495
rect 675496 574394 675524 574903
rect 675484 574388 675536 574394
rect 675484 574330 675536 574336
rect 675300 574252 675352 574258
rect 675300 574194 675352 574200
rect 675482 574152 675538 574161
rect 675482 574087 675484 574096
rect 675536 574087 675538 574096
rect 675484 574058 675536 574064
rect 675298 573744 675354 573753
rect 675298 573679 675354 573688
rect 675312 572762 675340 573679
rect 675482 572928 675538 572937
rect 675482 572863 675484 572872
rect 675536 572863 675538 572872
rect 675484 572834 675536 572840
rect 675300 572756 675352 572762
rect 675300 572698 675352 572704
rect 683500 571985 683528 591398
rect 684132 591320 684184 591326
rect 684132 591262 684184 591268
rect 684144 572801 684172 591262
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 684130 572792 684186 572801
rect 684130 572727 684186 572736
rect 683486 571976 683542 571985
rect 683486 571911 683542 571920
rect 675298 571296 675354 571305
rect 675298 571231 675300 571240
rect 675352 571231 675354 571240
rect 675300 571202 675352 571208
rect 676218 570752 676274 570761
rect 676218 570687 676274 570696
rect 675852 570104 675904 570110
rect 675496 570052 675852 570058
rect 675496 570046 675904 570052
rect 675496 570042 675892 570046
rect 675484 570036 675892 570042
rect 675536 570030 675892 570036
rect 675484 569978 675536 569984
rect 675482 569664 675538 569673
rect 675482 569599 675484 569608
rect 675536 569599 675538 569608
rect 675484 569570 675536 569576
rect 676232 565214 676260 570687
rect 683118 570344 683174 570353
rect 683118 570279 683174 570288
rect 683132 570110 683160 570279
rect 683120 570104 683172 570110
rect 683120 570046 683172 570052
rect 675852 565208 675904 565214
rect 675852 565150 675904 565156
rect 676220 565208 676272 565214
rect 676220 565150 676272 565156
rect 675300 564596 675352 564602
rect 675300 564538 675352 564544
rect 675312 564482 675340 564538
rect 675220 564454 675340 564482
rect 675484 564460 675536 564466
rect 675220 562306 675248 564454
rect 675484 564402 675536 564408
rect 675496 564346 675524 564402
rect 675312 564318 675524 564346
rect 675312 563054 675340 564318
rect 675864 563961 675892 565150
rect 675850 563952 675906 563961
rect 675850 563887 675906 563896
rect 675312 563026 675432 563054
rect 675404 562904 675432 563026
rect 675220 562278 675418 562306
rect 675390 561912 675446 561921
rect 675390 561847 675446 561856
rect 675404 561612 675432 561847
rect 675496 559473 675524 559776
rect 675482 559464 675538 559473
rect 675482 559399 675538 559408
rect 675772 559065 675800 559232
rect 675758 559056 675814 559065
rect 675758 558991 675814 559000
rect 675404 558278 675432 558620
rect 675392 558272 675444 558278
rect 675392 558214 675444 558220
rect 675312 557926 675418 557954
rect 675312 557734 675340 557926
rect 675300 557728 675352 557734
rect 675300 557670 675352 557676
rect 675300 557592 675352 557598
rect 675300 557534 675352 557540
rect 674944 557506 675156 557534
rect 674944 547641 674972 557506
rect 675312 555370 675340 557534
rect 675404 555370 675432 555492
rect 675312 555342 675432 555370
rect 675128 554905 675418 554933
rect 675128 554810 675156 554905
rect 675116 554804 675168 554810
rect 675116 554746 675168 554752
rect 675128 554254 675418 554282
rect 675128 554198 675156 554254
rect 675116 554192 675168 554198
rect 675116 554134 675168 554140
rect 675116 554056 675168 554062
rect 675116 553998 675168 554004
rect 675128 551253 675156 553998
rect 675404 553489 675432 553656
rect 675390 553480 675446 553489
rect 675390 553415 675446 553424
rect 675772 552129 675800 552432
rect 675758 552120 675814 552129
rect 675758 552055 675814 552064
rect 675128 551225 675418 551253
rect 675128 550582 675418 550610
rect 675128 547890 675156 550582
rect 675312 549937 675418 549965
rect 675312 549778 675340 549937
rect 675300 549772 675352 549778
rect 675300 549714 675352 549720
rect 675482 549672 675538 549681
rect 675312 549630 675482 549658
rect 675128 547862 675248 547890
rect 674930 547632 674986 547641
rect 674930 547567 674986 547576
rect 675024 545488 675076 545494
rect 675024 545430 675076 545436
rect 675036 540974 675064 545430
rect 675036 540946 675156 540974
rect 674932 534608 674984 534614
rect 674932 534550 674984 534556
rect 674944 534041 674972 534550
rect 674930 534032 674986 534041
rect 674930 533967 674986 533976
rect 674930 531176 674986 531185
rect 674930 531111 674986 531120
rect 674944 529990 674972 531111
rect 674932 529984 674984 529990
rect 674932 529926 674984 529932
rect 675128 524414 675156 540946
rect 674944 524386 675156 524414
rect 674654 484392 674710 484401
rect 674654 484327 674710 484336
rect 674104 481908 674156 481914
rect 674104 481850 674156 481856
rect 673920 395684 673972 395690
rect 673920 395626 673972 395632
rect 673932 376825 673960 395626
rect 673918 376816 673974 376825
rect 673918 376751 673974 376760
rect 673920 357060 673972 357066
rect 673920 357002 673972 357008
rect 673932 312526 673960 357002
rect 673920 312520 673972 312526
rect 673920 312462 673972 312468
rect 673918 249656 673974 249665
rect 673918 249591 673974 249600
rect 673932 215665 673960 249591
rect 673918 215656 673974 215665
rect 673918 215591 673974 215600
rect 673920 215484 673972 215490
rect 673920 215426 673972 215432
rect 673734 215384 673790 215393
rect 673734 215319 673790 215328
rect 673736 215212 673788 215218
rect 673736 215154 673788 215160
rect 673748 200802 673776 215154
rect 673932 201482 673960 215426
rect 673920 201476 673972 201482
rect 673920 201418 673972 201424
rect 673736 200796 673788 200802
rect 673736 200738 673788 200744
rect 673552 177744 673604 177750
rect 673552 177686 673604 177692
rect 673920 176860 673972 176866
rect 673920 176802 673972 176808
rect 673368 175228 673420 175234
rect 673368 175170 673420 175176
rect 673000 174412 673052 174418
rect 673000 174354 673052 174360
rect 672816 133816 672868 133822
rect 672816 133758 672868 133764
rect 673012 129742 673040 174354
rect 673184 168700 673236 168706
rect 673184 168642 673236 168648
rect 673196 151774 673224 168642
rect 673184 151768 673236 151774
rect 673184 151710 673236 151716
rect 673380 130558 673408 175170
rect 673552 162104 673604 162110
rect 673552 162046 673604 162052
rect 673564 155854 673592 162046
rect 673552 155848 673604 155854
rect 673552 155790 673604 155796
rect 673932 132190 673960 176802
rect 674116 148238 674144 481850
rect 674944 481545 674972 524386
rect 675220 511994 675248 547862
rect 675128 511966 675248 511994
rect 675128 508881 675156 511966
rect 675114 508872 675170 508881
rect 675114 508807 675170 508816
rect 675312 500313 675340 549630
rect 675482 549607 675538 549616
rect 675496 548457 675524 548760
rect 675482 548448 675538 548457
rect 675482 548383 675538 548392
rect 675758 547904 675814 547913
rect 675758 547839 675814 547848
rect 675482 536072 675538 536081
rect 675482 536007 675538 536016
rect 675496 535702 675524 536007
rect 675484 535696 675536 535702
rect 675484 535638 675536 535644
rect 675482 535528 675538 535537
rect 675482 535463 675484 535472
rect 675536 535463 675538 535472
rect 675484 535434 675536 535440
rect 675482 534848 675538 534857
rect 675482 534783 675538 534792
rect 675496 534478 675524 534783
rect 675484 534472 675536 534478
rect 675484 534414 675536 534420
rect 675482 534304 675538 534313
rect 675482 534239 675538 534248
rect 675496 534138 675524 534239
rect 675484 534132 675536 534138
rect 675484 534074 675536 534080
rect 675484 533384 675536 533390
rect 675482 533352 675484 533361
rect 675536 533352 675538 533361
rect 675482 533287 675538 533296
rect 675482 532808 675538 532817
rect 675482 532743 675484 532752
rect 675536 532743 675538 532752
rect 675484 532714 675536 532720
rect 675484 532568 675536 532574
rect 675482 532536 675484 532545
rect 675536 532536 675538 532545
rect 675482 532471 675538 532480
rect 675482 531584 675538 531593
rect 675482 531519 675538 531528
rect 675496 531418 675524 531519
rect 675484 531412 675536 531418
rect 675484 531354 675536 531360
rect 675484 530120 675536 530126
rect 675482 530088 675484 530097
rect 675536 530088 675538 530097
rect 675482 530023 675538 530032
rect 675482 529544 675538 529553
rect 675482 529479 675538 529488
rect 675496 528630 675524 529479
rect 675484 528624 675536 528630
rect 675484 528566 675536 528572
rect 675484 528488 675536 528494
rect 675482 528456 675484 528465
rect 675536 528456 675538 528465
rect 675482 528391 675538 528400
rect 675484 528080 675536 528086
rect 675482 528048 675484 528057
rect 675536 528048 675538 528057
rect 675482 527983 675538 527992
rect 675484 526856 675536 526862
rect 675482 526824 675484 526833
rect 675536 526824 675538 526833
rect 675482 526759 675538 526768
rect 675484 526448 675536 526454
rect 675482 526416 675484 526425
rect 675536 526416 675538 526425
rect 675482 526351 675538 526360
rect 675482 525872 675538 525881
rect 675482 525807 675484 525816
rect 675536 525807 675538 525816
rect 675484 525778 675536 525784
rect 675772 505094 675800 547839
rect 675942 547632 675998 547641
rect 675942 547567 675998 547576
rect 677506 547632 677562 547641
rect 677506 547567 677562 547576
rect 675956 546854 675984 547567
rect 676126 547360 676182 547369
rect 676126 547295 676182 547304
rect 675944 546848 675996 546854
rect 675944 546790 675996 546796
rect 676140 545766 676168 547295
rect 676128 545760 676180 545766
rect 676128 545702 676180 545708
rect 677520 529417 677548 547567
rect 683394 547088 683450 547097
rect 683394 547023 683450 547032
rect 681004 546848 681056 546854
rect 679622 546816 679678 546825
rect 681004 546790 681056 546796
rect 679622 546751 679678 546760
rect 679636 530641 679664 546751
rect 679622 530632 679678 530641
rect 679622 530567 679678 530576
rect 677506 529408 677562 529417
rect 677506 529343 677562 529352
rect 681016 525774 681044 546790
rect 683212 545760 683264 545766
rect 683212 545702 683264 545708
rect 683224 529009 683252 545702
rect 683408 531049 683436 547023
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683394 531040 683450 531049
rect 683394 530975 683450 530984
rect 683210 529000 683266 529009
rect 683210 528935 683266 528944
rect 681004 525768 681056 525774
rect 683120 525768 683172 525774
rect 681004 525710 681056 525716
rect 683118 525736 683120 525745
rect 683172 525736 683174 525745
rect 683118 525671 683174 525680
rect 676034 508872 676090 508881
rect 676034 508807 676090 508816
rect 675772 505066 675892 505094
rect 675298 500304 675354 500313
rect 675298 500239 675354 500248
rect 675298 492144 675354 492153
rect 675298 492079 675354 492088
rect 675312 491638 675340 492079
rect 675482 491736 675538 491745
rect 675482 491671 675538 491680
rect 675300 491632 675352 491638
rect 675300 491574 675352 491580
rect 675496 491502 675524 491671
rect 675484 491496 675536 491502
rect 675484 491438 675536 491444
rect 675484 491360 675536 491366
rect 675482 491328 675484 491337
rect 675536 491328 675538 491337
rect 675482 491263 675538 491272
rect 675482 490920 675538 490929
rect 675482 490855 675538 490864
rect 675496 490074 675524 490855
rect 675484 490068 675536 490074
rect 675484 490010 675536 490016
rect 675482 489288 675538 489297
rect 675482 489223 675538 489232
rect 675496 488714 675524 489223
rect 675666 488880 675722 488889
rect 675666 488815 675722 488824
rect 675484 488708 675536 488714
rect 675484 488650 675536 488656
rect 675298 486840 675354 486849
rect 675298 486775 675354 486784
rect 675312 485858 675340 486775
rect 675482 486024 675538 486033
rect 675482 485959 675484 485968
rect 675536 485959 675538 485968
rect 675484 485930 675536 485936
rect 675300 485852 675352 485858
rect 675300 485794 675352 485800
rect 675680 485774 675708 488815
rect 675864 487665 675892 505066
rect 676048 503538 676076 508807
rect 676036 503532 676088 503538
rect 676036 503474 676088 503480
rect 679624 503532 679676 503538
rect 679624 503474 679676 503480
rect 676034 500304 676090 500313
rect 676034 500239 676090 500248
rect 676048 498302 676076 500239
rect 676036 498296 676088 498302
rect 676036 498238 676088 498244
rect 676034 490512 676090 490521
rect 676090 490470 676260 490498
rect 676034 490447 676090 490456
rect 676232 490210 676260 490470
rect 676220 490204 676272 490210
rect 676220 490146 676272 490152
rect 677416 490204 677468 490210
rect 677416 490146 677468 490152
rect 676034 489696 676090 489705
rect 676090 489654 676260 489682
rect 676034 489631 676090 489640
rect 676232 488578 676260 489654
rect 676220 488572 676272 488578
rect 676220 488514 676272 488520
rect 677232 488572 677284 488578
rect 677232 488514 677284 488520
rect 676034 488064 676090 488073
rect 676034 487999 676090 488008
rect 675850 487656 675906 487665
rect 675850 487591 675906 487600
rect 675680 485746 675984 485774
rect 675484 485648 675536 485654
rect 675482 485616 675484 485625
rect 675536 485616 675538 485625
rect 675482 485551 675538 485560
rect 675482 485208 675538 485217
rect 675482 485143 675538 485152
rect 675496 484430 675524 485143
rect 675484 484424 675536 484430
rect 675484 484366 675536 484372
rect 675484 483608 675536 483614
rect 675482 483576 675484 483585
rect 675536 483576 675538 483585
rect 675482 483511 675538 483520
rect 675484 483200 675536 483206
rect 675482 483168 675484 483177
rect 675536 483168 675538 483177
rect 675482 483103 675538 483112
rect 675484 482792 675536 482798
rect 675482 482760 675484 482769
rect 675536 482760 675538 482769
rect 675482 482695 675538 482704
rect 675484 482384 675536 482390
rect 675482 482352 675484 482361
rect 675536 482352 675538 482361
rect 675482 482287 675538 482296
rect 675482 481944 675538 481953
rect 675482 481879 675484 481888
rect 675536 481879 675538 481888
rect 675484 481850 675536 481856
rect 674930 481536 674986 481545
rect 674930 481471 674986 481480
rect 675482 480720 675538 480729
rect 675482 480655 675484 480664
rect 675536 480655 675538 480664
rect 675484 480626 675536 480632
rect 675482 403880 675538 403889
rect 675482 403815 675538 403824
rect 675298 403472 675354 403481
rect 675298 403407 675300 403416
rect 675352 403407 675354 403416
rect 675300 403378 675352 403384
rect 675496 403306 675524 403815
rect 675484 403300 675536 403306
rect 675484 403242 675536 403248
rect 675484 403096 675536 403102
rect 675482 403064 675484 403073
rect 675536 403064 675538 403073
rect 675482 402999 675538 403008
rect 674654 402248 674710 402257
rect 674654 402183 674710 402192
rect 674470 401432 674526 401441
rect 674470 401367 674526 401376
rect 674286 393680 674342 393689
rect 674286 393615 674342 393624
rect 674104 148232 674156 148238
rect 674104 148174 674156 148180
rect 674300 144226 674328 393615
rect 674484 356697 674512 401367
rect 674668 357513 674696 402183
rect 675956 401033 675984 485746
rect 676048 470594 676076 487999
rect 676048 470566 676168 470594
rect 676140 412634 676168 470566
rect 676048 412606 676168 412634
rect 676048 408494 676076 412606
rect 676048 408466 676168 408494
rect 675942 401024 675998 401033
rect 675942 400959 675998 400968
rect 676140 400874 676168 408466
rect 677244 402121 677272 488514
rect 677428 402937 677456 490146
rect 679636 487257 679664 503474
rect 679808 498296 679860 498302
rect 679808 498238 679860 498244
rect 679622 487248 679678 487257
rect 679622 487183 679678 487192
rect 679820 486441 679848 498238
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 679806 486432 679862 486441
rect 679806 486367 679862 486376
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 677414 402928 677470 402937
rect 677414 402863 677470 402872
rect 677230 402112 677286 402121
rect 677230 402047 677286 402056
rect 675956 400846 676168 400874
rect 675482 400616 675538 400625
rect 675482 400551 675484 400560
rect 675536 400551 675538 400560
rect 675484 400522 675536 400528
rect 675956 400217 675984 400846
rect 675942 400208 675998 400217
rect 675942 400143 675998 400152
rect 675482 399800 675538 399809
rect 675482 399735 675484 399744
rect 675536 399735 675538 399744
rect 675484 399706 675536 399712
rect 674930 399392 674986 399401
rect 674930 399327 674986 399336
rect 674944 384810 674972 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675114 398168 675170 398177
rect 675114 398103 675170 398112
rect 674932 384804 674984 384810
rect 674932 384746 674984 384752
rect 675128 382582 675156 398103
rect 675482 397352 675538 397361
rect 675482 397287 675484 397296
rect 675536 397287 675538 397296
rect 675484 397258 675536 397264
rect 675482 396128 675538 396137
rect 675482 396063 675484 396072
rect 675536 396063 675538 396072
rect 675484 396034 675536 396040
rect 675482 395720 675538 395729
rect 675482 395655 675484 395664
rect 675536 395655 675538 395664
rect 675484 395626 675536 395632
rect 676232 394754 676260 398375
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 675312 394726 676260 394754
rect 675312 386186 675340 394726
rect 675482 394496 675538 394505
rect 675482 394431 675484 394440
rect 675536 394431 675538 394440
rect 675484 394402 675536 394408
rect 675482 394088 675538 394097
rect 675482 394023 675484 394032
rect 675536 394023 675538 394032
rect 675484 393994 675536 394000
rect 675482 392456 675538 392465
rect 675482 392391 675484 392400
rect 675536 392391 675538 392400
rect 675484 392362 675536 392368
rect 675852 392148 675904 392154
rect 675852 392090 675904 392096
rect 675864 389337 675892 392090
rect 675850 389328 675906 389337
rect 675850 389263 675906 389272
rect 681016 388521 681044 397559
rect 681186 396400 681242 396409
rect 681186 396335 681242 396344
rect 681002 388512 681058 388521
rect 681002 388447 681058 388456
rect 681200 387705 681228 396335
rect 683118 392728 683174 392737
rect 683118 392663 683174 392672
rect 683132 392154 683160 392663
rect 683120 392148 683172 392154
rect 683120 392090 683172 392096
rect 681186 387696 681242 387705
rect 681186 387631 681242 387640
rect 675312 386158 675432 386186
rect 675404 385696 675432 386158
rect 675312 385070 675418 385098
rect 675312 383625 675340 385070
rect 675484 384804 675536 384810
rect 675484 384746 675536 384752
rect 675496 384435 675524 384746
rect 675298 383616 675354 383625
rect 675298 383551 675354 383560
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675128 382554 675340 382582
rect 675404 382568 675432 382622
rect 675758 382256 675814 382265
rect 675758 382191 675814 382200
rect 675772 382024 675800 382191
rect 675128 381398 675418 381426
rect 675128 379506 675156 381398
rect 675772 380633 675800 380732
rect 675758 380624 675814 380633
rect 675758 380559 675814 380568
rect 675116 379500 675168 379506
rect 675116 379442 675168 379448
rect 675666 378584 675722 378593
rect 675666 378519 675722 378528
rect 675680 378284 675708 378519
rect 675300 377868 675352 377874
rect 675300 377810 675352 377816
rect 675312 377618 675340 377810
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 674930 376816 674986 376825
rect 674930 376751 674986 376760
rect 674944 375238 674972 376751
rect 675116 376644 675168 376650
rect 675116 376586 675168 376592
rect 675128 376462 675156 376586
rect 675128 376434 675340 376462
rect 675312 376394 675340 376434
rect 675404 376394 675432 376448
rect 675312 376366 675432 376394
rect 674944 375210 675418 375238
rect 675298 375048 675354 375057
rect 675298 374983 675354 374992
rect 675312 373402 675340 374983
rect 675312 373374 675418 373402
rect 675114 372600 675170 372609
rect 675404 372586 675432 372776
rect 675312 372570 675432 372586
rect 675114 372535 675170 372544
rect 675300 372564 675432 372570
rect 675128 371566 675156 372535
rect 675352 372558 675432 372564
rect 675300 372506 675352 372512
rect 675128 371538 675418 371566
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675298 358728 675354 358737
rect 675298 358663 675354 358672
rect 675114 358320 675170 358329
rect 675114 358255 675170 358264
rect 674654 357504 674710 357513
rect 675128 357474 675156 358255
rect 675312 357882 675340 358663
rect 675482 357912 675538 357921
rect 675300 357876 675352 357882
rect 675482 357847 675538 357856
rect 675300 357818 675352 357824
rect 675496 357610 675524 357847
rect 675484 357604 675536 357610
rect 675484 357546 675536 357552
rect 674654 357439 674710 357448
rect 675116 357468 675168 357474
rect 675116 357410 675168 357416
rect 675482 357096 675538 357105
rect 675482 357031 675484 357040
rect 675536 357031 675538 357040
rect 675484 357002 675536 357008
rect 674470 356688 674526 356697
rect 674470 356623 674526 356632
rect 674654 356280 674710 356289
rect 674654 356215 674710 356224
rect 674470 351384 674526 351393
rect 674470 351319 674526 351328
rect 674484 337958 674512 351319
rect 674472 337952 674524 337958
rect 674472 337894 674524 337900
rect 674668 311681 674696 356215
rect 675484 355904 675536 355910
rect 675482 355872 675484 355881
rect 675536 355872 675538 355881
rect 675482 355807 675538 355816
rect 675482 355464 675538 355473
rect 675482 355399 675484 355408
rect 675536 355399 675538 355408
rect 675484 355370 675536 355376
rect 675484 355088 675536 355094
rect 675482 355056 675484 355065
rect 675536 355056 675538 355065
rect 675482 354991 675538 355000
rect 675482 354648 675538 354657
rect 675482 354583 675484 354592
rect 675536 354583 675538 354592
rect 675484 354554 675536 354560
rect 675482 353832 675538 353841
rect 675482 353767 675538 353776
rect 675496 353666 675524 353767
rect 675484 353660 675536 353666
rect 675484 353602 675536 353608
rect 675482 353424 675538 353433
rect 675482 353359 675484 353368
rect 675536 353359 675538 353368
rect 675484 353330 675536 353336
rect 675482 352608 675538 352617
rect 675482 352543 675484 352552
rect 675536 352543 675538 352552
rect 675484 352514 675536 352520
rect 676034 350976 676090 350985
rect 676034 350911 676090 350920
rect 675850 350568 675906 350577
rect 675850 350503 675906 350512
rect 675482 350160 675538 350169
rect 675482 350095 675484 350104
rect 675536 350095 675538 350104
rect 675484 350066 675536 350072
rect 675482 349752 675538 349761
rect 675482 349687 675484 349696
rect 675536 349687 675538 349696
rect 675484 349658 675536 349664
rect 675482 349344 675538 349353
rect 675482 349279 675484 349288
rect 675536 349279 675538 349288
rect 675484 349250 675536 349256
rect 675482 348936 675538 348945
rect 675482 348871 675484 348880
rect 675536 348871 675538 348880
rect 675484 348842 675536 348848
rect 675482 348528 675538 348537
rect 675482 348463 675484 348472
rect 675536 348463 675538 348472
rect 675484 348434 675536 348440
rect 675864 347954 675892 350503
rect 675852 347948 675904 347954
rect 675852 347890 675904 347896
rect 675482 347304 675538 347313
rect 675482 347239 675484 347248
rect 675536 347239 675538 347248
rect 675484 347210 675536 347216
rect 676048 346633 676076 350911
rect 676588 347948 676640 347954
rect 676588 347890 676640 347896
rect 676034 346624 676090 346633
rect 676034 346559 676090 346568
rect 676600 346497 676628 347890
rect 683118 347712 683174 347721
rect 683118 347647 683174 347656
rect 676586 346488 676642 346497
rect 675852 346452 675904 346458
rect 683132 346458 683160 347647
rect 676586 346423 676642 346432
rect 683120 346452 683172 346458
rect 675852 346394 675904 346400
rect 683120 346394 683172 346400
rect 675864 342281 675892 346394
rect 675850 342272 675906 342281
rect 675850 342207 675906 342216
rect 675128 340530 675340 340558
rect 675128 338094 675156 340530
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340232 675814 340241
rect 675758 340167 675814 340176
rect 675772 339864 675800 340167
rect 675404 339017 675432 339252
rect 675390 339008 675446 339017
rect 675390 338943 675446 338952
rect 675116 338088 675168 338094
rect 675116 338030 675168 338036
rect 675116 337952 675168 337958
rect 675116 337894 675168 337900
rect 675128 336857 675156 337894
rect 675666 337784 675722 337793
rect 675666 337719 675722 337728
rect 675680 337416 675708 337719
rect 675128 336829 675418 336857
rect 675312 336178 675418 336206
rect 674932 336048 674984 336054
rect 675312 336002 675340 336178
rect 674932 335990 674984 335996
rect 674944 331889 674972 335990
rect 675220 335974 675340 336002
rect 675220 335354 675248 335974
rect 675392 335912 675444 335918
rect 675444 335860 675524 335866
rect 675392 335854 675524 335860
rect 675404 335838 675524 335854
rect 675496 335580 675524 335838
rect 675220 335345 675340 335354
rect 675220 335336 675354 335345
rect 675220 335326 675298 335336
rect 675298 335271 675354 335280
rect 675116 333940 675168 333946
rect 675116 333882 675168 333888
rect 675128 333078 675156 333882
rect 675128 333050 675418 333078
rect 675116 332648 675168 332654
rect 675116 332590 675168 332596
rect 675128 332534 675156 332590
rect 675128 332506 675418 332534
rect 674944 331861 675418 331889
rect 675116 331764 675168 331770
rect 675116 331706 675168 331712
rect 675128 331242 675156 331706
rect 675128 331214 675418 331242
rect 675298 331120 675354 331129
rect 675298 331055 675354 331064
rect 675312 330049 675340 331055
rect 675312 330021 675418 330049
rect 675312 328222 675432 328250
rect 675312 328182 675340 328222
rect 674944 328154 675340 328182
rect 675404 328168 675432 328222
rect 674944 325514 674972 328154
rect 675128 327542 675418 327570
rect 675128 325650 675156 327542
rect 675758 326904 675814 326913
rect 675758 326839 675814 326848
rect 675772 326332 675800 326839
rect 675116 325644 675168 325650
rect 675116 325586 675168 325592
rect 674932 325508 674984 325514
rect 674932 325450 674984 325456
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 675482 313712 675538 313721
rect 675482 313647 675538 313656
rect 675496 313478 675524 313647
rect 675484 313472 675536 313478
rect 675484 313414 675536 313420
rect 675484 313336 675536 313342
rect 675482 313304 675484 313313
rect 675536 313304 675538 313313
rect 675482 313239 675538 313248
rect 675298 312896 675354 312905
rect 675298 312831 675354 312840
rect 675312 312050 675340 312831
rect 675484 312520 675536 312526
rect 675482 312488 675484 312497
rect 675536 312488 675538 312497
rect 675482 312423 675538 312432
rect 675482 312080 675538 312089
rect 675300 312044 675352 312050
rect 675482 312015 675538 312024
rect 675300 311986 675352 311992
rect 675496 311914 675524 312015
rect 675484 311908 675536 311914
rect 675484 311850 675536 311856
rect 674654 311672 674710 311681
rect 674654 311607 674710 311616
rect 675482 311264 675538 311273
rect 675482 311199 675538 311208
rect 675496 310758 675524 311199
rect 675484 310752 675536 310758
rect 675484 310694 675536 310700
rect 675482 310448 675538 310457
rect 675482 310383 675484 310392
rect 675536 310383 675538 310392
rect 675484 310354 675536 310360
rect 675484 310072 675536 310078
rect 675482 310040 675484 310049
rect 675536 310040 675538 310049
rect 675482 309975 675538 309984
rect 675482 309632 675538 309641
rect 675482 309567 675538 309576
rect 675206 309224 675262 309233
rect 675496 309194 675524 309567
rect 675206 309159 675262 309168
rect 675484 309188 675536 309194
rect 675022 308000 675078 308009
rect 675022 307935 675078 307944
rect 674838 307592 674894 307601
rect 674838 307527 674894 307536
rect 674470 306368 674526 306377
rect 674470 306303 674526 306312
rect 674484 292330 674512 306303
rect 674654 304328 674710 304337
rect 674654 304263 674710 304272
rect 674472 292324 674524 292330
rect 674472 292266 674524 292272
rect 674668 287518 674696 304263
rect 674852 302234 674880 307527
rect 674852 302206 674972 302234
rect 674944 288062 674972 302206
rect 675036 292414 675064 307935
rect 675220 302234 675248 309159
rect 675484 309130 675536 309136
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 675482 305552 675538 305561
rect 675482 305487 675484 305496
rect 675536 305487 675538 305496
rect 675484 305458 675536 305464
rect 676232 305266 676260 308366
rect 678242 307184 678298 307193
rect 678242 307119 678298 307128
rect 675680 305238 676260 305266
rect 675482 303920 675538 303929
rect 675482 303855 675484 303864
rect 675536 303855 675538 303864
rect 675484 303826 675536 303832
rect 675482 303512 675538 303521
rect 675482 303447 675484 303456
rect 675536 303447 675538 303456
rect 675484 303418 675536 303424
rect 675128 302206 675248 302234
rect 675482 302288 675538 302297
rect 675482 302223 675484 302232
rect 675128 294250 675156 302206
rect 675536 302223 675538 302232
rect 675484 302194 675536 302200
rect 675680 299474 675708 305238
rect 675850 305144 675906 305153
rect 675850 305079 675906 305088
rect 675864 301617 675892 305079
rect 676034 304736 676090 304745
rect 676034 304671 676090 304680
rect 676048 302977 676076 304671
rect 676034 302968 676090 302977
rect 676034 302903 676090 302912
rect 675850 301608 675906 301617
rect 675850 301543 675906 301552
rect 675496 299446 675708 299474
rect 675496 296410 675524 299446
rect 678256 297401 678284 307119
rect 681002 306776 681058 306785
rect 681002 306711 681058 306720
rect 680360 302252 680412 302258
rect 680360 302194 680412 302200
rect 680372 299441 680400 302194
rect 680358 299432 680414 299441
rect 680358 299367 680414 299376
rect 678242 297392 678298 297401
rect 678242 297327 678298 297336
rect 681016 296954 681044 306711
rect 683118 302696 683174 302705
rect 683118 302631 683174 302640
rect 683132 302258 683160 302631
rect 683120 302252 683172 302258
rect 683120 302194 683172 302200
rect 675852 296948 675904 296954
rect 675852 296890 675904 296896
rect 681004 296948 681056 296954
rect 681004 296890 681056 296896
rect 675864 296562 675892 296890
rect 675680 296534 675892 296562
rect 675484 296404 675536 296410
rect 675484 296346 675536 296352
rect 675680 296290 675708 296534
rect 675220 296262 675708 296290
rect 675220 294893 675248 296262
rect 675484 295928 675536 295934
rect 675484 295870 675536 295876
rect 675496 295528 675524 295870
rect 675220 294865 675418 294893
rect 675128 294222 675418 294250
rect 675036 292386 675418 292414
rect 675116 292324 675168 292330
rect 675116 292266 675168 292272
rect 675128 291870 675156 292266
rect 675128 291842 675418 291870
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675758 291000 675814 291009
rect 675758 290935 675814 290944
rect 675772 290564 675800 290935
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674944 288034 675340 288062
rect 675404 288048 675432 288102
rect 674668 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 675298 268696 675354 268705
rect 675298 268631 675354 268640
rect 675312 268190 675340 268631
rect 675482 268288 675538 268297
rect 675482 268223 675538 268232
rect 675300 268184 675352 268190
rect 675300 268126 675352 268132
rect 675496 268054 675524 268223
rect 675484 268048 675536 268054
rect 675484 267990 675536 267996
rect 675482 267880 675538 267889
rect 675482 267815 675484 267824
rect 675536 267815 675538 267824
rect 675484 267786 675536 267792
rect 675114 267472 675170 267481
rect 675114 267407 675170 267416
rect 675128 266558 675156 267407
rect 675298 267064 675354 267073
rect 675298 266999 675354 267008
rect 675116 266552 675168 266558
rect 675116 266494 675168 266500
rect 675312 266422 675340 266999
rect 675484 266688 675536 266694
rect 675482 266656 675484 266665
rect 675536 266656 675538 266665
rect 675482 266591 675538 266600
rect 675300 266416 675352 266422
rect 675300 266358 675352 266364
rect 675482 266248 675538 266257
rect 675482 266183 675538 266192
rect 675300 265872 675352 265878
rect 675298 265840 675300 265849
rect 675352 265840 675354 265849
rect 675298 265775 675354 265784
rect 675496 265606 675524 266183
rect 675484 265600 675536 265606
rect 675484 265542 675536 265548
rect 675482 265432 675538 265441
rect 675482 265367 675538 265376
rect 675496 265266 675524 265367
rect 675484 265260 675536 265266
rect 675484 265202 675536 265208
rect 675484 265056 675536 265062
rect 675482 265024 675484 265033
rect 675536 265024 675538 265033
rect 675482 264959 675538 264968
rect 675482 264616 675538 264625
rect 675482 264551 675538 264560
rect 675022 264208 675078 264217
rect 675022 264143 675078 264152
rect 674470 262168 674526 262177
rect 674470 262103 674526 262112
rect 674484 247042 674512 262103
rect 674654 258904 674710 258913
rect 674654 258839 674710 258848
rect 674472 247036 674524 247042
rect 674472 246978 674524 246984
rect 674668 241466 674696 258839
rect 674838 254008 674894 254017
rect 674838 253943 674894 253952
rect 674852 247194 674880 253943
rect 675036 249778 675064 264143
rect 675496 263634 675524 264551
rect 675484 263628 675536 263634
rect 675484 263570 675536 263576
rect 676218 263256 676274 263265
rect 676218 263191 676274 263200
rect 675482 262984 675538 262993
rect 675482 262919 675484 262928
rect 675536 262919 675538 262928
rect 675484 262890 675536 262896
rect 675482 261352 675538 261361
rect 675482 261287 675484 261296
rect 675536 261287 675538 261296
rect 675484 261258 675536 261264
rect 675666 260536 675722 260545
rect 675666 260471 675722 260480
rect 675482 260128 675538 260137
rect 675482 260063 675538 260072
rect 675496 259758 675524 260063
rect 675484 259752 675536 259758
rect 675298 259720 675354 259729
rect 675484 259694 675536 259700
rect 675298 259655 675354 259664
rect 675312 259486 675340 259655
rect 675484 259616 675536 259622
rect 675680 259570 675708 260471
rect 676232 259570 676260 263191
rect 681002 262440 681058 262449
rect 681002 262375 681058 262384
rect 675536 259564 675708 259570
rect 675484 259558 675708 259564
rect 675496 259542 675708 259558
rect 675772 259542 676260 259570
rect 675300 259480 675352 259486
rect 675300 259422 675352 259428
rect 675482 259312 675538 259321
rect 675482 259247 675484 259256
rect 675536 259247 675538 259256
rect 675484 259218 675536 259224
rect 675482 258496 675538 258505
rect 675482 258431 675484 258440
rect 675536 258431 675538 258440
rect 675484 258402 675536 258408
rect 675482 257272 675538 257281
rect 675482 257207 675538 257216
rect 675496 256630 675524 257207
rect 675484 256624 675536 256630
rect 675484 256566 675536 256572
rect 675772 253934 675800 259542
rect 675944 256760 675996 256766
rect 675944 256702 675996 256708
rect 675956 254017 675984 256702
rect 675942 254008 675998 254017
rect 675942 253943 675998 253952
rect 675220 253906 675800 253934
rect 675220 250526 675248 253906
rect 681016 252657 681044 262375
rect 683118 257544 683174 257553
rect 683118 257479 683174 257488
rect 683132 256766 683160 257479
rect 683120 256760 683172 256766
rect 683120 256702 683172 256708
rect 681002 252648 681058 252657
rect 681002 252583 681058 252592
rect 675220 250498 675418 250526
rect 675758 250200 675814 250209
rect 675758 250135 675814 250144
rect 675772 249900 675800 250135
rect 675036 249750 675524 249778
rect 675114 249656 675170 249665
rect 675114 249591 675170 249600
rect 675298 249656 675354 249665
rect 675298 249591 675354 249600
rect 675128 249506 675156 249591
rect 675128 249478 675248 249506
rect 674852 247166 675064 247194
rect 674840 247036 674892 247042
rect 674840 246978 674892 246984
rect 674656 241460 674708 241466
rect 674656 241402 674708 241408
rect 674852 236382 674880 246978
rect 675036 246922 675064 247166
rect 674944 246894 675064 246922
rect 674944 237266 674972 246894
rect 675220 243522 675248 249478
rect 675312 245970 675340 249591
rect 675496 249220 675524 249750
rect 675482 247752 675538 247761
rect 675482 247687 675538 247696
rect 675496 247384 675524 247687
rect 675482 247072 675538 247081
rect 675482 247007 675538 247016
rect 675496 246840 675524 247007
rect 675758 246664 675814 246673
rect 675758 246599 675814 246608
rect 675772 246199 675800 246599
rect 675482 245984 675538 245993
rect 675312 245942 675482 245970
rect 675482 245919 675538 245928
rect 675404 245206 675432 245548
rect 675392 245200 675444 245206
rect 675392 245142 675444 245148
rect 675220 243494 675432 243522
rect 675404 243071 675432 243494
rect 675116 242888 675168 242894
rect 675116 242830 675168 242836
rect 675128 242533 675156 242830
rect 675128 242505 675418 242533
rect 675128 241862 675418 241890
rect 675128 241738 675156 241862
rect 675116 241732 675168 241738
rect 675116 241674 675168 241680
rect 675116 241460 675168 241466
rect 675116 241402 675168 241408
rect 675128 241245 675156 241402
rect 675128 241217 675418 241245
rect 675220 240026 675418 240054
rect 675220 237674 675248 240026
rect 675390 238640 675446 238649
rect 675390 238575 675446 238584
rect 675404 238204 675432 238575
rect 675220 237646 675340 237674
rect 675312 237386 675340 237646
rect 675300 237380 675352 237386
rect 675300 237322 675352 237328
rect 675496 237266 675524 237524
rect 674944 237238 675524 237266
rect 674852 236354 675418 236382
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 675114 223544 675170 223553
rect 675114 223479 675170 223488
rect 675128 222698 675156 223479
rect 675482 223136 675538 223145
rect 675482 223071 675538 223080
rect 675298 222728 675354 222737
rect 675116 222692 675168 222698
rect 675298 222663 675354 222672
rect 675116 222634 675168 222640
rect 675312 222426 675340 222663
rect 675496 222562 675524 223071
rect 675484 222556 675536 222562
rect 675484 222498 675536 222504
rect 675300 222420 675352 222426
rect 675300 222362 675352 222368
rect 675482 222320 675538 222329
rect 675482 222255 675484 222264
rect 675536 222255 675538 222264
rect 675484 222226 675536 222232
rect 675114 221912 675170 221921
rect 675114 221847 675170 221856
rect 675128 220998 675156 221847
rect 675482 221504 675538 221513
rect 675482 221439 675538 221448
rect 675496 221134 675524 221439
rect 675484 221128 675536 221134
rect 675298 221096 675354 221105
rect 675484 221070 675536 221076
rect 675298 221031 675354 221040
rect 675116 220992 675168 220998
rect 675116 220934 675168 220940
rect 675312 220862 675340 221031
rect 675300 220856 675352 220862
rect 675300 220798 675352 220804
rect 675298 220688 675354 220697
rect 675298 220623 675354 220632
rect 674654 220280 674710 220289
rect 674654 220215 674710 220224
rect 674470 219464 674526 219473
rect 674470 219399 674526 219408
rect 674484 198665 674512 219399
rect 674470 198656 674526 198665
rect 674470 198591 674526 198600
rect 674470 176080 674526 176089
rect 674470 176015 674526 176024
rect 674484 172122 674512 176015
rect 674668 175681 674696 220215
rect 675312 219774 675340 220623
rect 675482 219872 675538 219881
rect 675482 219807 675538 219816
rect 675300 219768 675352 219774
rect 675300 219710 675352 219716
rect 675496 219638 675524 219807
rect 675484 219632 675536 219638
rect 675484 219574 675536 219580
rect 674838 218240 674894 218249
rect 674838 218175 674894 218184
rect 674852 205766 674880 218175
rect 675298 217424 675354 217433
rect 675298 217359 675354 217368
rect 675312 216850 675340 217359
rect 675482 217016 675538 217025
rect 675482 216951 675538 216960
rect 675300 216844 675352 216850
rect 675300 216786 675352 216792
rect 675496 216714 675524 216951
rect 675484 216708 675536 216714
rect 675484 216650 675536 216656
rect 675114 216200 675170 216209
rect 675114 216135 675170 216144
rect 675128 212534 675156 216135
rect 675482 215792 675538 215801
rect 675482 215727 675538 215736
rect 675496 215490 675524 215727
rect 675484 215484 675536 215490
rect 675484 215426 675536 215432
rect 675298 215384 675354 215393
rect 675298 215319 675300 215328
rect 675352 215319 675354 215328
rect 675300 215290 675352 215296
rect 675482 214160 675538 214169
rect 675482 214095 675484 214104
rect 675536 214095 675538 214104
rect 675484 214066 675536 214072
rect 675482 213752 675538 213761
rect 675482 213687 675484 213696
rect 675536 213687 675538 213696
rect 675484 213658 675536 213664
rect 675482 213344 675538 213353
rect 675482 213279 675484 213288
rect 675536 213279 675538 213288
rect 675484 213250 675536 213256
rect 675036 212506 675156 212534
rect 683118 212528 683174 212537
rect 674840 205760 674892 205766
rect 674840 205702 674892 205708
rect 675036 202874 675064 212506
rect 683118 212463 683174 212472
rect 675482 212120 675538 212129
rect 675482 212055 675538 212064
rect 675496 208146 675524 212055
rect 683132 211818 683160 212463
rect 675852 211812 675904 211818
rect 675852 211754 675904 211760
rect 683120 211812 683172 211818
rect 683120 211754 683172 211760
rect 675864 209953 675892 211754
rect 675850 209944 675906 209953
rect 675850 209879 675906 209888
rect 675484 208140 675536 208146
rect 675484 208082 675536 208088
rect 675392 205760 675444 205766
rect 675392 205702 675444 205708
rect 675404 205323 675432 205702
rect 675758 205048 675814 205057
rect 675758 204983 675814 204992
rect 675772 204680 675800 204983
rect 675666 204232 675722 204241
rect 675666 204167 675722 204176
rect 675680 204035 675708 204167
rect 675036 202846 675156 202874
rect 675128 201634 675156 202846
rect 675390 202736 675446 202745
rect 675390 202671 675446 202680
rect 675404 202195 675432 202671
rect 675312 201742 675432 201770
rect 675312 201634 675340 201742
rect 675128 201606 675340 201634
rect 675404 201620 675432 201742
rect 675392 201476 675444 201482
rect 675392 201418 675444 201424
rect 675116 201272 675168 201278
rect 675116 201214 675168 201220
rect 674932 200796 674984 200802
rect 674932 200738 674984 200744
rect 674944 194834 674972 200738
rect 675128 196058 675156 201214
rect 675404 201008 675432 201418
rect 675772 200025 675800 200328
rect 675758 200016 675814 200025
rect 675758 199951 675814 199960
rect 675300 198688 675352 198694
rect 675300 198630 675352 198636
rect 675312 198370 675340 198630
rect 675312 198342 675432 198370
rect 675404 197880 675432 198342
rect 675300 197804 675352 197810
rect 675300 197746 675352 197752
rect 675312 197282 675340 197746
rect 675404 197282 675432 197336
rect 675312 197254 675432 197282
rect 675758 197160 675814 197169
rect 675758 197095 675814 197104
rect 675772 196656 675800 197095
rect 675128 196030 675418 196058
rect 674944 194806 675418 194834
rect 675758 193216 675814 193225
rect 675758 193151 675814 193160
rect 675772 192984 675800 193151
rect 675404 191978 675432 192372
rect 675312 191950 675432 191978
rect 675312 190330 675340 191950
rect 675482 191584 675538 191593
rect 675482 191519 675538 191528
rect 675496 191148 675524 191519
rect 675300 190324 675352 190330
rect 675300 190266 675352 190272
rect 676034 185872 676090 185881
rect 676034 185807 676090 185816
rect 675482 178528 675538 178537
rect 675482 178463 675538 178472
rect 675496 178294 675524 178463
rect 675484 178288 675536 178294
rect 675484 178230 675536 178236
rect 675484 178152 675536 178158
rect 675482 178120 675484 178129
rect 675536 178120 675538 178129
rect 675482 178055 675538 178064
rect 675484 177744 675536 177750
rect 675482 177712 675484 177721
rect 675536 177712 675538 177721
rect 675482 177647 675538 177656
rect 676048 177313 676076 185807
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 676034 177304 676090 177313
rect 676034 177239 676090 177248
rect 675482 176896 675538 176905
rect 675482 176831 675484 176840
rect 675536 176831 675538 176840
rect 675484 176802 675536 176808
rect 675482 176488 675538 176497
rect 675482 176423 675538 176432
rect 674654 175672 674710 175681
rect 674654 175607 674710 175616
rect 675496 175438 675524 176423
rect 675484 175432 675536 175438
rect 675484 175374 675536 175380
rect 675482 175264 675538 175273
rect 675482 175199 675484 175208
rect 675536 175199 675538 175208
rect 675484 175170 675536 175176
rect 675482 174448 675538 174457
rect 675482 174383 675484 174392
rect 675536 174383 675538 174392
rect 675484 174354 675536 174360
rect 675022 174040 675078 174049
rect 675022 173975 675078 173984
rect 674484 172094 674696 172122
rect 674470 172000 674526 172009
rect 674470 171935 674526 171944
rect 674484 148986 674512 171935
rect 674472 148980 674524 148986
rect 674472 148922 674524 148928
rect 674288 144220 674340 144226
rect 674288 144162 674340 144168
rect 673920 132184 673972 132190
rect 673920 132126 673972 132132
rect 674668 131345 674696 172094
rect 674838 162208 674894 162217
rect 674838 162143 674894 162152
rect 674852 157230 674880 162143
rect 675036 159066 675064 173975
rect 675850 173224 675906 173233
rect 675850 173159 675906 173168
rect 675206 171592 675262 171601
rect 675206 171527 675262 171536
rect 675220 159678 675248 171527
rect 675482 171184 675538 171193
rect 675482 171119 675484 171128
rect 675536 171119 675538 171128
rect 675484 171090 675536 171096
rect 675482 169552 675538 169561
rect 675482 169487 675484 169496
rect 675536 169487 675538 169496
rect 675484 169458 675536 169464
rect 675482 169144 675538 169153
rect 675482 169079 675484 169088
rect 675536 169079 675538 169088
rect 675484 169050 675536 169056
rect 675482 168736 675538 168745
rect 675482 168671 675484 168680
rect 675536 168671 675538 168680
rect 675484 168642 675536 168648
rect 675666 167920 675722 167929
rect 675666 167855 675722 167864
rect 675482 167104 675538 167113
rect 675482 167039 675484 167048
rect 675536 167039 675538 167048
rect 675484 167010 675536 167016
rect 675680 166954 675708 167855
rect 675864 166994 675892 173159
rect 676034 172816 676090 172825
rect 676090 172774 676260 172802
rect 676034 172751 676090 172760
rect 676232 169674 676260 172774
rect 678242 172408 678298 172417
rect 678242 172343 678298 172352
rect 676678 170776 676734 170785
rect 676678 170711 676734 170720
rect 676402 169960 676458 169969
rect 676402 169895 676458 169904
rect 675496 166926 675708 166954
rect 675772 166966 675892 166994
rect 676048 169646 676260 169674
rect 675496 166870 675524 166926
rect 675484 166864 675536 166870
rect 675484 166806 675536 166812
rect 675772 163690 675800 166966
rect 675312 163662 675800 163690
rect 675312 160290 675340 163662
rect 676048 162217 676076 169646
rect 676416 166433 676444 169895
rect 676402 166424 676458 166433
rect 676402 166359 676458 166368
rect 676692 166297 676720 170711
rect 676678 166288 676734 166297
rect 676678 166223 676734 166232
rect 676034 162208 676090 162217
rect 676034 162143 676090 162152
rect 678256 161945 678284 172343
rect 678242 161936 678298 161945
rect 678242 161871 678298 161880
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675220 159650 675418 159678
rect 675036 159038 675340 159066
rect 675312 158930 675340 159038
rect 675404 158930 675432 159052
rect 675312 158902 675432 158930
rect 674852 157202 675340 157230
rect 675312 157162 675340 157202
rect 675404 157162 675432 157216
rect 675312 157134 675432 157162
rect 675128 156629 675418 156657
rect 675128 154970 675156 156629
rect 675758 156360 675814 156369
rect 675758 156295 675814 156304
rect 675772 155992 675800 156295
rect 675392 155848 675444 155854
rect 675444 155796 675524 155802
rect 675392 155790 675524 155796
rect 675404 155774 675524 155790
rect 675496 155380 675524 155774
rect 675116 154964 675168 154970
rect 675116 154906 675168 154912
rect 675666 153096 675722 153105
rect 675666 153031 675722 153040
rect 675680 152864 675708 153031
rect 674944 152306 675418 152334
rect 674944 150414 674972 152306
rect 675116 151768 675168 151774
rect 675116 151710 675168 151716
rect 675128 151042 675156 151710
rect 675772 151473 675800 151675
rect 675758 151464 675814 151473
rect 675758 151399 675814 151408
rect 675128 151014 675418 151042
rect 674932 150408 674984 150414
rect 674932 150350 674984 150356
rect 675758 150376 675814 150385
rect 675758 150311 675814 150320
rect 675772 149835 675800 150311
rect 675300 148980 675352 148986
rect 675300 148922 675352 148928
rect 675312 146690 675340 148922
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675312 146662 675432 146690
rect 675404 146132 675432 146662
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 675484 133408 675536 133414
rect 675482 133376 675484 133385
rect 675536 133376 675538 133385
rect 675482 133311 675538 133320
rect 675482 132968 675538 132977
rect 675482 132903 675484 132912
rect 675536 132903 675538 132912
rect 675484 132874 675536 132880
rect 675484 132796 675536 132802
rect 675484 132738 675536 132744
rect 675496 132569 675524 132738
rect 675482 132560 675538 132569
rect 675482 132495 675538 132504
rect 675484 132184 675536 132190
rect 675482 132152 675484 132161
rect 675536 132152 675538 132161
rect 675482 132087 675538 132096
rect 675482 131744 675538 131753
rect 675482 131679 675538 131688
rect 674654 131336 674710 131345
rect 674654 131271 674710 131280
rect 675496 131238 675524 131679
rect 675484 131232 675536 131238
rect 675484 131174 675536 131180
rect 675482 130928 675538 130937
rect 675482 130863 675484 130872
rect 675536 130863 675538 130872
rect 675484 130834 675536 130840
rect 673368 130552 673420 130558
rect 675484 130552 675536 130558
rect 673368 130494 673420 130500
rect 675482 130520 675484 130529
rect 675536 130520 675538 130529
rect 675482 130455 675538 130464
rect 675482 130112 675538 130121
rect 675482 130047 675538 130056
rect 675496 129946 675524 130047
rect 675484 129940 675536 129946
rect 675484 129882 675536 129888
rect 673000 129736 673052 129742
rect 675484 129736 675536 129742
rect 673000 129678 673052 129684
rect 675482 129704 675484 129713
rect 675536 129704 675538 129713
rect 675482 129639 675538 129648
rect 675482 129296 675538 129305
rect 675482 129231 675538 129240
rect 675496 128382 675524 129231
rect 675484 128376 675536 128382
rect 675484 128318 675536 128324
rect 676218 128208 676274 128217
rect 676218 128143 676274 128152
rect 674838 127664 674894 127673
rect 674838 127599 674894 127608
rect 673184 125996 673236 126002
rect 673184 125938 673236 125944
rect 673000 125792 673052 125798
rect 673000 125734 673052 125740
rect 672632 115864 672684 115870
rect 672632 115806 672684 115812
rect 671528 111784 671580 111790
rect 671528 111726 671580 111732
rect 673012 111178 673040 125734
rect 673196 111790 673224 125938
rect 674378 125216 674434 125225
rect 674378 125151 674434 125160
rect 674194 124808 674250 124817
rect 674194 124743 674250 124752
rect 673368 123956 673420 123962
rect 673368 123898 673420 123904
rect 673184 111784 673236 111790
rect 673184 111726 673236 111732
rect 673000 111172 673052 111178
rect 673000 111114 673052 111120
rect 669136 108996 669188 109002
rect 669136 108938 669188 108944
rect 671344 108996 671396 109002
rect 671344 108938 671396 108944
rect 669148 107681 669176 108938
rect 669134 107672 669190 107681
rect 669134 107607 669190 107616
rect 673380 106554 673408 123898
rect 674012 123140 674064 123146
rect 674012 123082 674064 123088
rect 674024 114170 674052 123082
rect 674012 114164 674064 114170
rect 674012 114106 674064 114112
rect 674208 107030 674236 124743
rect 674196 107024 674248 107030
rect 674196 106966 674248 106972
rect 673368 106548 673420 106554
rect 673368 106490 673420 106496
rect 674392 104666 674420 125151
rect 674654 123584 674710 123593
rect 674654 123519 674710 123528
rect 674668 105822 674696 123519
rect 674852 112010 674880 127599
rect 675024 126200 675076 126206
rect 675024 126142 675076 126148
rect 675484 126200 675536 126206
rect 675852 126200 675904 126206
rect 675536 126160 675852 126188
rect 675484 126142 675536 126148
rect 675852 126142 675904 126148
rect 675036 115530 675064 126142
rect 675482 126032 675538 126041
rect 675482 125967 675484 125976
rect 675536 125967 675538 125976
rect 675484 125938 675536 125944
rect 675484 125792 675536 125798
rect 675484 125734 675536 125740
rect 675496 125633 675524 125734
rect 675482 125624 675538 125633
rect 675482 125559 675538 125568
rect 675482 123992 675538 124001
rect 675482 123927 675484 123936
rect 675536 123927 675538 123936
rect 675484 123898 675536 123904
rect 675482 123176 675538 123185
rect 675482 123111 675484 123120
rect 675536 123111 675538 123120
rect 675484 123082 675536 123088
rect 676232 122913 676260 128143
rect 676402 127800 676458 127809
rect 676402 127735 676458 127744
rect 676416 126206 676444 127735
rect 683118 126576 683174 126585
rect 683118 126511 683174 126520
rect 676404 126200 676456 126206
rect 676404 126142 676456 126148
rect 679622 126168 679678 126177
rect 679622 126103 679678 126112
rect 676218 122904 676274 122913
rect 676218 122839 676274 122848
rect 675482 122496 675538 122505
rect 675482 122431 675484 122440
rect 675536 122431 675538 122440
rect 675484 122402 675536 122408
rect 677598 122088 677654 122097
rect 677598 122023 677654 122032
rect 675482 121952 675538 121961
rect 675482 121887 675538 121896
rect 675496 121446 675524 121887
rect 675484 121440 675536 121446
rect 675484 121382 675536 121388
rect 675852 117292 675904 117298
rect 675852 117234 675904 117240
rect 675864 116090 675892 117234
rect 677612 116113 677640 122023
rect 679636 117298 679664 126103
rect 683132 124545 683160 126511
rect 683118 124536 683174 124545
rect 683118 124471 683174 124480
rect 679624 117292 679676 117298
rect 679624 117234 679676 117240
rect 675220 116062 675892 116090
rect 677598 116104 677654 116113
rect 675024 115524 675076 115530
rect 675024 115466 675076 115472
rect 675220 115274 675248 116062
rect 677598 116039 677654 116048
rect 675392 115524 675444 115530
rect 675392 115466 675444 115472
rect 675128 115246 675248 115274
rect 675128 114493 675156 115246
rect 675404 115124 675432 115466
rect 675128 114465 675418 114493
rect 675758 114200 675814 114209
rect 675758 114135 675814 114144
rect 675772 113832 675800 114135
rect 674852 111982 675418 112010
rect 675116 111784 675168 111790
rect 675116 111726 675168 111732
rect 675128 111466 675156 111726
rect 675128 111438 675418 111466
rect 675392 111172 675444 111178
rect 675392 111114 675444 111120
rect 675404 110772 675432 111114
rect 675758 110392 675814 110401
rect 675758 110327 675814 110336
rect 675772 110160 675800 110327
rect 675666 108080 675722 108089
rect 675666 108015 675722 108024
rect 675680 107644 675708 108015
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106554 675156 107086
rect 675300 107024 675352 107030
rect 675300 106966 675352 106972
rect 675116 106548 675168 106554
rect 675116 106490 675168 106496
rect 675312 106502 675340 106966
rect 675312 106474 675418 106502
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 674668 105794 675340 105822
rect 675404 105808 675432 105862
rect 674392 104638 675340 104666
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 668950 104408 669006 104417
rect 668950 104343 669006 104352
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 668582 102776 668638 102785
rect 668582 102711 668638 102720
rect 675666 102640 675722 102649
rect 675666 102575 675722 102584
rect 675680 102136 675708 102575
rect 580264 102128 580316 102134
rect 589464 102128 589516 102134
rect 580264 102070 580316 102076
rect 589462 102096 589464 102105
rect 589516 102096 589518 102105
rect 589462 102031 589518 102040
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 595272 100014 595608 100042
rect 596192 100014 596344 100042
rect 596560 100014 597080 100042
rect 597572 100014 597816 100042
rect 598032 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600424 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 577504 97980 577556 97986
rect 577504 97922 577556 97928
rect 594064 97980 594116 97986
rect 594064 97922 594116 97928
rect 592684 97708 592736 97714
rect 592684 97650 592736 97656
rect 578884 97300 578936 97306
rect 578884 97242 578936 97248
rect 577504 77308 577556 77314
rect 577504 77250 577556 77256
rect 145380 52964 145432 52970
rect 145380 52906 145432 52912
rect 78476 52686 78628 52714
rect 130824 52686 131068 52714
rect 78600 49745 78628 52686
rect 131040 50289 131068 52686
rect 145392 50810 145420 52906
rect 287868 52822 288204 52850
rect 392564 52822 392624 52850
rect 183172 52686 183508 52714
rect 235520 52686 235856 52714
rect 145084 50782 145420 50810
rect 183480 50386 183508 52686
rect 235828 51066 235856 52686
rect 288176 52426 288204 52822
rect 340216 52686 340552 52714
rect 288164 52420 288216 52426
rect 288164 52362 288216 52368
rect 288176 51066 288204 52362
rect 340524 51066 340552 52686
rect 392596 52290 392624 52822
rect 444912 52686 445248 52714
rect 497260 52686 497596 52714
rect 391940 52284 391992 52290
rect 391940 52226 391992 52232
rect 392584 52284 392636 52290
rect 392584 52226 392636 52232
rect 391952 51066 391980 52226
rect 235816 51060 235868 51066
rect 235816 51002 235868 51008
rect 288164 51060 288216 51066
rect 288164 51002 288216 51008
rect 340512 51060 340564 51066
rect 340512 51002 340564 51008
rect 391940 51060 391992 51066
rect 391940 51002 391992 51008
rect 405096 50516 405148 50522
rect 405096 50458 405148 50464
rect 183468 50380 183520 50386
rect 183468 50322 183520 50328
rect 131026 50280 131082 50289
rect 131026 50215 131082 50224
rect 78586 49736 78642 49745
rect 78586 49671 78642 49680
rect 151910 47288 151966 47297
rect 151910 47223 151966 47232
rect 142172 46702 142370 46730
rect 142172 43874 142200 46702
rect 151924 45937 151952 47223
rect 151910 45928 151966 45937
rect 151910 45863 151966 45872
rect 194048 44872 194100 44878
rect 194048 44814 194100 44820
rect 141896 43846 142200 43874
rect 141896 40202 141924 43846
rect 187514 42120 187570 42129
rect 187358 42078 187514 42106
rect 194060 42092 194088 44814
rect 315948 43444 316000 43450
rect 315948 43386 316000 43392
rect 306976 42392 307032 42401
rect 306976 42327 307032 42336
rect 306990 42092 307018 42327
rect 315960 42231 315988 43386
rect 315948 42225 316000 42231
rect 315948 42167 316000 42173
rect 310426 42120 310482 42129
rect 310132 42078 310426 42106
rect 187514 42055 187570 42064
rect 361946 42120 362002 42129
rect 361790 42078 361946 42106
rect 310426 42055 310482 42064
rect 365166 42120 365222 42129
rect 364918 42078 365166 42106
rect 361946 42055 362002 42064
rect 405108 42106 405136 50458
rect 406384 50380 406436 50386
rect 406384 50322 406436 50328
rect 406396 45121 406424 50322
rect 445220 50289 445248 52686
rect 497568 50561 497596 52686
rect 549272 52686 549608 52714
rect 497554 50552 497610 50561
rect 497554 50487 497610 50496
rect 549272 50289 549300 52686
rect 577516 52290 577544 77250
rect 577504 52284 577556 52290
rect 577504 52226 577556 52232
rect 578896 50522 578924 97242
rect 591304 77444 591356 77450
rect 591304 77386 591356 77392
rect 580264 75948 580316 75954
rect 580264 75890 580316 75896
rect 580276 53106 580304 75890
rect 580264 53100 580316 53106
rect 580264 53042 580316 53048
rect 578884 50516 578936 50522
rect 578884 50458 578936 50464
rect 445206 50280 445262 50289
rect 445206 50215 445262 50224
rect 549258 50280 549314 50289
rect 549258 50215 549314 50224
rect 415214 48104 415270 48113
rect 415214 48039 415270 48048
rect 406382 45112 406438 45121
rect 406382 45047 406438 45056
rect 411074 42800 411130 42809
rect 411074 42735 411130 42744
rect 411088 42500 411116 42735
rect 415228 42378 415256 48039
rect 591316 47569 591344 77386
rect 591302 47560 591358 47569
rect 591302 47495 591358 47504
rect 470612 47382 471008 47410
rect 470612 47297 470640 47382
rect 451278 47288 451334 47297
rect 451278 47223 451334 47232
rect 451462 47288 451518 47297
rect 451462 47223 451518 47232
rect 461030 47288 461086 47297
rect 461030 47223 461032 47232
rect 451292 46753 451320 47223
rect 451278 46744 451334 46753
rect 451278 46679 451334 46688
rect 451476 45937 451504 47223
rect 461084 47223 461086 47232
rect 461214 47288 461270 47297
rect 470598 47288 470654 47297
rect 461214 47223 461270 47232
rect 465908 47252 465960 47258
rect 461032 47194 461084 47200
rect 461228 46753 461256 47223
rect 470598 47223 470654 47232
rect 470782 47288 470838 47297
rect 470782 47223 470838 47232
rect 465908 47194 465960 47200
rect 461214 46744 461270 46753
rect 461214 46679 461270 46688
rect 465722 46744 465778 46753
rect 465722 46679 465778 46688
rect 451462 45928 451518 45937
rect 451462 45863 451518 45872
rect 465736 45801 465764 46679
rect 465920 45937 465948 47194
rect 470796 45937 470824 47223
rect 470980 45937 471008 47382
rect 499592 47382 499988 47410
rect 480442 47288 480498 47297
rect 480442 47223 480498 47232
rect 480626 47288 480682 47297
rect 480626 47223 480682 47232
rect 490010 47288 490066 47297
rect 490010 47223 490066 47232
rect 490194 47288 490250 47297
rect 490194 47223 490250 47232
rect 480456 45937 480484 47223
rect 465906 45928 465962 45937
rect 465906 45863 465962 45872
rect 470782 45928 470838 45937
rect 470782 45863 470838 45872
rect 470966 45928 471022 45937
rect 470966 45863 471022 45872
rect 480258 45928 480314 45937
rect 480258 45863 480314 45872
rect 480442 45928 480498 45937
rect 480442 45863 480498 45872
rect 465722 45792 465778 45801
rect 480272 45778 480300 45863
rect 480640 45778 480668 47223
rect 480272 45750 480668 45778
rect 490024 45778 490052 47223
rect 490208 45937 490236 47223
rect 499592 45937 499620 47382
rect 499960 47297 499988 47382
rect 499762 47288 499818 47297
rect 499762 47223 499818 47232
rect 499946 47288 500002 47297
rect 499946 47223 500002 47232
rect 513746 47288 513802 47297
rect 513746 47223 513802 47232
rect 499776 45937 499804 47223
rect 513760 47002 513788 47223
rect 514206 47016 514262 47025
rect 513760 46974 514206 47002
rect 514206 46951 514262 46960
rect 592696 46209 592724 97650
rect 594076 46481 594104 97922
rect 595272 97850 595300 100014
rect 596192 97986 596220 100014
rect 596180 97980 596232 97986
rect 596180 97922 596232 97928
rect 595260 97844 595312 97850
rect 595260 97786 595312 97792
rect 595628 97844 595680 97850
rect 595628 97786 595680 97792
rect 595444 97572 595496 97578
rect 595444 97514 595496 97520
rect 595456 48113 595484 97514
rect 595640 80714 595668 97786
rect 596560 84194 596588 100014
rect 597572 97714 597600 100014
rect 597560 97708 597612 97714
rect 597560 97650 597612 97656
rect 598032 84194 598060 100014
rect 598952 97306 598980 100014
rect 598940 97300 598992 97306
rect 598940 97242 598992 97248
rect 599504 84194 599532 100014
rect 600424 97578 600452 100014
rect 600412 97572 600464 97578
rect 600412 97514 600464 97520
rect 600884 84194 600912 100014
rect 601896 96966 601924 100014
rect 601056 96960 601108 96966
rect 601056 96902 601108 96908
rect 601884 96960 601936 96966
rect 601884 96902 601936 96908
rect 601068 84194 601096 96902
rect 602356 84194 602384 100014
rect 596192 84166 596588 84194
rect 597572 84166 598060 84194
rect 598952 84166 599532 84194
rect 600332 84166 600912 84194
rect 600976 84166 601096 84194
rect 601712 84166 602384 84194
rect 595628 80708 595680 80714
rect 595628 80650 595680 80656
rect 596192 48929 596220 84166
rect 596178 48920 596234 48929
rect 596178 48855 596234 48864
rect 595442 48104 595498 48113
rect 595442 48039 595498 48048
rect 597572 47841 597600 84166
rect 597558 47832 597614 47841
rect 597558 47767 597614 47776
rect 598952 47297 598980 84166
rect 600332 49201 600360 84166
rect 600318 49192 600374 49201
rect 600318 49127 600374 49136
rect 598938 47288 598994 47297
rect 598938 47223 598994 47232
rect 600976 46753 601004 84166
rect 600962 46744 601018 46753
rect 600962 46679 601018 46688
rect 594062 46472 594118 46481
rect 594062 46407 594118 46416
rect 592682 46200 592738 46209
rect 592682 46135 592738 46144
rect 490194 45928 490250 45937
rect 490194 45863 490250 45872
rect 490378 45928 490434 45937
rect 490378 45863 490434 45872
rect 499578 45928 499634 45937
rect 499578 45863 499634 45872
rect 499762 45928 499818 45937
rect 499762 45863 499818 45872
rect 490392 45778 490420 45863
rect 490024 45750 490420 45778
rect 465722 45727 465778 45736
rect 601712 44849 601740 84166
rect 603092 51785 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 607168 100042
rect 607384 100014 607720 100042
rect 608120 100014 608456 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613608 100042
rect 604426 99742 604500 99770
rect 603078 51776 603134 51785
rect 603078 51711 603134 51720
rect 601698 44840 601754 44849
rect 601698 44775 601754 44784
rect 604472 43489 604500 99742
rect 605484 97306 605512 100014
rect 605472 97300 605524 97306
rect 605472 97242 605524 97248
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606944 96960 606996 96966
rect 606944 96902 606996 96908
rect 606956 93854 606984 96902
rect 607140 96506 607168 100014
rect 607140 96478 607352 96506
rect 606956 93826 607168 93854
rect 607140 75206 607168 93826
rect 607324 88330 607352 96478
rect 607692 94518 607720 100014
rect 608428 95946 608456 100014
rect 609164 96898 609192 100014
rect 609152 96892 609204 96898
rect 609152 96834 609204 96840
rect 609704 96892 609756 96898
rect 609704 96834 609756 96840
rect 608416 95940 608468 95946
rect 608416 95882 608468 95888
rect 607680 94512 607732 94518
rect 607680 94454 607732 94460
rect 609716 93158 609744 96834
rect 609704 93152 609756 93158
rect 609704 93094 609756 93100
rect 607312 88324 607364 88330
rect 607312 88266 607364 88272
rect 609900 85542 609928 100014
rect 610636 96082 610664 100014
rect 610624 96076 610676 96082
rect 610624 96018 610676 96024
rect 611280 91050 611308 100014
rect 611912 97300 611964 97306
rect 611912 97242 611964 97248
rect 611924 93854 611952 97242
rect 612108 96762 612136 100014
rect 612660 96966 612688 100014
rect 612648 96960 612700 96966
rect 612648 96902 612700 96908
rect 613384 96960 613436 96966
rect 613384 96902 613436 96908
rect 612096 96756 612148 96762
rect 612096 96698 612148 96704
rect 612556 96756 612608 96762
rect 612556 96698 612608 96704
rect 611924 93826 612044 93854
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 607128 75200 607180 75206
rect 607128 75142 607180 75148
rect 612016 57254 612044 93826
rect 612568 80850 612596 96698
rect 612556 80844 612608 80850
rect 612556 80786 612608 80792
rect 613396 76566 613424 96902
rect 613580 96830 613608 100014
rect 613994 99770 614022 100028
rect 614744 100014 615080 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 617932 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613994 99742 614068 99770
rect 614040 96966 614068 99742
rect 614028 96960 614080 96966
rect 614028 96902 614080 96908
rect 614764 96960 614816 96966
rect 614764 96902 614816 96908
rect 613568 96824 613620 96830
rect 613568 96766 613620 96772
rect 614028 96824 614080 96830
rect 614028 96766 614080 96772
rect 614040 77994 614068 96766
rect 614028 77988 614080 77994
rect 614028 77930 614080 77936
rect 614776 76702 614804 96902
rect 615052 93854 615080 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 616524 95198 616552 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616512 95192 616564 95198
rect 616512 95134 616564 95140
rect 615052 93826 615448 93854
rect 614764 76696 614816 76702
rect 614764 76638 614816 76644
rect 613384 76560 613436 76566
rect 613384 76502 613436 76508
rect 615420 75342 615448 93826
rect 616800 79354 616828 96902
rect 617260 96762 617288 100014
rect 617248 96756 617300 96762
rect 617248 96698 617300 96704
rect 617904 92478 617932 100014
rect 618732 97442 618760 100014
rect 618720 97436 618772 97442
rect 618720 97378 618772 97384
rect 618076 96756 618128 96762
rect 618076 96698 618128 96704
rect 617892 92472 617944 92478
rect 617892 92414 617944 92420
rect 618088 91050 618116 96698
rect 619560 93838 619588 100014
rect 620204 97714 620232 100014
rect 620192 97708 620244 97714
rect 620192 97650 620244 97656
rect 620940 96286 620968 100014
rect 621676 98802 621704 100014
rect 621664 98796 621716 98802
rect 621664 98738 621716 98744
rect 622320 98666 622348 100014
rect 622308 98660 622360 98666
rect 622308 98602 622360 98608
rect 623148 97578 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 624620 97986 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628236 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 631916 100042
rect 632408 100014 632744 100042
rect 633144 100014 633388 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635688 100042
rect 625034 99742 625108 99770
rect 625080 99074 625108 99742
rect 625068 99068 625120 99074
rect 625068 99010 625120 99016
rect 624608 97980 624660 97986
rect 624608 97922 624660 97928
rect 626092 97850 626120 100014
rect 626080 97844 626132 97850
rect 626080 97786 626132 97792
rect 626080 97708 626132 97714
rect 626080 97650 626132 97656
rect 623136 97572 623188 97578
rect 623136 97514 623188 97520
rect 620928 96280 620980 96286
rect 620928 96222 620980 96228
rect 621664 96076 621716 96082
rect 621664 96018 621716 96024
rect 620284 95940 620336 95946
rect 620284 95882 620336 95888
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 618904 93152 618956 93158
rect 618904 93094 618956 93100
rect 617340 91044 617392 91050
rect 617340 90986 617392 90992
rect 618076 91044 618128 91050
rect 618076 90986 618128 90992
rect 617352 88194 617380 90986
rect 617340 88188 617392 88194
rect 617340 88130 617392 88136
rect 618916 84046 618944 93094
rect 620296 84182 620324 95882
rect 621676 86290 621704 96018
rect 623044 95192 623096 95198
rect 623044 95134 623096 95140
rect 623056 89690 623084 95134
rect 624976 94512 625028 94518
rect 626092 94489 626120 97650
rect 626264 97436 626316 97442
rect 626264 97378 626316 97384
rect 624976 94454 625028 94460
rect 626078 94480 626134 94489
rect 623044 89684 623096 89690
rect 623044 89626 623096 89632
rect 624988 88369 625016 94454
rect 626078 94415 626134 94424
rect 626276 92585 626304 97378
rect 626828 97170 626856 100014
rect 627564 97442 627592 100014
rect 627552 97436 627604 97442
rect 627552 97378 627604 97384
rect 628208 97306 628236 100014
rect 629036 98802 629064 100014
rect 629772 98938 629800 100014
rect 629760 98932 629812 98938
rect 629760 98874 629812 98880
rect 628380 98796 628432 98802
rect 628380 98738 628432 98744
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 628196 97300 628248 97306
rect 628196 97242 628248 97248
rect 626816 97164 626868 97170
rect 626816 97106 626868 97112
rect 626448 96280 626500 96286
rect 626448 96222 626500 96228
rect 626460 95441 626488 96222
rect 628392 95826 628420 98738
rect 630508 98666 630536 100014
rect 629484 98660 629536 98666
rect 629484 98602 629536 98608
rect 630496 98660 630548 98666
rect 630496 98602 630548 98608
rect 629496 95826 629524 98602
rect 630680 97572 630732 97578
rect 630680 97514 630732 97520
rect 630692 95826 630720 97514
rect 631244 96354 631272 100014
rect 631232 96348 631284 96354
rect 631232 96290 631284 96296
rect 631888 96218 631916 100014
rect 632152 99204 632204 99210
rect 632152 99146 632204 99152
rect 631876 96212 631928 96218
rect 631876 96154 631928 96160
rect 632164 95826 632192 99146
rect 632716 97578 632744 100014
rect 632980 97980 633032 97986
rect 632980 97922 633032 97928
rect 632704 97572 632756 97578
rect 632704 97514 632756 97520
rect 628392 95798 628728 95826
rect 629496 95798 629832 95826
rect 630692 95798 631028 95826
rect 632132 95798 632192 95826
rect 632992 95826 633020 97922
rect 633360 97714 633388 100014
rect 634188 97986 634216 100014
rect 634452 99068 634504 99074
rect 634452 99010 634504 99016
rect 634176 97980 634228 97986
rect 634176 97922 634228 97928
rect 633348 97708 633400 97714
rect 633348 97650 633400 97656
rect 634464 95826 634492 99010
rect 632992 95798 633328 95826
rect 634432 95798 634492 95826
rect 634740 95606 634768 100014
rect 635280 97844 635332 97850
rect 635280 97786 635332 97792
rect 635292 95826 635320 97786
rect 635660 96082 635688 100014
rect 635936 100014 636088 100042
rect 636824 100014 637068 100042
rect 637560 100014 637804 100042
rect 638296 100014 638632 100042
rect 639032 100014 639368 100042
rect 639768 100014 640104 100042
rect 640504 100014 640840 100042
rect 641240 100014 641576 100042
rect 641976 100014 642312 100042
rect 642712 100014 643048 100042
rect 643448 100014 643784 100042
rect 644184 100014 644336 100042
rect 644920 100014 645256 100042
rect 635648 96076 635700 96082
rect 635648 96018 635700 96024
rect 635292 95798 635628 95826
rect 635936 95713 635964 100014
rect 636384 97164 636436 97170
rect 636384 97106 636436 97112
rect 636396 95826 636424 97106
rect 637040 96937 637068 100014
rect 637580 97436 637632 97442
rect 637580 97378 637632 97384
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 95826 637620 97378
rect 637776 95946 637804 100014
rect 638604 96490 638632 100014
rect 639340 97714 639368 100014
rect 639880 98796 639932 98802
rect 639880 98738 639932 98744
rect 639328 97708 639380 97714
rect 639328 97650 639380 97656
rect 639052 97300 639104 97306
rect 639052 97242 639104 97248
rect 638592 96484 638644 96490
rect 638592 96426 638644 96432
rect 637764 95940 637816 95946
rect 637764 95882 637816 95888
rect 639064 95826 639092 97242
rect 636396 95798 636732 95826
rect 637592 95798 637928 95826
rect 639032 95798 639092 95826
rect 639892 95826 639920 98738
rect 640076 96082 640104 100014
rect 640064 96076 640116 96082
rect 640064 96018 640116 96024
rect 640812 95946 640840 100014
rect 640984 98932 641036 98938
rect 640984 98874 641036 98880
rect 640800 95940 640852 95946
rect 640800 95882 640852 95888
rect 640996 95826 641024 98874
rect 641548 96830 641576 100014
rect 642088 98660 642140 98666
rect 642088 98602 642140 98608
rect 641536 96824 641588 96830
rect 641536 96766 641588 96772
rect 639892 95798 640228 95826
rect 640996 95798 641332 95826
rect 635922 95704 635978 95713
rect 642100 95690 642128 98602
rect 642284 96626 642312 100014
rect 642824 96824 642876 96830
rect 642824 96766 642876 96772
rect 642272 96620 642324 96626
rect 642272 96562 642324 96568
rect 642836 96506 642864 96766
rect 643020 96762 643048 100014
rect 643376 97980 643428 97986
rect 643376 97922 643428 97928
rect 643008 96756 643060 96762
rect 643008 96698 643060 96704
rect 642836 96478 643048 96506
rect 642640 96348 642692 96354
rect 642640 96290 642692 96296
rect 642824 96348 642876 96354
rect 642824 96290 642876 96296
rect 642100 95662 642528 95690
rect 635922 95639 635978 95648
rect 634728 95600 634780 95606
rect 634728 95542 634780 95548
rect 626446 95432 626502 95441
rect 626446 95367 626502 95376
rect 642652 95169 642680 96290
rect 642836 95810 642864 96290
rect 642824 95804 642876 95810
rect 642824 95746 642876 95752
rect 643020 95690 643048 96478
rect 642928 95662 643048 95690
rect 642638 95160 642694 95169
rect 642638 95095 642694 95104
rect 642928 94518 642956 95662
rect 643100 95396 643152 95402
rect 643100 95338 643152 95344
rect 642916 94512 642968 94518
rect 642916 94454 642968 94460
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 626460 93537 626488 93774
rect 626446 93528 626502 93537
rect 626446 93463 626502 93472
rect 626262 92576 626318 92585
rect 626262 92511 626318 92520
rect 625436 92472 625488 92478
rect 625436 92414 625488 92420
rect 625448 91633 625476 92414
rect 625434 91624 625490 91633
rect 625434 91559 625490 91568
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90681 626488 90986
rect 626446 90672 626502 90681
rect 626446 90607 626502 90616
rect 626446 89720 626502 89729
rect 626446 89655 626448 89664
rect 626500 89655 626502 89664
rect 626448 89626 626500 89632
rect 624974 88360 625030 88369
rect 624974 88295 625030 88304
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 625620 88188 625672 88194
rect 625620 88130 625672 88136
rect 625632 87009 625660 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 625618 87000 625674 87009
rect 625618 86935 625674 86944
rect 621664 86284 621716 86290
rect 621664 86226 621716 86232
rect 626448 86284 626500 86290
rect 626448 86226 626500 86232
rect 626460 86057 626488 86226
rect 626446 86048 626502 86057
rect 626446 85983 626502 85992
rect 626448 85536 626500 85542
rect 626448 85478 626500 85484
rect 626460 85105 626488 85478
rect 626446 85096 626502 85105
rect 626446 85031 626502 85040
rect 620284 84176 620336 84182
rect 620284 84118 620336 84124
rect 626264 84176 626316 84182
rect 626264 84118 626316 84124
rect 626446 84144 626502 84153
rect 618904 84040 618956 84046
rect 618904 83982 618956 83988
rect 626276 83201 626304 84118
rect 626446 84079 626502 84088
rect 626460 83978 626488 84079
rect 626448 83972 626500 83978
rect 626448 83914 626500 83920
rect 626262 83192 626318 83201
rect 626262 83127 626318 83136
rect 643112 82793 643140 95338
rect 643388 84697 643416 97922
rect 643560 97844 643612 97850
rect 643560 97786 643612 97792
rect 643572 87145 643600 97786
rect 643756 94654 643784 100014
rect 644308 97578 644336 100014
rect 644296 97572 644348 97578
rect 644296 97514 644348 97520
rect 644756 97300 644808 97306
rect 644756 97242 644808 97248
rect 644112 96620 644164 96626
rect 644112 96562 644164 96568
rect 643744 94648 643796 94654
rect 643744 94590 643796 94596
rect 644124 93838 644152 96562
rect 644480 96212 644532 96218
rect 644480 96154 644532 96160
rect 644112 93832 644164 93838
rect 644112 93774 644164 93780
rect 644492 92177 644520 96154
rect 644478 92168 644534 92177
rect 644478 92103 644534 92112
rect 644768 89729 644796 97242
rect 645228 96966 645256 100014
rect 645642 99770 645670 100028
rect 646392 100014 646728 100042
rect 645596 99742 645670 99770
rect 645216 96960 645268 96966
rect 645216 96902 645268 96908
rect 645596 95674 645624 99742
rect 646504 97436 646556 97442
rect 646504 97378 646556 97384
rect 645768 96960 645820 96966
rect 645768 96902 645820 96908
rect 645584 95668 645636 95674
rect 645584 95610 645636 95616
rect 644754 89720 644810 89729
rect 644754 89655 644810 89664
rect 643558 87136 643614 87145
rect 643558 87071 643614 87080
rect 645780 87038 645808 96902
rect 646516 91050 646544 97378
rect 646700 96898 646728 100014
rect 647114 99770 647142 100028
rect 647864 100014 648200 100042
rect 648600 100014 649028 100042
rect 649336 100014 649672 100042
rect 650072 100014 650408 100042
rect 650808 100014 651144 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 647114 99742 647188 99770
rect 647160 97714 647188 99742
rect 647148 97708 647200 97714
rect 647148 97650 647200 97656
rect 646688 96892 646740 96898
rect 646688 96834 646740 96840
rect 647148 96892 647200 96898
rect 647148 96834 647200 96840
rect 646504 91044 646556 91050
rect 646504 90986 646556 90992
rect 647160 89010 647188 96834
rect 647148 89004 647200 89010
rect 647148 88946 647200 88952
rect 648172 87174 648200 100014
rect 649000 96354 649028 100014
rect 648804 96348 648856 96354
rect 648804 96290 648856 96296
rect 648988 96348 649040 96354
rect 648988 96290 649040 96296
rect 648160 87168 648212 87174
rect 648160 87110 648212 87116
rect 645768 87032 645820 87038
rect 645768 86974 645820 86980
rect 643374 84688 643430 84697
rect 643374 84623 643430 84632
rect 643098 82784 643154 82793
rect 643098 82719 643154 82728
rect 628562 81696 628618 81705
rect 628562 81631 628618 81640
rect 628576 80986 628604 81631
rect 628564 80980 628616 80986
rect 628564 80922 628616 80928
rect 631520 80974 631856 81002
rect 638972 80974 639308 81002
rect 642456 80980 642508 80986
rect 629206 80880 629262 80889
rect 629206 80815 629262 80824
rect 629220 79490 629248 80815
rect 629208 79484 629260 79490
rect 629208 79426 629260 79432
rect 616788 79348 616840 79354
rect 616788 79290 616840 79296
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 631060 77722 631088 78066
rect 631048 77716 631100 77722
rect 631048 77658 631100 77664
rect 628288 77580 628340 77586
rect 628288 77522 628340 77528
rect 625804 77444 625856 77450
rect 625804 77386 625856 77392
rect 615408 75336 615460 75342
rect 615408 75278 615460 75284
rect 612004 57248 612056 57254
rect 612004 57190 612056 57196
rect 625816 52426 625844 77386
rect 628300 75954 628328 77522
rect 628288 75948 628340 75954
rect 628288 75890 628340 75896
rect 628300 75290 628328 75890
rect 631060 75290 631088 77658
rect 631520 77586 631548 80974
rect 636108 80708 636160 80714
rect 636108 80650 636160 80656
rect 633898 77752 633954 77761
rect 633898 77687 633954 77696
rect 631508 77580 631560 77586
rect 631508 77522 631560 77528
rect 633912 77450 633940 77687
rect 633900 77444 633952 77450
rect 633900 77386 633952 77392
rect 633912 75290 633940 77386
rect 636120 77294 636148 80650
rect 637488 79484 637540 79490
rect 637488 79426 637540 79432
rect 637118 78568 637174 78577
rect 637118 78503 637174 78512
rect 637132 77314 637160 78503
rect 637500 78266 637528 79426
rect 637488 78260 637540 78266
rect 637488 78202 637540 78208
rect 638972 78130 639000 80974
rect 642456 80922 642508 80928
rect 638960 78124 639012 78130
rect 638960 78066 639012 78072
rect 637120 77308 637172 77314
rect 636120 77266 636332 77294
rect 628176 75262 628328 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636304 75154 636332 77266
rect 637120 77250 637172 77256
rect 639604 77308 639656 77314
rect 639604 77250 639656 77256
rect 639616 75290 639644 77250
rect 642468 75290 642496 80922
rect 645860 80844 645912 80850
rect 645860 80786 645912 80792
rect 645308 78260 645360 78266
rect 645308 78202 645360 78208
rect 645320 75290 645348 78202
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 636304 75126 636732 75154
rect 645872 66042 645900 80786
rect 647424 79348 647476 79354
rect 647424 79290 647476 79296
rect 646320 76696 646372 76702
rect 646320 76638 646372 76644
rect 646136 75336 646188 75342
rect 646136 75278 646188 75284
rect 646148 71777 646176 75278
rect 646134 71768 646190 71777
rect 646134 71703 646190 71712
rect 646332 70417 646360 76638
rect 646872 75200 646924 75206
rect 646872 75142 646924 75148
rect 646884 74497 646912 75142
rect 646870 74488 646926 74497
rect 646870 74423 646926 74432
rect 647436 73001 647464 79290
rect 647608 77988 647660 77994
rect 647608 77930 647660 77936
rect 647422 72992 647478 73001
rect 647422 72927 647478 72936
rect 646318 70408 646374 70417
rect 646318 70343 646374 70352
rect 647620 68513 647648 77930
rect 647606 68504 647662 68513
rect 647606 68439 647662 68448
rect 646134 66056 646190 66065
rect 645872 66014 646134 66042
rect 646134 65991 646190 66000
rect 648816 64025 648844 96290
rect 649264 96076 649316 96082
rect 649264 96018 649316 96024
rect 649276 95538 649304 96018
rect 649264 95532 649316 95538
rect 649264 95474 649316 95480
rect 649644 95198 649672 100014
rect 650380 97034 650408 100014
rect 651116 97238 651144 100014
rect 651852 97714 651880 100014
rect 651840 97708 651892 97714
rect 651840 97650 651892 97656
rect 651104 97232 651156 97238
rect 651104 97174 651156 97180
rect 650368 97028 650420 97034
rect 650368 96970 650420 96976
rect 652588 96626 652616 100014
rect 651288 96620 651340 96626
rect 651288 96562 651340 96568
rect 652576 96620 652628 96626
rect 652576 96562 652628 96568
rect 649632 95192 649684 95198
rect 649632 95134 649684 95140
rect 650644 95192 650696 95198
rect 650644 95134 650696 95140
rect 650656 86494 650684 95134
rect 651300 92478 651328 96562
rect 653324 96490 653352 100014
rect 653312 96484 653364 96490
rect 653312 96426 653364 96432
rect 652024 96212 652076 96218
rect 652024 96154 652076 96160
rect 651288 92472 651340 92478
rect 651288 92414 651340 92420
rect 652036 86766 652064 96154
rect 653404 94648 653456 94654
rect 653404 94590 653456 94596
rect 652024 86760 652076 86766
rect 652024 86702 652076 86708
rect 653416 86630 653444 94590
rect 653968 94217 653996 100014
rect 654324 97232 654376 97238
rect 654324 97174 654376 97180
rect 653954 94208 654010 94217
rect 653954 94143 654010 94152
rect 654140 93764 654192 93770
rect 654140 93706 654192 93712
rect 654152 92585 654180 93706
rect 654336 93401 654364 97174
rect 654796 96898 654824 100014
rect 655440 97850 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97844 655480 97850
rect 655428 97786 655480 97792
rect 654784 96892 654836 96898
rect 654784 96834 654836 96840
rect 655244 96892 655296 96898
rect 655244 96834 655296 96840
rect 654968 96620 655020 96626
rect 654968 96562 655020 96568
rect 654980 96354 655008 96562
rect 654968 96348 655020 96354
rect 654968 96290 655020 96296
rect 654322 93392 654378 93401
rect 654322 93327 654378 93336
rect 654138 92576 654194 92585
rect 654138 92511 654194 92520
rect 654324 92472 654376 92478
rect 654324 92414 654376 92420
rect 654336 91497 654364 92414
rect 654322 91488 654378 91497
rect 654322 91423 654378 91432
rect 654140 91044 654192 91050
rect 654140 90986 654192 90992
rect 654152 90681 654180 90986
rect 654138 90672 654194 90681
rect 654138 90607 654194 90616
rect 655256 88330 655284 96834
rect 655808 89865 655836 100014
rect 656820 97306 656848 100014
rect 656808 97300 656860 97306
rect 656808 97242 656860 97248
rect 656716 96892 656768 96898
rect 656716 96834 656768 96840
rect 656164 95668 656216 95674
rect 656164 95610 656216 95616
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 656176 88806 656204 95610
rect 656164 88800 656216 88806
rect 656164 88742 656216 88748
rect 656728 88670 656756 96834
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 658154 99742 658228 99770
rect 658200 97442 658228 99742
rect 658832 97572 658884 97578
rect 658832 97514 658884 97520
rect 658188 97436 658240 97442
rect 658188 97378 658240 97384
rect 658280 97028 658332 97034
rect 658280 96970 658332 96976
rect 658292 95132 658320 96970
rect 658844 95132 658872 97514
rect 659212 95674 659240 100014
rect 659948 97986 659976 100014
rect 660132 100014 660376 100042
rect 659752 97980 659804 97986
rect 659752 97922 659804 97928
rect 659936 97980 659988 97986
rect 659936 97922 659988 97928
rect 659764 97714 659792 97922
rect 659568 97708 659620 97714
rect 659568 97650 659620 97656
rect 659752 97708 659804 97714
rect 659752 97650 659804 97656
rect 659200 95668 659252 95674
rect 659200 95610 659252 95616
rect 659580 95132 659608 97650
rect 660132 96966 660160 100014
rect 665180 97980 665232 97986
rect 665180 97922 665232 97928
rect 662512 97844 662564 97850
rect 662512 97786 662564 97792
rect 661960 97708 662012 97714
rect 661960 97650 662012 97656
rect 661408 97300 661460 97306
rect 661408 97242 661460 97248
rect 660120 96960 660172 96966
rect 660120 96902 660172 96908
rect 660120 96756 660172 96762
rect 660120 96698 660172 96704
rect 660132 95132 660160 96698
rect 660672 96076 660724 96082
rect 660672 96018 660724 96024
rect 660684 95132 660712 96018
rect 661420 95132 661448 97242
rect 661972 95132 662000 97650
rect 662524 95132 662552 97786
rect 663064 97436 663116 97442
rect 663064 97378 663116 97384
rect 663076 95132 663104 97378
rect 663984 96484 664036 96490
rect 663984 96426 664036 96432
rect 663800 96212 663852 96218
rect 663800 96154 663852 96160
rect 663248 94512 663300 94518
rect 663248 94454 663300 94460
rect 663260 93129 663288 94454
rect 663246 93120 663302 93129
rect 663246 93055 663302 93064
rect 663812 90409 663840 96154
rect 663798 90400 663854 90409
rect 663798 90335 663854 90344
rect 663996 89049 664024 96426
rect 664168 95668 664220 95674
rect 664168 95610 664220 95616
rect 663982 89040 664038 89049
rect 656900 89004 656952 89010
rect 663982 88975 664038 88984
rect 656900 88946 656952 88952
rect 656912 88890 656940 88946
rect 656912 88862 657202 88890
rect 664180 88806 664208 95610
rect 665192 93401 665220 97922
rect 665548 96348 665600 96354
rect 665548 96290 665600 96296
rect 665364 95940 665416 95946
rect 665364 95882 665416 95888
rect 665178 93392 665234 93401
rect 665178 93327 665234 93336
rect 665376 91769 665404 95882
rect 665362 91760 665418 91769
rect 665362 91695 665418 91704
rect 665560 90681 665588 96290
rect 665546 90672 665602 90681
rect 665546 90607 665602 90616
rect 657452 88800 657504 88806
rect 662328 88800 662380 88806
rect 657504 88748 657754 88754
rect 657452 88742 657754 88748
rect 657464 88726 657754 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 664168 88800 664220 88806
rect 664168 88742 664220 88748
rect 661986 88726 662368 88742
rect 656716 88664 656768 88670
rect 656716 88606 656768 88612
rect 659292 88664 659344 88670
rect 659344 88612 659594 88618
rect 659292 88606 659594 88612
rect 659304 88590 659594 88606
rect 658306 88330 658504 88346
rect 655244 88324 655296 88330
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 655244 88266 655296 88272
rect 658464 88266 658516 88272
rect 653404 86624 653456 86630
rect 653404 86566 653456 86572
rect 658844 86494 658872 88196
rect 660132 86766 660160 88196
rect 660684 87038 660712 88196
rect 660672 87032 660724 87038
rect 660672 86974 660724 86980
rect 660120 86760 660172 86766
rect 660120 86702 660172 86708
rect 661420 86630 661448 88196
rect 662524 87174 662552 88196
rect 662512 87168 662564 87174
rect 662512 87110 662564 87116
rect 661408 86624 661460 86630
rect 661408 86566 661460 86572
rect 650644 86488 650696 86494
rect 650644 86430 650696 86436
rect 658832 86488 658884 86494
rect 658832 86430 658884 86436
rect 649172 76560 649224 76566
rect 649172 76502 649224 76508
rect 649184 67017 649212 76502
rect 649170 67008 649226 67017
rect 649170 66943 649226 66952
rect 648802 64016 648858 64025
rect 648802 63951 648858 63960
rect 662420 57248 662472 57254
rect 662420 57190 662472 57196
rect 625804 52420 625856 52426
rect 625804 52362 625856 52368
rect 661222 48240 661278 48249
rect 661222 48175 661278 48184
rect 661236 45554 661264 48175
rect 661590 47789 661646 47798
rect 661590 47724 661646 47733
rect 661144 45526 661264 45554
rect 474462 43480 474518 43489
rect 474462 43415 474518 43424
rect 604458 43480 604514 43489
rect 661144 43450 661172 45526
rect 661604 44878 661632 47724
rect 662432 47433 662460 57190
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661592 44872 661644 44878
rect 661592 44814 661644 44820
rect 604458 43415 604514 43424
rect 661132 43444 661184 43450
rect 416594 42800 416650 42809
rect 416594 42735 416650 42744
rect 464894 42800 464950 42809
rect 464894 42735 464950 42744
rect 415228 42350 415426 42378
rect 405108 42078 405582 42106
rect 416608 42092 416636 42735
rect 464908 42386 464936 42735
rect 474476 42500 474504 43415
rect 661132 43386 661184 43392
rect 518530 42392 518586 42401
rect 464896 42380 464948 42386
rect 464896 42322 464948 42328
rect 518586 42350 518834 42378
rect 518530 42327 518586 42336
rect 460570 42120 460626 42129
rect 460368 42078 460570 42106
rect 365166 42055 365222 42064
rect 471610 42120 471666 42129
rect 471408 42078 471610 42106
rect 460570 42055 460626 42064
rect 471610 42055 471666 42064
rect 514942 42120 514998 42129
rect 520462 42120 520518 42129
rect 514998 42078 515154 42106
rect 514942 42055 514998 42064
rect 525798 42120 525854 42129
rect 520518 42078 520674 42106
rect 520462 42055 520518 42064
rect 529570 42120 529626 42129
rect 525854 42078 526194 42106
rect 529322 42078 529570 42106
rect 525798 42055 525854 42064
rect 529570 42055 529626 42064
rect 521658 41984 521714 41993
rect 521714 41942 521870 41970
rect 521658 41919 521714 41928
rect 141758 40174 141924 40202
rect 141758 39984 141786 40174
<< via2 >>
rect 357714 1007140 357770 1007176
rect 505006 1007156 505008 1007176
rect 505008 1007156 505060 1007176
rect 505060 1007156 505062 1007176
rect 357714 1007120 357716 1007140
rect 357716 1007120 357768 1007140
rect 357768 1007120 357770 1007140
rect 505006 1007120 505062 1007156
rect 357714 1006884 357716 1006904
rect 357716 1006884 357768 1006904
rect 357768 1006884 357770 1006904
rect 357714 1006848 357770 1006884
rect 358542 1006748 358544 1006768
rect 358544 1006748 358596 1006768
rect 358596 1006748 358598 1006768
rect 358542 1006712 358598 1006748
rect 103150 1006596 103206 1006632
rect 103150 1006576 103152 1006596
rect 103152 1006576 103204 1006596
rect 103204 1006576 103206 1006596
rect 153750 1006596 153806 1006632
rect 153750 1006576 153752 1006596
rect 153752 1006576 153804 1006596
rect 153804 1006576 153806 1006596
rect 306930 1006596 306986 1006632
rect 306930 1006576 306932 1006596
rect 306932 1006576 306984 1006596
rect 306984 1006576 306986 1006596
rect 85946 995696 86002 995752
rect 80702 994472 80758 994528
rect 84658 995424 84714 995480
rect 86590 995424 86646 995480
rect 85026 995152 85082 995208
rect 90178 995424 90234 995480
rect 89350 994744 89406 994800
rect 93306 996376 93362 996432
rect 93490 995696 93546 995752
rect 93490 995016 93546 995072
rect 103978 1006460 104034 1006496
rect 103978 1006440 103980 1006460
rect 103980 1006440 104032 1006460
rect 104032 1006440 104034 1006460
rect 100298 1006324 100354 1006360
rect 100298 1006304 100300 1006324
rect 100300 1006304 100352 1006324
rect 100352 1006304 100354 1006324
rect 101954 1006188 102010 1006224
rect 101954 1006168 101956 1006188
rect 101956 1006168 102008 1006188
rect 102008 1006168 102010 1006188
rect 98274 1006052 98330 1006088
rect 98274 1006032 98276 1006052
rect 98276 1006032 98328 1006052
rect 98328 1006032 98330 1006052
rect 94502 994336 94558 994392
rect 87510 994064 87566 994120
rect 92662 994064 92718 994120
rect 41786 968768 41842 968824
rect 41970 967136 42026 967192
rect 41786 962104 41842 962160
rect 41786 959112 41842 959168
rect 41786 956528 41842 956584
rect 41786 955440 41842 955496
rect 39302 952448 39358 952504
rect 37922 952176 37978 952232
rect 35162 938406 35218 938462
rect 40038 951632 40094 951688
rect 41510 951632 41566 951688
rect 39302 937352 39358 937408
rect 37922 936944 37978 937000
rect 41326 941840 41382 941896
rect 40958 941024 41014 941080
rect 41142 939392 41198 939448
rect 40958 938406 41014 938462
rect 40038 935720 40094 935776
rect 40682 881864 40738 881920
rect 39946 819032 40002 819088
rect 35622 817944 35678 818000
rect 35806 817264 35862 817320
rect 40314 817944 40370 818000
rect 35254 816856 35310 816912
rect 35438 816448 35494 816504
rect 35806 816040 35862 816096
rect 35622 815632 35678 815688
rect 35438 815224 35494 815280
rect 35622 814816 35678 814872
rect 35806 814408 35862 814464
rect 41142 814000 41198 814056
rect 41142 812776 41198 812832
rect 42062 940208 42118 940264
rect 42246 937760 42302 937816
rect 42798 935312 42854 935368
rect 43074 934904 43130 934960
rect 43534 943472 43590 943528
rect 43442 942248 43498 942304
rect 43626 941332 43628 941352
rect 43628 941332 43680 941352
rect 43680 941332 43682 941352
rect 43626 941296 43682 941332
rect 43442 939820 43498 939856
rect 43442 939800 43444 939820
rect 43444 939800 43496 939820
rect 43496 939800 43498 939820
rect 43258 934496 43314 934552
rect 44638 943064 44694 943120
rect 47582 942656 47638 942712
rect 46202 940616 46258 940672
rect 97078 997228 97080 997248
rect 97080 997228 97132 997248
rect 97132 997228 97134 997248
rect 97078 997192 97134 997228
rect 98274 1001972 98330 1002008
rect 98274 1001952 98276 1001972
rect 98276 1001952 98328 1001972
rect 98328 1001952 98330 1001972
rect 97446 995560 97502 995616
rect 97262 995288 97318 995344
rect 100298 1002652 100354 1002688
rect 100298 1002632 100300 1002652
rect 100300 1002632 100352 1002652
rect 100352 1002632 100354 1002652
rect 101126 1002516 101182 1002552
rect 101126 1002496 101128 1002516
rect 101128 1002496 101180 1002516
rect 101180 1002496 101182 1002516
rect 99102 1002380 99158 1002416
rect 99102 1002360 99104 1002380
rect 99104 1002360 99156 1002380
rect 99156 1002360 99158 1002380
rect 101126 1002244 101182 1002280
rect 101126 1002224 101128 1002244
rect 101128 1002224 101180 1002244
rect 101180 1002224 101182 1002244
rect 99470 1002108 99526 1002144
rect 99470 1002088 99472 1002108
rect 99472 1002088 99524 1002108
rect 99524 1002088 99526 1002108
rect 100022 995016 100078 995072
rect 101954 1002788 102010 1002824
rect 101954 1002768 101956 1002788
rect 101956 1002768 102008 1002788
rect 102008 1002768 102010 1002788
rect 102322 1001972 102378 1002008
rect 102322 1001952 102324 1001972
rect 102324 1001952 102376 1001972
rect 102376 1001952 102378 1001972
rect 106830 1006188 106886 1006224
rect 106830 1006168 106832 1006188
rect 106832 1006168 106884 1006188
rect 106884 1006168 106886 1006188
rect 103978 1006052 104034 1006088
rect 103978 1006032 103980 1006052
rect 103980 1006032 104032 1006052
rect 104032 1006032 104034 1006052
rect 107658 1006052 107714 1006088
rect 107658 1006032 107660 1006052
rect 107660 1006032 107712 1006052
rect 107712 1006032 107714 1006052
rect 108486 1004692 108542 1004728
rect 108486 1004672 108488 1004692
rect 108488 1004672 108540 1004692
rect 108540 1004672 108542 1004692
rect 106002 1002516 106058 1002552
rect 106002 1002496 106004 1002516
rect 106004 1002496 106056 1002516
rect 106056 1002496 106058 1002516
rect 105634 1002380 105690 1002416
rect 105634 1002360 105636 1002380
rect 105636 1002360 105688 1002380
rect 105688 1002360 105690 1002380
rect 104806 1002244 104862 1002280
rect 104806 1002224 104808 1002244
rect 104808 1002224 104860 1002244
rect 104860 1002224 104862 1002244
rect 103150 1002108 103206 1002144
rect 103150 1002088 103152 1002108
rect 103152 1002088 103204 1002108
rect 103204 1002088 103206 1002108
rect 104806 1001952 104862 1002008
rect 106002 1001972 106058 1002008
rect 106002 1001952 106004 1001972
rect 106004 1001952 106056 1001972
rect 106056 1001952 106058 1001972
rect 108026 1002380 108082 1002416
rect 108026 1002360 108028 1002380
rect 108028 1002360 108080 1002380
rect 108080 1002360 108082 1002380
rect 106830 1002108 106886 1002144
rect 106830 1002088 106832 1002108
rect 106832 1002088 106884 1002108
rect 106884 1002088 106886 1002108
rect 106462 994744 106518 994800
rect 108486 1002244 108542 1002280
rect 108486 1002224 108488 1002244
rect 108488 1002224 108540 1002244
rect 108540 1002224 108542 1002244
rect 108854 1001972 108910 1002008
rect 108854 1001952 108856 1001972
rect 108856 1001952 108908 1001972
rect 108908 1001952 108910 1001972
rect 109682 1002108 109738 1002144
rect 109682 1002088 109684 1002108
rect 109684 1002088 109736 1002108
rect 109736 1002088 109738 1002108
rect 133050 995696 133106 995752
rect 137374 995696 137430 995752
rect 139122 995696 139178 995752
rect 140962 995696 141018 995752
rect 141790 995696 141846 995752
rect 143722 995696 143778 995752
rect 144274 996920 144330 996976
rect 129094 994744 129150 994800
rect 132406 995288 132462 995344
rect 129738 994472 129794 994528
rect 136638 995424 136694 995480
rect 135902 995016 135958 995072
rect 144826 996376 144882 996432
rect 152922 1006460 152978 1006496
rect 152922 1006440 152924 1006460
rect 152924 1006440 152976 1006460
rect 152976 1006440 152978 1006460
rect 152094 1006324 152150 1006360
rect 152094 1006304 152096 1006324
rect 152096 1006304 152148 1006324
rect 152148 1006304 152150 1006324
rect 158258 1006324 158314 1006360
rect 210422 1006340 210424 1006360
rect 210424 1006340 210476 1006360
rect 210476 1006340 210478 1006360
rect 158258 1006304 158260 1006324
rect 158260 1006304 158312 1006324
rect 158312 1006304 158314 1006324
rect 210422 1006304 210478 1006340
rect 159454 1006188 159510 1006224
rect 159454 1006168 159456 1006188
rect 159456 1006168 159508 1006188
rect 159508 1006168 159510 1006188
rect 160282 1006188 160338 1006224
rect 160282 1006168 160284 1006188
rect 160284 1006168 160336 1006188
rect 160336 1006168 160338 1006188
rect 146942 1006032 146998 1006088
rect 148874 1006052 148930 1006088
rect 148874 1006032 148876 1006052
rect 148876 1006032 148928 1006052
rect 148928 1006032 148930 1006052
rect 150070 1006052 150126 1006088
rect 150070 1006032 150072 1006052
rect 150072 1006032 150124 1006052
rect 150124 1006032 150126 1006052
rect 155774 1006052 155830 1006088
rect 155774 1006032 155776 1006052
rect 155776 1006032 155828 1006052
rect 155828 1006032 155830 1006052
rect 158626 1006052 158682 1006088
rect 158626 1006032 158628 1006052
rect 158628 1006032 158680 1006052
rect 158680 1006032 158682 1006052
rect 145746 996648 145802 996704
rect 133142 993928 133198 993984
rect 142802 993928 142858 993984
rect 148322 995424 148378 995480
rect 149242 1001972 149298 1002008
rect 149242 1001952 149244 1001972
rect 149244 1001952 149296 1001972
rect 149296 1001952 149298 1001972
rect 150898 1002380 150954 1002416
rect 150898 1002360 150900 1002380
rect 150900 1002360 150952 1002380
rect 150952 1002360 150954 1002380
rect 150898 1002108 150954 1002144
rect 150898 1002088 150900 1002108
rect 150900 1002088 150952 1002108
rect 150952 1002088 150954 1002108
rect 151726 1004692 151782 1004728
rect 151726 1004672 151728 1004692
rect 151728 1004672 151780 1004692
rect 151780 1004672 151782 1004692
rect 151726 1002244 151782 1002280
rect 151726 1002224 151728 1002244
rect 151728 1002224 151780 1002244
rect 151780 1002224 151782 1002244
rect 152922 1005372 152978 1005408
rect 152922 1005352 152924 1005372
rect 152924 1005352 152976 1005372
rect 152976 1005352 152978 1005372
rect 153750 1004964 153806 1005000
rect 153750 1004944 153752 1004964
rect 153752 1004944 153804 1004964
rect 153804 1004944 153806 1004964
rect 160650 1004964 160706 1005000
rect 160650 1004944 160652 1004964
rect 160652 1004944 160704 1004964
rect 160704 1004944 160706 1004964
rect 154118 1004828 154174 1004864
rect 154118 1004808 154120 1004828
rect 154120 1004808 154172 1004828
rect 154172 1004808 154174 1004828
rect 159454 1004828 159510 1004864
rect 159454 1004808 159456 1004828
rect 159456 1004808 159508 1004828
rect 159508 1004808 159510 1004828
rect 160650 1004692 160706 1004728
rect 160650 1004672 160652 1004692
rect 160652 1004672 160704 1004692
rect 160704 1004672 160706 1004692
rect 157430 1002652 157486 1002688
rect 157430 1002632 157432 1002652
rect 157432 1002632 157484 1002652
rect 157484 1002632 157486 1002652
rect 158626 1002516 158682 1002552
rect 158626 1002496 158628 1002516
rect 158628 1002496 158680 1002516
rect 158680 1002496 158682 1002516
rect 156602 1002380 156658 1002416
rect 156602 1002360 156604 1002380
rect 156604 1002360 156656 1002380
rect 156656 1002360 156658 1002380
rect 155774 1002244 155830 1002280
rect 155774 1002224 155776 1002244
rect 155776 1002224 155828 1002244
rect 155828 1002224 155830 1002244
rect 156602 1002108 156658 1002144
rect 156602 1002088 156604 1002108
rect 156604 1002088 156656 1002108
rect 156656 1002088 156658 1002108
rect 154578 1001988 154580 1002008
rect 154580 1001988 154632 1002008
rect 154632 1001988 154634 1002008
rect 154578 1001952 154634 1001988
rect 154946 1001972 155002 1002008
rect 154946 1001952 154948 1001972
rect 154948 1001952 155000 1001972
rect 155000 1001952 155002 1001972
rect 152462 995016 152518 995072
rect 151082 994744 151138 994800
rect 157798 1001972 157854 1002008
rect 157798 1001952 157800 1001972
rect 157800 1001952 157852 1001972
rect 157852 1001952 157854 1001972
rect 155222 994472 155278 994528
rect 208398 1006204 208400 1006224
rect 208400 1006204 208452 1006224
rect 208452 1006204 208454 1006224
rect 208398 1006168 208454 1006204
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 195242 996648 195298 996704
rect 188066 995696 188122 995752
rect 189354 995696 189410 995752
rect 192482 995696 192538 995752
rect 193126 995696 193182 995752
rect 195058 995696 195114 995752
rect 183834 995424 183890 995480
rect 187606 994880 187662 994936
rect 188802 994608 188858 994664
rect 184846 994336 184902 994392
rect 194690 994608 194746 994664
rect 202694 1005252 202696 1005272
rect 202696 1005252 202748 1005272
rect 202748 1005252 202750 1005272
rect 202694 1005216 202750 1005252
rect 209226 1005100 209282 1005136
rect 209226 1005080 209228 1005100
rect 209228 1005080 209280 1005100
rect 209280 1005080 209282 1005100
rect 207570 1004964 207626 1005000
rect 207570 1004944 207572 1004964
rect 207572 1004944 207624 1004964
rect 207624 1004944 207626 1004964
rect 209226 1004692 209282 1004728
rect 209226 1004672 209228 1004692
rect 209228 1004672 209280 1004692
rect 209280 1004672 209282 1004692
rect 206374 1002244 206430 1002280
rect 206374 1002224 206376 1002244
rect 206376 1002224 206428 1002244
rect 206428 1002224 206430 1002244
rect 195702 997192 195758 997248
rect 195518 995968 195574 996024
rect 195058 994336 195114 994392
rect 196806 996376 196862 996432
rect 190366 994064 190422 994120
rect 200670 998164 200726 998200
rect 200670 998144 200672 998164
rect 200672 998144 200724 998164
rect 200724 998144 200726 998164
rect 202694 998300 202750 998336
rect 202694 998280 202696 998300
rect 202696 998280 202748 998300
rect 202748 998280 202750 998300
rect 201866 998028 201922 998064
rect 201866 998008 201868 998028
rect 201868 998008 201920 998028
rect 201920 998008 201922 998028
rect 200210 996412 200212 996432
rect 200212 996412 200264 996432
rect 200264 996412 200266 996432
rect 200210 996376 200266 996412
rect 202326 995424 202382 995480
rect 205546 1002108 205602 1002144
rect 205546 1002088 205548 1002108
rect 205548 1002088 205600 1002108
rect 205600 1002088 205602 1002108
rect 203522 998572 203578 998608
rect 203522 998552 203524 998572
rect 203524 998552 203576 998572
rect 203576 998552 203578 998572
rect 203522 997772 203524 997792
rect 203524 997772 203576 997792
rect 203576 997772 203578 997792
rect 203522 997736 203578 997772
rect 204350 998708 204406 998744
rect 204350 998688 204352 998708
rect 204352 998688 204404 998708
rect 204404 998688 204406 998708
rect 203890 998436 203946 998472
rect 203890 998416 203892 998436
rect 203892 998416 203944 998436
rect 203944 998416 203946 998436
rect 204718 997908 204720 997928
rect 204720 997908 204772 997928
rect 204772 997908 204774 997928
rect 204718 997872 204774 997908
rect 204074 995832 204130 995888
rect 203338 994880 203394 994936
rect 206374 1001952 206430 1002008
rect 206742 1001972 206798 1002008
rect 206742 1001952 206744 1001972
rect 206744 1001952 206796 1001972
rect 206796 1001952 206798 1001972
rect 207570 1001952 207626 1002008
rect 208398 1001952 208454 1002008
rect 210054 1002244 210110 1002280
rect 210054 1002224 210056 1002244
rect 210056 1002224 210108 1002244
rect 210108 1002224 210110 1002244
rect 210422 1001952 210478 1002008
rect 211250 1002380 211306 1002416
rect 211250 1002360 211252 1002380
rect 211252 1002360 211304 1002380
rect 211304 1002360 211306 1002380
rect 211250 1002108 211306 1002144
rect 211250 1002088 211252 1002108
rect 211252 1002088 211304 1002108
rect 211304 1002088 211306 1002108
rect 212538 1004692 212594 1004728
rect 212538 1004672 212540 1004692
rect 212540 1004672 212592 1004692
rect 212592 1004672 212594 1004692
rect 212078 1001972 212134 1002008
rect 212078 1001952 212080 1001972
rect 212080 1001952 212132 1001972
rect 212132 1001952 212134 1001972
rect 200762 994064 200818 994120
rect 256146 1006324 256202 1006360
rect 256146 1006304 256148 1006324
rect 256148 1006304 256200 1006324
rect 256200 1006304 256202 1006324
rect 229006 997192 229062 997248
rect 229190 997192 229246 997248
rect 238574 995696 238630 995752
rect 239586 995696 239642 995752
rect 242070 995696 242126 995752
rect 243266 995696 243322 995752
rect 243818 995560 243874 995616
rect 244094 995560 244150 995616
rect 235906 995424 235962 995480
rect 236550 994880 236606 994936
rect 245566 995288 245622 995344
rect 240874 994608 240930 994664
rect 246762 996376 246818 996432
rect 247222 997056 247278 997112
rect 247038 995560 247094 995616
rect 246578 995288 246634 995344
rect 247866 996104 247922 996160
rect 247682 994608 247738 994664
rect 252466 1006188 252522 1006224
rect 252466 1006168 252468 1006188
rect 252468 1006168 252520 1006188
rect 252520 1006168 252522 1006188
rect 262678 1006188 262734 1006224
rect 262678 1006168 262680 1006188
rect 262680 1006168 262732 1006188
rect 262732 1006168 262734 1006188
rect 254122 1006052 254178 1006088
rect 254122 1006032 254124 1006052
rect 254124 1006032 254176 1006052
rect 254176 1006032 254178 1006052
rect 261850 1006052 261906 1006088
rect 261850 1006032 261852 1006052
rect 261852 1006032 261904 1006052
rect 261904 1006032 261906 1006052
rect 263046 1005252 263048 1005272
rect 263048 1005252 263100 1005272
rect 263100 1005252 263102 1005272
rect 263046 1005216 263102 1005252
rect 256514 1004692 256570 1004728
rect 256514 1004672 256516 1004692
rect 256516 1004672 256568 1004692
rect 256568 1004672 256570 1004692
rect 249890 996784 249946 996840
rect 255318 1002788 255374 1002824
rect 255318 1002768 255320 1002788
rect 255320 1002768 255372 1002788
rect 255372 1002768 255374 1002788
rect 255318 1002532 255320 1002552
rect 255320 1002532 255372 1002552
rect 255372 1002532 255374 1002552
rect 255318 1002496 255374 1002532
rect 261022 1002516 261078 1002552
rect 261022 1002496 261024 1002516
rect 261024 1002496 261076 1002516
rect 261076 1002496 261078 1002516
rect 254490 1002244 254546 1002280
rect 254490 1002224 254492 1002244
rect 254492 1002224 254544 1002244
rect 254544 1002224 254546 1002244
rect 256146 1002108 256202 1002144
rect 256146 1002088 256148 1002108
rect 256148 1002088 256200 1002108
rect 256200 1002088 256202 1002108
rect 263506 1002108 263562 1002144
rect 263506 1002088 263508 1002108
rect 263508 1002088 263560 1002108
rect 263560 1002088 263562 1002108
rect 253294 998028 253350 998064
rect 253294 998008 253296 998028
rect 253296 998008 253348 998028
rect 253348 998008 253350 998028
rect 252466 997892 252522 997928
rect 252466 997872 252468 997892
rect 252468 997872 252520 997892
rect 252520 997872 252522 997892
rect 261022 1001972 261078 1002008
rect 261022 1001952 261024 1001972
rect 261024 1001952 261076 1001972
rect 261076 1001952 261078 1001972
rect 263874 1001972 263930 1002008
rect 263874 1001952 263876 1001972
rect 263876 1001952 263928 1001972
rect 263928 1001952 263930 1001972
rect 256974 1001172 256976 1001192
rect 256976 1001172 257028 1001192
rect 257028 1001172 257030 1001192
rect 256974 1001136 257030 1001172
rect 258998 998436 259054 998472
rect 258998 998416 259000 998436
rect 259000 998416 259052 998436
rect 259052 998416 259054 998436
rect 253662 998164 253718 998200
rect 257342 998180 257344 998200
rect 257344 998180 257396 998200
rect 257396 998180 257398 998200
rect 253662 998144 253664 998164
rect 253664 998144 253716 998164
rect 253716 998144 253718 998164
rect 257342 998144 257398 998180
rect 258170 998044 258172 998064
rect 258172 998044 258224 998064
rect 258224 998044 258226 998064
rect 253478 995832 253534 995888
rect 251822 994880 251878 994936
rect 258170 998008 258226 998044
rect 260194 998044 260196 998064
rect 260196 998044 260248 998064
rect 260248 998044 260250 998064
rect 260194 998008 260250 998044
rect 258998 997908 259000 997928
rect 259000 997908 259052 997928
rect 259052 997908 259054 997928
rect 258998 997872 259054 997908
rect 259826 997908 259828 997928
rect 259828 997908 259880 997928
rect 259880 997908 259882 997928
rect 259826 997872 259882 997908
rect 258170 997772 258172 997792
rect 258172 997772 258224 997792
rect 258224 997772 258226 997792
rect 258170 997736 258226 997772
rect 260194 997772 260196 997792
rect 260196 997772 260248 997792
rect 260248 997772 260250 997792
rect 260194 997736 260250 997772
rect 261850 997736 261906 997792
rect 298098 1002224 298154 1002280
rect 298282 997872 298338 997928
rect 292486 995696 292542 995752
rect 295062 995696 295118 995752
rect 296166 995696 296222 995752
rect 298098 995696 298154 995752
rect 280710 995560 280766 995616
rect 290278 995016 290334 995072
rect 287794 994744 287850 994800
rect 294878 995424 294934 995480
rect 307758 1006460 307814 1006496
rect 307758 1006440 307760 1006460
rect 307760 1006440 307812 1006460
rect 307812 1006440 307814 1006460
rect 360198 1006460 360254 1006496
rect 360198 1006440 360200 1006460
rect 360200 1006440 360252 1006460
rect 360252 1006440 360254 1006460
rect 299110 996376 299166 996432
rect 298926 995968 298982 996024
rect 291474 994200 291530 994256
rect 298650 995424 298706 995480
rect 314658 1006324 314714 1006360
rect 314658 1006304 314660 1006324
rect 314660 1006304 314712 1006324
rect 314712 1006304 314714 1006324
rect 360566 1006324 360622 1006360
rect 360566 1006304 360568 1006324
rect 360568 1006304 360620 1006324
rect 360620 1006304 360622 1006324
rect 306102 1006188 306158 1006224
rect 306102 1006168 306104 1006188
rect 306104 1006168 306156 1006188
rect 306156 1006168 306158 1006188
rect 304078 1006052 304134 1006088
rect 304078 1006032 304080 1006052
rect 304080 1006032 304132 1006052
rect 304132 1006032 304134 1006052
rect 311806 1006032 311862 1006088
rect 314658 1006052 314714 1006088
rect 314658 1006032 314660 1006052
rect 314660 1006032 314712 1006052
rect 314712 1006032 314714 1006052
rect 313830 1004828 313886 1004864
rect 313830 1004808 313832 1004828
rect 313832 1004808 313884 1004828
rect 313884 1004808 313886 1004828
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 302146 1002224 302202 1002280
rect 310978 1002108 311034 1002144
rect 310978 1002088 310980 1002108
rect 310980 1002088 311032 1002108
rect 311032 1002088 311034 1002108
rect 310150 1001972 310206 1002008
rect 310150 1001952 310152 1001972
rect 310152 1001952 310204 1001972
rect 310204 1001952 310206 1001972
rect 312634 1001972 312690 1002008
rect 312634 1001952 312636 1001972
rect 312636 1001952 312688 1001972
rect 312688 1001952 312690 1001972
rect 305274 999132 305276 999152
rect 305276 999132 305328 999152
rect 305328 999132 305330 999152
rect 305274 999096 305330 999132
rect 308954 998572 309010 998608
rect 308954 998552 308956 998572
rect 308956 998552 309008 998572
rect 309008 998552 309010 998572
rect 302146 995560 302202 995616
rect 300122 994744 300178 994800
rect 287518 993928 287574 993984
rect 298006 993928 298062 993984
rect 307298 998436 307354 998472
rect 307298 998416 307300 998436
rect 307300 998416 307352 998436
rect 307352 998416 307354 998436
rect 303250 997872 303306 997928
rect 306102 998300 306158 998336
rect 306102 998280 306104 998300
rect 306104 998280 306156 998300
rect 306156 998280 306158 998300
rect 310610 998280 310666 998336
rect 308126 998164 308182 998200
rect 308126 998144 308128 998164
rect 308128 998144 308180 998164
rect 308180 998144 308182 998164
rect 304906 997892 304962 997928
rect 304906 997872 304908 997892
rect 304908 997872 304960 997892
rect 304960 997872 304962 997892
rect 306930 998028 306986 998064
rect 306930 998008 306932 998028
rect 306932 998008 306984 998028
rect 306984 998008 306986 998028
rect 307022 995016 307078 995072
rect 308954 997892 309010 997928
rect 308954 997872 308956 997892
rect 308956 997872 309008 997892
rect 309008 997872 309010 997892
rect 309782 997736 309838 997792
rect 310610 998028 310666 998064
rect 310610 998008 310612 998028
rect 310612 998008 310664 998028
rect 310664 998008 310666 998028
rect 354862 1006052 354918 1006088
rect 354862 1006032 354864 1006052
rect 354864 1006032 354916 1006052
rect 354916 1006032 354918 1006052
rect 355690 1006052 355746 1006088
rect 355690 1006032 355692 1006052
rect 355692 1006032 355744 1006052
rect 355744 1006032 355746 1006052
rect 361394 1006052 361450 1006088
rect 361394 1006032 361396 1006052
rect 361396 1006032 361448 1006052
rect 361448 1006032 361450 1006052
rect 365074 1006052 365130 1006088
rect 365074 1006032 365076 1006052
rect 365076 1006032 365128 1006052
rect 365128 1006032 365130 1006052
rect 304262 994200 304318 994256
rect 355690 1004828 355746 1004864
rect 355690 1004808 355692 1004828
rect 355692 1004808 355744 1004828
rect 355744 1004808 355746 1004828
rect 356518 1003892 356520 1003912
rect 356520 1003892 356572 1003912
rect 356572 1003892 356574 1003912
rect 356518 1003856 356574 1003892
rect 354034 1001972 354090 1002008
rect 354034 1001952 354036 1001972
rect 354036 1001952 354088 1001972
rect 354088 1001952 354090 1001972
rect 358542 1002108 358598 1002144
rect 358542 1002088 358544 1002108
rect 358544 1002088 358596 1002108
rect 358596 1002088 358598 1002108
rect 356518 1001972 356574 1002008
rect 356518 1001952 356520 1001972
rect 356520 1001952 356572 1001972
rect 356572 1001952 356574 1001972
rect 357346 1001972 357402 1002008
rect 357346 1001952 357348 1001972
rect 357348 1001952 357400 1001972
rect 357400 1001952 357402 1001972
rect 359370 1001952 359426 1002008
rect 360566 1005252 360568 1005272
rect 360568 1005252 360620 1005272
rect 360620 1005252 360622 1005272
rect 360566 1005216 360622 1005252
rect 363418 1005100 363474 1005136
rect 363418 1005080 363420 1005100
rect 363420 1005080 363472 1005100
rect 363472 1005080 363474 1005100
rect 365074 1004964 365130 1005000
rect 365074 1004944 365076 1004964
rect 365076 1004944 365128 1004964
rect 365128 1004944 365130 1004964
rect 362590 1004828 362646 1004864
rect 362590 1004808 362592 1004828
rect 362592 1004808 362644 1004828
rect 362644 1004808 362646 1004828
rect 364246 1004692 364302 1004728
rect 364246 1004672 364248 1004692
rect 364248 1004672 364300 1004692
rect 364300 1004672 364302 1004692
rect 359738 1002108 359794 1002144
rect 359738 1002088 359740 1002108
rect 359740 1002088 359792 1002108
rect 359792 1002088 359794 1002108
rect 361394 1001972 361450 1002008
rect 361394 1001952 361396 1001972
rect 361396 1001952 361448 1001972
rect 361448 1001952 361450 1001972
rect 425518 1007004 425574 1007040
rect 505374 1007020 505376 1007040
rect 505376 1007020 505428 1007040
rect 505428 1007020 505430 1007040
rect 425518 1006984 425520 1007004
rect 425520 1006984 425572 1007004
rect 425572 1006984 425574 1007004
rect 505374 1006984 505430 1007020
rect 365902 1001972 365958 1002008
rect 365902 1001952 365904 1001972
rect 365904 1001952 365956 1001972
rect 365956 1001952 365958 1001972
rect 427542 1006868 427598 1006904
rect 427542 1006848 427544 1006868
rect 427544 1006848 427596 1006868
rect 427596 1006848 427598 1006868
rect 430854 1006732 430910 1006768
rect 430854 1006712 430856 1006732
rect 430856 1006712 430908 1006732
rect 430908 1006712 430910 1006732
rect 372342 996376 372398 996432
rect 374642 995016 374698 995072
rect 376022 996920 376078 996976
rect 375562 994744 375618 994800
rect 383290 997600 383346 997656
rect 383474 997192 383530 997248
rect 383106 995696 383162 995752
rect 381450 995288 381506 995344
rect 385038 995696 385094 995752
rect 385774 995696 385830 995752
rect 387890 995696 387946 995752
rect 388718 995696 388774 995752
rect 389362 995696 389418 995752
rect 392398 995696 392454 995752
rect 396538 995696 396594 995752
rect 392306 995288 392362 995344
rect 388350 995016 388406 995072
rect 393502 995288 393558 995344
rect 395158 994744 395214 994800
rect 429198 1006596 429254 1006632
rect 429198 1006576 429200 1006596
rect 429200 1006576 429252 1006596
rect 429252 1006576 429254 1006596
rect 425150 1006324 425206 1006360
rect 425150 1006304 425152 1006324
rect 425152 1006304 425204 1006324
rect 425204 1006304 425206 1006324
rect 423494 1006188 423550 1006224
rect 423494 1006168 423496 1006188
rect 423496 1006168 423548 1006188
rect 423548 1006168 423550 1006188
rect 422666 1006052 422722 1006088
rect 422666 1006032 422668 1006052
rect 422668 1006032 422720 1006052
rect 422720 1006032 422722 1006052
rect 430026 1006052 430082 1006088
rect 430026 1006032 430028 1006052
rect 430028 1006032 430080 1006052
rect 430080 1006032 430082 1006052
rect 423494 1005660 423496 1005680
rect 423496 1005660 423548 1005680
rect 423548 1005660 423550 1005680
rect 423494 1005624 423550 1005660
rect 428370 1005524 428372 1005544
rect 428372 1005524 428424 1005544
rect 428424 1005524 428426 1005544
rect 428370 1005488 428426 1005524
rect 427174 1005372 427230 1005408
rect 427174 1005352 427176 1005372
rect 427176 1005352 427228 1005372
rect 427228 1005352 427230 1005372
rect 429198 1004964 429254 1005000
rect 429198 1004944 429200 1004964
rect 429200 1004944 429252 1004964
rect 429252 1004944 429254 1004964
rect 421470 1001972 421526 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 421010 996412 421012 996432
rect 421012 996412 421064 996432
rect 421064 996412 421066 996432
rect 421010 996376 421066 996412
rect 422666 1004672 422722 1004728
rect 424690 1002668 424692 1002688
rect 424692 1002668 424744 1002688
rect 424744 1002668 424746 1002688
rect 424690 1002632 424746 1002668
rect 426346 1002532 426348 1002552
rect 426348 1002532 426400 1002552
rect 426400 1002532 426402 1002552
rect 426346 1002496 426402 1002532
rect 428002 1002244 428058 1002280
rect 428002 1002224 428004 1002244
rect 428004 1002224 428056 1002244
rect 428056 1002224 428058 1002244
rect 425150 1002108 425206 1002144
rect 425150 1002088 425152 1002108
rect 425152 1002088 425204 1002108
rect 425204 1002088 425206 1002108
rect 428370 1002108 428426 1002144
rect 428370 1002088 428372 1002108
rect 428372 1002088 428424 1002108
rect 428424 1002088 428426 1002108
rect 424322 1001972 424378 1002008
rect 424322 1001952 424324 1001972
rect 424324 1001952 424376 1001972
rect 424376 1001952 424378 1001972
rect 426346 1001972 426402 1002008
rect 426346 1001952 426348 1001972
rect 426348 1001952 426400 1001972
rect 426400 1001952 426402 1001972
rect 432050 1005796 432052 1005816
rect 432052 1005796 432104 1005816
rect 432104 1005796 432106 1005816
rect 432050 1005760 432106 1005796
rect 430854 1005236 430910 1005272
rect 430854 1005216 430856 1005236
rect 430856 1005216 430908 1005236
rect 430908 1005216 430910 1005236
rect 432050 1005116 432052 1005136
rect 432052 1005116 432104 1005136
rect 432104 1005116 432106 1005136
rect 432050 1005080 432106 1005116
rect 431682 1004828 431738 1004864
rect 431682 1004808 431684 1004828
rect 431684 1004808 431736 1004828
rect 431736 1004808 431738 1004828
rect 430026 1004692 430082 1004728
rect 430026 1004672 430028 1004692
rect 430028 1004672 430080 1004692
rect 430080 1004672 430082 1004692
rect 433338 1002108 433394 1002144
rect 433338 1002088 433340 1002108
rect 433340 1002088 433392 1002108
rect 433392 1002088 433394 1002108
rect 432878 1001972 432934 1002008
rect 432878 1001952 432880 1001972
rect 432880 1001952 432932 1001972
rect 432932 1001952 432934 1001972
rect 503350 1006884 503352 1006904
rect 503352 1006884 503404 1006904
rect 503404 1006884 503406 1006904
rect 503350 1006848 503406 1006884
rect 506202 1006612 506204 1006632
rect 506204 1006612 506256 1006632
rect 506256 1006612 506258 1006632
rect 506202 1006576 506258 1006612
rect 439686 998280 439742 998336
rect 439686 996648 439742 996704
rect 439870 996376 439926 996432
rect 449162 996104 449218 996160
rect 446862 994880 446918 994936
rect 462318 995832 462374 995888
rect 452290 994608 452346 994664
rect 505374 1006476 505376 1006496
rect 505376 1006476 505428 1006496
rect 505428 1006476 505430 1006496
rect 505374 1006440 505430 1006476
rect 502154 1006324 502210 1006360
rect 502154 1006304 502156 1006324
rect 502156 1006304 502208 1006324
rect 502208 1006304 502210 1006324
rect 508226 1006188 508282 1006224
rect 508226 1006168 508228 1006188
rect 508228 1006168 508280 1006188
rect 508280 1006168 508282 1006188
rect 498842 1006052 498898 1006088
rect 498842 1006032 498844 1006052
rect 498844 1006032 498896 1006052
rect 498896 1006032 498898 1006052
rect 501326 1006052 501382 1006088
rect 501326 1006032 501328 1006052
rect 501328 1006032 501380 1006052
rect 501380 1006032 501382 1006052
rect 509054 1006052 509110 1006088
rect 509054 1006032 509056 1006052
rect 509056 1006032 509108 1006052
rect 509108 1006032 509110 1006052
rect 472070 995152 472126 995208
rect 473358 995696 473414 995752
rect 475934 995696 475990 995752
rect 476486 995696 476542 995752
rect 477038 995696 477094 995752
rect 485686 995696 485742 995752
rect 488906 995696 488962 995752
rect 480810 995424 480866 995480
rect 478234 995152 478290 995208
rect 478786 995152 478842 995208
rect 475750 994880 475806 994936
rect 466458 994336 466514 994392
rect 481546 995152 481602 995208
rect 487802 994880 487858 994936
rect 484122 994608 484178 994664
rect 482926 994336 482982 994392
rect 475750 994064 475806 994120
rect 499670 1004828 499726 1004864
rect 499670 1004808 499672 1004828
rect 499672 1004808 499724 1004828
rect 499724 1004808 499726 1004828
rect 500498 1004692 500554 1004728
rect 500498 1004672 500500 1004692
rect 500500 1004672 500552 1004692
rect 500552 1004672 500554 1004692
rect 498474 1001972 498530 1002008
rect 498474 1001952 498476 1001972
rect 498476 1001952 498528 1001972
rect 498528 1001952 498530 1001972
rect 504546 1004436 504548 1004456
rect 504548 1004436 504600 1004456
rect 504600 1004436 504602 1004456
rect 504546 1004400 504602 1004436
rect 501694 1002516 501750 1002552
rect 501694 1002496 501696 1002516
rect 501696 1002496 501748 1002516
rect 501748 1002496 501750 1002516
rect 502154 1002380 502210 1002416
rect 502154 1002360 502156 1002380
rect 502156 1002360 502208 1002380
rect 502208 1002360 502210 1002380
rect 500498 1002244 500554 1002280
rect 500498 1002224 500500 1002244
rect 500500 1002224 500552 1002244
rect 500552 1002224 500554 1002244
rect 502522 1002108 502578 1002144
rect 502522 1002088 502524 1002108
rect 502524 1002088 502576 1002108
rect 502576 1002088 502578 1002108
rect 503350 1001972 503406 1002008
rect 503350 1001952 503352 1001972
rect 503352 1001952 503404 1001972
rect 503404 1001952 503406 1001972
rect 504178 1001972 504234 1002008
rect 504178 1001952 504180 1001972
rect 504180 1001952 504232 1001972
rect 504232 1001952 504234 1001972
rect 506202 1001972 506258 1002008
rect 506202 1001952 506204 1001972
rect 506204 1001952 506256 1001972
rect 506256 1001952 506258 1001972
rect 507030 1005236 507086 1005272
rect 507030 1005216 507032 1005236
rect 507032 1005216 507084 1005236
rect 507084 1005216 507086 1005236
rect 508226 1005100 508282 1005136
rect 508226 1005080 508228 1005100
rect 508228 1005080 508280 1005100
rect 508280 1005080 508282 1005100
rect 507858 1004964 507914 1005000
rect 507858 1004944 507860 1004964
rect 507860 1004944 507912 1004964
rect 507912 1004944 507914 1004964
rect 507398 1004828 507454 1004864
rect 507398 1004808 507400 1004828
rect 507400 1004808 507452 1004828
rect 507452 1004808 507454 1004828
rect 509054 1004692 509110 1004728
rect 509054 1004672 509056 1004692
rect 509056 1004672 509108 1004692
rect 509108 1004672 509110 1004692
rect 509882 1002244 509938 1002280
rect 509882 1002224 509884 1002244
rect 509884 1002224 509936 1002244
rect 509936 1002224 509938 1002244
rect 510342 1002108 510398 1002144
rect 510342 1002088 510344 1002108
rect 510344 1002088 510396 1002108
rect 510396 1002088 510398 1002108
rect 551098 1007004 551154 1007040
rect 551098 1006984 551100 1007004
rect 551100 1006984 551152 1007004
rect 551152 1006984 551154 1007004
rect 517242 998552 517298 998608
rect 516874 996376 516930 996432
rect 516690 996104 516746 996160
rect 518162 994744 518218 994800
rect 559654 1006868 559710 1006904
rect 559654 1006848 559656 1006868
rect 559656 1006848 559708 1006868
rect 559708 1006848 559710 1006868
rect 553122 1006460 553178 1006496
rect 553122 1006440 553124 1006460
rect 553124 1006440 553176 1006460
rect 553176 1006440 553178 1006460
rect 553950 1005388 553952 1005408
rect 553952 1005388 554004 1005408
rect 554004 1005388 554006 1005408
rect 553950 1005352 554006 1005388
rect 552294 1005252 552296 1005272
rect 552296 1005252 552348 1005272
rect 552348 1005252 552350 1005272
rect 552294 1005216 552350 1005252
rect 523130 995152 523186 995208
rect 523498 998552 523554 998608
rect 523682 995696 523738 995752
rect 551098 998028 551154 998064
rect 551098 998008 551100 998028
rect 551100 998008 551152 998028
rect 551152 998008 551154 998028
rect 524050 996648 524106 996704
rect 524786 995696 524842 995752
rect 529846 995696 529902 995752
rect 536562 995696 536618 995752
rect 537206 995696 537262 995752
rect 523498 995424 523554 995480
rect 527914 995424 527970 995480
rect 526258 995172 526314 995208
rect 526258 995152 526260 995172
rect 526260 995152 526312 995172
rect 526312 995152 526314 995172
rect 533434 995424 533490 995480
rect 537850 995424 537906 995480
rect 535550 994744 535606 994800
rect 538218 995424 538274 995480
rect 550270 997892 550326 997928
rect 550270 997872 550272 997892
rect 550272 997872 550324 997892
rect 550324 997872 550326 997892
rect 551466 997736 551522 997792
rect 552294 997736 552350 997792
rect 553306 997892 553362 997928
rect 553306 997872 553308 997892
rect 553308 997872 553360 997892
rect 553360 997872 553362 997892
rect 555974 1006732 556030 1006768
rect 555974 1006712 555976 1006732
rect 555976 1006712 556028 1006732
rect 556028 1006712 556030 1006732
rect 556802 1006324 556858 1006360
rect 556802 1006304 556804 1006324
rect 556804 1006304 556856 1006324
rect 556856 1006304 556858 1006324
rect 557170 1006188 557226 1006224
rect 557170 1006168 557172 1006188
rect 557172 1006168 557224 1006188
rect 557224 1006168 557226 1006188
rect 555146 1005524 555148 1005544
rect 555148 1005524 555200 1005544
rect 555200 1005524 555202 1005544
rect 555146 1005488 555202 1005524
rect 555974 1004828 556030 1004864
rect 555974 1004808 555976 1004828
rect 555976 1004808 556028 1004828
rect 556028 1004808 556030 1004828
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 557998 1002380 558054 1002416
rect 557998 1002360 558000 1002380
rect 558000 1002360 558052 1002380
rect 558052 1002360 558054 1002380
rect 554318 1002244 554374 1002280
rect 554318 1002224 554320 1002244
rect 554320 1002224 554372 1002244
rect 554372 1002224 554374 1002244
rect 555146 1002108 555202 1002144
rect 555146 1002088 555148 1002108
rect 555148 1002088 555200 1002108
rect 555200 1002088 555202 1002108
rect 557998 1002108 558054 1002144
rect 557998 1002088 558000 1002108
rect 558000 1002088 558052 1002108
rect 558052 1002088 558054 1002108
rect 554318 1001972 554374 1002008
rect 554318 1001952 554320 1001972
rect 554320 1001952 554372 1001972
rect 554372 1001952 554374 1001972
rect 558826 1002516 558882 1002552
rect 558826 1002496 558828 1002516
rect 558828 1002496 558880 1002516
rect 558880 1002496 558882 1002516
rect 558826 1001972 558882 1002008
rect 558826 1001952 558828 1001972
rect 558828 1001952 558880 1001972
rect 558880 1001952 558882 1001972
rect 560850 1005660 560852 1005680
rect 560852 1005660 560904 1005680
rect 560904 1005660 560906 1005680
rect 560850 1005624 560906 1005660
rect 560482 1002380 560538 1002416
rect 560482 1002360 560484 1002380
rect 560484 1002360 560536 1002380
rect 560536 1002360 560538 1002380
rect 560022 1002244 560078 1002280
rect 560022 1002224 560024 1002244
rect 560024 1002224 560076 1002244
rect 560076 1002224 560078 1002244
rect 560850 1002108 560906 1002144
rect 560850 1002088 560852 1002108
rect 560852 1002088 560904 1002108
rect 560904 1002088 560906 1002108
rect 561678 1001972 561734 1002008
rect 561678 1001952 561680 1001972
rect 561680 1001952 561732 1001972
rect 561732 1001952 561734 1001972
rect 567842 993656 567898 993712
rect 590566 996668 590622 996704
rect 590566 996648 590568 996668
rect 590568 996648 590620 996668
rect 590620 996648 590622 996668
rect 590566 996376 590622 996432
rect 625434 995968 625490 996024
rect 623686 995696 623742 995752
rect 617338 995016 617394 995072
rect 626538 995696 626594 995752
rect 627182 995696 627238 995752
rect 631506 995696 631562 995752
rect 625618 995424 625674 995480
rect 630218 995424 630274 995480
rect 630862 995424 630918 995480
rect 629666 995016 629722 995072
rect 625434 994744 625490 994800
rect 576306 989440 576362 989496
rect 634726 994744 634782 994800
rect 633990 993656 634046 993712
rect 62118 975976 62174 976032
rect 62118 962920 62174 962976
rect 62118 949864 62174 949920
rect 62118 936980 62120 937000
rect 62120 936980 62172 937000
rect 62172 936980 62174 937000
rect 62118 936944 62174 936980
rect 44822 936128 44878 936184
rect 44454 934088 44510 934144
rect 44178 933680 44234 933736
rect 43442 933272 43498 933328
rect 42522 932864 42578 932920
rect 42798 932048 42854 932104
rect 42430 881864 42486 881920
rect 42062 817944 42118 818000
rect 41878 814680 41934 814736
rect 42890 814680 42946 814736
rect 41786 812776 41842 812832
rect 35162 812368 35218 812424
rect 32402 811144 32458 811200
rect 31666 809920 31722 809976
rect 33782 809512 33838 809568
rect 40958 811960 41014 812016
rect 36542 809104 36598 809160
rect 35162 803800 35218 803856
rect 41326 811588 41328 811608
rect 41328 811588 41380 811608
rect 41380 811588 41382 811608
rect 41326 811552 41382 811588
rect 40958 804752 41014 804808
rect 39762 801896 39818 801952
rect 39854 800944 39910 801000
rect 41970 810328 42026 810384
rect 42062 806656 42118 806712
rect 41786 805296 41842 805352
rect 41234 800808 41290 800864
rect 40038 800672 40094 800728
rect 42614 801896 42670 801952
rect 42338 801080 42394 801136
rect 42338 800808 42394 800864
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 42154 797272 42210 797328
rect 41786 796184 41842 796240
rect 42062 794960 42118 795016
rect 41786 794416 41842 794472
rect 41786 793464 41842 793520
rect 42154 792920 42210 792976
rect 42430 791968 42486 792024
rect 42614 790064 42670 790120
rect 42338 789112 42394 789168
rect 42246 788160 42302 788216
rect 42522 787888 42578 787944
rect 39762 775240 39818 775296
rect 35806 774324 35808 774344
rect 35808 774324 35860 774344
rect 35860 774324 35862 774344
rect 35806 774288 35862 774324
rect 35806 773880 35862 773936
rect 35346 773472 35402 773528
rect 35530 773064 35586 773120
rect 35806 773100 35808 773120
rect 35808 773100 35860 773120
rect 35860 773100 35862 773120
rect 35806 773064 35862 773100
rect 40866 773064 40922 773120
rect 35346 772248 35402 772304
rect 35530 771840 35586 771896
rect 35806 771840 35862 771896
rect 35806 771024 35862 771080
rect 35622 770616 35678 770672
rect 43258 813592 43314 813648
rect 43074 808696 43130 808752
rect 43074 773064 43130 773120
rect 39854 770616 39910 770672
rect 42890 770616 42946 770672
rect 35806 770208 35862 770264
rect 39854 770208 39910 770264
rect 35622 769392 35678 769448
rect 35806 768984 35862 769040
rect 35806 768168 35862 768224
rect 35622 767760 35678 767816
rect 32402 767352 32458 767408
rect 35162 766944 35218 767000
rect 32402 759600 32458 759656
rect 35806 766536 35862 766592
rect 35806 766128 35862 766184
rect 35806 764496 35862 764552
rect 35622 764088 35678 764144
rect 35806 763308 35808 763328
rect 35808 763308 35860 763328
rect 35860 763308 35862 763328
rect 35806 763272 35862 763308
rect 35806 762864 35862 762920
rect 39118 763680 39174 763736
rect 42522 768712 42578 768768
rect 39762 764496 39818 764552
rect 41694 763292 41750 763328
rect 41694 763272 41696 763292
rect 41696 763272 41748 763292
rect 41748 763272 41750 763292
rect 39302 757696 39358 757752
rect 42246 758376 42302 758432
rect 40222 758104 40278 758160
rect 41970 757832 42026 757888
rect 42430 757832 42486 757888
rect 39946 757424 40002 757480
rect 42246 757424 42302 757480
rect 41786 757016 41842 757072
rect 41970 755384 42026 755440
rect 42154 754840 42210 754896
rect 42062 754024 42118 754080
rect 42246 752120 42302 752176
rect 42062 751712 42118 751768
rect 41786 751032 41842 751088
rect 42246 749400 42302 749456
rect 42246 746544 42302 746600
rect 42062 746000 42118 746056
rect 42062 745456 42118 745512
rect 42430 746272 42486 746328
rect 42614 746000 42670 746056
rect 42706 745456 42762 745512
rect 42614 745048 42670 745104
rect 43258 764496 43314 764552
rect 43626 807200 43682 807256
rect 43626 797272 43682 797328
rect 44454 812776 44510 812832
rect 44638 807880 44694 807936
rect 44638 794960 44694 795016
rect 46202 819032 46258 819088
rect 46202 806248 46258 806304
rect 44822 775240 44878 775296
rect 44270 770208 44326 770264
rect 43442 754024 43498 754080
rect 43442 751712 43498 751768
rect 43258 730904 43314 730960
rect 43442 730496 43498 730552
rect 43074 730088 43130 730144
rect 42890 729272 42946 729328
rect 40866 728626 40922 728682
rect 41326 728680 41382 728682
rect 41326 728628 41328 728680
rect 41328 728628 41380 728680
rect 41380 728628 41382 728680
rect 41326 728626 41382 728628
rect 42890 728048 42946 728104
rect 41050 727456 41106 727458
rect 41050 727404 41052 727456
rect 41052 727404 41104 727456
rect 41104 727404 41106 727456
rect 41050 727402 41106 727404
rect 41326 726824 41382 726880
rect 42522 726416 42578 726472
rect 40958 726178 41014 726234
rect 37922 725192 37978 725248
rect 35162 724784 35218 724840
rect 33046 724376 33102 724432
rect 31758 720316 31814 720352
rect 31758 720296 31760 720316
rect 31760 720296 31812 720316
rect 31812 720296 31814 720316
rect 33782 723730 33838 723786
rect 33046 716760 33102 716816
rect 40682 723152 40738 723208
rect 40314 714856 40370 714912
rect 41786 725736 41842 725792
rect 41326 725600 41382 725656
rect 41142 721712 41198 721768
rect 41786 722336 41842 722392
rect 42338 719888 42394 719944
rect 41786 718528 41842 718584
rect 41326 718256 41382 718312
rect 42338 718256 42394 718312
rect 42522 715128 42578 715184
rect 42338 714856 42394 714912
rect 40682 714176 40738 714232
rect 41786 713904 41842 713960
rect 41786 713496 41842 713552
rect 42154 711592 42210 711648
rect 41786 709824 41842 709880
rect 41786 708464 41842 708520
rect 41878 707104 41934 707160
rect 42246 706152 42302 706208
rect 42246 703704 42302 703760
rect 42062 703432 42118 703488
rect 42062 703024 42118 703080
rect 43258 723560 43314 723616
rect 42706 703024 42762 703080
rect 42614 702344 42670 702400
rect 42430 701800 42486 701856
rect 40958 688336 41014 688392
rect 41142 686840 41198 686896
rect 40866 685854 40922 685910
rect 41326 685908 41382 685910
rect 41326 685856 41328 685908
rect 41328 685856 41380 685908
rect 41380 685856 41382 685908
rect 41326 685854 41382 685856
rect 41142 685208 41198 685264
rect 42706 684800 42762 684856
rect 40958 683576 41014 683632
rect 40774 682760 40830 682816
rect 40590 682352 40646 682408
rect 37922 681944 37978 682000
rect 36542 681536 36598 681592
rect 32402 681128 32458 681184
rect 33782 680720 33838 680776
rect 32402 672696 32458 672752
rect 41326 683168 41382 683224
rect 41786 682352 41842 682408
rect 41786 678816 41842 678872
rect 41142 677048 41198 677104
rect 41142 672424 41198 672480
rect 42246 672152 42302 672208
rect 39486 671472 39542 671528
rect 40038 671236 40040 671256
rect 40040 671236 40092 671256
rect 40092 671236 40094 671256
rect 40038 671200 40094 671236
rect 43166 703432 43222 703488
rect 43258 687656 43314 687712
rect 43442 687248 43498 687304
rect 43074 684392 43130 684448
rect 43258 683984 43314 684040
rect 42706 671472 42762 671528
rect 42706 671200 42762 671256
rect 41786 669024 41842 669080
rect 42062 667664 42118 667720
rect 42430 667392 42486 667448
rect 42062 665080 42118 665136
rect 41786 664128 41842 664184
rect 42154 662768 42210 662824
rect 42614 660320 42670 660376
rect 42430 658824 42486 658880
rect 42246 658552 42302 658608
rect 39394 646040 39450 646096
rect 35530 644680 35586 644736
rect 35806 644716 35808 644736
rect 35808 644716 35860 644736
rect 35860 644716 35862 644736
rect 35806 644680 35862 644716
rect 39762 644680 39818 644736
rect 35346 643864 35402 643920
rect 39854 643864 39910 643920
rect 35530 643456 35586 643512
rect 35806 643492 35808 643512
rect 35808 643492 35860 643512
rect 35860 643492 35862 643512
rect 35806 643456 35862 643492
rect 39670 643492 39672 643512
rect 39672 643492 39724 643512
rect 39724 643492 39726 643512
rect 39670 643456 39726 643492
rect 39578 643048 39634 643104
rect 35438 642640 35494 642696
rect 35622 642232 35678 642288
rect 38934 642252 38990 642288
rect 38934 642232 38936 642252
rect 38936 642232 38988 642252
rect 38988 642232 38990 642252
rect 35806 641824 35862 641880
rect 35806 641416 35862 641472
rect 35622 641008 35678 641064
rect 35806 640600 35862 640656
rect 43442 680312 43498 680368
rect 43258 678272 43314 678328
rect 43258 665080 43314 665136
rect 44454 729680 44510 729736
rect 44178 722744 44234 722800
rect 43626 667664 43682 667720
rect 43074 643864 43130 643920
rect 42890 642232 42946 642288
rect 39670 640192 39726 640248
rect 35346 639784 35402 639840
rect 33782 638560 33838 638616
rect 32402 638152 32458 638208
rect 35530 639376 35586 639432
rect 35806 639376 35862 639432
rect 35530 637744 35586 637800
rect 35806 637764 35862 637800
rect 35806 637744 35808 637764
rect 35808 637744 35860 637764
rect 35860 637744 35862 637764
rect 40038 637336 40094 637392
rect 35806 636520 35862 636576
rect 41510 638152 41566 638208
rect 40958 637744 41014 637800
rect 35622 635296 35678 635352
rect 40222 635296 40278 635352
rect 35806 634888 35862 634944
rect 39578 634888 39634 634944
rect 35806 634480 35862 634536
rect 35806 633664 35862 633720
rect 40682 634480 40738 634536
rect 42338 633800 42394 633856
rect 40498 632032 40554 632088
rect 42338 625368 42394 625424
rect 42154 624552 42210 624608
rect 42154 623328 42210 623384
rect 42062 620880 42118 620936
rect 42890 624552 42946 624608
rect 43258 640192 43314 640248
rect 42062 620200 42118 620256
rect 42706 620200 42762 620256
rect 42246 619792 42302 619848
rect 42430 618976 42486 619032
rect 42706 618704 42762 618760
rect 42246 615984 42302 616040
rect 41786 612720 41842 612776
rect 35806 601724 35862 601760
rect 35806 601704 35808 601724
rect 35808 601704 35860 601724
rect 35860 601704 35862 601724
rect 41326 599256 41382 599312
rect 40866 598848 40922 598904
rect 42706 598440 42762 598496
rect 41050 597848 41106 597850
rect 41050 597796 41052 597848
rect 41052 597796 41104 597848
rect 41104 597796 41106 597848
rect 41050 597794 41106 597796
rect 41326 597794 41382 597850
rect 41142 597216 41198 597272
rect 42246 596808 42302 596864
rect 42062 595992 42118 596048
rect 41694 595720 41750 595776
rect 33046 595584 33102 595640
rect 31022 594360 31078 594416
rect 35162 595176 35218 595232
rect 34426 594768 34482 594824
rect 34426 587152 34482 587208
rect 36542 593544 36598 593600
rect 41694 592884 41750 592920
rect 41694 592864 41696 592884
rect 41696 592864 41748 592884
rect 41748 592864 41750 592884
rect 39946 590688 40002 590744
rect 39578 586608 39634 586664
rect 39578 585792 39634 585848
rect 41786 592320 41842 592376
rect 40774 589600 40830 589656
rect 41786 589464 41842 589520
rect 39946 585520 40002 585576
rect 42982 593136 43038 593192
rect 42430 585384 42486 585440
rect 40498 584704 40554 584760
rect 42062 584704 42118 584760
rect 39670 584568 39726 584624
rect 41786 582528 41842 582584
rect 42430 581576 42486 581632
rect 42246 581440 42302 581496
rect 42062 581168 42118 581224
rect 42246 580080 42302 580136
rect 42062 578856 42118 578912
rect 42154 578176 42210 578232
rect 42154 576952 42210 577008
rect 42246 575592 42302 575648
rect 42062 574640 42118 574696
rect 42614 579808 42670 579864
rect 42614 572736 42670 572792
rect 42522 572056 42578 572112
rect 41786 570152 41842 570208
rect 40590 556008 40646 556064
rect 40866 555600 40922 555656
rect 43258 591504 43314 591560
rect 44270 686432 44326 686488
rect 45006 763680 45062 763736
rect 44822 758104 44878 758160
rect 44638 727640 44694 727696
rect 43994 676640 44050 676696
rect 43810 644680 43866 644736
rect 44638 679496 44694 679552
rect 44638 643456 44694 643512
rect 44270 643048 44326 643104
rect 43626 637744 43682 637800
rect 43810 634888 43866 634944
rect 43994 634480 44050 634536
rect 43994 623328 44050 623384
rect 43442 581168 43498 581224
rect 43166 578856 43222 578912
rect 42982 578176 43038 578232
rect 43258 558456 43314 558512
rect 43442 558048 43498 558104
rect 43442 557640 43498 557696
rect 42982 555192 43038 555248
rect 40038 553352 40094 553408
rect 40866 553352 40922 553408
rect 34426 551928 34482 551984
rect 31758 547460 31814 547496
rect 31758 547440 31760 547460
rect 31760 547440 31812 547460
rect 31812 547440 31814 547460
rect 41878 550568 41934 550624
rect 42154 549888 42210 549944
rect 41970 549480 42026 549536
rect 41142 548140 41198 548142
rect 41142 548088 41144 548140
rect 41144 548088 41196 548140
rect 41196 548088 41198 548140
rect 41142 548086 41198 548088
rect 41694 547712 41750 547768
rect 40866 545808 40922 545864
rect 42154 545536 42210 545592
rect 41970 545264 42026 545320
rect 39762 542172 39764 542192
rect 39764 542172 39816 542192
rect 39816 542172 39818 542192
rect 39762 542136 39818 542172
rect 42338 542136 42394 542192
rect 39486 541864 39542 541920
rect 42062 541864 42118 541920
rect 43350 551520 43406 551576
rect 42338 538192 42394 538248
rect 42154 537920 42210 537976
rect 42706 537920 42762 537976
rect 41786 535200 41842 535256
rect 42246 533296 42302 533352
rect 42614 530168 42670 530224
rect 42706 529760 42762 529816
rect 41786 529352 41842 529408
rect 40682 522688 40738 522744
rect 40682 431160 40738 431216
rect 41326 430480 41382 430536
rect 41142 430072 41198 430128
rect 40958 429426 41014 429482
rect 41326 429480 41382 429482
rect 41326 429428 41328 429480
rect 41328 429428 41380 429480
rect 41380 429428 41382 429480
rect 41326 429426 41382 429428
rect 41142 428848 41198 428904
rect 42706 428440 42762 428496
rect 43442 547712 43498 547768
rect 43442 547032 43498 547088
rect 43258 522688 43314 522744
rect 41326 427794 41382 427850
rect 40958 427624 41014 427680
rect 41142 427216 41198 427272
rect 41326 425992 41382 426048
rect 40774 425176 40830 425232
rect 42614 424360 42670 424416
rect 41786 421096 41842 421152
rect 41878 419872 41934 419928
rect 42430 420688 42486 420744
rect 42062 412936 42118 412992
rect 42614 412936 42670 412992
rect 41786 407496 41842 407552
rect 41786 403824 41842 403880
rect 41786 401920 41842 401976
rect 41786 400016 41842 400072
rect 41878 398792 41934 398848
rect 35438 387504 35494 387560
rect 35806 387540 35808 387560
rect 35808 387540 35860 387560
rect 35860 387540 35862 387560
rect 35806 387504 35862 387540
rect 39946 387096 40002 387152
rect 35806 386688 35862 386744
rect 40130 386708 40186 386744
rect 40130 386688 40132 386708
rect 40132 386688 40184 386708
rect 40184 386688 40186 386708
rect 35622 386280 35678 386336
rect 35346 385872 35402 385928
rect 35530 385464 35586 385520
rect 35806 385484 35862 385520
rect 35806 385464 35808 385484
rect 35808 385464 35860 385484
rect 35860 385464 35862 385484
rect 39946 385056 40002 385112
rect 35622 384648 35678 384704
rect 35806 384240 35862 384296
rect 35806 383832 35862 383888
rect 39762 383832 39818 383888
rect 43074 421504 43130 421560
rect 43810 600888 43866 600944
rect 44362 638152 44418 638208
rect 44546 600480 44602 600536
rect 44362 600072 44418 600128
rect 44178 599664 44234 599720
rect 44270 557232 44326 557288
rect 44638 591912 44694 591968
rect 44638 556824 44694 556880
rect 44454 556416 44510 556472
rect 43810 554784 43866 554840
rect 43810 554376 43866 554432
rect 43994 549072 44050 549128
rect 44178 548664 44234 548720
rect 43442 422728 43498 422784
rect 43258 387096 43314 387152
rect 42798 383832 42854 383888
rect 35254 383424 35310 383480
rect 40130 383424 40186 383480
rect 35438 383016 35494 383072
rect 35806 382644 35808 382664
rect 35808 382644 35860 382664
rect 35860 382644 35862 382664
rect 35806 382608 35862 382644
rect 35622 382200 35678 382256
rect 40038 382200 40094 382256
rect 35622 381792 35678 381848
rect 39026 381792 39082 381848
rect 32402 381384 32458 381440
rect 28814 376488 28870 376544
rect 35806 380976 35862 381032
rect 35622 380568 35678 380624
rect 35806 380160 35862 380216
rect 40038 380160 40094 380216
rect 35806 379752 35862 379808
rect 35806 378936 35862 378992
rect 35622 377712 35678 377768
rect 41418 380976 41474 381032
rect 40222 378936 40278 378992
rect 41510 378528 41566 378584
rect 41234 378120 41290 378176
rect 39946 377712 40002 377768
rect 35806 377304 35862 377360
rect 39578 377304 39634 377360
rect 41694 376932 41696 376952
rect 41696 376932 41748 376952
rect 41748 376932 41750 376952
rect 41694 376896 41750 376932
rect 35806 376080 35862 376136
rect 42062 369688 42118 369744
rect 41786 365608 41842 365664
rect 41786 363704 41842 363760
rect 41786 360576 41842 360632
rect 41878 358672 41934 358728
rect 41786 356904 41842 356960
rect 41970 355680 42026 355736
rect 39210 345888 39266 345944
rect 35806 344256 35862 344312
rect 35622 343848 35678 343904
rect 35806 343440 35862 343496
rect 35622 343032 35678 343088
rect 40038 343032 40094 343088
rect 35806 342660 35808 342680
rect 35808 342660 35860 342680
rect 35860 342660 35862 342680
rect 35806 342624 35862 342660
rect 40314 342660 40316 342680
rect 40316 342660 40368 342680
rect 40368 342660 40370 342680
rect 40314 342624 40370 342660
rect 35622 342252 35624 342272
rect 35624 342252 35676 342272
rect 35676 342252 35678 342272
rect 35622 342216 35678 342252
rect 35806 341808 35862 341864
rect 42982 377712 43038 377768
rect 43258 377304 43314 377360
rect 43258 342624 43314 342680
rect 35346 341400 35402 341456
rect 35622 341400 35678 341456
rect 35806 341028 35808 341048
rect 35808 341028 35860 341048
rect 35860 341028 35862 341048
rect 35806 340992 35862 341028
rect 35806 340176 35862 340232
rect 35622 338952 35678 339008
rect 41418 338952 41474 339008
rect 35806 338544 35862 338600
rect 41786 338680 41842 338736
rect 41694 338136 41750 338192
rect 35806 337728 35862 337784
rect 35530 336912 35586 336968
rect 35806 336932 35862 336968
rect 35806 336912 35808 336932
rect 35808 336912 35860 336932
rect 35860 336912 35862 336932
rect 35622 335688 35678 335744
rect 35806 335588 35808 335608
rect 35808 335588 35860 335608
rect 35860 335588 35862 335608
rect 35806 335552 35862 335588
rect 35622 334872 35678 334928
rect 35438 334464 35494 334520
rect 35806 334464 35862 334520
rect 35806 333240 35862 333296
rect 35806 332832 35862 332888
rect 40314 335688 40370 335744
rect 40222 334872 40278 334928
rect 39854 332832 39910 332888
rect 40314 333648 40370 333704
rect 40866 332424 40922 332480
rect 40130 331200 40186 331256
rect 39302 330656 39358 330712
rect 41786 324808 41842 324864
rect 41786 322768 41842 322824
rect 41786 315560 41842 315616
rect 41786 313656 41842 313712
rect 41786 312976 41842 313032
rect 40958 300464 41014 300520
rect 41142 300056 41198 300112
rect 41142 299240 41198 299296
rect 40958 298424 41014 298480
rect 42706 298832 42762 298888
rect 40958 298016 41014 298072
rect 41142 297608 41198 297664
rect 40774 295568 40830 295624
rect 37922 294752 37978 294808
rect 40498 292544 40500 292588
rect 40500 292544 40552 292588
rect 40552 292544 40554 292588
rect 41786 295160 41842 295216
rect 41786 294480 41842 294536
rect 41326 294344 41382 294400
rect 41786 293528 41842 293584
rect 40498 292532 40554 292544
rect 41786 292032 41842 292088
rect 41142 291896 41198 291952
rect 40958 291080 41014 291136
rect 41142 290264 41198 290320
rect 43074 332424 43130 332480
rect 43074 301280 43130 301336
rect 43074 299648 43130 299704
rect 42982 293120 43038 293176
rect 41970 289584 42026 289640
rect 41970 281424 42026 281480
rect 42522 278704 42578 278760
rect 41786 277344 41842 277400
rect 41786 272992 41842 273048
rect 41786 272312 41842 272368
rect 41786 270408 41842 270464
rect 39946 259528 40002 259584
rect 35806 258032 35862 258088
rect 35622 257488 35678 257544
rect 39578 257488 39634 257544
rect 35438 257080 35494 257136
rect 35806 257116 35808 257136
rect 35808 257116 35860 257136
rect 35860 257116 35862 257136
rect 35806 257080 35862 257116
rect 35438 256264 35494 256320
rect 35622 255856 35678 255912
rect 35806 255448 35862 255504
rect 35438 255040 35494 255096
rect 35806 255040 35862 255096
rect 35622 254632 35678 254688
rect 35806 254260 35808 254280
rect 35808 254260 35860 254280
rect 35860 254260 35862 254280
rect 35806 254224 35862 254260
rect 35530 253000 35586 253056
rect 35806 253000 35862 253056
rect 40038 253816 40094 253872
rect 44546 426808 44602 426864
rect 43994 423952 44050 424008
rect 43810 423136 43866 423192
rect 43626 386688 43682 386744
rect 44362 385056 44418 385112
rect 44638 383424 44694 383480
rect 43626 381792 43682 381848
rect 44178 380976 44234 381032
rect 43810 378120 43866 378176
rect 44362 378528 44418 378584
rect 44178 369688 44234 369744
rect 44270 338952 44326 339008
rect 43810 335688 43866 335744
rect 43994 334872 44050 334928
rect 43626 300872 43682 300928
rect 43626 290672 43682 290728
rect 43166 257488 43222 257544
rect 41234 254224 41290 254280
rect 42890 253816 42946 253872
rect 42430 253544 42486 253600
rect 40406 253000 40462 253056
rect 39762 252592 39818 252648
rect 31022 252184 31078 252240
rect 35530 251776 35586 251832
rect 35806 251776 35862 251832
rect 35438 250960 35494 251016
rect 35622 250552 35678 250608
rect 35806 250180 35808 250200
rect 35808 250180 35860 250200
rect 35860 250180 35862 250200
rect 35806 250144 35862 250180
rect 39394 250180 39396 250200
rect 39396 250180 39448 250200
rect 39448 250180 39450 250200
rect 39394 250144 39450 250180
rect 35438 249328 35494 249384
rect 35622 248920 35678 248976
rect 35806 248512 35862 248568
rect 39118 248548 39120 248568
rect 39120 248548 39172 248568
rect 39172 248548 39174 248568
rect 39118 248512 39174 248548
rect 35806 248104 35862 248160
rect 35622 247696 35678 247752
rect 35806 247288 35862 247344
rect 41694 252184 41750 252240
rect 41510 251776 41566 251832
rect 41694 251368 41750 251424
rect 39854 245656 39910 245712
rect 40406 247288 40462 247344
rect 40130 245112 40186 245168
rect 42062 240080 42118 240136
rect 41786 238448 41842 238504
rect 42062 238312 42118 238368
rect 42246 237632 42302 237688
rect 43442 252592 43498 252648
rect 43258 250144 43314 250200
rect 43074 245112 43130 245168
rect 42614 238312 42670 238368
rect 42430 237360 42486 237416
rect 41786 236544 41842 236600
rect 41970 228928 42026 228984
rect 42062 227296 42118 227352
rect 28538 223896 28594 223952
rect 41694 223624 41750 223680
rect 40682 222264 40738 222320
rect 40314 216688 40370 216744
rect 35806 215056 35862 215112
rect 33046 214240 33102 214296
rect 35806 214240 35862 214296
rect 39946 214240 40002 214296
rect 39946 213832 40002 213888
rect 35438 213424 35494 213480
rect 28538 212608 28594 212664
rect 35622 213016 35678 213072
rect 35806 212608 35862 212664
rect 41510 217252 41566 217288
rect 41510 217232 41512 217252
rect 41512 217232 41564 217252
rect 41564 217232 41566 217252
rect 41510 215056 41566 215112
rect 40958 212200 41014 212256
rect 35806 211792 35862 211848
rect 35622 211384 35678 211440
rect 39670 211404 39726 211440
rect 39670 211384 39672 211404
rect 39672 211384 39724 211404
rect 39724 211384 39726 211404
rect 35806 210976 35862 211032
rect 41510 210976 41566 211032
rect 35622 210568 35678 210624
rect 35806 210160 35862 210216
rect 35806 209344 35862 209400
rect 30286 208936 30342 208992
rect 42062 217268 42064 217288
rect 42064 217268 42116 217288
rect 42116 217268 42118 217288
rect 42062 217232 42118 217268
rect 43166 215056 43222 215112
rect 44638 330656 44694 330712
rect 44362 297200 44418 297256
rect 44178 291488 44234 291544
rect 44270 254224 44326 254280
rect 44546 251776 44602 251832
rect 43810 248512 43866 248568
rect 44178 247288 44234 247344
rect 44546 240080 44602 240136
rect 45190 679904 45246 679960
rect 45006 677864 45062 677920
rect 45190 632032 45246 632088
rect 45190 620880 45246 620936
rect 45374 552336 45430 552392
rect 45190 551112 45246 551168
rect 45558 424768 45614 424824
rect 45190 423544 45246 423600
rect 45374 421232 45430 421288
rect 45742 419464 45798 419520
rect 45190 376896 45246 376952
rect 45006 276664 45062 276720
rect 45374 343032 45430 343088
rect 45558 338680 45614 338736
rect 45374 338136 45430 338192
rect 46018 333648 46074 333704
rect 45834 332832 45890 332888
rect 45558 295976 45614 296032
rect 45374 293936 45430 293992
rect 43626 214240 43682 214296
rect 45374 253000 45430 253056
rect 45558 252184 45614 252240
rect 45742 245656 45798 245712
rect 47582 763272 47638 763328
rect 46386 721112 46442 721168
rect 46570 345888 46626 345944
rect 46754 331200 46810 331256
rect 47030 294480 47086 294536
rect 46570 259528 46626 259584
rect 47030 251368 47086 251424
rect 46386 228792 46442 228848
rect 47766 731312 47822 731368
rect 47766 646040 47822 646096
rect 47766 601296 47822 601352
rect 47766 590280 47822 590336
rect 49146 228520 49202 228576
rect 47766 228248 47822 228304
rect 47582 222536 47638 222592
rect 45282 216688 45338 216744
rect 45006 213832 45062 213888
rect 43350 212200 43406 212256
rect 42890 211384 42946 211440
rect 42338 210976 42394 211032
rect 40038 208936 40094 208992
rect 35806 208528 35862 208584
rect 35530 207304 35586 207360
rect 35806 207324 35862 207360
rect 35806 207304 35808 207324
rect 35808 207304 35860 207324
rect 35860 207304 35862 207324
rect 35806 206488 35862 206544
rect 35806 205692 35862 205728
rect 35806 205672 35808 205692
rect 35808 205672 35860 205692
rect 35860 205672 35862 205692
rect 35622 205264 35678 205320
rect 35806 204892 35808 204912
rect 35808 204892 35860 204912
rect 35860 204892 35862 204912
rect 35806 204856 35862 204892
rect 35530 204448 35586 204504
rect 35806 204484 35808 204504
rect 35808 204484 35860 204504
rect 35860 204484 35862 204504
rect 35806 204448 35862 204484
rect 40130 206896 40186 206952
rect 39946 205672 40002 205728
rect 42890 206896 42946 206952
rect 40958 205264 41014 205320
rect 40774 204448 40830 204504
rect 39762 204040 39818 204096
rect 35622 203632 35678 203688
rect 35806 203224 35862 203280
rect 40038 203224 40094 203280
rect 41786 202952 41842 203008
rect 30286 202136 30342 202192
rect 41786 197104 41842 197160
rect 44178 205672 44234 205728
rect 43258 205264 43314 205320
rect 41786 195200 41842 195256
rect 41786 191528 41842 191584
rect 43810 204040 43866 204096
rect 43626 202952 43682 203008
rect 41786 185816 41842 185872
rect 41786 184048 41842 184104
rect 44546 204448 44602 204504
rect 50710 265512 50766 265568
rect 62118 923752 62174 923808
rect 62118 910696 62174 910752
rect 62118 897776 62174 897832
rect 62118 884740 62174 884776
rect 62118 884720 62120 884740
rect 62120 884720 62172 884740
rect 62172 884720 62174 884740
rect 62118 871664 62174 871720
rect 62118 858608 62174 858664
rect 62118 845552 62174 845608
rect 62118 832496 62174 832552
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 62118 793620 62174 793656
rect 62118 793600 62120 793620
rect 62120 793600 62172 793620
rect 62172 793600 62174 793620
rect 62118 780408 62174 780464
rect 54482 278024 54538 278080
rect 53470 276936 53526 276992
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 62118 741240 62174 741296
rect 62118 728184 62174 728240
rect 62118 715264 62174 715320
rect 62118 702208 62174 702264
rect 62118 689152 62174 689208
rect 62118 676096 62174 676152
rect 62118 663040 62174 663096
rect 62118 649984 62174 650040
rect 62118 637064 62174 637120
rect 62118 624008 62174 624064
rect 62118 610952 62174 611008
rect 62118 597896 62174 597952
rect 62118 584840 62174 584896
rect 62118 571784 62174 571840
rect 62118 558728 62174 558784
rect 62118 545808 62174 545864
rect 62762 532752 62818 532808
rect 62118 519696 62174 519752
rect 62118 506640 62174 506696
rect 62118 493584 62174 493640
rect 62118 480528 62174 480584
rect 62118 467472 62174 467528
rect 62118 454552 62174 454608
rect 62118 441496 62174 441552
rect 62118 428440 62174 428496
rect 62118 415420 62120 415440
rect 62120 415420 62172 415440
rect 62172 415420 62174 415440
rect 62118 415384 62174 415420
rect 62118 402328 62174 402384
rect 62118 389292 62174 389328
rect 62118 389272 62120 389292
rect 62120 389272 62172 389292
rect 62172 389272 62174 389292
rect 62118 376216 62174 376272
rect 62118 363296 62174 363352
rect 62118 350240 62174 350296
rect 62118 337184 62174 337240
rect 62762 324128 62818 324184
rect 62762 311072 62818 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 56046 230016 56102 230072
rect 54666 229744 54722 229800
rect 53286 227432 53342 227488
rect 50342 227160 50398 227216
rect 62118 285096 62174 285152
rect 61382 230288 61438 230344
rect 60002 226888 60058 226944
rect 59266 226616 59322 226672
rect 56874 226072 56930 226128
rect 50342 221992 50398 222048
rect 51722 221720 51778 221776
rect 56506 219952 56562 220008
rect 60002 221992 60058 222048
rect 60002 221448 60058 221504
rect 366638 267280 366694 267336
rect 369122 270136 369178 270192
rect 369306 266756 369362 266792
rect 369306 266736 369308 266756
rect 369308 266736 369360 266756
rect 369360 266736 369362 266756
rect 370502 267300 370558 267336
rect 370502 267280 370504 267300
rect 370504 267280 370556 267300
rect 370556 267280 370558 267300
rect 371790 266736 371846 266792
rect 373722 269456 373778 269512
rect 375194 269492 375196 269512
rect 375196 269492 375248 269512
rect 375248 269492 375250 269512
rect 375194 269456 375250 269492
rect 376942 270172 376944 270192
rect 376944 270172 376996 270192
rect 376996 270172 376998 270192
rect 376942 270136 376998 270172
rect 377126 270000 377182 270056
rect 379150 270308 379152 270328
rect 379152 270308 379204 270328
rect 379204 270308 379206 270328
rect 379150 270272 379206 270308
rect 379518 270272 379574 270328
rect 380530 270272 380586 270328
rect 379334 270000 379390 270056
rect 379334 267572 379390 267608
rect 379334 267552 379336 267572
rect 379336 267552 379388 267572
rect 379388 267552 379390 267572
rect 381358 267572 381414 267608
rect 381358 267552 381360 267572
rect 381360 267552 381412 267572
rect 381412 267552 381414 267572
rect 383566 270308 383568 270328
rect 383568 270308 383620 270328
rect 383620 270308 383622 270328
rect 383566 270272 383622 270308
rect 383658 270000 383714 270056
rect 383382 269592 383438 269648
rect 383750 269592 383806 269648
rect 384118 269492 384120 269512
rect 384120 269492 384172 269512
rect 384172 269492 384174 269512
rect 384118 269456 384174 269492
rect 386970 270000 387026 270056
rect 388166 267280 388222 267336
rect 388994 269492 388996 269512
rect 388996 269492 389048 269512
rect 389048 269492 389050 269512
rect 388994 269456 389050 269492
rect 390466 267300 390522 267336
rect 390466 267280 390468 267300
rect 390468 267280 390520 267300
rect 390520 267280 390522 267300
rect 391754 271532 391756 271552
rect 391756 271532 391808 271552
rect 391808 271532 391810 271552
rect 391754 271496 391810 271532
rect 392582 267572 392638 267608
rect 392582 267552 392584 267572
rect 392584 267552 392636 267572
rect 392636 267552 392638 267572
rect 393686 269356 393688 269376
rect 393688 269356 393740 269376
rect 393740 269356 393742 269376
rect 393686 269320 393742 269356
rect 393410 267552 393466 267608
rect 396262 266484 396318 266520
rect 396262 266464 396264 266484
rect 396264 266464 396316 266484
rect 396316 266464 396318 266484
rect 399666 275732 399722 275768
rect 399666 275712 399668 275732
rect 399668 275712 399720 275732
rect 399720 275712 399722 275732
rect 397918 269628 397920 269648
rect 397920 269628 397972 269648
rect 397972 269628 397974 269648
rect 397918 269592 397974 269628
rect 398930 269592 398986 269648
rect 398470 266464 398526 266520
rect 400770 275732 400826 275768
rect 400770 275712 400772 275732
rect 400772 275712 400824 275732
rect 400824 275712 400826 275732
rect 400126 269728 400182 269784
rect 401598 269320 401654 269376
rect 402610 271496 402666 271552
rect 402978 270952 403034 271008
rect 402794 270580 402796 270600
rect 402796 270580 402848 270600
rect 402848 270580 402850 270600
rect 402794 270544 402850 270580
rect 403070 270544 403126 270600
rect 404174 270544 404230 270600
rect 405922 270580 405924 270600
rect 405924 270580 405976 270600
rect 405976 270580 405978 270600
rect 405922 270544 405978 270580
rect 406750 270172 406752 270192
rect 406752 270172 406804 270192
rect 406804 270172 406806 270192
rect 406750 270136 406806 270172
rect 408774 270172 408776 270192
rect 408776 270172 408828 270192
rect 408828 270172 408830 270192
rect 408774 270136 408830 270172
rect 408498 269048 408554 269104
rect 409694 271632 409750 271688
rect 411258 270952 411314 271008
rect 410798 266328 410854 266384
rect 412914 271088 412970 271144
rect 412822 266892 412878 266928
rect 412822 266872 412824 266892
rect 412824 266872 412876 266892
rect 412876 266872 412878 266892
rect 413926 271088 413982 271144
rect 415858 269456 415914 269512
rect 414662 266872 414718 266928
rect 417698 270852 417700 270872
rect 417700 270852 417752 270872
rect 417752 270852 417754 270872
rect 417698 270816 417754 270852
rect 416778 269048 416834 269104
rect 416686 268116 416742 268152
rect 416686 268096 416688 268116
rect 416688 268096 416740 268116
rect 416740 268096 416742 268116
rect 417698 267824 417754 267880
rect 418158 270852 418160 270872
rect 418160 270852 418212 270872
rect 418212 270852 418214 270872
rect 418158 270816 418214 270852
rect 418066 268096 418122 268152
rect 417422 266364 417424 266384
rect 417424 266364 417476 266384
rect 417476 266364 417478 266384
rect 417422 266328 417478 266364
rect 420734 266600 420790 266656
rect 424506 272348 424508 272368
rect 424508 272348 424560 272368
rect 424560 272348 424562 272368
rect 424506 272312 424562 272348
rect 422666 267824 422722 267880
rect 423862 266600 423918 266656
rect 425242 268232 425298 268288
rect 424874 267980 424930 268016
rect 424874 267960 424876 267980
rect 424876 267960 424928 267980
rect 424928 267960 424930 267980
rect 426254 273536 426310 273592
rect 427266 272312 427322 272368
rect 426898 267028 426954 267064
rect 427358 267572 427414 267608
rect 427358 267552 427360 267572
rect 427360 267552 427412 267572
rect 427412 267552 427414 267572
rect 426898 267008 426900 267028
rect 426900 267008 426952 267028
rect 426952 267008 426954 267028
rect 428002 267572 428058 267608
rect 428002 267552 428004 267572
rect 428004 267552 428056 267572
rect 428056 267552 428058 267572
rect 428094 267280 428150 267336
rect 429290 272176 429346 272232
rect 429106 270680 429162 270736
rect 428462 267980 428518 268016
rect 428462 267960 428464 267980
rect 428464 267960 428516 267980
rect 428516 267960 428518 267980
rect 432050 273536 432106 273592
rect 431866 272448 431922 272504
rect 431498 271088 431554 271144
rect 429934 269184 429990 269240
rect 429290 268232 429346 268288
rect 434350 274080 434406 274136
rect 432970 271360 433026 271416
rect 432786 269184 432842 269240
rect 432602 267008 432658 267064
rect 433614 271088 433670 271144
rect 641994 278024 642050 278080
rect 436282 270716 436284 270736
rect 436284 270716 436336 270736
rect 436336 270716 436338 270736
rect 436282 270680 436338 270716
rect 436006 267708 436062 267744
rect 436006 267688 436008 267708
rect 436008 267688 436060 267708
rect 436060 267688 436062 267708
rect 436926 272856 436982 272912
rect 437938 272856 437994 272912
rect 437570 272448 437626 272504
rect 437110 272176 437166 272232
rect 437386 272212 437388 272232
rect 437388 272212 437440 272232
rect 437440 272212 437442 272232
rect 437386 272176 437442 272212
rect 438674 270000 438730 270056
rect 437018 269048 437074 269104
rect 437386 267708 437442 267744
rect 437386 267688 437388 267708
rect 437388 267688 437440 267708
rect 437440 267688 437442 267708
rect 437386 266756 437442 266792
rect 437386 266736 437388 266756
rect 437388 266736 437440 266756
rect 437440 266736 437442 266756
rect 442446 272176 442502 272232
rect 441526 271904 441582 271960
rect 438858 269048 438914 269104
rect 441342 268932 441398 268968
rect 441342 268912 441344 268932
rect 441344 268912 441396 268932
rect 441396 268912 441398 268932
rect 442446 266736 442502 266792
rect 444194 271904 444250 271960
rect 446218 275440 446274 275496
rect 445390 272176 445446 272232
rect 443550 270272 443606 270328
rect 443182 268912 443238 268968
rect 445114 270000 445170 270056
rect 447874 272212 447876 272232
rect 447876 272212 447928 272232
rect 447928 272212 447930 272232
rect 447874 272176 447930 272212
rect 446034 271360 446090 271416
rect 446310 271360 446366 271416
rect 447046 268504 447102 268560
rect 446862 266192 446918 266248
rect 448334 271904 448390 271960
rect 449714 273128 449770 273184
rect 448518 268504 448574 268560
rect 449070 266212 449126 266248
rect 449070 266192 449072 266212
rect 449072 266192 449124 266212
rect 449124 266192 449126 266212
rect 450542 272856 450598 272912
rect 450174 267008 450230 267064
rect 451002 273164 451004 273184
rect 451004 273164 451056 273184
rect 451056 273164 451058 273184
rect 451002 273128 451058 273164
rect 452106 272856 452162 272912
rect 452106 272448 452162 272504
rect 451094 271904 451150 271960
rect 451370 271360 451426 271416
rect 451554 271360 451610 271416
rect 453762 272856 453818 272912
rect 454866 273808 454922 273864
rect 454682 272892 454684 272912
rect 454684 272892 454736 272912
rect 454736 272892 454738 272912
rect 454682 272856 454738 272892
rect 454406 272484 454408 272504
rect 454408 272484 454460 272504
rect 454460 272484 454462 272504
rect 454406 272448 454462 272484
rect 455142 269184 455198 269240
rect 454866 267008 454922 267064
rect 454958 266328 455014 266384
rect 456890 271360 456946 271416
rect 456752 271124 456754 271144
rect 456754 271124 456806 271144
rect 456806 271124 456808 271144
rect 456752 271088 456808 271124
rect 456798 269184 456854 269240
rect 458638 272176 458694 272232
rect 457902 268096 457958 268152
rect 456890 266328 456946 266384
rect 457166 266328 457222 266384
rect 459374 270000 459430 270056
rect 460938 274352 460994 274408
rect 461030 273828 461086 273864
rect 461030 273808 461032 273828
rect 461032 273808 461084 273828
rect 461084 273808 461086 273828
rect 460846 272448 460902 272504
rect 460110 268368 460166 268424
rect 461766 272484 461768 272504
rect 461768 272484 461820 272504
rect 461820 272484 461822 272504
rect 461766 272448 461822 272484
rect 461766 271088 461822 271144
rect 461766 270000 461822 270056
rect 462502 271224 462558 271280
rect 461582 268640 461638 268696
rect 461030 266056 461086 266112
rect 462318 268388 462374 268424
rect 462318 268368 462320 268388
rect 462320 268368 462372 268388
rect 462372 268368 462374 268388
rect 461950 268096 462006 268152
rect 463606 266736 463662 266792
rect 462502 266328 462558 266384
rect 461766 266076 461822 266112
rect 461766 266056 461768 266076
rect 461768 266056 461820 266076
rect 461820 266056 461822 266076
rect 462686 265784 462742 265840
rect 464894 272448 464950 272504
rect 464710 268096 464766 268152
rect 466274 272720 466330 272776
rect 466274 272176 466330 272232
rect 466458 271360 466514 271416
rect 465354 271260 465356 271280
rect 465356 271260 465408 271280
rect 465408 271260 465410 271280
rect 465354 271224 465410 271260
rect 465998 271088 466054 271144
rect 466550 271124 466552 271144
rect 466552 271124 466604 271144
rect 466604 271124 466606 271144
rect 466550 271088 466606 271124
rect 465814 265240 465870 265296
rect 466458 268912 466514 268968
rect 466366 268368 466422 268424
rect 466182 267552 466238 267608
rect 466182 266464 466238 266520
rect 466734 268388 466790 268424
rect 466734 268368 466736 268388
rect 466736 268368 466788 268388
rect 466788 268368 466790 268388
rect 467010 267552 467066 267608
rect 466826 267008 466882 267064
rect 466918 265240 466974 265296
rect 468022 268912 468078 268968
rect 468206 267688 468262 267744
rect 470230 274644 470286 274680
rect 470230 274624 470232 274644
rect 470232 274624 470284 274644
rect 470284 274624 470286 274644
rect 470414 274352 470470 274408
rect 472162 274624 472218 274680
rect 470506 270000 470562 270056
rect 469218 268096 469274 268152
rect 470046 267008 470102 267064
rect 472254 270544 472310 270600
rect 471426 267708 471482 267744
rect 471426 267688 471428 267708
rect 471428 267688 471480 267708
rect 471480 267688 471482 267708
rect 473726 268096 473782 268152
rect 475842 274352 475898 274408
rect 475658 272176 475714 272232
rect 474922 270000 474978 270056
rect 475566 268368 475622 268424
rect 474002 266736 474058 266792
rect 474646 266736 474702 266792
rect 476026 272720 476082 272776
rect 476026 269184 476082 269240
rect 480166 275712 480222 275768
rect 480350 275712 480406 275768
rect 479798 274352 479854 274408
rect 477498 269184 477554 269240
rect 481454 275168 481510 275224
rect 480074 272720 480130 272776
rect 480994 272720 481050 272776
rect 480074 272176 480130 272232
rect 480994 272176 481050 272232
rect 480534 271360 480590 271416
rect 480442 271088 480498 271144
rect 480074 270000 480130 270056
rect 480258 268912 480314 268968
rect 480350 268388 480406 268424
rect 480350 268368 480352 268388
rect 480352 268368 480404 268388
rect 480404 268368 480406 268388
rect 479890 266756 479946 266792
rect 479890 266736 479892 266756
rect 479892 266736 479944 266756
rect 479944 266736 479946 266756
rect 479614 265784 479670 265840
rect 483018 275984 483074 276040
rect 482558 274352 482614 274408
rect 483018 270000 483074 270056
rect 483110 267552 483166 267608
rect 485594 270816 485650 270872
rect 485778 270544 485834 270600
rect 487802 272992 487858 273048
rect 487618 272720 487674 272776
rect 487618 271904 487674 271960
rect 489918 276004 489974 276040
rect 489918 275984 489920 276004
rect 489920 275984 489972 276004
rect 489972 275984 489974 276004
rect 490102 275984 490158 276040
rect 489734 275712 489790 275768
rect 490010 275732 490066 275768
rect 490010 275712 490012 275732
rect 490012 275712 490064 275732
rect 490064 275712 490066 275732
rect 491850 276120 491906 276176
rect 491482 275984 491538 276040
rect 489918 274896 489974 274952
rect 490470 274488 490526 274544
rect 489734 274352 489790 274408
rect 489458 273808 489514 273864
rect 489274 271360 489330 271416
rect 488170 269900 488172 269920
rect 488172 269900 488224 269920
rect 488224 269900 488226 269920
rect 488170 269864 488226 269900
rect 487986 269728 488042 269784
rect 488078 266736 488134 266792
rect 489734 273536 489790 273592
rect 490102 273536 490158 273592
rect 490010 272176 490066 272232
rect 489642 271904 489698 271960
rect 490010 271768 490066 271824
rect 490102 271360 490158 271416
rect 489642 271088 489698 271144
rect 490286 271088 490342 271144
rect 489734 269864 489790 269920
rect 489734 269184 489790 269240
rect 490654 272992 490710 273048
rect 491206 272992 491262 273048
rect 489734 267552 489790 267608
rect 490470 267572 490526 267608
rect 490470 267552 490472 267572
rect 490472 267552 490524 267572
rect 490524 267552 490526 267572
rect 489734 266464 489790 266520
rect 490194 266736 490250 266792
rect 490470 266736 490526 266792
rect 491390 267552 491446 267608
rect 493046 271088 493102 271144
rect 492126 267552 492182 267608
rect 494978 274896 495034 274952
rect 493690 270000 493746 270056
rect 495070 270544 495126 270600
rect 494150 267824 494206 267880
rect 494886 266736 494942 266792
rect 494518 266464 494574 266520
rect 497462 276392 497518 276448
rect 497186 274508 497242 274544
rect 497186 274488 497188 274508
rect 497188 274488 497240 274508
rect 497240 274488 497242 274508
rect 496726 271088 496782 271144
rect 496542 266736 496598 266792
rect 495438 264288 495494 264344
rect 499578 277344 499634 277400
rect 499210 276120 499266 276176
rect 499394 275984 499450 276040
rect 499762 275984 499818 276040
rect 497646 273536 497702 273592
rect 499210 272720 499266 272776
rect 497462 267008 497518 267064
rect 498014 266464 498070 266520
rect 498842 272176 498898 272232
rect 499854 272176 499910 272232
rect 499394 271768 499450 271824
rect 499762 271632 499818 271688
rect 499670 270580 499672 270600
rect 499672 270580 499724 270600
rect 499724 270580 499726 270600
rect 499670 270544 499726 270580
rect 499394 270036 499396 270056
rect 499396 270036 499448 270056
rect 499448 270036 499450 270056
rect 499394 270000 499450 270036
rect 502338 277344 502394 277400
rect 501142 275712 501198 275768
rect 500222 271904 500278 271960
rect 500038 270000 500094 270056
rect 499210 269184 499266 269240
rect 499762 269184 499818 269240
rect 499210 268912 499266 268968
rect 499394 268912 499450 268968
rect 499026 267008 499082 267064
rect 499210 266736 499266 266792
rect 499394 266484 499450 266520
rect 499394 266464 499396 266484
rect 499396 266464 499448 266484
rect 499448 266464 499450 266484
rect 503626 274624 503682 274680
rect 504730 275712 504786 275768
rect 505282 273536 505338 273592
rect 504546 270816 504602 270872
rect 503626 269456 503682 269512
rect 501142 268912 501198 268968
rect 508870 276392 508926 276448
rect 509238 275712 509294 275768
rect 509330 274624 509386 274680
rect 507858 272176 507914 272232
rect 509422 271632 509478 271688
rect 509238 270680 509294 270736
rect 512182 275712 512238 275768
rect 514114 272720 514170 272776
rect 509054 269184 509110 269240
rect 510618 269184 510674 269240
rect 508870 267824 508926 267880
rect 518346 270680 518402 270736
rect 532974 267280 533030 267336
rect 541070 275440 541126 275496
rect 543462 274080 543518 274136
rect 557906 270272 557962 270328
rect 578882 267552 578938 267608
rect 587898 268640 587954 268696
rect 589278 266056 589334 266112
rect 593142 272448 593198 272504
rect 607218 268368 607274 268424
rect 619086 275168 619142 275224
rect 614762 265784 614818 265840
rect 626170 271360 626226 271416
rect 632150 273808 632206 273864
rect 637578 270000 637634 270056
rect 640706 269728 640762 269784
rect 636198 267008 636254 267064
rect 499762 264288 499818 264344
rect 511538 262656 511594 262712
rect 511354 260208 511410 260264
rect 511446 257760 511502 257816
rect 511170 255312 511226 255368
rect 510618 250416 510674 250472
rect 511906 252864 511962 252920
rect 511078 247968 511134 248024
rect 66718 221992 66774 222048
rect 71686 224168 71742 224224
rect 72882 221176 72938 221232
rect 111062 229472 111118 229528
rect 130382 245656 130438 245712
rect 129186 230832 129242 230888
rect 510710 240624 510766 240680
rect 507490 237904 507546 237960
rect 132590 230852 132646 230888
rect 132590 230832 132592 230852
rect 132592 230832 132644 230852
rect 132644 230832 132646 230852
rect 144642 230832 144698 230888
rect 132498 230560 132554 230616
rect 145838 230288 145894 230344
rect 146022 230288 146078 230344
rect 130382 225800 130438 225856
rect 129002 225528 129058 225584
rect 130198 220360 130254 220416
rect 136546 222808 136602 222864
rect 145838 229200 145894 229256
rect 142894 227976 142950 228032
rect 142158 227704 142214 227760
rect 142342 226500 142398 226502
rect 142342 226448 142344 226500
rect 142344 226448 142396 226500
rect 142396 226448 142398 226500
rect 142342 226446 142398 226448
rect 141698 226380 141700 226400
rect 141700 226380 141752 226400
rect 141752 226380 141754 226400
rect 141698 226344 141754 226380
rect 142158 223080 142214 223136
rect 142618 222808 142674 222864
rect 142066 219544 142122 219600
rect 142250 219544 142306 219600
rect 147034 224440 147090 224496
rect 143078 219700 143134 219736
rect 143078 219680 143080 219700
rect 143080 219680 143132 219700
rect 143132 219680 143134 219700
rect 147678 220632 147734 220688
rect 149150 226072 149206 226128
rect 148322 223080 148378 223136
rect 148966 222808 149022 222864
rect 148046 219952 148102 220008
rect 147770 219680 147826 219736
rect 150530 230288 150586 230344
rect 150806 227976 150862 228032
rect 151910 229200 151966 229256
rect 151358 226616 151414 226672
rect 151450 225256 151506 225312
rect 150162 223352 150218 223408
rect 150346 220088 150402 220144
rect 151634 225020 151636 225040
rect 151636 225020 151688 225040
rect 151688 225020 151690 225040
rect 151634 224984 151690 225020
rect 153842 230832 153898 230888
rect 153750 230288 153806 230344
rect 153290 227704 153346 227760
rect 152738 225256 152794 225312
rect 152186 224984 152242 225040
rect 151910 224440 151966 224496
rect 151634 221176 151690 221232
rect 154302 226616 154358 226672
rect 152094 220632 152150 220688
rect 152830 219680 152886 219736
rect 155038 224476 155040 224496
rect 155040 224476 155092 224496
rect 155092 224476 155094 224496
rect 155038 224440 155094 224476
rect 154762 221992 154818 222048
rect 154670 219700 154726 219736
rect 154670 219680 154672 219700
rect 154672 219680 154724 219700
rect 154724 219680 154726 219700
rect 155590 223352 155646 223408
rect 156602 227976 156658 228032
rect 157430 227704 157486 227760
rect 157798 226616 157854 226672
rect 157338 224712 157394 224768
rect 157430 224476 157432 224496
rect 157432 224476 157484 224496
rect 157484 224476 157486 224496
rect 157430 224440 157486 224476
rect 157798 224440 157854 224496
rect 157154 223080 157210 223136
rect 157430 223116 157432 223136
rect 157432 223116 157484 223136
rect 157484 223116 157486 223136
rect 157430 223080 157486 223116
rect 157338 222844 157340 222864
rect 157340 222844 157392 222864
rect 157392 222844 157394 222864
rect 157338 222808 157394 222844
rect 157522 222808 157578 222864
rect 156234 221176 156290 221232
rect 157982 224168 158038 224224
rect 157982 223080 158038 223136
rect 156878 220632 156934 220688
rect 157798 220632 157854 220688
rect 158442 229064 158498 229120
rect 158350 222844 158352 222864
rect 158352 222844 158404 222864
rect 158404 222844 158406 222864
rect 158350 222808 158406 222844
rect 160466 230288 160522 230344
rect 160190 227976 160246 228032
rect 158902 220904 158958 220960
rect 159914 224476 159916 224496
rect 159916 224476 159968 224496
rect 159968 224476 159970 224496
rect 159914 224440 159970 224476
rect 161478 230288 161534 230344
rect 161478 224712 161534 224768
rect 159822 221176 159878 221232
rect 160926 221176 160982 221232
rect 161110 221176 161166 221232
rect 160926 219564 160982 219600
rect 160926 219544 160928 219564
rect 160928 219544 160980 219564
rect 160980 219544 160982 219564
rect 164330 230560 164386 230616
rect 165158 229472 165214 229528
rect 163778 229064 163834 229120
rect 166814 230832 166870 230888
rect 166998 230288 167054 230344
rect 166538 227704 166594 227760
rect 166998 226244 167000 226264
rect 167000 226244 167052 226264
rect 167052 226244 167054 226264
rect 166998 226208 167054 226244
rect 165710 223080 165766 223136
rect 165986 220380 166042 220416
rect 165986 220360 165988 220380
rect 165988 220360 166040 220380
rect 166040 220360 166042 220380
rect 165618 219544 165674 219600
rect 166630 221176 166686 221232
rect 166814 221040 166870 221096
rect 169298 230832 169354 230888
rect 168838 230288 168894 230344
rect 170034 229472 170090 229528
rect 169022 220360 169078 220416
rect 171138 221992 171194 222048
rect 171230 221060 171286 221096
rect 171230 221040 171232 221060
rect 171232 221040 171284 221060
rect 171284 221040 171286 221060
rect 171046 219816 171102 219872
rect 172058 230288 172114 230344
rect 172334 227976 172390 228032
rect 173622 226244 173624 226264
rect 173624 226244 173676 226264
rect 173676 226244 173678 226264
rect 173622 226208 173678 226244
rect 173070 222944 173126 223000
rect 173438 220360 173494 220416
rect 173254 219816 173310 219872
rect 174082 222980 174084 223000
rect 174084 222980 174136 223000
rect 174136 222980 174138 223000
rect 174082 222944 174138 222980
rect 175002 229472 175058 229528
rect 174818 221992 174874 222048
rect 175830 220360 175886 220416
rect 176474 226108 176476 226128
rect 176476 226108 176528 226128
rect 176528 226108 176530 226128
rect 176474 226072 176530 226108
rect 176750 226072 176806 226128
rect 178130 225292 178132 225312
rect 178132 225292 178184 225312
rect 178184 225292 178186 225312
rect 178130 225256 178186 225292
rect 176566 220768 176622 220824
rect 177854 220496 177910 220552
rect 179878 225256 179934 225312
rect 180798 226072 180854 226128
rect 180522 219564 180578 219600
rect 180522 219544 180524 219564
rect 180524 219544 180576 219564
rect 180576 219544 180578 219564
rect 181350 226108 181352 226128
rect 181352 226108 181404 226128
rect 181404 226108 181406 226128
rect 181350 226072 181406 226108
rect 182362 227976 182418 228032
rect 181166 222944 181222 223000
rect 181442 220768 181498 220824
rect 181166 220360 181222 220416
rect 181994 222012 182050 222048
rect 181994 221992 181996 222012
rect 181996 221992 182048 222012
rect 182048 221992 182050 222012
rect 182178 219544 182234 219600
rect 183282 219564 183338 219600
rect 183282 219544 183284 219564
rect 183284 219544 183336 219564
rect 183336 219544 183338 219564
rect 185030 223352 185086 223408
rect 185950 226616 186006 226672
rect 185582 223352 185638 223408
rect 187054 224984 187110 225040
rect 187974 226616 188030 226672
rect 187790 221992 187846 222048
rect 187974 219564 188030 219600
rect 187974 219544 187976 219564
rect 187976 219544 188028 219564
rect 188028 219544 188030 219564
rect 190274 230444 190330 230480
rect 190274 230424 190276 230444
rect 190276 230424 190328 230444
rect 190328 230424 190330 230444
rect 190458 230444 190514 230480
rect 190458 230424 190460 230444
rect 190460 230424 190512 230444
rect 190512 230424 190514 230444
rect 190918 229492 190974 229528
rect 190918 229472 190920 229492
rect 190920 229472 190972 229492
rect 190972 229472 190974 229492
rect 190642 229200 190698 229256
rect 190274 226244 190276 226264
rect 190276 226244 190328 226264
rect 190328 226244 190330 226264
rect 190274 226208 190330 226244
rect 189998 224984 190054 225040
rect 189630 222944 189686 223000
rect 191562 229200 191618 229256
rect 191378 226208 191434 226264
rect 190366 224712 190422 224768
rect 190642 224712 190698 224768
rect 189906 220360 189962 220416
rect 192298 221196 192354 221232
rect 192298 221176 192300 221196
rect 192300 221176 192352 221196
rect 192352 221176 192354 221196
rect 192482 220652 192538 220688
rect 192482 220632 192484 220652
rect 192484 220632 192536 220652
rect 192536 220632 192538 220652
rect 193494 224168 193550 224224
rect 194046 220632 194102 220688
rect 196070 229472 196126 229528
rect 196346 221176 196402 221232
rect 199198 224168 199254 224224
rect 200118 221992 200174 222048
rect 199474 221040 199530 221096
rect 200302 221040 200358 221096
rect 199658 220788 199714 220824
rect 199658 220768 199660 220788
rect 199660 220768 199712 220788
rect 199712 220768 199714 220788
rect 202602 229356 202658 229392
rect 202602 229336 202604 229356
rect 202604 229336 202656 229356
rect 202656 229336 202658 229356
rect 201958 220768 202014 220824
rect 202326 219700 202382 219736
rect 202326 219680 202328 219700
rect 202328 219680 202380 219700
rect 202380 219680 202382 219700
rect 204534 229336 204590 229392
rect 204350 220088 204406 220144
rect 204994 219408 205050 219464
rect 206834 224340 206836 224360
rect 206836 224340 206888 224360
rect 206888 224340 206890 224360
rect 206834 224304 206890 224340
rect 205914 221992 205970 222048
rect 205914 219700 205970 219736
rect 205914 219680 205916 219700
rect 205916 219680 205968 219700
rect 205968 219680 205970 219700
rect 205638 219408 205694 219464
rect 208766 224304 208822 224360
rect 209686 219836 209742 219872
rect 209686 219816 209688 219836
rect 209688 219816 209740 219836
rect 209740 219816 209742 219836
rect 209870 219836 209926 219872
rect 209870 219816 209872 219836
rect 209872 219816 209924 219836
rect 209924 219816 209926 219836
rect 212354 225256 212410 225312
rect 213366 222808 213422 222864
rect 214102 229472 214158 229528
rect 214654 229472 214710 229528
rect 214746 225292 214748 225312
rect 214748 225292 214800 225312
rect 214800 225292 214802 225312
rect 214746 225256 214802 225292
rect 214378 224848 214434 224904
rect 214746 222808 214802 222864
rect 215574 224848 215630 224904
rect 219346 220108 219402 220144
rect 219346 220088 219348 220108
rect 219348 220088 219400 220108
rect 219400 220088 219402 220108
rect 220082 220088 220138 220144
rect 437294 221176 437350 221232
rect 442906 220088 442962 220144
rect 449898 220360 449954 220416
rect 458086 221992 458142 222048
rect 459374 225256 459430 225312
rect 462778 222808 462834 222864
rect 467562 226072 467618 226128
rect 474462 219544 474518 219600
rect 476578 219564 476634 219600
rect 476578 219544 476580 219564
rect 476580 219544 476632 219564
rect 476632 219544 476634 219564
rect 481086 224576 481142 224632
rect 479982 224304 480038 224360
rect 481086 224304 481142 224360
rect 483294 230324 483296 230344
rect 483296 230324 483348 230344
rect 483348 230324 483350 230344
rect 483294 230288 483350 230324
rect 483294 229472 483350 229528
rect 481454 224576 481510 224632
rect 481454 221176 481510 221232
rect 480350 219544 480406 219600
rect 483386 223080 483442 223136
rect 484766 230560 484822 230616
rect 486422 227704 486478 227760
rect 511814 245520 511870 245576
rect 511262 243072 511318 243128
rect 510894 235728 510950 235784
rect 510618 233280 510674 233336
rect 491390 230560 491446 230616
rect 488446 230288 488502 230344
rect 489182 229472 489238 229528
rect 486790 224984 486846 225040
rect 485226 224440 485282 224496
rect 485870 223116 485872 223136
rect 485872 223116 485924 223136
rect 485924 223116 485926 223136
rect 485870 223080 485926 223116
rect 485870 221176 485926 221232
rect 485870 220632 485926 220688
rect 485870 219564 485926 219600
rect 485870 219544 485872 219564
rect 485872 219544 485924 219564
rect 485924 219544 485926 219564
rect 484858 216688 484914 216744
rect 489090 224440 489146 224496
rect 488538 220632 488594 220688
rect 489918 226616 489974 226672
rect 489550 226344 489606 226400
rect 490010 226344 490066 226400
rect 489734 224984 489790 225040
rect 489918 224984 489974 225040
rect 490930 226616 490986 226672
rect 489274 223080 489330 223136
rect 490838 223352 490894 223408
rect 491574 227704 491630 227760
rect 490286 220360 490342 220416
rect 490286 218048 490342 218104
rect 491666 220904 491722 220960
rect 492770 224984 492826 225040
rect 493322 220088 493378 220144
rect 495254 223080 495310 223136
rect 495254 221176 495310 221232
rect 495254 220496 495310 220552
rect 494794 218320 494850 218376
rect 495070 218320 495126 218376
rect 493322 217776 493378 217832
rect 496818 220496 496874 220552
rect 497462 218592 497518 218648
rect 499578 224576 499634 224632
rect 499302 224304 499358 224360
rect 499670 224304 499726 224360
rect 499532 223352 499588 223408
rect 499302 223080 499358 223136
rect 499670 223080 499726 223136
rect 499762 221176 499818 221232
rect 499946 221176 500002 221232
rect 488170 217232 488226 217288
rect 485778 216960 485834 217016
rect 486882 216960 486938 217016
rect 505190 224576 505246 224632
rect 504730 223352 504786 223408
rect 502338 219952 502394 220008
rect 504730 221176 504786 221232
rect 505098 219836 505154 219872
rect 505098 219816 505100 219836
rect 505100 219816 505152 219836
rect 505152 219816 505154 219836
rect 504178 217776 504234 217832
rect 507766 219408 507822 219464
rect 510066 223352 510122 223408
rect 511998 220244 512054 220280
rect 511998 220224 512000 220244
rect 512000 220224 512052 220244
rect 512052 220224 512054 220244
rect 512642 220224 512698 220280
rect 504178 217232 504234 217288
rect 514574 223352 514630 223408
rect 517426 223352 517482 223408
rect 513838 216416 513894 216472
rect 521658 221992 521714 222048
rect 525062 225256 525118 225312
rect 524234 224612 524236 224632
rect 524236 224612 524288 224632
rect 524288 224612 524290 224632
rect 524234 224576 524290 224612
rect 524234 223352 524290 223408
rect 526350 224576 526406 224632
rect 525062 219952 525118 220008
rect 530398 222808 530454 222864
rect 520646 216436 520702 216472
rect 520646 216416 520648 216436
rect 520648 216416 520700 216436
rect 520700 216416 520702 216436
rect 526074 216436 526130 216472
rect 526074 216416 526076 216436
rect 526076 216416 526128 216436
rect 526128 216416 526130 216436
rect 531226 216436 531282 216472
rect 533526 219952 533582 220008
rect 533066 219680 533122 219736
rect 537482 226072 537538 226128
rect 535366 218864 535422 218920
rect 531226 216416 531228 216436
rect 531228 216416 531280 216436
rect 531280 216416 531282 216436
rect 537390 216436 537446 216472
rect 541162 217504 541218 217560
rect 542082 217606 542138 217662
rect 542542 219136 542598 219192
rect 542496 217504 542552 217560
rect 543462 219136 543518 219192
rect 543646 217504 543702 217560
rect 545762 220768 545818 220824
rect 544382 219136 544438 219192
rect 546130 217504 546186 217560
rect 548154 220516 548210 220552
rect 548154 220496 548156 220516
rect 548156 220496 548208 220516
rect 548208 220496 548210 220516
rect 547970 217504 548026 217560
rect 549350 220768 549406 220824
rect 548890 220496 548946 220552
rect 552662 219136 552718 219192
rect 550638 217776 550694 217832
rect 537390 216416 537392 216436
rect 537392 216416 537444 216436
rect 537444 216416 537446 216436
rect 545670 216436 545726 216472
rect 545670 216416 545672 216436
rect 545672 216416 545724 216436
rect 545724 216416 545726 216436
rect 546774 216436 546830 216472
rect 546774 216416 546776 216436
rect 546776 216416 546828 216436
rect 546828 216416 546830 216436
rect 549442 216416 549498 216472
rect 553490 219136 553546 219192
rect 554962 220496 555018 220552
rect 556986 219136 557042 219192
rect 556802 217796 556858 217832
rect 556802 217776 556804 217796
rect 556804 217776 556856 217796
rect 556856 217776 556858 217796
rect 560114 217776 560170 217832
rect 560574 220768 560630 220824
rect 561034 217776 561090 217832
rect 562322 221040 562378 221096
rect 562138 220768 562194 220824
rect 562966 220652 563022 220654
rect 562966 220600 562968 220652
rect 562968 220600 563020 220652
rect 563020 220600 563022 220652
rect 562966 220598 563022 220600
rect 562506 219136 562562 219192
rect 563426 219136 563482 219192
rect 564070 221040 564126 221096
rect 563150 217776 563206 217832
rect 563426 217776 563482 217832
rect 563702 217776 563758 217832
rect 572442 220768 572498 220824
rect 572626 220768 572682 220824
rect 575110 220768 575166 220824
rect 572534 220516 572590 220552
rect 572534 220496 572536 220516
rect 572536 220496 572588 220516
rect 572588 220496 572590 220516
rect 572258 220360 572314 220416
rect 572442 220224 572498 220280
rect 572442 219680 572498 219736
rect 572166 219136 572222 219192
rect 573730 219136 573786 219192
rect 572626 217776 572682 217832
rect 553950 216436 554006 216472
rect 553950 216416 553952 216436
rect 553952 216416 554004 216436
rect 554004 216416 554006 216436
rect 556986 216416 557042 216472
rect 574650 218320 574706 218376
rect 574466 217776 574522 217832
rect 574466 217504 574522 217560
rect 574006 216144 574062 216200
rect 574466 216144 574522 216200
rect 574558 215872 574614 215928
rect 575846 220496 575902 220552
rect 576030 220224 576086 220280
rect 575478 216144 575534 216200
rect 576766 216416 576822 216472
rect 576582 215736 576638 215792
rect 576030 215328 576086 215384
rect 47582 203224 47638 203280
rect 41786 183368 41842 183424
rect 578698 216008 578754 216064
rect 578514 212744 578570 212800
rect 579250 214240 579306 214296
rect 586702 215484 586758 215520
rect 586702 215464 586704 215484
rect 586704 215464 586756 215484
rect 586756 215464 586758 215484
rect 586610 215192 586666 215248
rect 594062 215192 594118 215248
rect 578882 211148 578884 211168
rect 578884 211148 578936 211168
rect 578936 211148 578938 211168
rect 578882 211112 578938 211148
rect 579250 209788 579252 209808
rect 579252 209788 579304 209808
rect 579304 209788 579306 209808
rect 579250 209752 579306 209788
rect 578422 208256 578478 208312
rect 578698 206760 578754 206816
rect 579066 205284 579122 205320
rect 579066 205264 579068 205284
rect 579068 205264 579120 205284
rect 579120 205264 579122 205284
rect 578698 203768 578754 203824
rect 578238 202272 578294 202328
rect 578514 200776 578570 200832
rect 578882 199280 578938 199336
rect 578330 197784 578386 197840
rect 579250 196288 579306 196344
rect 578882 194792 578938 194848
rect 578514 193452 578570 193488
rect 578514 193432 578516 193452
rect 578516 193432 578568 193452
rect 578568 193432 578570 193452
rect 578238 190304 578294 190360
rect 578514 187312 578570 187368
rect 579526 191836 579528 191856
rect 579528 191836 579580 191856
rect 579580 191836 579582 191856
rect 579526 191800 579582 191836
rect 579250 188828 579306 188864
rect 579250 188808 579252 188828
rect 579252 188808 579304 188828
rect 579304 188808 579306 188828
rect 596270 215872 596326 215928
rect 595810 215736 595866 215792
rect 595994 215600 596050 215656
rect 596638 215620 596694 215656
rect 596638 215600 596640 215620
rect 596640 215600 596692 215620
rect 596692 215600 596694 215620
rect 600502 215872 600558 215928
rect 614026 219952 614082 220008
rect 613382 218864 613438 218920
rect 612278 218048 612334 218104
rect 611726 216960 611782 217016
rect 612830 217232 612886 217288
rect 614946 219680 615002 219736
rect 615498 219408 615554 219464
rect 631046 218592 631102 218648
rect 631598 216688 631654 216744
rect 642730 271088 642786 271144
rect 648710 276664 648766 276720
rect 647330 228792 647386 228848
rect 648066 227160 648122 227216
rect 651102 227432 651158 227488
rect 651562 975840 651618 975896
rect 651562 962512 651618 962568
rect 651562 949320 651618 949376
rect 651562 936128 651618 936184
rect 651562 922664 651618 922720
rect 651562 909492 651618 909528
rect 651562 909472 651564 909492
rect 651564 909472 651616 909492
rect 651616 909472 651618 909492
rect 651562 896144 651618 896200
rect 651562 869624 651618 869680
rect 651562 856296 651618 856352
rect 651562 842968 651618 843024
rect 651562 829776 651618 829832
rect 651562 816448 651618 816504
rect 651562 803276 651618 803312
rect 651562 803256 651564 803276
rect 651564 803256 651616 803276
rect 651616 803256 651618 803276
rect 651562 789928 651618 789984
rect 651562 776600 651618 776656
rect 651562 763292 651618 763328
rect 651562 763272 651564 763292
rect 651564 763272 651616 763292
rect 651616 763272 651618 763292
rect 651562 750080 651618 750136
rect 651562 736752 651618 736808
rect 651562 723424 651618 723480
rect 651562 710232 651618 710288
rect 651562 696940 651564 696960
rect 651564 696940 651616 696960
rect 651616 696940 651618 696960
rect 651562 696904 651618 696940
rect 651562 683576 651618 683632
rect 651562 670384 651618 670440
rect 651562 657056 651618 657112
rect 651562 643728 651618 643784
rect 651562 630536 651618 630592
rect 651562 617208 651618 617264
rect 651562 590708 651618 590744
rect 651562 590688 651564 590708
rect 651564 590688 651616 590708
rect 651616 590688 651618 590708
rect 651562 577360 651618 577416
rect 651562 550840 651618 550896
rect 651562 537512 651618 537568
rect 651562 524184 651618 524240
rect 651562 510992 651618 511048
rect 651562 497664 651618 497720
rect 651562 484492 651618 484528
rect 651562 484472 651564 484492
rect 651564 484472 651616 484492
rect 651616 484472 651618 484492
rect 651562 471144 651618 471200
rect 651562 457816 651618 457872
rect 651562 444508 651618 444544
rect 651562 444488 651564 444508
rect 651564 444488 651616 444508
rect 651616 444488 651618 444508
rect 651562 431296 651618 431352
rect 651562 417968 651618 418024
rect 651562 404640 651618 404696
rect 651562 391448 651618 391504
rect 651562 378156 651564 378176
rect 651564 378156 651616 378176
rect 651616 378156 651618 378176
rect 651562 378120 651618 378156
rect 651562 364792 651618 364848
rect 651562 324944 651618 325000
rect 651562 311752 651618 311808
rect 651562 285232 651618 285288
rect 651562 228248 651618 228304
rect 652390 882816 652446 882872
rect 652574 603880 652630 603936
rect 652390 564032 652446 564088
rect 652022 351600 652078 351656
rect 652206 338272 652262 338328
rect 652206 298424 652262 298480
rect 589462 208120 589518 208176
rect 589462 206488 589518 206544
rect 589462 204856 589518 204912
rect 589462 203224 589518 203280
rect 589370 201592 589426 201648
rect 589462 199996 589464 200016
rect 589464 199996 589516 200016
rect 589516 199996 589518 200016
rect 589462 199960 589518 199996
rect 590382 198328 590438 198384
rect 589462 196696 589518 196752
rect 589462 195064 589518 195120
rect 589462 193432 589518 193488
rect 578330 185816 578386 185872
rect 579526 184320 579582 184376
rect 578882 182824 578938 182880
rect 578514 181348 578570 181384
rect 578514 181328 578516 181348
rect 578516 181328 578568 181348
rect 578568 181328 578570 181348
rect 578974 179832 579030 179888
rect 578606 178356 578662 178392
rect 578606 178336 578608 178356
rect 578608 178336 578660 178356
rect 578660 178336 578662 178356
rect 579526 176860 579582 176896
rect 579526 176840 579528 176860
rect 579528 176840 579580 176860
rect 579580 176840 579582 176860
rect 579434 175480 579490 175536
rect 578330 173848 578386 173904
rect 579066 172352 579122 172408
rect 579526 170856 579582 170912
rect 578238 169360 578294 169416
rect 579434 167864 579490 167920
rect 579066 166368 579122 166424
rect 579526 164348 579582 164384
rect 579526 164328 579528 164348
rect 579528 164328 579580 164348
rect 579580 164328 579582 164348
rect 578698 163376 578754 163432
rect 578882 161880 578938 161936
rect 578514 160384 578570 160440
rect 578698 152904 578754 152960
rect 579526 158888 579582 158944
rect 579434 157392 579490 157448
rect 579250 155896 579306 155952
rect 579250 154400 579306 154456
rect 579158 151408 579214 151464
rect 578882 149912 578938 149968
rect 579526 148416 579582 148472
rect 589646 191664 589702 191720
rect 589462 190168 589518 190224
rect 589462 188536 589518 188592
rect 589370 186904 589426 186960
rect 589462 185272 589518 185328
rect 590382 183504 590438 183560
rect 588542 182008 588598 182064
rect 589462 180376 589518 180432
rect 589554 178744 589610 178800
rect 589462 177112 589518 177168
rect 589462 175480 589518 175536
rect 589278 173868 589334 173904
rect 589278 173848 589280 173868
rect 589280 173848 589332 173868
rect 589332 173848 589334 173868
rect 589370 172216 589426 172272
rect 589462 170584 589518 170640
rect 589462 168952 589518 169008
rect 589462 167320 589518 167376
rect 589462 165572 589518 165608
rect 589462 165552 589464 165572
rect 589464 165552 589516 165572
rect 589516 165552 589518 165572
rect 589922 164056 589978 164112
rect 589462 162424 589518 162480
rect 589462 160792 589518 160848
rect 588726 159160 588782 159216
rect 579250 146920 579306 146976
rect 579434 145424 579490 145480
rect 578514 143928 578570 143984
rect 579526 142432 579582 142488
rect 578882 140936 578938 140992
rect 578238 134952 578294 135008
rect 578514 133456 578570 133512
rect 578422 131960 578478 132016
rect 578606 130464 578662 130520
rect 579526 139460 579582 139496
rect 579526 139440 579528 139460
rect 579528 139440 579580 139460
rect 579580 139440 579582 139460
rect 579250 137964 579306 138000
rect 579250 137944 579252 137964
rect 579252 137944 579304 137964
rect 579304 137944 579306 137964
rect 579066 136448 579122 136504
rect 589462 157528 589518 157584
rect 589370 154264 589426 154320
rect 589462 152632 589518 152688
rect 589462 151000 589518 151056
rect 589462 149368 589518 149424
rect 588542 146104 588598 146160
rect 579434 128968 579490 129024
rect 578330 127472 578386 127528
rect 578514 125976 578570 126032
rect 578882 124480 578938 124536
rect 578882 122984 578938 123040
rect 578330 117020 578386 117056
rect 578330 117000 578332 117020
rect 578332 117000 578384 117020
rect 578384 117000 578386 117020
rect 579526 121508 579582 121544
rect 579526 121488 579528 121508
rect 579528 121488 579580 121508
rect 579580 121488 579582 121508
rect 579250 119992 579306 120048
rect 579066 118496 579122 118552
rect 589462 147600 589518 147656
rect 590382 155896 590438 155952
rect 656898 276936 656954 276992
rect 654138 230016 654194 230072
rect 653034 228520 653090 228576
rect 654322 229744 654378 229800
rect 658462 265512 658518 265568
rect 659842 226888 659898 226944
rect 661498 225800 661554 225856
rect 662418 225528 662474 225584
rect 662878 222536 662934 222592
rect 663798 221448 663854 221504
rect 665178 273672 665234 273728
rect 665730 273672 665786 273728
rect 665546 273400 665602 273456
rect 666742 245656 666798 245712
rect 666742 245384 666798 245440
rect 666742 223896 666798 223952
rect 666558 184184 666614 184240
rect 589922 144472 589978 144528
rect 590014 142840 590070 142896
rect 589462 141208 589518 141264
rect 589462 139576 589518 139632
rect 589462 137964 589518 138000
rect 589462 137944 589464 137964
rect 589464 137944 589516 137964
rect 589516 137944 589518 137964
rect 589370 136312 589426 136368
rect 588726 134680 588782 134736
rect 589462 131416 589518 131472
rect 589462 129684 589464 129704
rect 589464 129684 589516 129704
rect 589516 129684 589518 129704
rect 589462 129648 589518 129684
rect 589462 128188 589464 128208
rect 589464 128188 589516 128208
rect 589516 128188 589518 128208
rect 589462 128152 589518 128188
rect 589738 126520 589794 126576
rect 590382 133048 590438 133104
rect 589922 124888 589978 124944
rect 589462 123256 589518 123312
rect 590382 121624 590438 121680
rect 589462 120028 589464 120048
rect 589464 120028 589516 120048
rect 589516 120028 589518 120048
rect 589462 119992 589518 120028
rect 588542 118360 588598 118416
rect 589462 116728 589518 116784
rect 589278 115096 589334 115152
rect 589462 113464 589518 113520
rect 589462 111732 589464 111752
rect 589464 111732 589516 111752
rect 589516 111732 589518 111752
rect 589462 111696 589518 111732
rect 589922 110200 589978 110256
rect 667846 684936 667902 684992
rect 667846 615848 667902 615904
rect 667018 187584 667074 187640
rect 668030 245656 668086 245712
rect 675390 966456 675446 966512
rect 672998 959112 673054 959168
rect 668582 773744 668638 773800
rect 669226 752936 669282 752992
rect 669042 730088 669098 730144
rect 669042 663448 669098 663504
rect 668398 245792 668454 245848
rect 668398 222264 668454 222320
rect 668214 197376 668270 197432
rect 668030 163104 668086 163160
rect 668214 135360 668270 135416
rect 669226 572056 669282 572112
rect 668766 563896 668822 563952
rect 668582 182688 668638 182744
rect 668582 177792 668638 177848
rect 668950 223624 669006 223680
rect 668766 158208 668822 158264
rect 668766 148416 668822 148472
rect 668766 145152 668822 145208
rect 668766 143520 668822 143576
rect 668766 140256 668822 140312
rect 668766 138624 668822 138680
rect 668306 130464 668362 130520
rect 668214 125568 668270 125624
rect 668030 123936 668086 123992
rect 668306 112512 668362 112568
rect 666742 109316 666798 109372
rect 589462 108568 589518 108624
rect 589370 106936 589426 106992
rect 589278 105304 589334 105360
rect 589370 103672 589426 103728
rect 669134 221720 669190 221776
rect 669318 209888 669374 209944
rect 669226 133764 669228 133784
rect 669228 133764 669280 133784
rect 669280 133764 669282 133784
rect 669226 133728 669282 133764
rect 670422 872208 670478 872264
rect 670054 774968 670110 775024
rect 670054 710640 670110 710696
rect 670422 752664 670478 752720
rect 669594 208256 669650 208312
rect 670146 607144 670202 607200
rect 670330 606872 670386 606928
rect 670238 548392 670294 548448
rect 670238 342216 670294 342272
rect 671802 867992 671858 868048
rect 671710 733624 671766 733680
rect 675758 965096 675814 965152
rect 675206 963328 675262 963384
rect 674102 952176 674158 952232
rect 674102 933408 674158 933464
rect 674286 932184 674342 932240
rect 675758 961968 675814 962024
rect 674930 959384 674986 959440
rect 675114 959112 675170 959168
rect 675758 958296 675814 958352
rect 675758 956392 675814 956448
rect 674930 948912 674986 948968
rect 675482 952176 675538 952232
rect 677506 951496 677562 951552
rect 674930 941840 674986 941896
rect 674930 939528 674986 939584
rect 674930 937896 674986 937952
rect 675850 941840 675906 941896
rect 675482 939936 675538 939992
rect 675298 939120 675354 939176
rect 675482 938732 675538 938768
rect 675482 938712 675484 938732
rect 675484 938712 675536 938732
rect 675536 938712 675538 938732
rect 675482 938304 675538 938360
rect 675298 937488 675354 937544
rect 675482 937080 675538 937136
rect 675666 936672 675722 936728
rect 675482 936264 675538 936320
rect 675298 935856 675354 935912
rect 675850 934632 675906 934688
rect 675114 934088 675170 934144
rect 675482 933816 675538 933872
rect 675482 933020 675538 933056
rect 675482 933000 675484 933020
rect 675484 933000 675536 933020
rect 675536 933000 675538 933020
rect 674654 932592 674710 932648
rect 674470 931368 674526 931424
rect 683302 950000 683358 950056
rect 677506 931096 677562 931152
rect 675482 930164 675538 930200
rect 675482 930144 675484 930164
rect 675484 930144 675536 930164
rect 675536 930144 675538 930164
rect 683302 935584 683358 935640
rect 682382 935176 682438 935232
rect 675482 929736 675538 929792
rect 683118 929464 683174 929520
rect 675482 928512 675538 928568
rect 675758 877104 675814 877160
rect 675298 876424 675354 876480
rect 675390 873976 675446 874032
rect 672630 873568 672686 873624
rect 675390 873568 675446 873624
rect 672354 751304 672410 751360
rect 671710 643456 671766 643512
rect 671158 377712 671214 377768
rect 671066 212608 671122 212664
rect 670882 210432 670938 210488
rect 670790 209616 670846 209672
rect 669962 169632 670018 169688
rect 669226 128832 669282 128888
rect 669686 120672 669742 120728
rect 669226 119040 669282 119096
rect 670606 193568 670662 193624
rect 672538 734168 672594 734224
rect 672170 625096 672226 625152
rect 672722 688608 672778 688664
rect 672538 645360 672594 645416
rect 671986 553424 672042 553480
rect 671250 155080 671306 155136
rect 671802 247016 671858 247072
rect 672354 586200 672410 586256
rect 673458 732672 673514 732728
rect 675390 872208 675446 872264
rect 675666 869624 675722 869680
rect 674838 869488 674894 869544
rect 675482 867992 675538 868048
rect 675298 784216 675354 784272
rect 675114 783944 675170 784000
rect 674654 772384 674710 772440
rect 674654 772112 674710 772168
rect 675482 774968 675538 775024
rect 675482 773744 675538 773800
rect 675114 770616 675170 770672
rect 674930 766536 674986 766592
rect 679622 772656 679678 772712
rect 676034 772384 676090 772440
rect 675850 772132 675906 772168
rect 675850 772112 675852 772132
rect 675852 772112 675904 772132
rect 675904 772112 675906 772132
rect 675850 770616 675906 770672
rect 675482 761504 675538 761560
rect 675298 761096 675354 761152
rect 675482 760688 675538 760744
rect 675298 760300 675354 760336
rect 675298 760280 675300 760300
rect 675300 760280 675352 760300
rect 675352 760280 675354 760300
rect 675482 759892 675538 759928
rect 675482 759872 675484 759892
rect 675484 759872 675536 759892
rect 675536 759872 675538 759892
rect 675482 759500 675484 759520
rect 675484 759500 675536 759520
rect 675536 759500 675538 759520
rect 675482 759464 675538 759500
rect 675482 759076 675538 759112
rect 675482 759056 675484 759076
rect 675484 759056 675536 759076
rect 675536 759056 675538 759076
rect 675482 758684 675484 758704
rect 675484 758684 675536 758704
rect 675536 758684 675538 758704
rect 675482 758648 675538 758684
rect 675482 758260 675538 758296
rect 675482 758240 675484 758260
rect 675484 758240 675536 758260
rect 675536 758240 675538 758260
rect 675482 757868 675484 757888
rect 675484 757868 675536 757888
rect 675536 757868 675538 757888
rect 675482 757832 675538 757868
rect 675482 757444 675538 757480
rect 675482 757424 675484 757444
rect 675484 757424 675536 757444
rect 675536 757424 675538 757444
rect 682382 768712 682438 768768
rect 679622 756200 679678 756256
rect 675850 755792 675906 755848
rect 682382 755384 682438 755440
rect 675482 755012 675484 755032
rect 675484 755012 675536 755032
rect 675536 755012 675538 755032
rect 675482 754976 675538 755012
rect 675482 754604 675484 754624
rect 675484 754604 675536 754624
rect 675536 754604 675538 754624
rect 675482 754568 675538 754604
rect 675482 754196 675484 754216
rect 675484 754196 675536 754216
rect 675536 754196 675538 754216
rect 675482 754160 675538 754196
rect 675114 753752 675170 753808
rect 675482 753380 675484 753400
rect 675484 753380 675536 753400
rect 675536 753380 675538 753400
rect 675482 753344 675538 753380
rect 684130 756608 684186 756664
rect 675850 752936 675906 752992
rect 683302 752936 683358 752992
rect 674930 752392 674986 752448
rect 675482 752156 675484 752176
rect 675484 752156 675536 752176
rect 675536 752156 675538 752176
rect 675482 752120 675538 752156
rect 675482 751748 675484 751768
rect 675484 751748 675536 751768
rect 675536 751748 675538 751768
rect 675482 751712 675538 751748
rect 683118 750692 683174 750748
rect 675482 750100 675538 750136
rect 675482 750080 675484 750100
rect 675484 750080 675536 750100
rect 675536 750080 675538 750100
rect 674194 727504 674250 727560
rect 674010 683032 674066 683088
rect 674654 728048 674710 728104
rect 675114 738112 675170 738168
rect 675114 732944 675170 733000
rect 675482 734168 675538 734224
rect 675482 733624 675538 733680
rect 675482 732672 675538 732728
rect 675114 730088 675170 730144
rect 675850 728048 675906 728104
rect 677506 728048 677562 728104
rect 676034 727504 676090 727560
rect 674838 721520 674894 721576
rect 675482 716524 675484 716544
rect 675484 716524 675536 716544
rect 675536 716524 675538 716544
rect 675482 716488 675538 716524
rect 675298 716080 675354 716136
rect 675114 715300 675116 715320
rect 675116 715300 675168 715320
rect 675168 715300 675170 715320
rect 675114 715264 675170 715300
rect 675482 715672 675538 715728
rect 675482 714876 675538 714912
rect 675482 714856 675484 714876
rect 675484 714856 675536 714876
rect 675536 714856 675538 714876
rect 675482 714484 675484 714504
rect 675484 714484 675536 714504
rect 675536 714484 675538 714504
rect 675482 714448 675538 714484
rect 675482 714060 675538 714096
rect 675482 714040 675484 714060
rect 675484 714040 675536 714060
rect 675536 714040 675538 714060
rect 675482 713668 675484 713688
rect 675484 713668 675536 713688
rect 675536 713668 675538 713688
rect 675482 713632 675538 713668
rect 676770 713432 676826 713488
rect 675482 713244 675538 713280
rect 675482 713224 675484 713244
rect 675484 713224 675536 713244
rect 675536 713224 675538 713244
rect 675482 712852 675484 712872
rect 675484 712852 675536 712872
rect 675536 712852 675538 712872
rect 675482 712816 675538 712852
rect 675482 712428 675538 712464
rect 675482 712408 675484 712428
rect 675484 712408 675536 712428
rect 675536 712408 675538 712428
rect 676034 712000 676090 712056
rect 683394 727776 683450 727832
rect 676034 711592 676090 711648
rect 675482 711220 675484 711240
rect 675484 711220 675536 711240
rect 675536 711220 675538 711240
rect 675482 711184 675538 711220
rect 675850 710640 675906 710696
rect 675298 710368 675354 710424
rect 675482 709960 675538 710016
rect 675482 709588 675484 709608
rect 675484 709588 675536 709608
rect 675536 709588 675538 709608
rect 675482 709552 675538 709588
rect 675482 707956 675484 707976
rect 675484 707956 675536 707976
rect 675536 707956 675538 707976
rect 675482 707920 675538 707956
rect 675482 707548 675484 707568
rect 675484 707548 675536 707568
rect 675536 707548 675538 707568
rect 675482 707512 675538 707548
rect 675482 707140 675484 707160
rect 675484 707140 675536 707160
rect 675536 707140 675538 707160
rect 675482 707104 675538 707140
rect 675482 706732 675484 706752
rect 675484 706732 675536 706752
rect 675536 706732 675538 706752
rect 675482 706696 675538 706732
rect 684222 710776 684278 710832
rect 683394 709144 683450 709200
rect 683210 708328 683266 708384
rect 683118 705472 683174 705528
rect 675482 705084 675538 705120
rect 675482 705064 675484 705084
rect 675484 705064 675536 705084
rect 675536 705064 675538 705084
rect 675390 698536 675446 698592
rect 675390 696768 675446 696824
rect 675666 694320 675722 694376
rect 674470 663992 674526 664048
rect 674102 644272 674158 644328
rect 674010 640464 674066 640520
rect 673642 637064 673698 637120
rect 672722 598440 672778 598496
rect 673826 618568 673882 618624
rect 673458 592864 673514 592920
rect 673918 599120 673974 599176
rect 674470 644680 674526 644736
rect 674286 617752 674342 617808
rect 673826 597352 673882 597408
rect 675482 688608 675538 688664
rect 675022 685208 675078 685264
rect 675482 684936 675538 684992
rect 675850 683032 675906 683088
rect 674838 669296 674894 669352
rect 674838 649188 674894 649224
rect 674838 649168 674840 649188
rect 674840 649168 674892 649188
rect 674892 649168 674894 649188
rect 674838 643048 674894 643104
rect 674838 639376 674894 639432
rect 678242 678272 678298 678328
rect 675298 671336 675354 671392
rect 675482 670928 675538 670984
rect 675666 670520 675722 670576
rect 675298 670112 675354 670168
rect 675482 669704 675538 669760
rect 675298 668888 675354 668944
rect 675482 668516 675484 668536
rect 675484 668516 675536 668536
rect 675536 668516 675538 668536
rect 675482 668480 675538 668516
rect 675482 668092 675538 668128
rect 675482 668072 675484 668092
rect 675484 668072 675536 668092
rect 675536 668072 675538 668092
rect 675482 667700 675484 667720
rect 675484 667700 675536 667720
rect 675536 667700 675538 667720
rect 675482 667664 675538 667700
rect 675482 667276 675538 667312
rect 675482 667256 675484 667276
rect 675484 667256 675536 667276
rect 675536 667256 675538 667276
rect 683210 674056 683266 674112
rect 678242 666984 678298 667040
rect 675298 666440 675354 666496
rect 675482 666068 675484 666088
rect 675484 666068 675536 666088
rect 675536 666068 675538 666088
rect 675482 666032 675538 666068
rect 675482 665624 675538 665680
rect 675482 664844 675484 664864
rect 675484 664844 675536 664864
rect 675536 664844 675538 664864
rect 675482 664808 675538 664844
rect 675482 664400 675538 664456
rect 675850 663448 675906 663504
rect 675482 663212 675484 663232
rect 675484 663212 675536 663232
rect 675536 663212 675538 663232
rect 675482 663176 675538 663212
rect 675482 662804 675484 662824
rect 675484 662804 675536 662824
rect 675536 662804 675538 662824
rect 675482 662768 675538 662804
rect 675482 661988 675484 662008
rect 675484 661988 675536 662008
rect 675536 661988 675538 662008
rect 675482 661952 675538 661988
rect 675482 661580 675484 661600
rect 675484 661580 675536 661600
rect 675536 661580 675538 661600
rect 675482 661544 675538 661580
rect 675482 661156 675538 661192
rect 675482 661136 675484 661156
rect 675484 661136 675536 661156
rect 675536 661136 675538 661156
rect 675482 659948 675484 659968
rect 675484 659948 675536 659968
rect 675536 659948 675538 659968
rect 675482 659912 675538 659948
rect 683394 663720 683450 663776
rect 683210 662496 683266 662552
rect 683118 660048 683174 660104
rect 675574 652840 675630 652896
rect 675482 649168 675538 649224
rect 675574 648624 675630 648680
rect 675298 645768 675354 645824
rect 675482 645360 675538 645416
rect 675390 644680 675446 644736
rect 675390 644272 675446 644328
rect 675482 643456 675538 643512
rect 675482 643048 675538 643104
rect 675482 640464 675538 640520
rect 675390 639376 675446 639432
rect 675206 638152 675262 638208
rect 675758 638152 675814 638208
rect 675298 637744 675354 637800
rect 675574 637608 675630 637664
rect 675022 637336 675078 637392
rect 675114 625912 675170 625968
rect 674838 623872 674894 623928
rect 676034 637336 676090 637392
rect 676034 637064 676090 637120
rect 675574 631352 675630 631408
rect 675482 626320 675538 626376
rect 675482 625504 675538 625560
rect 675482 625096 675538 625152
rect 675482 624708 675538 624744
rect 675482 624688 675484 624708
rect 675484 624688 675536 624708
rect 675536 624688 675538 624708
rect 675482 624316 675484 624336
rect 675484 624316 675536 624336
rect 675536 624316 675538 624336
rect 675482 624280 675538 624316
rect 675482 623500 675484 623520
rect 675484 623500 675536 623520
rect 675536 623500 675538 623520
rect 675482 623464 675538 623500
rect 675482 623076 675538 623112
rect 675482 623056 675484 623076
rect 675484 623056 675536 623076
rect 675536 623056 675538 623076
rect 675482 622684 675484 622704
rect 675484 622684 675536 622704
rect 675536 622684 675538 622704
rect 675482 622648 675538 622684
rect 675482 622260 675538 622296
rect 675482 622240 675484 622260
rect 675484 622240 675536 622260
rect 675536 622240 675538 622260
rect 682566 621968 682622 622024
rect 682382 621560 682438 621616
rect 675022 619828 675024 619848
rect 675024 619828 675076 619848
rect 675076 619828 675078 619848
rect 675022 619792 675078 619828
rect 674654 617344 674710 617400
rect 683302 620744 683358 620800
rect 675482 620200 675538 620256
rect 675482 619384 675538 619440
rect 675666 618160 675722 618216
rect 675482 616972 675484 616992
rect 675484 616972 675536 616992
rect 675536 616972 675538 616992
rect 675482 616936 675538 616972
rect 675482 616564 675484 616584
rect 675484 616564 675536 616584
rect 675536 616564 675538 616584
rect 675482 616528 675538 616564
rect 675482 616140 675538 616176
rect 675482 616120 675484 616140
rect 675484 616120 675536 616140
rect 675536 616120 675538 616140
rect 675850 615848 675906 615904
rect 683118 615440 683174 615496
rect 675482 614916 675538 614952
rect 675482 614896 675484 614916
rect 675484 614896 675536 614916
rect 675536 614896 675538 614916
rect 674838 601160 674894 601216
rect 675390 607824 675446 607880
rect 675758 607280 675814 607336
rect 674930 597624 674986 597680
rect 675298 602928 675354 602984
rect 675390 601160 675446 601216
rect 675482 599120 675538 599176
rect 675482 598440 675538 598496
rect 675482 597352 675538 597408
rect 675022 594496 675078 594552
rect 674470 592184 674526 592240
rect 674194 591232 674250 591288
rect 675482 594768 675538 594824
rect 675850 592864 675906 592920
rect 675850 592492 675852 592512
rect 675852 592492 675904 592512
rect 675904 592492 675906 592512
rect 675850 592456 675906 592492
rect 675850 592184 675906 592240
rect 675850 591268 675852 591288
rect 675852 591268 675904 591288
rect 675904 591268 675906 591288
rect 675850 591232 675906 591268
rect 674930 580624 674986 580680
rect 674930 579400 674986 579456
rect 674194 547304 674250 547360
rect 674470 535064 674526 535120
rect 674286 533568 674342 533624
rect 674010 527584 674066 527640
rect 672630 474816 672686 474872
rect 672354 393216 672410 393272
rect 672814 389272 672870 389328
rect 672722 310800 672778 310856
rect 672630 217368 672686 217424
rect 672078 168272 672134 168328
rect 671986 168000 672042 168056
rect 669962 117408 670018 117464
rect 669226 115812 669228 115832
rect 669228 115812 669280 115832
rect 669280 115812 669282 115832
rect 669226 115776 669282 115812
rect 669226 114164 669282 114200
rect 669226 114144 669228 114164
rect 669228 114144 669280 114164
rect 669280 114144 669282 114164
rect 669042 110880 669098 110936
rect 668766 105984 668822 106040
rect 673090 286456 673146 286512
rect 673274 285504 673330 285560
rect 673090 278704 673146 278760
rect 673274 247696 673330 247752
rect 673090 214512 673146 214568
rect 672538 183504 672594 183560
rect 673274 200776 673330 200832
rect 674470 531936 674526 531992
rect 674286 490048 674342 490104
rect 674470 488416 674526 488472
rect 675298 586200 675354 586256
rect 675482 581052 675538 581088
rect 675482 581032 675484 581052
rect 675484 581032 675536 581052
rect 675536 581032 675538 581052
rect 675298 580216 675354 580272
rect 675482 579808 675538 579864
rect 675298 578992 675354 579048
rect 675482 578584 675538 578640
rect 675482 578176 675538 578232
rect 675298 577768 675354 577824
rect 675482 577360 675538 577416
rect 675482 576972 675538 577008
rect 675482 576952 675484 576972
rect 675484 576952 675536 576972
rect 675536 576952 675538 576972
rect 675482 576544 675538 576600
rect 682382 589192 682438 589248
rect 683302 576408 683358 576464
rect 682382 576000 682438 576056
rect 678242 575592 678298 575648
rect 675482 574912 675538 574968
rect 675298 574504 675354 574560
rect 675482 574116 675538 574152
rect 675482 574096 675484 574116
rect 675484 574096 675536 574116
rect 675536 574096 675538 574116
rect 675298 573688 675354 573744
rect 675482 572892 675538 572928
rect 675482 572872 675484 572892
rect 675484 572872 675536 572892
rect 675536 572872 675538 572892
rect 684130 572736 684186 572792
rect 683486 571920 683542 571976
rect 675298 571260 675354 571296
rect 675298 571240 675300 571260
rect 675300 571240 675352 571260
rect 675352 571240 675354 571260
rect 676218 570696 676274 570752
rect 675482 569628 675538 569664
rect 675482 569608 675484 569628
rect 675484 569608 675536 569628
rect 675536 569608 675538 569628
rect 683118 570288 683174 570344
rect 675850 563896 675906 563952
rect 675390 561856 675446 561912
rect 675482 559408 675538 559464
rect 675758 559000 675814 559056
rect 675390 553424 675446 553480
rect 675758 552064 675814 552120
rect 674930 547576 674986 547632
rect 674930 533976 674986 534032
rect 674930 531120 674986 531176
rect 674654 484336 674710 484392
rect 673918 376760 673974 376816
rect 673918 249600 673974 249656
rect 673918 215600 673974 215656
rect 673734 215328 673790 215384
rect 675114 508816 675170 508872
rect 675482 549616 675538 549672
rect 675482 548392 675538 548448
rect 675758 547848 675814 547904
rect 675482 536016 675538 536072
rect 675482 535492 675538 535528
rect 675482 535472 675484 535492
rect 675484 535472 675536 535492
rect 675536 535472 675538 535492
rect 675482 534792 675538 534848
rect 675482 534248 675538 534304
rect 675482 533332 675484 533352
rect 675484 533332 675536 533352
rect 675536 533332 675538 533352
rect 675482 533296 675538 533332
rect 675482 532772 675538 532808
rect 675482 532752 675484 532772
rect 675484 532752 675536 532772
rect 675536 532752 675538 532772
rect 675482 532516 675484 532536
rect 675484 532516 675536 532536
rect 675536 532516 675538 532536
rect 675482 532480 675538 532516
rect 675482 531528 675538 531584
rect 675482 530068 675484 530088
rect 675484 530068 675536 530088
rect 675536 530068 675538 530088
rect 675482 530032 675538 530068
rect 675482 529488 675538 529544
rect 675482 528436 675484 528456
rect 675484 528436 675536 528456
rect 675536 528436 675538 528456
rect 675482 528400 675538 528436
rect 675482 528028 675484 528048
rect 675484 528028 675536 528048
rect 675536 528028 675538 528048
rect 675482 527992 675538 528028
rect 675482 526804 675484 526824
rect 675484 526804 675536 526824
rect 675536 526804 675538 526824
rect 675482 526768 675538 526804
rect 675482 526396 675484 526416
rect 675484 526396 675536 526416
rect 675536 526396 675538 526416
rect 675482 526360 675538 526396
rect 675482 525836 675538 525872
rect 675482 525816 675484 525836
rect 675484 525816 675536 525836
rect 675536 525816 675538 525836
rect 675942 547576 675998 547632
rect 677506 547576 677562 547632
rect 676126 547304 676182 547360
rect 683394 547032 683450 547088
rect 679622 546760 679678 546816
rect 679622 530576 679678 530632
rect 677506 529352 677562 529408
rect 683394 530984 683450 531040
rect 683210 528944 683266 529000
rect 683118 525716 683120 525736
rect 683120 525716 683172 525736
rect 683172 525716 683174 525736
rect 683118 525680 683174 525716
rect 676034 508816 676090 508872
rect 675298 500248 675354 500304
rect 675298 492088 675354 492144
rect 675482 491680 675538 491736
rect 675482 491308 675484 491328
rect 675484 491308 675536 491328
rect 675536 491308 675538 491328
rect 675482 491272 675538 491308
rect 675482 490864 675538 490920
rect 675482 489232 675538 489288
rect 675666 488824 675722 488880
rect 675298 486784 675354 486840
rect 675482 485988 675538 486024
rect 675482 485968 675484 485988
rect 675484 485968 675536 485988
rect 675536 485968 675538 485988
rect 676034 500248 676090 500304
rect 676034 490456 676090 490512
rect 676034 489640 676090 489696
rect 676034 488008 676090 488064
rect 675850 487600 675906 487656
rect 675482 485596 675484 485616
rect 675484 485596 675536 485616
rect 675536 485596 675538 485616
rect 675482 485560 675538 485596
rect 675482 485152 675538 485208
rect 675482 483556 675484 483576
rect 675484 483556 675536 483576
rect 675536 483556 675538 483576
rect 675482 483520 675538 483556
rect 675482 483148 675484 483168
rect 675484 483148 675536 483168
rect 675536 483148 675538 483168
rect 675482 483112 675538 483148
rect 675482 482740 675484 482760
rect 675484 482740 675536 482760
rect 675536 482740 675538 482760
rect 675482 482704 675538 482740
rect 675482 482332 675484 482352
rect 675484 482332 675536 482352
rect 675536 482332 675538 482352
rect 675482 482296 675538 482332
rect 675482 481908 675538 481944
rect 675482 481888 675484 481908
rect 675484 481888 675536 481908
rect 675536 481888 675538 481908
rect 674930 481480 674986 481536
rect 675482 480684 675538 480720
rect 675482 480664 675484 480684
rect 675484 480664 675536 480684
rect 675536 480664 675538 480684
rect 675482 403824 675538 403880
rect 675298 403436 675354 403472
rect 675298 403416 675300 403436
rect 675300 403416 675352 403436
rect 675352 403416 675354 403436
rect 675482 403044 675484 403064
rect 675484 403044 675536 403064
rect 675536 403044 675538 403064
rect 675482 403008 675538 403044
rect 674654 402192 674710 402248
rect 674470 401376 674526 401432
rect 674286 393624 674342 393680
rect 675942 400968 675998 401024
rect 679622 487192 679678 487248
rect 679806 486376 679862 486432
rect 677414 402872 677470 402928
rect 677230 402056 677286 402112
rect 675482 400580 675538 400616
rect 675482 400560 675484 400580
rect 675484 400560 675536 400580
rect 675536 400560 675538 400580
rect 675942 400152 675998 400208
rect 675482 399764 675538 399800
rect 675482 399744 675484 399764
rect 675484 399744 675536 399764
rect 675536 399744 675538 399764
rect 674930 399336 674986 399392
rect 676218 398384 676274 398440
rect 675114 398112 675170 398168
rect 675482 397316 675538 397352
rect 675482 397296 675484 397316
rect 675484 397296 675536 397316
rect 675536 397296 675538 397316
rect 675482 396092 675538 396128
rect 675482 396072 675484 396092
rect 675484 396072 675536 396092
rect 675536 396072 675538 396092
rect 675482 395684 675538 395720
rect 675482 395664 675484 395684
rect 675484 395664 675536 395684
rect 675536 395664 675538 395684
rect 681002 397568 681058 397624
rect 675482 394460 675538 394496
rect 675482 394440 675484 394460
rect 675484 394440 675536 394460
rect 675536 394440 675538 394460
rect 675482 394052 675538 394088
rect 675482 394032 675484 394052
rect 675484 394032 675536 394052
rect 675536 394032 675538 394052
rect 675482 392420 675538 392456
rect 675482 392400 675484 392420
rect 675484 392400 675536 392420
rect 675536 392400 675538 392420
rect 675850 389272 675906 389328
rect 681186 396344 681242 396400
rect 681002 388456 681058 388512
rect 683118 392672 683174 392728
rect 681186 387640 681242 387696
rect 675298 383560 675354 383616
rect 675758 382200 675814 382256
rect 675758 380568 675814 380624
rect 675666 378528 675722 378584
rect 675758 377304 675814 377360
rect 674930 376760 674986 376816
rect 675298 374992 675354 375048
rect 675114 372544 675170 372600
rect 675298 358672 675354 358728
rect 675114 358264 675170 358320
rect 674654 357448 674710 357504
rect 675482 357856 675538 357912
rect 675482 357060 675538 357096
rect 675482 357040 675484 357060
rect 675484 357040 675536 357060
rect 675536 357040 675538 357060
rect 674470 356632 674526 356688
rect 674654 356224 674710 356280
rect 674470 351328 674526 351384
rect 675482 355852 675484 355872
rect 675484 355852 675536 355872
rect 675536 355852 675538 355872
rect 675482 355816 675538 355852
rect 675482 355428 675538 355464
rect 675482 355408 675484 355428
rect 675484 355408 675536 355428
rect 675536 355408 675538 355428
rect 675482 355036 675484 355056
rect 675484 355036 675536 355056
rect 675536 355036 675538 355056
rect 675482 355000 675538 355036
rect 675482 354612 675538 354648
rect 675482 354592 675484 354612
rect 675484 354592 675536 354612
rect 675536 354592 675538 354612
rect 675482 353776 675538 353832
rect 675482 353388 675538 353424
rect 675482 353368 675484 353388
rect 675484 353368 675536 353388
rect 675536 353368 675538 353388
rect 675482 352572 675538 352608
rect 675482 352552 675484 352572
rect 675484 352552 675536 352572
rect 675536 352552 675538 352572
rect 676034 350920 676090 350976
rect 675850 350512 675906 350568
rect 675482 350124 675538 350160
rect 675482 350104 675484 350124
rect 675484 350104 675536 350124
rect 675536 350104 675538 350124
rect 675482 349716 675538 349752
rect 675482 349696 675484 349716
rect 675484 349696 675536 349716
rect 675536 349696 675538 349716
rect 675482 349308 675538 349344
rect 675482 349288 675484 349308
rect 675484 349288 675536 349308
rect 675536 349288 675538 349308
rect 675482 348900 675538 348936
rect 675482 348880 675484 348900
rect 675484 348880 675536 348900
rect 675536 348880 675538 348900
rect 675482 348492 675538 348528
rect 675482 348472 675484 348492
rect 675484 348472 675536 348492
rect 675536 348472 675538 348492
rect 675482 347268 675538 347304
rect 675482 347248 675484 347268
rect 675484 347248 675536 347268
rect 675536 347248 675538 347268
rect 676034 346568 676090 346624
rect 683118 347656 683174 347712
rect 676586 346432 676642 346488
rect 675850 342216 675906 342272
rect 675758 340176 675814 340232
rect 675390 338952 675446 339008
rect 675666 337728 675722 337784
rect 675298 335280 675354 335336
rect 675298 331064 675354 331120
rect 675758 326848 675814 326904
rect 675482 313656 675538 313712
rect 675482 313284 675484 313304
rect 675484 313284 675536 313304
rect 675536 313284 675538 313304
rect 675482 313248 675538 313284
rect 675298 312840 675354 312896
rect 675482 312468 675484 312488
rect 675484 312468 675536 312488
rect 675536 312468 675538 312488
rect 675482 312432 675538 312468
rect 675482 312024 675538 312080
rect 674654 311616 674710 311672
rect 675482 311208 675538 311264
rect 675482 310412 675538 310448
rect 675482 310392 675484 310412
rect 675484 310392 675536 310412
rect 675536 310392 675538 310412
rect 675482 310020 675484 310040
rect 675484 310020 675536 310040
rect 675536 310020 675538 310040
rect 675482 309984 675538 310020
rect 675482 309576 675538 309632
rect 675206 309168 675262 309224
rect 675022 307944 675078 308000
rect 674838 307536 674894 307592
rect 674470 306312 674526 306368
rect 674654 304272 674710 304328
rect 676034 308352 676090 308408
rect 675482 305516 675538 305552
rect 675482 305496 675484 305516
rect 675484 305496 675536 305516
rect 675536 305496 675538 305516
rect 678242 307128 678298 307184
rect 675482 303884 675538 303920
rect 675482 303864 675484 303884
rect 675484 303864 675536 303884
rect 675536 303864 675538 303884
rect 675482 303476 675538 303512
rect 675482 303456 675484 303476
rect 675484 303456 675536 303476
rect 675536 303456 675538 303476
rect 675482 302252 675538 302288
rect 675482 302232 675484 302252
rect 675484 302232 675536 302252
rect 675536 302232 675538 302252
rect 675850 305088 675906 305144
rect 676034 304680 676090 304736
rect 676034 302912 676090 302968
rect 675850 301552 675906 301608
rect 681002 306720 681058 306776
rect 680358 299376 680414 299432
rect 678242 297336 678298 297392
rect 683118 302640 683174 302696
rect 675758 291488 675814 291544
rect 675758 290944 675814 291000
rect 675758 287000 675814 287056
rect 675390 286456 675446 286512
rect 675114 285504 675170 285560
rect 675758 283600 675814 283656
rect 675666 282784 675722 282840
rect 675666 281560 675722 281616
rect 675298 268640 675354 268696
rect 675482 268232 675538 268288
rect 675482 267844 675538 267880
rect 675482 267824 675484 267844
rect 675484 267824 675536 267844
rect 675536 267824 675538 267844
rect 675114 267416 675170 267472
rect 675298 267008 675354 267064
rect 675482 266636 675484 266656
rect 675484 266636 675536 266656
rect 675536 266636 675538 266656
rect 675482 266600 675538 266636
rect 675482 266192 675538 266248
rect 675298 265820 675300 265840
rect 675300 265820 675352 265840
rect 675352 265820 675354 265840
rect 675298 265784 675354 265820
rect 675482 265376 675538 265432
rect 675482 265004 675484 265024
rect 675484 265004 675536 265024
rect 675536 265004 675538 265024
rect 675482 264968 675538 265004
rect 675482 264560 675538 264616
rect 675022 264152 675078 264208
rect 674470 262112 674526 262168
rect 674654 258848 674710 258904
rect 674838 253952 674894 254008
rect 676218 263200 676274 263256
rect 675482 262948 675538 262984
rect 675482 262928 675484 262948
rect 675484 262928 675536 262948
rect 675536 262928 675538 262948
rect 675482 261316 675538 261352
rect 675482 261296 675484 261316
rect 675484 261296 675536 261316
rect 675536 261296 675538 261316
rect 675666 260480 675722 260536
rect 675482 260072 675538 260128
rect 675298 259664 675354 259720
rect 681002 262384 681058 262440
rect 675482 259276 675538 259312
rect 675482 259256 675484 259276
rect 675484 259256 675536 259276
rect 675536 259256 675538 259276
rect 675482 258460 675538 258496
rect 675482 258440 675484 258460
rect 675484 258440 675536 258460
rect 675536 258440 675538 258460
rect 675482 257216 675538 257272
rect 675942 253952 675998 254008
rect 683118 257488 683174 257544
rect 681002 252592 681058 252648
rect 675758 250144 675814 250200
rect 675114 249600 675170 249656
rect 675298 249600 675354 249656
rect 675482 247696 675538 247752
rect 675482 247016 675538 247072
rect 675758 246608 675814 246664
rect 675482 245928 675538 245984
rect 675390 238584 675446 238640
rect 675114 223488 675170 223544
rect 675482 223080 675538 223136
rect 675298 222672 675354 222728
rect 675482 222284 675538 222320
rect 675482 222264 675484 222284
rect 675484 222264 675536 222284
rect 675536 222264 675538 222284
rect 675114 221856 675170 221912
rect 675482 221448 675538 221504
rect 675298 221040 675354 221096
rect 675298 220632 675354 220688
rect 674654 220224 674710 220280
rect 674470 219408 674526 219464
rect 674470 198600 674526 198656
rect 674470 176024 674526 176080
rect 675482 219816 675538 219872
rect 674838 218184 674894 218240
rect 675298 217368 675354 217424
rect 675482 216960 675538 217016
rect 675114 216144 675170 216200
rect 675482 215736 675538 215792
rect 675298 215348 675354 215384
rect 675298 215328 675300 215348
rect 675300 215328 675352 215348
rect 675352 215328 675354 215348
rect 675482 214124 675538 214160
rect 675482 214104 675484 214124
rect 675484 214104 675536 214124
rect 675536 214104 675538 214124
rect 675482 213716 675538 213752
rect 675482 213696 675484 213716
rect 675484 213696 675536 213716
rect 675536 213696 675538 213716
rect 675482 213308 675538 213344
rect 675482 213288 675484 213308
rect 675484 213288 675536 213308
rect 675536 213288 675538 213308
rect 683118 212472 683174 212528
rect 675482 212064 675538 212120
rect 675850 209888 675906 209944
rect 675758 204992 675814 205048
rect 675666 204176 675722 204232
rect 675390 202680 675446 202736
rect 675758 199960 675814 200016
rect 675758 197104 675814 197160
rect 675758 193160 675814 193216
rect 675482 191528 675538 191584
rect 676034 185816 676090 185872
rect 675482 178472 675538 178528
rect 675482 178100 675484 178120
rect 675484 178100 675536 178120
rect 675536 178100 675538 178120
rect 675482 178064 675538 178100
rect 675482 177692 675484 177712
rect 675484 177692 675536 177712
rect 675536 177692 675538 177712
rect 675482 177656 675538 177692
rect 676034 177248 676090 177304
rect 675482 176860 675538 176896
rect 675482 176840 675484 176860
rect 675484 176840 675536 176860
rect 675536 176840 675538 176860
rect 675482 176432 675538 176488
rect 674654 175616 674710 175672
rect 675482 175228 675538 175264
rect 675482 175208 675484 175228
rect 675484 175208 675536 175228
rect 675536 175208 675538 175228
rect 675482 174412 675538 174448
rect 675482 174392 675484 174412
rect 675484 174392 675536 174412
rect 675536 174392 675538 174412
rect 675022 173984 675078 174040
rect 674470 171944 674526 172000
rect 674838 162152 674894 162208
rect 675850 173168 675906 173224
rect 675206 171536 675262 171592
rect 675482 171148 675538 171184
rect 675482 171128 675484 171148
rect 675484 171128 675536 171148
rect 675536 171128 675538 171148
rect 675482 169516 675538 169552
rect 675482 169496 675484 169516
rect 675484 169496 675536 169516
rect 675536 169496 675538 169516
rect 675482 169108 675538 169144
rect 675482 169088 675484 169108
rect 675484 169088 675536 169108
rect 675536 169088 675538 169108
rect 675482 168700 675538 168736
rect 675482 168680 675484 168700
rect 675484 168680 675536 168700
rect 675536 168680 675538 168700
rect 675666 167864 675722 167920
rect 675482 167068 675538 167104
rect 675482 167048 675484 167068
rect 675484 167048 675536 167068
rect 675536 167048 675538 167068
rect 676034 172760 676090 172816
rect 678242 172352 678298 172408
rect 676678 170720 676734 170776
rect 676402 169904 676458 169960
rect 676402 166368 676458 166424
rect 676678 166232 676734 166288
rect 676034 162152 676090 162208
rect 678242 161880 678298 161936
rect 675758 156304 675814 156360
rect 675666 153040 675722 153096
rect 675758 151408 675814 151464
rect 675758 150320 675814 150376
rect 675758 148416 675814 148472
rect 675666 147600 675722 147656
rect 675482 133356 675484 133376
rect 675484 133356 675536 133376
rect 675536 133356 675538 133376
rect 675482 133320 675538 133356
rect 675482 132932 675538 132968
rect 675482 132912 675484 132932
rect 675484 132912 675536 132932
rect 675536 132912 675538 132932
rect 675482 132504 675538 132560
rect 675482 132132 675484 132152
rect 675484 132132 675536 132152
rect 675536 132132 675538 132152
rect 675482 132096 675538 132132
rect 675482 131688 675538 131744
rect 674654 131280 674710 131336
rect 675482 130892 675538 130928
rect 675482 130872 675484 130892
rect 675484 130872 675536 130892
rect 675536 130872 675538 130892
rect 675482 130500 675484 130520
rect 675484 130500 675536 130520
rect 675536 130500 675538 130520
rect 675482 130464 675538 130500
rect 675482 130056 675538 130112
rect 675482 129684 675484 129704
rect 675484 129684 675536 129704
rect 675536 129684 675538 129704
rect 675482 129648 675538 129684
rect 675482 129240 675538 129296
rect 676218 128152 676274 128208
rect 674838 127608 674894 127664
rect 674378 125160 674434 125216
rect 674194 124752 674250 124808
rect 669134 107616 669190 107672
rect 674654 123528 674710 123584
rect 675482 125996 675538 126032
rect 675482 125976 675484 125996
rect 675484 125976 675536 125996
rect 675536 125976 675538 125996
rect 675482 125568 675538 125624
rect 675482 123956 675538 123992
rect 675482 123936 675484 123956
rect 675484 123936 675536 123956
rect 675536 123936 675538 123956
rect 675482 123140 675538 123176
rect 675482 123120 675484 123140
rect 675484 123120 675536 123140
rect 675536 123120 675538 123140
rect 676402 127744 676458 127800
rect 683118 126520 683174 126576
rect 679622 126112 679678 126168
rect 676218 122848 676274 122904
rect 675482 122460 675538 122496
rect 675482 122440 675484 122460
rect 675484 122440 675536 122460
rect 675536 122440 675538 122460
rect 677598 122032 677654 122088
rect 675482 121896 675538 121952
rect 683118 124480 683174 124536
rect 677598 116048 677654 116104
rect 675758 114144 675814 114200
rect 675758 110336 675814 110392
rect 675666 108024 675722 108080
rect 668950 104352 669006 104408
rect 675758 103128 675814 103184
rect 668582 102720 668638 102776
rect 675666 102584 675722 102640
rect 589462 102076 589464 102096
rect 589464 102076 589516 102096
rect 589516 102076 589518 102096
rect 589462 102040 589518 102076
rect 675758 101360 675814 101416
rect 131026 50224 131082 50280
rect 78586 49680 78642 49736
rect 151910 47232 151966 47288
rect 151910 45872 151966 45928
rect 187514 42064 187570 42120
rect 306976 42336 307032 42392
rect 310426 42064 310482 42120
rect 361946 42064 362002 42120
rect 365166 42064 365222 42120
rect 497554 50496 497610 50552
rect 445206 50224 445262 50280
rect 549258 50224 549314 50280
rect 415214 48048 415270 48104
rect 406382 45056 406438 45112
rect 411074 42744 411130 42800
rect 591302 47504 591358 47560
rect 451278 47232 451334 47288
rect 451462 47232 451518 47288
rect 461030 47252 461086 47288
rect 461030 47232 461032 47252
rect 461032 47232 461084 47252
rect 461084 47232 461086 47252
rect 451278 46688 451334 46744
rect 461214 47232 461270 47288
rect 470598 47232 470654 47288
rect 470782 47232 470838 47288
rect 461214 46688 461270 46744
rect 465722 46688 465778 46744
rect 451462 45872 451518 45928
rect 480442 47232 480498 47288
rect 480626 47232 480682 47288
rect 490010 47232 490066 47288
rect 490194 47232 490250 47288
rect 465906 45872 465962 45928
rect 470782 45872 470838 45928
rect 470966 45872 471022 45928
rect 480258 45872 480314 45928
rect 480442 45872 480498 45928
rect 465722 45736 465778 45792
rect 499762 47232 499818 47288
rect 499946 47232 500002 47288
rect 513746 47232 513802 47288
rect 514206 46960 514262 47016
rect 596178 48864 596234 48920
rect 595442 48048 595498 48104
rect 597558 47776 597614 47832
rect 600318 49136 600374 49192
rect 598938 47232 598994 47288
rect 600962 46688 601018 46744
rect 594062 46416 594118 46472
rect 592682 46144 592738 46200
rect 490194 45872 490250 45928
rect 490378 45872 490434 45928
rect 499578 45872 499634 45928
rect 499762 45872 499818 45928
rect 603078 51720 603134 51776
rect 601698 44784 601754 44840
rect 626078 94424 626134 94480
rect 637026 96872 637082 96928
rect 635922 95648 635978 95704
rect 626446 95376 626502 95432
rect 642638 95104 642694 95160
rect 626446 93472 626502 93528
rect 626262 92520 626318 92576
rect 625434 91568 625490 91624
rect 626446 90616 626502 90672
rect 626446 89684 626502 89720
rect 626446 89664 626448 89684
rect 626448 89664 626500 89684
rect 626500 89664 626502 89684
rect 624974 88304 625030 88360
rect 626446 87896 626502 87952
rect 625618 86944 625674 87000
rect 626446 85992 626502 86048
rect 626446 85040 626502 85096
rect 626446 84088 626502 84144
rect 626262 83136 626318 83192
rect 644478 92112 644534 92168
rect 644754 89664 644810 89720
rect 643558 87080 643614 87136
rect 643374 84632 643430 84688
rect 643098 82728 643154 82784
rect 628562 81640 628618 81696
rect 629206 80824 629262 80880
rect 633898 77696 633954 77752
rect 637118 78512 637174 78568
rect 646134 71712 646190 71768
rect 646870 74432 646926 74488
rect 647422 72936 647478 72992
rect 646318 70352 646374 70408
rect 647606 68448 647662 68504
rect 646134 66000 646190 66056
rect 653954 94152 654010 94208
rect 654322 93336 654378 93392
rect 654138 92520 654194 92576
rect 654322 91432 654378 91488
rect 654138 90616 654194 90672
rect 655794 89800 655850 89856
rect 663246 93064 663302 93120
rect 663798 90344 663854 90400
rect 663982 88984 664038 89040
rect 665178 93336 665234 93392
rect 665362 91704 665418 91760
rect 665546 90616 665602 90672
rect 649170 66952 649226 67008
rect 648802 63960 648858 64016
rect 661222 48184 661278 48240
rect 661590 47733 661646 47789
rect 474462 43424 474518 43480
rect 604458 43424 604514 43480
rect 662418 47368 662474 47424
rect 416594 42744 416650 42800
rect 464894 42744 464950 42800
rect 518530 42336 518586 42392
rect 460570 42064 460626 42120
rect 471610 42064 471666 42120
rect 514942 42064 514998 42120
rect 520462 42064 520518 42120
rect 525798 42064 525854 42120
rect 529570 42064 529626 42120
rect 521658 41928 521714 41984
<< metal3 >>
rect 357709 1007178 357775 1007181
rect 505001 1007178 505067 1007181
rect 357709 1007176 357972 1007178
rect 357709 1007120 357714 1007176
rect 357770 1007120 357972 1007176
rect 357709 1007118 357972 1007120
rect 504804 1007176 505067 1007178
rect 504804 1007120 505006 1007176
rect 505062 1007120 505067 1007176
rect 504804 1007118 505067 1007120
rect 357709 1007115 357775 1007118
rect 505001 1007115 505067 1007118
rect 425513 1007042 425579 1007045
rect 505369 1007042 505435 1007045
rect 551093 1007042 551159 1007045
rect 425513 1007040 425776 1007042
rect 425513 1006984 425518 1007040
rect 425574 1006984 425776 1007040
rect 425513 1006982 425776 1006984
rect 505172 1007040 505435 1007042
rect 505172 1006984 505374 1007040
rect 505430 1006984 505435 1007040
rect 505172 1006982 505435 1006984
rect 550436 1007040 551159 1007042
rect 550436 1006984 551098 1007040
rect 551154 1006984 551159 1007040
rect 550436 1006982 551159 1006984
rect 425513 1006979 425579 1006982
rect 505369 1006979 505435 1006982
rect 551093 1006979 551159 1006982
rect 357709 1006906 357775 1006909
rect 427537 1006906 427603 1006909
rect 503345 1006906 503411 1006909
rect 559649 1006906 559715 1006909
rect 357604 1006904 357775 1006906
rect 357604 1006848 357714 1006904
rect 357770 1006848 357775 1006904
rect 357604 1006846 357775 1006848
rect 427340 1006904 427603 1006906
rect 427340 1006848 427542 1006904
rect 427598 1006848 427603 1006904
rect 427340 1006846 427603 1006848
rect 503148 1006904 503411 1006906
rect 503148 1006848 503350 1006904
rect 503406 1006848 503411 1006904
rect 503148 1006846 503411 1006848
rect 559452 1006904 559715 1006906
rect 559452 1006848 559654 1006904
rect 559710 1006848 559715 1006904
rect 559452 1006846 559715 1006848
rect 357709 1006843 357775 1006846
rect 427537 1006843 427603 1006846
rect 503345 1006843 503411 1006846
rect 559649 1006843 559715 1006846
rect 358537 1006770 358603 1006773
rect 358340 1006768 358603 1006770
rect 358340 1006712 358542 1006768
rect 358598 1006712 358603 1006768
rect 358340 1006710 358603 1006712
rect 358537 1006707 358603 1006710
rect 430849 1006770 430915 1006773
rect 555969 1006770 556035 1006773
rect 430849 1006768 431020 1006770
rect 430849 1006712 430854 1006768
rect 430910 1006712 431020 1006768
rect 430849 1006710 431020 1006712
rect 555969 1006768 556232 1006770
rect 555969 1006712 555974 1006768
rect 556030 1006712 556232 1006768
rect 555969 1006710 556232 1006712
rect 430849 1006707 430915 1006710
rect 555969 1006707 556035 1006710
rect 103145 1006634 103211 1006637
rect 153745 1006634 153811 1006637
rect 102948 1006632 103211 1006634
rect 102948 1006576 103150 1006632
rect 103206 1006576 103211 1006632
rect 102948 1006574 103211 1006576
rect 153548 1006632 153811 1006634
rect 153548 1006576 153750 1006632
rect 153806 1006576 153811 1006632
rect 153548 1006574 153811 1006576
rect 103145 1006571 103211 1006574
rect 153745 1006571 153811 1006574
rect 306925 1006634 306991 1006637
rect 429193 1006634 429259 1006637
rect 506197 1006634 506263 1006637
rect 306925 1006632 307188 1006634
rect 306925 1006576 306930 1006632
rect 306986 1006576 307188 1006632
rect 306925 1006574 307188 1006576
rect 428996 1006632 429259 1006634
rect 428996 1006576 429198 1006632
rect 429254 1006576 429259 1006632
rect 428996 1006574 429259 1006576
rect 506000 1006632 506263 1006634
rect 506000 1006576 506202 1006632
rect 506258 1006576 506263 1006632
rect 506000 1006574 506263 1006576
rect 306925 1006571 306991 1006574
rect 429193 1006571 429259 1006574
rect 506197 1006571 506263 1006574
rect 103973 1006498 104039 1006501
rect 152917 1006498 152983 1006501
rect 103973 1006496 104236 1006498
rect 103973 1006440 103978 1006496
rect 104034 1006440 104236 1006496
rect 103973 1006438 104236 1006440
rect 152720 1006496 152983 1006498
rect 152720 1006440 152922 1006496
rect 152978 1006440 152983 1006496
rect 152720 1006438 152983 1006440
rect 103973 1006435 104039 1006438
rect 152917 1006435 152983 1006438
rect 307753 1006498 307819 1006501
rect 360193 1006498 360259 1006501
rect 307753 1006496 307924 1006498
rect 307753 1006440 307758 1006496
rect 307814 1006440 307924 1006496
rect 307753 1006438 307924 1006440
rect 359996 1006496 360259 1006498
rect 359996 1006440 360198 1006496
rect 360254 1006440 360259 1006496
rect 359996 1006438 360259 1006440
rect 307753 1006435 307819 1006438
rect 360193 1006435 360259 1006438
rect 505369 1006498 505435 1006501
rect 553117 1006498 553183 1006501
rect 505369 1006496 505632 1006498
rect 505369 1006440 505374 1006496
rect 505430 1006440 505632 1006496
rect 505369 1006438 505632 1006440
rect 552920 1006496 553183 1006498
rect 552920 1006440 553122 1006496
rect 553178 1006440 553183 1006496
rect 552920 1006438 553183 1006440
rect 505369 1006435 505435 1006438
rect 553117 1006435 553183 1006438
rect 100293 1006362 100359 1006365
rect 152089 1006362 152155 1006365
rect 158253 1006362 158319 1006365
rect 210417 1006362 210483 1006365
rect 100293 1006360 100556 1006362
rect 100293 1006304 100298 1006360
rect 100354 1006304 100556 1006360
rect 100293 1006302 100556 1006304
rect 152089 1006360 152352 1006362
rect 152089 1006304 152094 1006360
rect 152150 1006304 152352 1006360
rect 152089 1006302 152352 1006304
rect 158056 1006360 158319 1006362
rect 158056 1006304 158258 1006360
rect 158314 1006304 158319 1006360
rect 158056 1006302 158319 1006304
rect 210220 1006360 210483 1006362
rect 210220 1006304 210422 1006360
rect 210478 1006304 210483 1006360
rect 210220 1006302 210483 1006304
rect 100293 1006299 100359 1006302
rect 152089 1006299 152155 1006302
rect 158253 1006299 158319 1006302
rect 210417 1006299 210483 1006302
rect 256141 1006362 256207 1006365
rect 314653 1006362 314719 1006365
rect 360561 1006362 360627 1006365
rect 425145 1006362 425211 1006365
rect 502149 1006362 502215 1006365
rect 556797 1006362 556863 1006365
rect 256141 1006360 256404 1006362
rect 256141 1006304 256146 1006360
rect 256202 1006304 256404 1006360
rect 256141 1006302 256404 1006304
rect 314653 1006360 314916 1006362
rect 314653 1006304 314658 1006360
rect 314714 1006304 314916 1006360
rect 314653 1006302 314916 1006304
rect 360561 1006360 360824 1006362
rect 360561 1006304 360566 1006360
rect 360622 1006304 360824 1006360
rect 360561 1006302 360824 1006304
rect 424948 1006360 425211 1006362
rect 424948 1006304 425150 1006360
rect 425206 1006304 425211 1006360
rect 424948 1006302 425211 1006304
rect 501952 1006360 502215 1006362
rect 501952 1006304 502154 1006360
rect 502210 1006304 502215 1006360
rect 501952 1006302 502215 1006304
rect 556600 1006360 556863 1006362
rect 556600 1006304 556802 1006360
rect 556858 1006304 556863 1006360
rect 556600 1006302 556863 1006304
rect 256141 1006299 256207 1006302
rect 314653 1006299 314719 1006302
rect 360561 1006299 360627 1006302
rect 425145 1006299 425211 1006302
rect 502149 1006299 502215 1006302
rect 556797 1006299 556863 1006302
rect 101949 1006226 102015 1006229
rect 106825 1006226 106891 1006229
rect 159449 1006226 159515 1006229
rect 160277 1006226 160343 1006229
rect 101949 1006224 102212 1006226
rect 101949 1006168 101954 1006224
rect 102010 1006168 102212 1006224
rect 101949 1006166 102212 1006168
rect 106628 1006224 106891 1006226
rect 106628 1006168 106830 1006224
rect 106886 1006168 106891 1006224
rect 106628 1006166 106891 1006168
rect 159252 1006224 159515 1006226
rect 159252 1006168 159454 1006224
rect 159510 1006168 159515 1006224
rect 159252 1006166 159515 1006168
rect 160080 1006224 160343 1006226
rect 160080 1006168 160282 1006224
rect 160338 1006168 160343 1006224
rect 160080 1006166 160343 1006168
rect 101949 1006163 102015 1006166
rect 106825 1006163 106891 1006166
rect 159449 1006163 159515 1006166
rect 160277 1006163 160343 1006166
rect 208393 1006226 208459 1006229
rect 252461 1006226 252527 1006229
rect 262673 1006226 262739 1006229
rect 208393 1006224 208656 1006226
rect 208393 1006168 208398 1006224
rect 208454 1006168 208656 1006224
rect 208393 1006166 208656 1006168
rect 252461 1006224 252724 1006226
rect 252461 1006168 252466 1006224
rect 252522 1006196 252724 1006224
rect 262476 1006224 262739 1006226
rect 252522 1006168 252754 1006196
rect 252461 1006166 252754 1006168
rect 262476 1006168 262678 1006224
rect 262734 1006168 262739 1006224
rect 262476 1006166 262739 1006168
rect 208393 1006163 208459 1006166
rect 252461 1006163 252527 1006166
rect 98269 1006090 98335 1006093
rect 103973 1006090 104039 1006093
rect 107653 1006090 107719 1006093
rect 98269 1006088 98900 1006090
rect 98269 1006032 98274 1006088
rect 98330 1006032 98900 1006088
rect 98269 1006030 98900 1006032
rect 103776 1006088 104039 1006090
rect 103776 1006032 103978 1006088
rect 104034 1006032 104039 1006088
rect 103776 1006030 104039 1006032
rect 107456 1006088 107719 1006090
rect 107456 1006032 107658 1006088
rect 107714 1006032 107719 1006088
rect 107456 1006030 107719 1006032
rect 98269 1006027 98335 1006030
rect 103973 1006027 104039 1006030
rect 107653 1006027 107719 1006030
rect 146937 1006090 147003 1006093
rect 148869 1006090 148935 1006093
rect 150065 1006090 150131 1006093
rect 155769 1006090 155835 1006093
rect 158621 1006090 158687 1006093
rect 201033 1006090 201099 1006093
rect 252694 1006090 252754 1006166
rect 262673 1006163 262739 1006166
rect 306097 1006226 306163 1006229
rect 423489 1006226 423555 1006229
rect 508221 1006226 508287 1006229
rect 557165 1006226 557231 1006229
rect 306097 1006224 306360 1006226
rect 306097 1006168 306102 1006224
rect 306158 1006168 306360 1006224
rect 306097 1006166 306360 1006168
rect 423489 1006224 423752 1006226
rect 423489 1006168 423494 1006224
rect 423550 1006168 423752 1006224
rect 423489 1006166 423752 1006168
rect 508221 1006224 508484 1006226
rect 508221 1006168 508226 1006224
rect 508282 1006168 508484 1006224
rect 508221 1006166 508484 1006168
rect 557060 1006224 557231 1006226
rect 557060 1006168 557170 1006224
rect 557226 1006168 557231 1006224
rect 557060 1006166 557231 1006168
rect 306097 1006163 306163 1006166
rect 423489 1006163 423555 1006166
rect 508221 1006163 508287 1006166
rect 557165 1006163 557231 1006166
rect 254117 1006090 254183 1006093
rect 261845 1006090 261911 1006093
rect 146937 1006088 148935 1006090
rect 146937 1006032 146942 1006088
rect 146998 1006032 148874 1006088
rect 148930 1006032 148935 1006088
rect 146937 1006030 148935 1006032
rect 149868 1006088 150328 1006090
rect 149868 1006032 150070 1006088
rect 150126 1006032 150328 1006088
rect 149868 1006030 150328 1006032
rect 155769 1006088 156032 1006090
rect 155769 1006032 155774 1006088
rect 155830 1006032 156032 1006088
rect 155769 1006030 156032 1006032
rect 158621 1006088 158884 1006090
rect 158621 1006032 158626 1006088
rect 158682 1006032 158884 1006088
rect 158621 1006030 158884 1006032
rect 201033 1006088 201756 1006090
rect 201033 1006032 201038 1006088
rect 201094 1006032 201756 1006088
rect 252694 1006060 253092 1006090
rect 201033 1006030 201756 1006032
rect 252724 1006030 253092 1006060
rect 254117 1006088 254380 1006090
rect 254117 1006032 254122 1006088
rect 254178 1006032 254380 1006088
rect 254117 1006030 254380 1006032
rect 261648 1006088 261911 1006090
rect 261648 1006032 261850 1006088
rect 261906 1006032 261911 1006088
rect 261648 1006030 261911 1006032
rect 146937 1006027 147003 1006030
rect 148869 1006027 148935 1006030
rect 150065 1006027 150131 1006030
rect 155769 1006027 155835 1006030
rect 158621 1006027 158687 1006030
rect 201033 1006027 201099 1006030
rect 254117 1006027 254183 1006030
rect 261845 1006027 261911 1006030
rect 304073 1006090 304139 1006093
rect 311801 1006090 311867 1006093
rect 314653 1006090 314719 1006093
rect 354857 1006090 354923 1006093
rect 355685 1006090 355751 1006093
rect 361389 1006090 361455 1006093
rect 365069 1006090 365135 1006093
rect 422661 1006090 422727 1006093
rect 430021 1006090 430087 1006093
rect 304073 1006088 304704 1006090
rect 304073 1006032 304078 1006088
rect 304134 1006032 304704 1006088
rect 304073 1006030 304704 1006032
rect 311801 1006088 312064 1006090
rect 311801 1006032 311806 1006088
rect 311862 1006032 312064 1006088
rect 311801 1006030 312064 1006032
rect 314548 1006088 314719 1006090
rect 314548 1006032 314658 1006088
rect 314714 1006032 314719 1006088
rect 314548 1006030 314719 1006032
rect 354660 1006088 355120 1006090
rect 354660 1006032 354862 1006088
rect 354918 1006032 355120 1006088
rect 354660 1006030 355120 1006032
rect 355685 1006088 355948 1006090
rect 355685 1006032 355690 1006088
rect 355746 1006032 355948 1006088
rect 355685 1006030 355948 1006032
rect 361389 1006088 361652 1006090
rect 361389 1006032 361394 1006088
rect 361450 1006032 361652 1006088
rect 361389 1006030 361652 1006032
rect 364872 1006088 365135 1006090
rect 364872 1006032 365074 1006088
rect 365130 1006032 365135 1006088
rect 364872 1006030 365135 1006032
rect 422096 1006088 422727 1006090
rect 422096 1006032 422666 1006088
rect 422722 1006032 422727 1006088
rect 422096 1006030 422727 1006032
rect 429824 1006088 430087 1006090
rect 429824 1006032 430026 1006088
rect 430082 1006032 430087 1006088
rect 429824 1006030 430087 1006032
rect 304073 1006027 304139 1006030
rect 311801 1006027 311867 1006030
rect 314653 1006027 314719 1006030
rect 354857 1006027 354923 1006030
rect 355685 1006027 355751 1006030
rect 361389 1006027 361455 1006030
rect 365069 1006027 365135 1006030
rect 422661 1006027 422727 1006030
rect 430021 1006027 430087 1006030
rect 498837 1006090 498903 1006093
rect 501321 1006090 501387 1006093
rect 498837 1006088 499468 1006090
rect 498837 1006032 498842 1006088
rect 498898 1006032 499468 1006088
rect 498837 1006030 499468 1006032
rect 501124 1006088 501387 1006090
rect 501124 1006032 501326 1006088
rect 501382 1006032 501387 1006088
rect 501124 1006030 501387 1006032
rect 498837 1006027 498903 1006030
rect 501321 1006027 501387 1006030
rect 509049 1006090 509115 1006093
rect 509049 1006088 509312 1006090
rect 509049 1006032 509054 1006088
rect 509110 1006032 509312 1006088
rect 509049 1006030 509312 1006032
rect 509049 1006027 509115 1006030
rect 432045 1005818 432111 1005821
rect 431940 1005816 432111 1005818
rect 431940 1005760 432050 1005816
rect 432106 1005760 432111 1005816
rect 431940 1005758 432111 1005760
rect 432045 1005755 432111 1005758
rect 423489 1005682 423555 1005685
rect 423292 1005680 423555 1005682
rect 423292 1005624 423494 1005680
rect 423550 1005624 423555 1005680
rect 423292 1005622 423555 1005624
rect 423489 1005619 423555 1005622
rect 560845 1005682 560911 1005685
rect 560845 1005680 561108 1005682
rect 560845 1005624 560850 1005680
rect 560906 1005624 561108 1005680
rect 560845 1005622 561108 1005624
rect 560845 1005619 560911 1005622
rect 428365 1005546 428431 1005549
rect 428260 1005544 428431 1005546
rect 428260 1005488 428370 1005544
rect 428426 1005488 428431 1005544
rect 428260 1005486 428431 1005488
rect 428365 1005483 428431 1005486
rect 555141 1005546 555207 1005549
rect 555141 1005544 555404 1005546
rect 555141 1005488 555146 1005544
rect 555202 1005488 555404 1005544
rect 555141 1005486 555404 1005488
rect 555141 1005483 555207 1005486
rect 152917 1005410 152983 1005413
rect 427169 1005410 427235 1005413
rect 553945 1005410 554011 1005413
rect 152917 1005408 153180 1005410
rect 152917 1005352 152922 1005408
rect 152978 1005352 153180 1005408
rect 152917 1005350 153180 1005352
rect 426972 1005408 427235 1005410
rect 426972 1005352 427174 1005408
rect 427230 1005352 427235 1005408
rect 426972 1005350 427235 1005352
rect 553748 1005408 554011 1005410
rect 553748 1005352 553950 1005408
rect 554006 1005352 554011 1005408
rect 553748 1005350 554011 1005352
rect 152917 1005347 152983 1005350
rect 427169 1005347 427235 1005350
rect 553945 1005347 554011 1005350
rect 202689 1005274 202755 1005277
rect 263041 1005274 263107 1005277
rect 360561 1005274 360627 1005277
rect 430849 1005274 430915 1005277
rect 507025 1005274 507091 1005277
rect 202492 1005272 202755 1005274
rect 202492 1005216 202694 1005272
rect 202750 1005216 202755 1005272
rect 202492 1005214 202755 1005216
rect 262844 1005272 263107 1005274
rect 262844 1005216 263046 1005272
rect 263102 1005216 263107 1005272
rect 262844 1005214 263107 1005216
rect 360364 1005272 360627 1005274
rect 360364 1005216 360566 1005272
rect 360622 1005216 360627 1005272
rect 360364 1005214 360627 1005216
rect 430652 1005272 430915 1005274
rect 430652 1005216 430854 1005272
rect 430910 1005216 430915 1005272
rect 430652 1005214 430915 1005216
rect 506828 1005272 507091 1005274
rect 506828 1005216 507030 1005272
rect 507086 1005216 507091 1005272
rect 506828 1005214 507091 1005216
rect 202689 1005211 202755 1005214
rect 263041 1005211 263107 1005214
rect 360561 1005211 360627 1005214
rect 430849 1005211 430915 1005214
rect 507025 1005211 507091 1005214
rect 552289 1005274 552355 1005277
rect 552289 1005272 552552 1005274
rect 552289 1005216 552294 1005272
rect 552350 1005216 552552 1005272
rect 552289 1005214 552552 1005216
rect 552289 1005211 552355 1005214
rect 209221 1005138 209287 1005141
rect 363413 1005138 363479 1005141
rect 209221 1005136 209484 1005138
rect 209221 1005080 209226 1005136
rect 209282 1005080 209484 1005136
rect 209221 1005078 209484 1005080
rect 363308 1005136 363479 1005138
rect 363308 1005080 363418 1005136
rect 363474 1005080 363479 1005136
rect 363308 1005078 363479 1005080
rect 209221 1005075 209287 1005078
rect 363413 1005075 363479 1005078
rect 432045 1005138 432111 1005141
rect 508221 1005138 508287 1005141
rect 432045 1005136 432308 1005138
rect 432045 1005080 432050 1005136
rect 432106 1005080 432308 1005136
rect 432045 1005078 432308 1005080
rect 508116 1005136 508287 1005138
rect 508116 1005080 508226 1005136
rect 508282 1005080 508287 1005136
rect 508116 1005078 508287 1005080
rect 432045 1005075 432111 1005078
rect 508221 1005075 508287 1005078
rect 153745 1005002 153811 1005005
rect 160645 1005002 160711 1005005
rect 207565 1005002 207631 1005005
rect 153745 1005000 153916 1005002
rect 153745 1004944 153750 1005000
rect 153806 1004944 153916 1005000
rect 153745 1004942 153916 1004944
rect 160645 1005000 160908 1005002
rect 160645 1004944 160650 1005000
rect 160706 1004944 160908 1005000
rect 160645 1004942 160908 1004944
rect 207460 1005000 207631 1005002
rect 207460 1004944 207570 1005000
rect 207626 1004944 207631 1005000
rect 207460 1004942 207631 1004944
rect 153745 1004939 153811 1004942
rect 160645 1004939 160711 1004942
rect 207565 1004939 207631 1004942
rect 365069 1005002 365135 1005005
rect 429193 1005002 429259 1005005
rect 507853 1005002 507919 1005005
rect 365069 1005000 365332 1005002
rect 365069 1004944 365074 1005000
rect 365130 1004944 365332 1005000
rect 365069 1004942 365332 1004944
rect 429193 1005000 429456 1005002
rect 429193 1004944 429198 1005000
rect 429254 1004944 429456 1005000
rect 429193 1004942 429456 1004944
rect 507656 1005000 507919 1005002
rect 507656 1004944 507858 1005000
rect 507914 1004944 507919 1005000
rect 507656 1004942 507919 1004944
rect 365069 1004939 365135 1004942
rect 429193 1004939 429259 1004942
rect 507853 1004939 507919 1004942
rect 154113 1004866 154179 1004869
rect 159449 1004866 159515 1004869
rect 313825 1004866 313891 1004869
rect 355685 1004866 355751 1004869
rect 362585 1004866 362651 1004869
rect 431677 1004866 431743 1004869
rect 154113 1004864 154376 1004866
rect 154113 1004808 154118 1004864
rect 154174 1004808 154376 1004864
rect 154113 1004806 154376 1004808
rect 159449 1004864 159712 1004866
rect 159449 1004808 159454 1004864
rect 159510 1004808 159712 1004864
rect 159449 1004806 159712 1004808
rect 313628 1004864 313891 1004866
rect 313628 1004808 313830 1004864
rect 313886 1004808 313891 1004864
rect 313628 1004806 313891 1004808
rect 355488 1004864 355751 1004866
rect 355488 1004808 355690 1004864
rect 355746 1004808 355751 1004864
rect 355488 1004806 355751 1004808
rect 362388 1004864 362651 1004866
rect 362388 1004808 362590 1004864
rect 362646 1004808 362651 1004864
rect 362388 1004806 362651 1004808
rect 431480 1004864 431743 1004866
rect 431480 1004808 431682 1004864
rect 431738 1004808 431743 1004864
rect 431480 1004806 431743 1004808
rect 154113 1004803 154179 1004806
rect 159449 1004803 159515 1004806
rect 313825 1004803 313891 1004806
rect 355685 1004803 355751 1004806
rect 362585 1004803 362651 1004806
rect 431677 1004803 431743 1004806
rect 499665 1004866 499731 1004869
rect 507393 1004866 507459 1004869
rect 555969 1004866 556035 1004869
rect 499665 1004864 499928 1004866
rect 499665 1004808 499670 1004864
rect 499726 1004808 499928 1004864
rect 499665 1004806 499928 1004808
rect 507196 1004864 507459 1004866
rect 507196 1004808 507398 1004864
rect 507454 1004808 507459 1004864
rect 507196 1004806 507459 1004808
rect 555772 1004864 556035 1004866
rect 555772 1004808 555974 1004864
rect 556030 1004808 556035 1004864
rect 555772 1004806 556035 1004808
rect 499665 1004803 499731 1004806
rect 507393 1004803 507459 1004806
rect 555969 1004803 556035 1004806
rect 108481 1004730 108547 1004733
rect 151721 1004730 151787 1004733
rect 160645 1004730 160711 1004733
rect 209221 1004730 209287 1004733
rect 212533 1004730 212599 1004733
rect 108481 1004728 108652 1004730
rect 108481 1004672 108486 1004728
rect 108542 1004672 108652 1004728
rect 108481 1004670 108652 1004672
rect 151721 1004728 151892 1004730
rect 151721 1004672 151726 1004728
rect 151782 1004672 151892 1004728
rect 151721 1004670 151892 1004672
rect 160540 1004728 160711 1004730
rect 160540 1004672 160650 1004728
rect 160706 1004672 160711 1004728
rect 160540 1004670 160711 1004672
rect 209024 1004728 209287 1004730
rect 209024 1004672 209226 1004728
rect 209282 1004672 209287 1004728
rect 209024 1004670 209287 1004672
rect 212336 1004728 212599 1004730
rect 212336 1004672 212538 1004728
rect 212594 1004672 212599 1004728
rect 212336 1004670 212599 1004672
rect 108481 1004667 108547 1004670
rect 151721 1004667 151787 1004670
rect 160645 1004667 160711 1004670
rect 209221 1004667 209287 1004670
rect 212533 1004667 212599 1004670
rect 256509 1004730 256575 1004733
rect 315481 1004730 315547 1004733
rect 364241 1004730 364307 1004733
rect 256509 1004728 256772 1004730
rect 256509 1004672 256514 1004728
rect 256570 1004672 256772 1004728
rect 256509 1004670 256772 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 364044 1004728 364307 1004730
rect 364044 1004672 364246 1004728
rect 364302 1004672 364307 1004728
rect 364044 1004670 364307 1004672
rect 256509 1004667 256575 1004670
rect 315481 1004667 315547 1004670
rect 364241 1004667 364307 1004670
rect 422661 1004730 422727 1004733
rect 430021 1004730 430087 1004733
rect 500493 1004730 500559 1004733
rect 509049 1004730 509115 1004733
rect 557625 1004730 557691 1004733
rect 422661 1004728 422924 1004730
rect 422661 1004672 422666 1004728
rect 422722 1004672 422924 1004728
rect 422661 1004670 422924 1004672
rect 430021 1004728 430284 1004730
rect 430021 1004672 430026 1004728
rect 430082 1004672 430284 1004728
rect 430021 1004670 430284 1004672
rect 500296 1004728 500559 1004730
rect 500296 1004672 500498 1004728
rect 500554 1004672 500559 1004728
rect 500296 1004670 500559 1004672
rect 508852 1004728 509115 1004730
rect 508852 1004672 509054 1004728
rect 509110 1004672 509115 1004728
rect 508852 1004670 509115 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 422661 1004667 422727 1004670
rect 430021 1004667 430087 1004670
rect 500493 1004667 500559 1004670
rect 509049 1004667 509115 1004670
rect 557625 1004667 557691 1004670
rect 504541 1004458 504607 1004461
rect 504436 1004456 504607 1004458
rect 504436 1004400 504546 1004456
rect 504602 1004400 504607 1004456
rect 504436 1004398 504607 1004400
rect 504541 1004395 504607 1004398
rect 356513 1003914 356579 1003917
rect 356316 1003912 356579 1003914
rect 356316 1003856 356518 1003912
rect 356574 1003856 356579 1003912
rect 356316 1003854 356579 1003856
rect 356513 1003851 356579 1003854
rect 101949 1002826 102015 1002829
rect 255313 1002826 255379 1002829
rect 101752 1002824 102015 1002826
rect 101752 1002768 101954 1002824
rect 102010 1002768 102015 1002824
rect 101752 1002766 102015 1002768
rect 255116 1002824 255379 1002826
rect 255116 1002768 255318 1002824
rect 255374 1002768 255379 1002824
rect 255116 1002766 255379 1002768
rect 101949 1002763 102015 1002766
rect 255313 1002763 255379 1002766
rect 100293 1002690 100359 1002693
rect 157425 1002690 157491 1002693
rect 424685 1002690 424751 1002693
rect 100096 1002688 100359 1002690
rect 100096 1002632 100298 1002688
rect 100354 1002632 100359 1002688
rect 100096 1002630 100359 1002632
rect 157228 1002688 157491 1002690
rect 157228 1002632 157430 1002688
rect 157486 1002632 157491 1002688
rect 157228 1002630 157491 1002632
rect 424580 1002688 424751 1002690
rect 424580 1002632 424690 1002688
rect 424746 1002632 424751 1002688
rect 424580 1002630 424751 1002632
rect 100293 1002627 100359 1002630
rect 157425 1002627 157491 1002630
rect 424685 1002627 424751 1002630
rect 101121 1002554 101187 1002557
rect 105997 1002554 106063 1002557
rect 158621 1002554 158687 1002557
rect 100924 1002552 101187 1002554
rect 100924 1002496 101126 1002552
rect 101182 1002496 101187 1002552
rect 100924 1002494 101187 1002496
rect 105892 1002552 106063 1002554
rect 105892 1002496 106002 1002552
rect 106058 1002496 106063 1002552
rect 105892 1002494 106063 1002496
rect 158516 1002552 158687 1002554
rect 158516 1002496 158626 1002552
rect 158682 1002496 158687 1002552
rect 158516 1002494 158687 1002496
rect 101121 1002491 101187 1002494
rect 105997 1002491 106063 1002494
rect 158621 1002491 158687 1002494
rect 255313 1002554 255379 1002557
rect 261017 1002554 261083 1002557
rect 426341 1002554 426407 1002557
rect 501689 1002554 501755 1002557
rect 255313 1002552 255576 1002554
rect 255313 1002496 255318 1002552
rect 255374 1002496 255576 1002552
rect 255313 1002494 255576 1002496
rect 260820 1002552 261083 1002554
rect 260820 1002496 261022 1002552
rect 261078 1002496 261083 1002552
rect 260820 1002494 261083 1002496
rect 426144 1002552 426407 1002554
rect 426144 1002496 426346 1002552
rect 426402 1002496 426407 1002552
rect 426144 1002494 426407 1002496
rect 501492 1002552 501755 1002554
rect 501492 1002496 501694 1002552
rect 501750 1002496 501755 1002552
rect 501492 1002494 501755 1002496
rect 255313 1002491 255379 1002494
rect 261017 1002491 261083 1002494
rect 426341 1002491 426407 1002494
rect 501689 1002491 501755 1002494
rect 558821 1002554 558887 1002557
rect 558821 1002552 559084 1002554
rect 558821 1002496 558826 1002552
rect 558882 1002496 559084 1002552
rect 558821 1002494 559084 1002496
rect 558821 1002491 558887 1002494
rect 99097 1002418 99163 1002421
rect 105629 1002418 105695 1002421
rect 108021 1002418 108087 1002421
rect 99097 1002416 99268 1002418
rect 99097 1002360 99102 1002416
rect 99158 1002360 99268 1002416
rect 99097 1002358 99268 1002360
rect 105432 1002416 105695 1002418
rect 105432 1002360 105634 1002416
rect 105690 1002360 105695 1002416
rect 105432 1002358 105695 1002360
rect 107916 1002416 108087 1002418
rect 107916 1002360 108026 1002416
rect 108082 1002360 108087 1002416
rect 107916 1002358 108087 1002360
rect 99097 1002355 99163 1002358
rect 105629 1002355 105695 1002358
rect 108021 1002355 108087 1002358
rect 150893 1002418 150959 1002421
rect 156597 1002418 156663 1002421
rect 211245 1002418 211311 1002421
rect 502149 1002418 502215 1002421
rect 557993 1002418 558059 1002421
rect 560477 1002418 560543 1002421
rect 150893 1002416 151156 1002418
rect 150893 1002360 150898 1002416
rect 150954 1002360 151156 1002416
rect 150893 1002358 151156 1002360
rect 156597 1002416 156860 1002418
rect 156597 1002360 156602 1002416
rect 156658 1002360 156860 1002416
rect 156597 1002358 156860 1002360
rect 211245 1002416 211508 1002418
rect 211245 1002360 211250 1002416
rect 211306 1002360 211508 1002416
rect 211245 1002358 211508 1002360
rect 502149 1002416 502412 1002418
rect 502149 1002360 502154 1002416
rect 502210 1002360 502412 1002416
rect 502149 1002358 502412 1002360
rect 557796 1002416 558059 1002418
rect 557796 1002360 557998 1002416
rect 558054 1002360 558059 1002416
rect 557796 1002358 558059 1002360
rect 560280 1002416 560543 1002418
rect 560280 1002360 560482 1002416
rect 560538 1002360 560543 1002416
rect 560280 1002358 560543 1002360
rect 150893 1002355 150959 1002358
rect 156597 1002355 156663 1002358
rect 211245 1002355 211311 1002358
rect 502149 1002355 502215 1002358
rect 557993 1002355 558059 1002358
rect 560477 1002355 560543 1002358
rect 101121 1002282 101187 1002285
rect 104801 1002282 104867 1002285
rect 108481 1002282 108547 1002285
rect 151721 1002282 151787 1002285
rect 155769 1002282 155835 1002285
rect 206369 1002282 206435 1002285
rect 210049 1002282 210115 1002285
rect 101121 1002280 101292 1002282
rect 101121 1002224 101126 1002280
rect 101182 1002224 101292 1002280
rect 101121 1002222 101292 1002224
rect 104604 1002280 104867 1002282
rect 104604 1002224 104806 1002280
rect 104862 1002224 104867 1002280
rect 104604 1002222 104867 1002224
rect 108284 1002280 108547 1002282
rect 108284 1002224 108486 1002280
rect 108542 1002224 108547 1002280
rect 108284 1002222 108547 1002224
rect 151524 1002280 151787 1002282
rect 151524 1002224 151726 1002280
rect 151782 1002224 151787 1002280
rect 151524 1002222 151787 1002224
rect 155572 1002280 155835 1002282
rect 155572 1002224 155774 1002280
rect 155830 1002224 155835 1002280
rect 155572 1002222 155835 1002224
rect 206172 1002280 206435 1002282
rect 206172 1002224 206374 1002280
rect 206430 1002224 206435 1002280
rect 206172 1002222 206435 1002224
rect 209852 1002280 210115 1002282
rect 209852 1002224 210054 1002280
rect 210110 1002224 210115 1002280
rect 209852 1002222 210115 1002224
rect 101121 1002219 101187 1002222
rect 104801 1002219 104867 1002222
rect 108481 1002219 108547 1002222
rect 151721 1002219 151787 1002222
rect 155769 1002219 155835 1002222
rect 206369 1002219 206435 1002222
rect 210049 1002219 210115 1002222
rect 254485 1002282 254551 1002285
rect 298093 1002282 298159 1002285
rect 302141 1002282 302207 1002285
rect 427997 1002282 428063 1002285
rect 254485 1002280 254748 1002282
rect 254485 1002224 254490 1002280
rect 254546 1002224 254748 1002280
rect 254485 1002222 254748 1002224
rect 298093 1002280 302207 1002282
rect 298093 1002224 298098 1002280
rect 298154 1002224 302146 1002280
rect 302202 1002224 302207 1002280
rect 298093 1002222 302207 1002224
rect 427800 1002280 428063 1002282
rect 427800 1002224 428002 1002280
rect 428058 1002224 428063 1002280
rect 427800 1002222 428063 1002224
rect 254485 1002219 254551 1002222
rect 298093 1002219 298159 1002222
rect 302141 1002219 302207 1002222
rect 427997 1002219 428063 1002222
rect 500493 1002282 500559 1002285
rect 509877 1002282 509943 1002285
rect 500493 1002280 500756 1002282
rect 500493 1002224 500498 1002280
rect 500554 1002224 500756 1002280
rect 500493 1002222 500756 1002224
rect 509680 1002280 509943 1002282
rect 509680 1002224 509882 1002280
rect 509938 1002224 509943 1002280
rect 509680 1002222 509943 1002224
rect 500493 1002219 500559 1002222
rect 509877 1002219 509943 1002222
rect 554313 1002282 554379 1002285
rect 560017 1002282 560083 1002285
rect 554313 1002280 554576 1002282
rect 554313 1002224 554318 1002280
rect 554374 1002224 554576 1002280
rect 554313 1002222 554576 1002224
rect 559820 1002280 560083 1002282
rect 559820 1002224 560022 1002280
rect 560078 1002224 560083 1002280
rect 559820 1002222 560083 1002224
rect 554313 1002219 554379 1002222
rect 560017 1002219 560083 1002222
rect 99465 1002146 99531 1002149
rect 103145 1002146 103211 1002149
rect 106825 1002146 106891 1002149
rect 109677 1002146 109743 1002149
rect 150893 1002146 150959 1002149
rect 156597 1002146 156663 1002149
rect 99465 1002144 99728 1002146
rect 99465 1002088 99470 1002144
rect 99526 1002088 99728 1002144
rect 99465 1002086 99728 1002088
rect 103145 1002144 103408 1002146
rect 103145 1002088 103150 1002144
rect 103206 1002088 103408 1002144
rect 103145 1002086 103408 1002088
rect 106825 1002144 107088 1002146
rect 106825 1002088 106830 1002144
rect 106886 1002088 107088 1002144
rect 106825 1002086 107088 1002088
rect 109480 1002144 109743 1002146
rect 109480 1002088 109682 1002144
rect 109738 1002088 109743 1002144
rect 109480 1002086 109743 1002088
rect 150696 1002144 150959 1002146
rect 150696 1002088 150898 1002144
rect 150954 1002088 150959 1002144
rect 150696 1002086 150959 1002088
rect 156400 1002144 156663 1002146
rect 156400 1002088 156602 1002144
rect 156658 1002088 156663 1002144
rect 156400 1002086 156663 1002088
rect 99465 1002083 99531 1002086
rect 103145 1002083 103211 1002086
rect 106825 1002083 106891 1002086
rect 109677 1002083 109743 1002086
rect 150893 1002083 150959 1002086
rect 156597 1002083 156663 1002086
rect 205541 1002146 205607 1002149
rect 211245 1002146 211311 1002149
rect 256141 1002146 256207 1002149
rect 263501 1002146 263567 1002149
rect 205541 1002144 205804 1002146
rect 205541 1002088 205546 1002144
rect 205602 1002088 205804 1002144
rect 205541 1002086 205804 1002088
rect 211140 1002144 211311 1002146
rect 211140 1002088 211250 1002144
rect 211306 1002088 211311 1002144
rect 211140 1002086 211311 1002088
rect 255944 1002144 256207 1002146
rect 255944 1002088 256146 1002144
rect 256202 1002088 256207 1002144
rect 255944 1002086 256207 1002088
rect 263304 1002144 263567 1002146
rect 263304 1002088 263506 1002144
rect 263562 1002088 263567 1002144
rect 263304 1002086 263567 1002088
rect 205541 1002083 205607 1002086
rect 211245 1002083 211311 1002086
rect 256141 1002083 256207 1002086
rect 263501 1002083 263567 1002086
rect 310973 1002146 311039 1002149
rect 358537 1002146 358603 1002149
rect 359733 1002146 359799 1002149
rect 310973 1002144 311236 1002146
rect 310973 1002088 310978 1002144
rect 311034 1002088 311236 1002144
rect 310973 1002086 311236 1002088
rect 358537 1002144 358800 1002146
rect 358537 1002088 358542 1002144
rect 358598 1002088 358800 1002144
rect 358537 1002086 358800 1002088
rect 359628 1002144 359799 1002146
rect 359628 1002088 359738 1002144
rect 359794 1002088 359799 1002144
rect 359628 1002086 359799 1002088
rect 310973 1002083 311039 1002086
rect 358537 1002083 358603 1002086
rect 359733 1002083 359799 1002086
rect 425145 1002146 425211 1002149
rect 428365 1002146 428431 1002149
rect 433333 1002146 433399 1002149
rect 425145 1002144 425316 1002146
rect 425145 1002088 425150 1002144
rect 425206 1002088 425316 1002144
rect 425145 1002086 425316 1002088
rect 428365 1002144 428628 1002146
rect 428365 1002088 428370 1002144
rect 428426 1002088 428628 1002144
rect 428365 1002086 428628 1002088
rect 433136 1002144 433399 1002146
rect 433136 1002088 433338 1002144
rect 433394 1002088 433399 1002144
rect 433136 1002086 433399 1002088
rect 425145 1002083 425211 1002086
rect 428365 1002083 428431 1002086
rect 433333 1002083 433399 1002086
rect 502517 1002146 502583 1002149
rect 510337 1002146 510403 1002149
rect 555141 1002146 555207 1002149
rect 502517 1002144 502780 1002146
rect 502517 1002088 502522 1002144
rect 502578 1002088 502780 1002144
rect 502517 1002086 502780 1002088
rect 510140 1002144 510403 1002146
rect 510140 1002088 510342 1002144
rect 510398 1002088 510403 1002144
rect 510140 1002086 510403 1002088
rect 555036 1002144 555207 1002146
rect 555036 1002088 555146 1002144
rect 555202 1002088 555207 1002144
rect 555036 1002086 555207 1002088
rect 502517 1002083 502583 1002086
rect 510337 1002083 510403 1002086
rect 555141 1002083 555207 1002086
rect 557993 1002146 558059 1002149
rect 560845 1002146 560911 1002149
rect 557993 1002144 558256 1002146
rect 557993 1002088 557998 1002144
rect 558054 1002088 558256 1002144
rect 557993 1002086 558256 1002088
rect 560740 1002144 560911 1002146
rect 560740 1002088 560850 1002144
rect 560906 1002088 560911 1002144
rect 560740 1002086 560911 1002088
rect 557993 1002083 558059 1002086
rect 560845 1002083 560911 1002086
rect 98269 1002010 98335 1002013
rect 98072 1002008 98335 1002010
rect 98072 1001952 98274 1002008
rect 98330 1001952 98335 1002008
rect 98072 1001950 98335 1001952
rect 98269 1001947 98335 1001950
rect 102317 1002010 102383 1002013
rect 104801 1002010 104867 1002013
rect 105997 1002010 106063 1002013
rect 108849 1002010 108915 1002013
rect 149237 1002010 149303 1002013
rect 154573 1002010 154639 1002013
rect 154941 1002010 155007 1002013
rect 157793 1002010 157859 1002013
rect 102317 1002008 102580 1002010
rect 102317 1001952 102322 1002008
rect 102378 1001952 102580 1002008
rect 102317 1001950 102580 1001952
rect 104801 1002008 104972 1002010
rect 104801 1001952 104806 1002008
rect 104862 1001952 104972 1002008
rect 104801 1001950 104972 1001952
rect 105997 1002008 106260 1002010
rect 105997 1001952 106002 1002008
rect 106058 1001952 106260 1002008
rect 105997 1001950 106260 1001952
rect 108849 1002008 109112 1002010
rect 108849 1001952 108854 1002008
rect 108910 1001952 109112 1002008
rect 108849 1001950 109112 1001952
rect 149237 1002008 149500 1002010
rect 149237 1001952 149242 1002008
rect 149298 1001952 149500 1002008
rect 149237 1001950 149500 1001952
rect 154573 1002008 154836 1002010
rect 154573 1001952 154578 1002008
rect 154634 1001952 154836 1002008
rect 154573 1001950 154836 1001952
rect 154941 1002008 155204 1002010
rect 154941 1001952 154946 1002008
rect 155002 1001952 155204 1002008
rect 154941 1001950 155204 1001952
rect 157596 1002008 157859 1002010
rect 157596 1001952 157798 1002008
rect 157854 1001952 157859 1002008
rect 157596 1001950 157859 1001952
rect 102317 1001947 102383 1001950
rect 104801 1001947 104867 1001950
rect 105997 1001947 106063 1001950
rect 108849 1001947 108915 1001950
rect 149237 1001947 149303 1001950
rect 154573 1001947 154639 1001950
rect 154941 1001947 155007 1001950
rect 157793 1001947 157859 1001950
rect 206369 1002010 206435 1002013
rect 206737 1002010 206803 1002013
rect 207565 1002010 207631 1002013
rect 208393 1002010 208459 1002013
rect 206369 1002008 206540 1002010
rect 206369 1001952 206374 1002008
rect 206430 1001952 206540 1002008
rect 206369 1001950 206540 1001952
rect 206737 1002008 207000 1002010
rect 206737 1001952 206742 1002008
rect 206798 1001952 207000 1002008
rect 206737 1001950 207000 1001952
rect 207565 1002008 207828 1002010
rect 207565 1001952 207570 1002008
rect 207626 1001952 207828 1002008
rect 207565 1001950 207828 1001952
rect 208196 1002008 208459 1002010
rect 208196 1001952 208398 1002008
rect 208454 1001952 208459 1002008
rect 208196 1001950 208459 1001952
rect 206369 1001947 206435 1001950
rect 206737 1001947 206803 1001950
rect 207565 1001947 207631 1001950
rect 208393 1001947 208459 1001950
rect 210417 1002010 210483 1002013
rect 212073 1002010 212139 1002013
rect 210417 1002008 210680 1002010
rect 210417 1001952 210422 1002008
rect 210478 1001952 210680 1002008
rect 210417 1001950 210680 1001952
rect 211876 1002008 212139 1002010
rect 211876 1001952 212078 1002008
rect 212134 1001952 212139 1002008
rect 211876 1001950 212139 1001952
rect 210417 1001947 210483 1001950
rect 212073 1001947 212139 1001950
rect 261017 1002010 261083 1002013
rect 263869 1002010 263935 1002013
rect 310145 1002010 310211 1002013
rect 261017 1002008 261280 1002010
rect 261017 1001952 261022 1002008
rect 261078 1001952 261280 1002008
rect 261017 1001950 261280 1001952
rect 263764 1002008 263935 1002010
rect 263764 1001952 263874 1002008
rect 263930 1001952 263935 1002008
rect 263764 1001950 263935 1001952
rect 309948 1002008 310211 1002010
rect 309948 1001952 310150 1002008
rect 310206 1001952 310211 1002008
rect 309948 1001950 310211 1001952
rect 261017 1001947 261083 1001950
rect 263869 1001947 263935 1001950
rect 310145 1001947 310211 1001950
rect 312629 1002010 312695 1002013
rect 354029 1002010 354095 1002013
rect 356513 1002010 356579 1002013
rect 357341 1002010 357407 1002013
rect 359365 1002010 359431 1002013
rect 361389 1002010 361455 1002013
rect 365897 1002010 365963 1002013
rect 312629 1002008 312892 1002010
rect 312629 1001952 312634 1002008
rect 312690 1001952 312892 1002008
rect 312629 1001950 312892 1001952
rect 354029 1002008 354292 1002010
rect 354029 1001952 354034 1002008
rect 354090 1001952 354292 1002008
rect 354029 1001950 354292 1001952
rect 356513 1002008 356684 1002010
rect 356513 1001952 356518 1002008
rect 356574 1001952 356684 1002008
rect 356513 1001950 356684 1001952
rect 357144 1002008 357407 1002010
rect 357144 1001952 357346 1002008
rect 357402 1001952 357407 1002008
rect 357144 1001950 357407 1001952
rect 359168 1002008 359431 1002010
rect 359168 1001952 359370 1002008
rect 359426 1001952 359431 1002008
rect 359168 1001950 359431 1001952
rect 361192 1002008 361455 1002010
rect 361192 1001952 361394 1002008
rect 361450 1001952 361455 1002008
rect 361192 1001950 361455 1001952
rect 365700 1002008 365963 1002010
rect 365700 1001952 365902 1002008
rect 365958 1001952 365963 1002008
rect 365700 1001950 365963 1001952
rect 312629 1001947 312695 1001950
rect 354029 1001947 354095 1001950
rect 356513 1001947 356579 1001950
rect 357341 1001947 357407 1001950
rect 359365 1001947 359431 1001950
rect 361389 1001947 361455 1001950
rect 365897 1001947 365963 1001950
rect 421465 1002010 421531 1002013
rect 424317 1002010 424383 1002013
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 424120 1002008 424383 1002010
rect 424120 1001952 424322 1002008
rect 424378 1001952 424383 1002008
rect 424120 1001950 424383 1001952
rect 421465 1001947 421531 1001950
rect 424317 1001947 424383 1001950
rect 426341 1002010 426407 1002013
rect 432873 1002010 432939 1002013
rect 426341 1002008 426604 1002010
rect 426341 1001952 426346 1002008
rect 426402 1001952 426604 1002008
rect 426341 1001950 426604 1001952
rect 432676 1002008 432939 1002010
rect 432676 1001952 432878 1002008
rect 432934 1001952 432939 1002008
rect 432676 1001950 432939 1001952
rect 426341 1001947 426407 1001950
rect 432873 1001947 432939 1001950
rect 498469 1002010 498535 1002013
rect 503345 1002010 503411 1002013
rect 504173 1002010 504239 1002013
rect 498469 1002008 498732 1002010
rect 498469 1001952 498474 1002008
rect 498530 1001952 498732 1002008
rect 498469 1001950 498732 1001952
rect 503345 1002008 503608 1002010
rect 503345 1001952 503350 1002008
rect 503406 1001952 503608 1002008
rect 503345 1001950 503608 1001952
rect 503976 1002008 504239 1002010
rect 503976 1001952 504178 1002008
rect 504234 1001952 504239 1002008
rect 503976 1001950 504239 1001952
rect 498469 1001947 498535 1001950
rect 503345 1001947 503411 1001950
rect 504173 1001947 504239 1001950
rect 506197 1002010 506263 1002013
rect 554313 1002010 554379 1002013
rect 558821 1002010 558887 1002013
rect 561673 1002010 561739 1002013
rect 506197 1002008 506460 1002010
rect 506197 1001952 506202 1002008
rect 506258 1001952 506460 1002008
rect 506197 1001950 506460 1001952
rect 554116 1002008 554379 1002010
rect 554116 1001952 554318 1002008
rect 554374 1001952 554379 1002008
rect 554116 1001950 554379 1001952
rect 558624 1002008 558887 1002010
rect 558624 1001952 558826 1002008
rect 558882 1001952 558887 1002008
rect 558624 1001950 558887 1001952
rect 561476 1002008 561739 1002010
rect 561476 1001952 561678 1002008
rect 561734 1001952 561739 1002008
rect 561476 1001950 561739 1001952
rect 506197 1001947 506263 1001950
rect 554313 1001947 554379 1001950
rect 558821 1001947 558887 1001950
rect 561673 1001947 561739 1001950
rect 256969 1001194 257035 1001197
rect 256969 1001192 257140 1001194
rect 256969 1001136 256974 1001192
rect 257030 1001136 257140 1001192
rect 256969 1001134 257140 1001136
rect 256969 1001131 257035 1001134
rect 305269 999154 305335 999157
rect 305269 999152 305532 999154
rect 305269 999096 305274 999152
rect 305330 999096 305532 999152
rect 305269 999094 305532 999096
rect 305269 999091 305335 999094
rect 204345 998746 204411 998749
rect 204345 998744 204516 998746
rect 204345 998688 204350 998744
rect 204406 998688 204516 998744
rect 204345 998686 204516 998688
rect 204345 998683 204411 998686
rect 203517 998610 203583 998613
rect 308949 998610 309015 998613
rect 203517 998608 203780 998610
rect 203517 998552 203522 998608
rect 203578 998552 203780 998608
rect 203517 998550 203780 998552
rect 308752 998608 309015 998610
rect 308752 998552 308954 998608
rect 309010 998552 309015 998608
rect 308752 998550 309015 998552
rect 203517 998547 203583 998550
rect 308949 998547 309015 998550
rect 517237 998610 517303 998613
rect 523493 998610 523559 998613
rect 517237 998608 523559 998610
rect 517237 998552 517242 998608
rect 517298 998552 523498 998608
rect 523554 998552 523559 998608
rect 517237 998550 523559 998552
rect 517237 998547 517303 998550
rect 523493 998547 523559 998550
rect 203885 998474 203951 998477
rect 258993 998474 259059 998477
rect 203885 998472 204148 998474
rect 203885 998416 203890 998472
rect 203946 998416 204148 998472
rect 203885 998414 204148 998416
rect 258796 998472 259059 998474
rect 258796 998416 258998 998472
rect 259054 998416 259059 998472
rect 258796 998414 259059 998416
rect 203885 998411 203951 998414
rect 258993 998411 259059 998414
rect 307293 998474 307359 998477
rect 307293 998472 307556 998474
rect 307293 998416 307298 998472
rect 307354 998416 307556 998472
rect 307293 998414 307556 998416
rect 307293 998411 307359 998414
rect 202689 998338 202755 998341
rect 306097 998338 306163 998341
rect 310605 998338 310671 998341
rect 202689 998336 202952 998338
rect 202689 998280 202694 998336
rect 202750 998280 202952 998336
rect 202689 998278 202952 998280
rect 305900 998336 306163 998338
rect 305900 998280 306102 998336
rect 306158 998280 306163 998336
rect 305900 998278 306163 998280
rect 310408 998336 310671 998338
rect 310408 998280 310610 998336
rect 310666 998280 310671 998336
rect 310408 998278 310671 998280
rect 202689 998275 202755 998278
rect 306097 998275 306163 998278
rect 310605 998275 310671 998278
rect 439681 998338 439747 998341
rect 439681 998336 451290 998338
rect 439681 998280 439686 998336
rect 439742 998280 451290 998336
rect 439681 998278 451290 998280
rect 439681 998275 439747 998278
rect 200665 998202 200731 998205
rect 253657 998202 253723 998205
rect 257337 998202 257403 998205
rect 308121 998202 308187 998205
rect 451230 998202 451290 998278
rect 200665 998200 200836 998202
rect 200665 998144 200670 998200
rect 200726 998144 200836 998200
rect 200665 998142 200836 998144
rect 253657 998200 253920 998202
rect 253657 998144 253662 998200
rect 253718 998144 253920 998200
rect 253657 998142 253920 998144
rect 257337 998200 257600 998202
rect 257337 998144 257342 998200
rect 257398 998144 257600 998200
rect 257337 998142 257600 998144
rect 308121 998200 308384 998202
rect 308121 998144 308126 998200
rect 308182 998144 308384 998200
rect 308121 998142 308384 998144
rect 451230 998142 470610 998202
rect 200665 998139 200731 998142
rect 253657 998139 253723 998142
rect 257337 998139 257403 998142
rect 308121 998139 308187 998142
rect 201861 998066 201927 998069
rect 253289 998066 253355 998069
rect 258165 998066 258231 998069
rect 260189 998066 260255 998069
rect 306925 998066 306991 998069
rect 201861 998064 202124 998066
rect 201861 998008 201866 998064
rect 201922 998008 202124 998064
rect 201861 998006 202124 998008
rect 253289 998064 253460 998066
rect 253289 998008 253294 998064
rect 253350 998008 253460 998064
rect 253289 998006 253460 998008
rect 258165 998064 258428 998066
rect 258165 998008 258170 998064
rect 258226 998008 258428 998064
rect 258165 998006 258428 998008
rect 260084 998064 260255 998066
rect 260084 998008 260194 998064
rect 260250 998008 260255 998064
rect 260084 998006 260255 998008
rect 306728 998064 306991 998066
rect 306728 998008 306930 998064
rect 306986 998008 306991 998064
rect 306728 998006 306991 998008
rect 201861 998003 201927 998006
rect 253289 998003 253355 998006
rect 258165 998003 258231 998006
rect 260189 998003 260255 998006
rect 306925 998003 306991 998006
rect 310605 998066 310671 998069
rect 310605 998064 310868 998066
rect 310605 998008 310610 998064
rect 310666 998008 310868 998064
rect 310605 998006 310868 998008
rect 310605 998003 310671 998006
rect 204713 997930 204779 997933
rect 252461 997930 252527 997933
rect 204713 997928 204976 997930
rect 204713 997872 204718 997928
rect 204774 997872 204976 997928
rect 204713 997870 204976 997872
rect 252264 997928 252527 997930
rect 252264 997872 252466 997928
rect 252522 997872 252527 997928
rect 252264 997870 252527 997872
rect 204713 997867 204779 997870
rect 252461 997867 252527 997870
rect 258993 997930 259059 997933
rect 259821 997930 259887 997933
rect 258993 997928 259164 997930
rect 258993 997872 258998 997928
rect 259054 997872 259164 997928
rect 258993 997870 259164 997872
rect 259624 997928 259887 997930
rect 259624 997872 259826 997928
rect 259882 997872 259887 997928
rect 259624 997870 259887 997872
rect 258993 997867 259059 997870
rect 259821 997867 259887 997870
rect 298277 997930 298343 997933
rect 303245 997930 303311 997933
rect 298277 997928 303311 997930
rect 298277 997872 298282 997928
rect 298338 997872 303250 997928
rect 303306 997872 303311 997928
rect 298277 997870 303311 997872
rect 298277 997867 298343 997870
rect 303245 997867 303311 997870
rect 304901 997930 304967 997933
rect 308949 997930 309015 997933
rect 304901 997928 305164 997930
rect 304901 997872 304906 997928
rect 304962 997872 305164 997928
rect 304901 997870 305164 997872
rect 308949 997928 309212 997930
rect 308949 997872 308954 997928
rect 309010 997872 309212 997928
rect 308949 997870 309212 997872
rect 304901 997867 304967 997870
rect 308949 997867 309015 997870
rect 203517 997794 203583 997797
rect 258165 997794 258231 997797
rect 203320 997792 203583 997794
rect 203320 997736 203522 997792
rect 203578 997736 203583 997792
rect 203320 997734 203583 997736
rect 257968 997792 258231 997794
rect 257968 997736 258170 997792
rect 258226 997736 258231 997792
rect 257968 997734 258231 997736
rect 203517 997731 203583 997734
rect 258165 997731 258231 997734
rect 260189 997794 260255 997797
rect 261845 997794 261911 997797
rect 309777 997794 309843 997797
rect 260189 997792 260452 997794
rect 260189 997736 260194 997792
rect 260250 997736 260452 997792
rect 260189 997734 260452 997736
rect 261845 997792 262108 997794
rect 261845 997736 261850 997792
rect 261906 997736 262108 997792
rect 261845 997734 262108 997736
rect 309580 997792 309843 997794
rect 309580 997736 309782 997792
rect 309838 997736 309843 997792
rect 309580 997734 309843 997736
rect 260189 997731 260255 997734
rect 261845 997731 261911 997734
rect 309777 997731 309843 997734
rect 383285 997660 383351 997661
rect 383285 997658 383332 997660
rect 383240 997656 383332 997658
rect 383240 997600 383290 997656
rect 383240 997598 383332 997600
rect 383285 997596 383332 997598
rect 383396 997596 383402 997660
rect 383285 997595 383351 997596
rect 97073 997250 97139 997253
rect 93810 997248 97139 997250
rect 93810 997192 97078 997248
rect 97134 997192 97139 997248
rect 93810 997190 97139 997192
rect 93810 996978 93870 997190
rect 97073 997187 97139 997190
rect 194358 997188 194364 997252
rect 194428 997250 194434 997252
rect 195697 997250 195763 997253
rect 194428 997248 195763 997250
rect 194428 997192 195702 997248
rect 195758 997192 195763 997248
rect 194428 997190 195763 997192
rect 194428 997188 194434 997190
rect 195697 997187 195763 997190
rect 229001 997250 229067 997253
rect 229185 997250 229251 997253
rect 229001 997248 229251 997250
rect 229001 997192 229006 997248
rect 229062 997192 229190 997248
rect 229246 997192 229251 997248
rect 229001 997190 229251 997192
rect 229001 997187 229067 997190
rect 229185 997187 229251 997190
rect 383469 997250 383535 997253
rect 389030 997250 389036 997252
rect 383469 997248 389036 997250
rect 383469 997192 383474 997248
rect 383530 997192 389036 997248
rect 383469 997190 389036 997192
rect 383469 997187 383535 997190
rect 389030 997188 389036 997190
rect 389100 997188 389106 997252
rect 247217 997114 247283 997117
rect 238526 997112 247283 997114
rect 238526 997056 247222 997112
rect 247278 997056 247283 997112
rect 238526 997054 247283 997056
rect 85990 996918 93870 996978
rect 85990 995757 86050 996918
rect 138054 996916 138060 996980
rect 138124 996978 138130 996980
rect 144269 996978 144335 996981
rect 138124 996976 144335 996978
rect 138124 996920 144274 996976
rect 144330 996920 144335 996976
rect 138124 996918 144335 996920
rect 138124 996916 138130 996918
rect 144269 996915 144335 996918
rect 145741 996706 145807 996709
rect 139166 996704 145807 996706
rect 139166 996648 145746 996704
rect 145802 996648 145807 996704
rect 139166 996646 145807 996648
rect 90214 996372 90220 996436
rect 90284 996434 90290 996436
rect 93301 996434 93367 996437
rect 90284 996432 93367 996434
rect 90284 996376 93306 996432
rect 93362 996376 93367 996432
rect 90284 996374 93367 996376
rect 90284 996372 90290 996374
rect 93301 996371 93367 996374
rect 86902 995964 86908 996028
rect 86972 996026 86978 996028
rect 86972 995966 93870 996026
rect 86972 995964 86978 995966
rect 85941 995752 86050 995757
rect 93485 995754 93551 995757
rect 85941 995696 85946 995752
rect 86002 995696 86050 995752
rect 85941 995694 86050 995696
rect 86358 995752 93551 995754
rect 86358 995696 93490 995752
rect 93546 995696 93551 995752
rect 86358 995694 93551 995696
rect 85941 995691 86007 995694
rect 84653 995482 84719 995485
rect 86358 995482 86418 995694
rect 93485 995691 93551 995694
rect 93810 995618 93870 995966
rect 139166 995757 139226 996646
rect 145741 996643 145807 996646
rect 195237 996706 195303 996709
rect 195237 996704 197186 996706
rect 195237 996648 195242 996704
rect 195298 996648 197186 996704
rect 195237 996646 197186 996648
rect 195237 996643 195303 996646
rect 144821 996434 144887 996437
rect 196801 996434 196867 996437
rect 141006 996432 144887 996434
rect 141006 996376 144826 996432
rect 144882 996376 144887 996432
rect 141006 996374 144887 996376
rect 141006 995757 141066 996374
rect 144821 996371 144887 996374
rect 188110 996432 196867 996434
rect 188110 996376 196806 996432
rect 196862 996376 196867 996432
rect 188110 996374 196867 996376
rect 197126 996434 197186 996646
rect 200205 996434 200271 996437
rect 197126 996432 200271 996434
rect 197126 996376 200210 996432
rect 200266 996376 200271 996432
rect 197126 996374 200271 996376
rect 188110 995757 188170 996374
rect 196801 996371 196867 996374
rect 200205 996371 200271 996374
rect 195513 996026 195579 996029
rect 192710 996024 195579 996026
rect 192710 995968 195518 996024
rect 195574 995968 195579 996024
rect 192710 995966 195579 995968
rect 133045 995754 133111 995757
rect 132450 995752 133111 995754
rect 132450 995696 133050 995752
rect 133106 995696 133111 995752
rect 132450 995694 133111 995696
rect 97441 995618 97507 995621
rect 93810 995616 97507 995618
rect 93810 995560 97446 995616
rect 97502 995560 97507 995616
rect 93810 995558 97507 995560
rect 97441 995555 97507 995558
rect 84653 995480 86418 995482
rect 84653 995424 84658 995480
rect 84714 995424 86418 995480
rect 84653 995422 86418 995424
rect 86585 995482 86651 995485
rect 90173 995484 90239 995485
rect 86902 995482 86908 995484
rect 86585 995480 86908 995482
rect 86585 995424 86590 995480
rect 86646 995424 86908 995480
rect 86585 995422 86908 995424
rect 84653 995419 84719 995422
rect 86585 995419 86651 995422
rect 86902 995420 86908 995422
rect 86972 995420 86978 995484
rect 90173 995482 90220 995484
rect 90128 995480 90220 995482
rect 90128 995424 90178 995480
rect 90128 995422 90220 995424
rect 90173 995420 90220 995422
rect 90284 995420 90290 995484
rect 90173 995419 90239 995420
rect 132450 995349 132510 995694
rect 133045 995691 133111 995694
rect 137369 995754 137435 995757
rect 138054 995754 138060 995756
rect 137369 995752 138060 995754
rect 137369 995696 137374 995752
rect 137430 995696 138060 995752
rect 137369 995694 138060 995696
rect 137369 995691 137435 995694
rect 138054 995692 138060 995694
rect 138124 995692 138130 995756
rect 139117 995752 139226 995757
rect 139117 995696 139122 995752
rect 139178 995696 139226 995752
rect 139117 995694 139226 995696
rect 140957 995752 141066 995757
rect 140957 995696 140962 995752
rect 141018 995696 141066 995752
rect 140957 995694 141066 995696
rect 141785 995754 141851 995757
rect 143717 995754 143783 995757
rect 141785 995752 143783 995754
rect 141785 995696 141790 995752
rect 141846 995696 143722 995752
rect 143778 995696 143783 995752
rect 141785 995694 143783 995696
rect 139117 995691 139183 995694
rect 140957 995691 141023 995694
rect 141785 995691 141851 995694
rect 143717 995691 143783 995694
rect 188061 995752 188170 995757
rect 189349 995756 189415 995757
rect 189349 995754 189396 995756
rect 188061 995696 188066 995752
rect 188122 995696 188170 995752
rect 188061 995694 188170 995696
rect 189304 995752 189396 995754
rect 189304 995696 189354 995752
rect 189304 995694 189396 995696
rect 188061 995691 188127 995694
rect 189349 995692 189396 995694
rect 189460 995692 189466 995756
rect 192477 995754 192543 995757
rect 192710 995754 192770 995966
rect 195513 995963 195579 995966
rect 204069 995890 204135 995893
rect 205314 995890 205374 996132
rect 204069 995888 205374 995890
rect 204069 995832 204074 995888
rect 204130 995832 205374 995888
rect 204069 995830 205374 995832
rect 204069 995827 204135 995830
rect 238526 995757 238586 997054
rect 247217 997051 247283 997054
rect 376017 996978 376083 996981
rect 470550 996978 470610 998142
rect 551093 998066 551159 998069
rect 551093 998064 551356 998066
rect 551093 998008 551098 998064
rect 551154 998008 551356 998064
rect 551093 998006 551356 998008
rect 551093 998003 551159 998006
rect 550265 997930 550331 997933
rect 550068 997928 550331 997930
rect 550068 997872 550270 997928
rect 550326 997872 550331 997928
rect 550068 997870 550331 997872
rect 550265 997867 550331 997870
rect 553301 997930 553367 997933
rect 553301 997928 553380 997930
rect 553301 997872 553306 997928
rect 553362 997872 553380 997928
rect 553301 997870 553380 997872
rect 553301 997867 553367 997870
rect 551461 997794 551527 997797
rect 552289 997794 552355 997797
rect 551461 997792 551724 997794
rect 551461 997736 551466 997792
rect 551522 997736 551724 997792
rect 551461 997734 551724 997736
rect 552092 997792 552355 997794
rect 552092 997736 552294 997792
rect 552350 997736 552355 997792
rect 552092 997734 552355 997736
rect 551461 997731 551527 997734
rect 552289 997731 552355 997734
rect 376017 996976 387994 996978
rect 376017 996920 376022 996976
rect 376078 996920 387994 996976
rect 376017 996918 387994 996920
rect 470550 996918 477050 996978
rect 376017 996915 376083 996918
rect 242566 996780 242572 996844
rect 242636 996842 242642 996844
rect 249885 996842 249951 996845
rect 242636 996840 249951 996842
rect 242636 996784 249890 996840
rect 249946 996784 249951 996840
rect 242636 996782 249951 996784
rect 242636 996780 242642 996782
rect 249885 996779 249951 996782
rect 246757 996434 246823 996437
rect 243126 996432 246823 996434
rect 243126 996376 246762 996432
rect 246818 996376 246823 996432
rect 243126 996374 246823 996376
rect 243126 995890 243186 996374
rect 246757 996371 246823 996374
rect 295006 996372 295012 996436
rect 295076 996434 295082 996436
rect 299105 996434 299171 996437
rect 295076 996432 299171 996434
rect 295076 996376 299110 996432
rect 299166 996376 299171 996432
rect 295076 996374 299171 996376
rect 295076 996372 295082 996374
rect 299105 996371 299171 996374
rect 372337 996434 372403 996437
rect 372337 996432 385786 996434
rect 372337 996376 372342 996432
rect 372398 996376 385786 996432
rect 372337 996374 385786 996376
rect 372337 996371 372403 996374
rect 243854 996100 243860 996164
rect 243924 996162 243930 996164
rect 247861 996162 247927 996165
rect 243924 996160 247927 996162
rect 243924 996104 247866 996160
rect 247922 996104 247927 996160
rect 243924 996102 247927 996104
rect 243924 996100 243930 996102
rect 247861 996099 247927 996102
rect 298921 996026 298987 996029
rect 294462 996024 298987 996026
rect 294462 995968 298926 996024
rect 298982 995968 298987 996024
rect 294462 995966 298987 995968
rect 253473 995890 253539 995893
rect 242942 995830 243186 995890
rect 243494 995888 253539 995890
rect 243494 995832 253478 995888
rect 253534 995832 253539 995888
rect 243494 995830 253539 995832
rect 192477 995752 192770 995754
rect 192477 995696 192482 995752
rect 192538 995696 192770 995752
rect 192477 995694 192770 995696
rect 193121 995754 193187 995757
rect 195053 995754 195119 995757
rect 193121 995752 195119 995754
rect 193121 995696 193126 995752
rect 193182 995696 195058 995752
rect 195114 995696 195119 995752
rect 193121 995694 195119 995696
rect 238526 995752 238635 995757
rect 239581 995756 239647 995757
rect 239581 995754 239628 995756
rect 238526 995696 238574 995752
rect 238630 995696 238635 995752
rect 238526 995694 238635 995696
rect 239536 995752 239628 995754
rect 239536 995696 239586 995752
rect 239536 995694 239628 995696
rect 189349 995691 189415 995692
rect 192477 995691 192543 995694
rect 193121 995691 193187 995694
rect 195053 995691 195119 995694
rect 238569 995691 238635 995694
rect 239581 995692 239628 995694
rect 239692 995692 239698 995756
rect 242065 995754 242131 995757
rect 242942 995754 243002 995830
rect 243261 995756 243327 995757
rect 243261 995754 243308 995756
rect 242065 995752 243002 995754
rect 242065 995696 242070 995752
rect 242126 995696 243002 995752
rect 242065 995694 243002 995696
rect 243216 995752 243308 995754
rect 243216 995696 243266 995752
rect 243216 995694 243308 995696
rect 239581 995691 239647 995692
rect 242065 995691 242131 995694
rect 243261 995692 243308 995694
rect 243372 995692 243378 995756
rect 243261 995691 243327 995692
rect 136633 995482 136699 995485
rect 148317 995482 148383 995485
rect 136633 995480 148383 995482
rect 136633 995424 136638 995480
rect 136694 995424 148322 995480
rect 148378 995424 148383 995480
rect 136633 995422 148383 995424
rect 136633 995419 136699 995422
rect 148317 995419 148383 995422
rect 183829 995482 183895 995485
rect 202321 995482 202387 995485
rect 183829 995480 202387 995482
rect 183829 995424 183834 995480
rect 183890 995424 202326 995480
rect 202382 995424 202387 995480
rect 183829 995422 202387 995424
rect 183829 995419 183895 995422
rect 202321 995419 202387 995422
rect 235901 995482 235967 995485
rect 243494 995482 243554 995830
rect 253473 995827 253539 995830
rect 292481 995754 292547 995757
rect 294462 995754 294522 995966
rect 298921 995963 298987 995966
rect 295057 995756 295123 995757
rect 292481 995752 294522 995754
rect 292481 995696 292486 995752
rect 292542 995696 294522 995752
rect 292481 995694 294522 995696
rect 292481 995691 292547 995694
rect 295006 995692 295012 995756
rect 295076 995754 295123 995756
rect 296161 995754 296227 995757
rect 298093 995754 298159 995757
rect 295076 995752 295168 995754
rect 295118 995696 295168 995752
rect 295076 995694 295168 995696
rect 296161 995752 298159 995754
rect 296161 995696 296166 995752
rect 296222 995696 298098 995752
rect 298154 995696 298159 995752
rect 296161 995694 298159 995696
rect 295076 995692 295123 995694
rect 295057 995691 295123 995692
rect 296161 995691 296227 995694
rect 298093 995691 298159 995694
rect 243813 995620 243879 995621
rect 243813 995618 243860 995620
rect 243768 995616 243860 995618
rect 243768 995560 243818 995616
rect 243768 995558 243860 995560
rect 243813 995556 243860 995558
rect 243924 995556 243930 995620
rect 244089 995618 244155 995621
rect 247033 995618 247099 995621
rect 244089 995616 247099 995618
rect 244089 995560 244094 995616
rect 244150 995560 247038 995616
rect 247094 995560 247099 995616
rect 244089 995558 247099 995560
rect 243813 995555 243879 995556
rect 244089 995555 244155 995558
rect 247033 995555 247099 995558
rect 274582 995556 274588 995620
rect 274652 995618 274658 995620
rect 280705 995618 280771 995621
rect 274652 995616 280771 995618
rect 274652 995560 280710 995616
rect 280766 995560 280771 995616
rect 274652 995558 280771 995560
rect 274652 995556 274658 995558
rect 280705 995555 280771 995558
rect 302141 995618 302207 995621
rect 303846 995618 303906 996132
rect 385726 995757 385786 996374
rect 387934 995757 387994 996918
rect 439681 996706 439747 996709
rect 473302 996706 473308 996708
rect 439681 996704 473308 996706
rect 439681 996648 439686 996704
rect 439742 996648 473308 996704
rect 439681 996646 473308 996648
rect 439681 996643 439747 996646
rect 473302 996644 473308 996646
rect 473372 996644 473378 996708
rect 421005 996434 421071 996437
rect 396582 996432 421071 996434
rect 396582 996376 421010 996432
rect 421066 996376 421071 996432
rect 396582 996374 421071 996376
rect 396582 995757 396642 996374
rect 421005 996371 421071 996374
rect 439865 996434 439931 996437
rect 439865 996432 476498 996434
rect 439865 996376 439870 996432
rect 439926 996376 476498 996432
rect 439865 996374 476498 996376
rect 439865 996371 439931 996374
rect 449157 996162 449223 996165
rect 449157 996160 475394 996162
rect 449157 996104 449162 996160
rect 449218 996104 475394 996160
rect 449157 996102 475394 996104
rect 449157 996099 449223 996102
rect 462313 995890 462379 995893
rect 462313 995888 470610 995890
rect 462313 995832 462318 995888
rect 462374 995832 470610 995888
rect 462313 995830 470610 995832
rect 462313 995827 462379 995830
rect 383101 995754 383167 995757
rect 385033 995754 385099 995757
rect 383101 995752 385099 995754
rect 383101 995696 383106 995752
rect 383162 995696 385038 995752
rect 385094 995696 385099 995752
rect 383101 995694 385099 995696
rect 385726 995752 385835 995757
rect 385726 995696 385774 995752
rect 385830 995696 385835 995752
rect 385726 995694 385835 995696
rect 383101 995691 383167 995694
rect 385033 995691 385099 995694
rect 385769 995691 385835 995694
rect 387885 995752 387994 995757
rect 387885 995696 387890 995752
rect 387946 995696 387994 995752
rect 387885 995694 387994 995696
rect 387885 995691 387951 995694
rect 388110 995692 388116 995756
rect 388180 995754 388186 995756
rect 388713 995754 388779 995757
rect 388180 995752 388779 995754
rect 388180 995696 388718 995752
rect 388774 995696 388779 995752
rect 388180 995694 388779 995696
rect 388180 995692 388186 995694
rect 388713 995691 388779 995694
rect 389030 995692 389036 995756
rect 389100 995754 389106 995756
rect 389357 995754 389423 995757
rect 389100 995752 389423 995754
rect 389100 995696 389362 995752
rect 389418 995696 389423 995752
rect 389100 995694 389423 995696
rect 389100 995692 389106 995694
rect 389357 995691 389423 995694
rect 392393 995754 392459 995757
rect 392393 995752 393514 995754
rect 392393 995696 392398 995752
rect 392454 995696 393514 995752
rect 392393 995694 393514 995696
rect 392393 995691 392459 995694
rect 302141 995616 303906 995618
rect 302141 995560 302146 995616
rect 302202 995560 303906 995616
rect 302141 995558 303906 995560
rect 302141 995555 302207 995558
rect 235901 995480 243554 995482
rect 235901 995424 235906 995480
rect 235962 995424 243554 995480
rect 235901 995422 243554 995424
rect 294873 995482 294939 995485
rect 298645 995482 298711 995485
rect 294873 995480 298711 995482
rect 294873 995424 294878 995480
rect 294934 995424 298650 995480
rect 298706 995424 298711 995480
rect 294873 995422 298711 995424
rect 235901 995419 235967 995422
rect 294873 995419 294939 995422
rect 298645 995419 298711 995422
rect 393454 995349 393514 995694
rect 396533 995752 396642 995757
rect 396533 995696 396538 995752
rect 396594 995696 396642 995752
rect 396533 995694 396642 995696
rect 396533 995691 396599 995694
rect 470550 995482 470610 995830
rect 473353 995756 473419 995757
rect 473302 995692 473308 995756
rect 473372 995754 473419 995756
rect 475334 995754 475394 996102
rect 476438 995757 476498 996374
rect 476990 995757 477050 996918
rect 524045 996706 524111 996709
rect 529606 996706 529612 996708
rect 524045 996704 529612 996706
rect 524045 996648 524050 996704
rect 524106 996648 529612 996704
rect 524045 996646 529612 996648
rect 524045 996643 524111 996646
rect 529606 996644 529612 996646
rect 529676 996644 529682 996708
rect 590561 996706 590627 996709
rect 627126 996706 627132 996708
rect 590561 996704 627132 996706
rect 590561 996648 590566 996704
rect 590622 996648 627132 996704
rect 590561 996646 627132 996648
rect 590561 996643 590627 996646
rect 627126 996644 627132 996646
rect 627196 996644 627202 996708
rect 516869 996434 516935 996437
rect 590561 996434 590627 996437
rect 630806 996434 630812 996436
rect 516869 996432 537218 996434
rect 516869 996376 516874 996432
rect 516930 996376 537218 996432
rect 516869 996374 537218 996376
rect 516869 996371 516935 996374
rect 516685 996162 516751 996165
rect 516685 996160 528570 996162
rect 516685 996104 516690 996160
rect 516746 996104 528570 996160
rect 516685 996102 528570 996104
rect 516685 996099 516751 996102
rect 475929 995754 475995 995757
rect 473372 995752 473464 995754
rect 473414 995696 473464 995752
rect 473372 995694 473464 995696
rect 475334 995752 475995 995754
rect 475334 995696 475934 995752
rect 475990 995696 475995 995752
rect 475334 995694 475995 995696
rect 476438 995752 476547 995757
rect 476438 995696 476486 995752
rect 476542 995696 476547 995752
rect 476438 995694 476547 995696
rect 476990 995752 477099 995757
rect 476990 995696 477038 995752
rect 477094 995696 477099 995752
rect 476990 995694 477099 995696
rect 473372 995692 473419 995694
rect 473353 995691 473419 995692
rect 475929 995691 475995 995694
rect 476481 995691 476547 995694
rect 477033 995691 477099 995694
rect 485681 995754 485747 995757
rect 488901 995754 488967 995757
rect 485681 995752 488967 995754
rect 485681 995696 485686 995752
rect 485742 995696 488906 995752
rect 488962 995696 488967 995752
rect 485681 995694 488967 995696
rect 485681 995691 485747 995694
rect 488901 995691 488967 995694
rect 523677 995754 523743 995757
rect 524781 995754 524847 995757
rect 523677 995752 524847 995754
rect 523677 995696 523682 995752
rect 523738 995696 524786 995752
rect 524842 995696 524847 995752
rect 523677 995694 524847 995696
rect 523677 995691 523743 995694
rect 524781 995691 524847 995694
rect 480805 995482 480871 995485
rect 470550 995480 480871 995482
rect 470550 995424 480810 995480
rect 480866 995424 480871 995480
rect 470550 995422 480871 995424
rect 480805 995419 480871 995422
rect 523493 995482 523559 995485
rect 527909 995482 527975 995485
rect 523493 995480 527975 995482
rect 523493 995424 523498 995480
rect 523554 995424 527914 995480
rect 527970 995424 527975 995480
rect 523493 995422 527975 995424
rect 528510 995482 528570 996102
rect 537158 995757 537218 996374
rect 590561 996432 630812 996434
rect 590561 996376 590566 996432
rect 590622 996376 630812 996432
rect 590561 996374 630812 996376
rect 590561 996371 590627 996374
rect 630806 996372 630812 996374
rect 630876 996372 630882 996436
rect 625429 996026 625495 996029
rect 625429 996024 630690 996026
rect 625429 995968 625434 996024
rect 625490 995968 630690 996024
rect 625429 995966 630690 995968
rect 625429 995963 625495 995966
rect 529606 995692 529612 995756
rect 529676 995754 529682 995756
rect 529841 995754 529907 995757
rect 536557 995756 536623 995757
rect 536557 995754 536604 995756
rect 529676 995752 529907 995754
rect 529676 995696 529846 995752
rect 529902 995696 529907 995752
rect 529676 995694 529907 995696
rect 536512 995752 536604 995754
rect 536512 995696 536562 995752
rect 536512 995694 536604 995696
rect 529676 995692 529682 995694
rect 529841 995691 529907 995694
rect 536557 995692 536604 995694
rect 536668 995692 536674 995756
rect 537158 995752 537267 995757
rect 537158 995696 537206 995752
rect 537262 995696 537267 995752
rect 537158 995694 537267 995696
rect 536557 995691 536623 995692
rect 537201 995691 537267 995694
rect 623681 995754 623747 995757
rect 626533 995754 626599 995757
rect 627177 995756 627243 995757
rect 623681 995752 626599 995754
rect 623681 995696 623686 995752
rect 623742 995696 626538 995752
rect 626594 995696 626599 995752
rect 623681 995694 626599 995696
rect 623681 995691 623747 995694
rect 626533 995691 626599 995694
rect 627126 995692 627132 995756
rect 627196 995754 627243 995756
rect 630630 995754 630690 995966
rect 631501 995754 631567 995757
rect 627196 995752 627288 995754
rect 627238 995696 627288 995752
rect 627196 995694 627288 995696
rect 630630 995752 631567 995754
rect 630630 995696 631506 995752
rect 631562 995696 631567 995752
rect 630630 995694 631567 995696
rect 627196 995692 627243 995694
rect 627177 995691 627243 995692
rect 631501 995691 631567 995694
rect 533429 995482 533495 995485
rect 528510 995480 533495 995482
rect 528510 995424 533434 995480
rect 533490 995424 533495 995480
rect 528510 995422 533495 995424
rect 523493 995419 523559 995422
rect 527909 995419 527975 995422
rect 533429 995419 533495 995422
rect 537845 995482 537911 995485
rect 538213 995482 538279 995485
rect 537845 995480 538279 995482
rect 537845 995424 537850 995480
rect 537906 995424 538218 995480
rect 538274 995424 538279 995480
rect 537845 995422 538279 995424
rect 537845 995419 537911 995422
rect 538213 995419 538279 995422
rect 625613 995482 625679 995485
rect 630213 995482 630279 995485
rect 630857 995484 630923 995485
rect 625613 995480 630279 995482
rect 625613 995424 625618 995480
rect 625674 995424 630218 995480
rect 630274 995424 630279 995480
rect 625613 995422 630279 995424
rect 625613 995419 625679 995422
rect 630213 995419 630279 995422
rect 630806 995420 630812 995484
rect 630876 995482 630923 995484
rect 630876 995480 630968 995482
rect 630918 995424 630968 995480
rect 630876 995422 630968 995424
rect 630876 995420 630923 995422
rect 630857 995419 630923 995420
rect 97257 995346 97323 995349
rect 93350 995344 97323 995346
rect 93350 995288 97262 995344
rect 97318 995288 97323 995344
rect 93350 995286 97323 995288
rect 85021 995210 85087 995213
rect 93350 995210 93410 995286
rect 97257 995283 97323 995286
rect 132401 995344 132510 995349
rect 132401 995288 132406 995344
rect 132462 995288 132510 995344
rect 132401 995286 132510 995288
rect 245561 995346 245627 995349
rect 246573 995346 246639 995349
rect 245561 995344 246639 995346
rect 245561 995288 245566 995344
rect 245622 995288 246578 995344
rect 246634 995288 246639 995344
rect 245561 995286 246639 995288
rect 132401 995283 132467 995286
rect 245561 995283 245627 995286
rect 246573 995283 246639 995286
rect 381445 995346 381511 995349
rect 392301 995346 392367 995349
rect 381445 995344 392367 995346
rect 381445 995288 381450 995344
rect 381506 995288 392306 995344
rect 392362 995288 392367 995344
rect 381445 995286 392367 995288
rect 393454 995344 393563 995349
rect 393454 995288 393502 995344
rect 393558 995288 393563 995344
rect 393454 995286 393563 995288
rect 381445 995283 381511 995286
rect 392301 995283 392367 995286
rect 393497 995283 393563 995286
rect 85021 995208 93410 995210
rect 85021 995152 85026 995208
rect 85082 995152 93410 995208
rect 85021 995150 93410 995152
rect 472065 995210 472131 995213
rect 478229 995210 478295 995213
rect 472065 995208 478295 995210
rect 472065 995152 472070 995208
rect 472126 995152 478234 995208
rect 478290 995152 478295 995208
rect 472065 995150 478295 995152
rect 85021 995147 85087 995150
rect 472065 995147 472131 995150
rect 478229 995147 478295 995150
rect 478781 995210 478847 995213
rect 481541 995210 481607 995213
rect 478781 995208 481607 995210
rect 478781 995152 478786 995208
rect 478842 995152 481546 995208
rect 481602 995152 481607 995208
rect 478781 995150 481607 995152
rect 478781 995147 478847 995150
rect 481541 995147 481607 995150
rect 523125 995210 523191 995213
rect 526253 995210 526319 995213
rect 523125 995208 526319 995210
rect 523125 995152 523130 995208
rect 523186 995152 526258 995208
rect 526314 995152 526319 995208
rect 523125 995150 526319 995152
rect 523125 995147 523191 995150
rect 526253 995147 526319 995150
rect 93485 995074 93551 995077
rect 100017 995074 100083 995077
rect 93485 995072 100083 995074
rect 93485 995016 93490 995072
rect 93546 995016 100022 995072
rect 100078 995016 100083 995072
rect 93485 995014 100083 995016
rect 93485 995011 93551 995014
rect 100017 995011 100083 995014
rect 135897 995074 135963 995077
rect 152457 995074 152523 995077
rect 135897 995072 152523 995074
rect 135897 995016 135902 995072
rect 135958 995016 152462 995072
rect 152518 995016 152523 995072
rect 135897 995014 152523 995016
rect 135897 995011 135963 995014
rect 152457 995011 152523 995014
rect 290273 995074 290339 995077
rect 307017 995074 307083 995077
rect 290273 995072 307083 995074
rect 290273 995016 290278 995072
rect 290334 995016 307022 995072
rect 307078 995016 307083 995072
rect 290273 995014 307083 995016
rect 290273 995011 290339 995014
rect 307017 995011 307083 995014
rect 374637 995074 374703 995077
rect 388345 995074 388411 995077
rect 374637 995072 388411 995074
rect 374637 995016 374642 995072
rect 374698 995016 388350 995072
rect 388406 995016 388411 995072
rect 374637 995014 388411 995016
rect 374637 995011 374703 995014
rect 388345 995011 388411 995014
rect 617333 995074 617399 995077
rect 629661 995074 629727 995077
rect 617333 995072 629727 995074
rect 617333 995016 617338 995072
rect 617394 995016 629666 995072
rect 629722 995016 629727 995072
rect 617333 995014 629727 995016
rect 617333 995011 617399 995014
rect 629661 995011 629727 995014
rect 187601 994938 187667 994941
rect 203333 994938 203399 994941
rect 187601 994936 203399 994938
rect 187601 994880 187606 994936
rect 187662 994880 203338 994936
rect 203394 994880 203399 994936
rect 187601 994878 203399 994880
rect 187601 994875 187667 994878
rect 203333 994875 203399 994878
rect 236545 994938 236611 994941
rect 251817 994938 251883 994941
rect 236545 994936 251883 994938
rect 236545 994880 236550 994936
rect 236606 994880 251822 994936
rect 251878 994880 251883 994936
rect 236545 994878 251883 994880
rect 236545 994875 236611 994878
rect 251817 994875 251883 994878
rect 446857 994938 446923 994941
rect 475745 994938 475811 994941
rect 487797 994938 487863 994941
rect 446857 994936 475578 994938
rect 446857 994880 446862 994936
rect 446918 994880 475578 994936
rect 446857 994878 475578 994880
rect 446857 994875 446923 994878
rect 89345 994802 89411 994805
rect 106457 994802 106523 994805
rect 89345 994800 106523 994802
rect 89345 994744 89350 994800
rect 89406 994744 106462 994800
rect 106518 994744 106523 994800
rect 89345 994742 106523 994744
rect 89345 994739 89411 994742
rect 106457 994739 106523 994742
rect 129089 994802 129155 994805
rect 151077 994802 151143 994805
rect 129089 994800 151143 994802
rect 129089 994744 129094 994800
rect 129150 994744 151082 994800
rect 151138 994744 151143 994800
rect 129089 994742 151143 994744
rect 129089 994739 129155 994742
rect 151077 994739 151143 994742
rect 287789 994802 287855 994805
rect 300117 994802 300183 994805
rect 287789 994800 300183 994802
rect 287789 994744 287794 994800
rect 287850 994744 300122 994800
rect 300178 994744 300183 994800
rect 287789 994742 300183 994744
rect 287789 994739 287855 994742
rect 300117 994739 300183 994742
rect 375557 994802 375623 994805
rect 395153 994802 395219 994805
rect 375557 994800 395219 994802
rect 375557 994744 375562 994800
rect 375618 994744 395158 994800
rect 395214 994744 395219 994800
rect 375557 994742 395219 994744
rect 375557 994739 375623 994742
rect 395153 994739 395219 994742
rect 188797 994666 188863 994669
rect 194685 994666 194751 994669
rect 188797 994664 194751 994666
rect 188797 994608 188802 994664
rect 188858 994608 194690 994664
rect 194746 994608 194751 994664
rect 188797 994606 194751 994608
rect 188797 994603 188863 994606
rect 194685 994603 194751 994606
rect 240869 994666 240935 994669
rect 247677 994666 247743 994669
rect 240869 994664 247743 994666
rect 240869 994608 240874 994664
rect 240930 994608 247682 994664
rect 247738 994608 247743 994664
rect 240869 994606 247743 994608
rect 240869 994603 240935 994606
rect 247677 994603 247743 994606
rect 452285 994666 452351 994669
rect 475518 994666 475578 994878
rect 475745 994936 487863 994938
rect 475745 994880 475750 994936
rect 475806 994880 487802 994936
rect 487858 994880 487863 994936
rect 475745 994878 487863 994880
rect 475745 994875 475811 994878
rect 487797 994875 487863 994878
rect 518157 994802 518223 994805
rect 535545 994802 535611 994805
rect 518157 994800 535611 994802
rect 518157 994744 518162 994800
rect 518218 994744 535550 994800
rect 535606 994744 535611 994800
rect 518157 994742 535611 994744
rect 518157 994739 518223 994742
rect 535545 994739 535611 994742
rect 625429 994802 625495 994805
rect 634721 994802 634787 994805
rect 625429 994800 634787 994802
rect 625429 994744 625434 994800
rect 625490 994744 634726 994800
rect 634782 994744 634787 994800
rect 625429 994742 634787 994744
rect 625429 994739 625495 994742
rect 634721 994739 634787 994742
rect 484117 994666 484183 994669
rect 452285 994664 475394 994666
rect 452285 994608 452290 994664
rect 452346 994608 475394 994664
rect 452285 994606 475394 994608
rect 475518 994664 484183 994666
rect 475518 994608 484122 994664
rect 484178 994608 484183 994664
rect 475518 994606 484183 994608
rect 452285 994603 452351 994606
rect 80697 994530 80763 994533
rect 129733 994530 129799 994533
rect 155217 994530 155283 994533
rect 80697 994528 84210 994530
rect 80697 994472 80702 994528
rect 80758 994472 84210 994528
rect 80697 994470 84210 994472
rect 80697 994467 80763 994470
rect 84150 994394 84210 994470
rect 129733 994528 155283 994530
rect 129733 994472 129738 994528
rect 129794 994472 155222 994528
rect 155278 994472 155283 994528
rect 129733 994470 155283 994472
rect 129733 994467 129799 994470
rect 155217 994467 155283 994470
rect 94497 994394 94563 994397
rect 84150 994392 94563 994394
rect 84150 994336 94502 994392
rect 94558 994336 94563 994392
rect 84150 994334 94563 994336
rect 94497 994331 94563 994334
rect 184841 994394 184907 994397
rect 195053 994394 195119 994397
rect 184841 994392 195119 994394
rect 184841 994336 184846 994392
rect 184902 994336 195058 994392
rect 195114 994336 195119 994392
rect 184841 994334 195119 994336
rect 184841 994331 184907 994334
rect 195053 994331 195119 994334
rect 466453 994394 466519 994397
rect 475334 994394 475394 994606
rect 484117 994603 484183 994606
rect 482921 994394 482987 994397
rect 466453 994392 470610 994394
rect 466453 994336 466458 994392
rect 466514 994336 470610 994392
rect 466453 994334 470610 994336
rect 475334 994392 482987 994394
rect 475334 994336 482926 994392
rect 482982 994336 482987 994392
rect 475334 994334 482987 994336
rect 466453 994331 466519 994334
rect 291469 994258 291535 994261
rect 304257 994258 304323 994261
rect 291469 994256 304323 994258
rect 291469 994200 291474 994256
rect 291530 994200 304262 994256
rect 304318 994200 304323 994256
rect 291469 994198 304323 994200
rect 291469 994195 291535 994198
rect 304257 994195 304323 994198
rect 87505 994122 87571 994125
rect 92657 994122 92723 994125
rect 87505 994120 92723 994122
rect 87505 994064 87510 994120
rect 87566 994064 92662 994120
rect 92718 994064 92723 994120
rect 87505 994062 92723 994064
rect 87505 994059 87571 994062
rect 92657 994059 92723 994062
rect 190361 994122 190427 994125
rect 200757 994122 200823 994125
rect 190361 994120 200823 994122
rect 190361 994064 190366 994120
rect 190422 994064 200762 994120
rect 200818 994064 200823 994120
rect 190361 994062 200823 994064
rect 470550 994122 470610 994334
rect 482921 994331 482987 994334
rect 475745 994122 475811 994125
rect 470550 994120 475811 994122
rect 470550 994064 475750 994120
rect 475806 994064 475811 994120
rect 470550 994062 475811 994064
rect 190361 994059 190427 994062
rect 200757 994059 200823 994062
rect 475745 994059 475811 994062
rect 133137 993986 133203 993989
rect 142797 993986 142863 993989
rect 133137 993984 142863 993986
rect 133137 993928 133142 993984
rect 133198 993928 142802 993984
rect 142858 993928 142863 993984
rect 133137 993926 142863 993928
rect 133137 993923 133203 993926
rect 142797 993923 142863 993926
rect 287513 993986 287579 993989
rect 298001 993986 298067 993989
rect 287513 993984 298067 993986
rect 287513 993928 287518 993984
rect 287574 993928 298006 993984
rect 298062 993928 298067 993984
rect 287513 993926 298067 993928
rect 287513 993923 287579 993926
rect 298001 993923 298067 993926
rect 567837 993714 567903 993717
rect 633985 993714 634051 993717
rect 567837 993712 634051 993714
rect 567837 993656 567842 993712
rect 567898 993656 633990 993712
rect 634046 993656 634051 993712
rect 567837 993654 634051 993656
rect 567837 993651 567903 993654
rect 633985 993651 634051 993654
rect 573214 989436 573220 989500
rect 573284 989498 573290 989500
rect 576301 989498 576367 989501
rect 573284 989496 576367 989498
rect 573284 989440 576306 989496
rect 576362 989440 576367 989496
rect 573284 989438 576367 989440
rect 573284 989436 573290 989438
rect 576301 989435 576367 989438
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651557 975898 651623 975901
rect 650164 975896 651623 975898
rect 650164 975840 651562 975896
rect 651618 975840 651623 975896
rect 650164 975838 651623 975840
rect 651557 975835 651623 975838
rect 41454 968764 41460 968828
rect 41524 968826 41530 968828
rect 41781 968826 41847 968829
rect 41524 968824 41847 968826
rect 41524 968768 41786 968824
rect 41842 968768 41847 968824
rect 41524 968766 41847 968768
rect 41524 968764 41530 968766
rect 41781 968763 41847 968766
rect 41965 967196 42031 967197
rect 41965 967192 42012 967196
rect 42076 967194 42082 967196
rect 41965 967136 41970 967192
rect 41965 967132 42012 967136
rect 42076 967134 42122 967194
rect 42076 967132 42082 967134
rect 41965 967131 42031 967132
rect 675385 966516 675451 966517
rect 675334 966514 675340 966516
rect 675294 966454 675340 966514
rect 675404 966512 675451 966516
rect 675446 966456 675451 966512
rect 675334 966452 675340 966454
rect 675404 966452 675451 966456
rect 675385 966451 675451 966452
rect 675753 965154 675819 965157
rect 676070 965154 676076 965156
rect 675753 965152 676076 965154
rect 675753 965096 675758 965152
rect 675814 965096 676076 965152
rect 675753 965094 676076 965096
rect 675753 965091 675819 965094
rect 676070 965092 676076 965094
rect 676140 965092 676146 965156
rect 675201 963388 675267 963389
rect 675150 963386 675156 963388
rect 675110 963326 675156 963386
rect 675220 963384 675267 963388
rect 675262 963328 675267 963384
rect 675150 963324 675156 963326
rect 675220 963324 675267 963328
rect 675201 963323 675267 963324
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 651557 962570 651623 962573
rect 650164 962568 651623 962570
rect 650164 962512 651562 962568
rect 651618 962512 651623 962568
rect 650164 962510 651623 962512
rect 651557 962507 651623 962510
rect 41781 962164 41847 962165
rect 41781 962160 41828 962164
rect 41892 962162 41898 962164
rect 41781 962104 41786 962160
rect 41781 962100 41828 962104
rect 41892 962102 41938 962162
rect 41892 962100 41898 962102
rect 41781 962099 41847 962100
rect 675753 962026 675819 962029
rect 676622 962026 676628 962028
rect 675753 962024 676628 962026
rect 675753 961968 675758 962024
rect 675814 961968 676628 962024
rect 675753 961966 676628 961968
rect 675753 961963 675819 961966
rect 676622 961964 676628 961966
rect 676692 961964 676698 962028
rect 674925 959442 674991 959445
rect 675150 959442 675156 959444
rect 674925 959440 675156 959442
rect 674925 959384 674930 959440
rect 674986 959384 675156 959440
rect 674925 959382 675156 959384
rect 674925 959379 674991 959382
rect 675150 959380 675156 959382
rect 675220 959380 675226 959444
rect 41270 959108 41276 959172
rect 41340 959170 41346 959172
rect 41781 959170 41847 959173
rect 41340 959168 41847 959170
rect 41340 959112 41786 959168
rect 41842 959112 41847 959168
rect 41340 959110 41847 959112
rect 41340 959108 41346 959110
rect 41781 959107 41847 959110
rect 672993 959170 673059 959173
rect 675109 959170 675175 959173
rect 672993 959168 675175 959170
rect 672993 959112 672998 959168
rect 673054 959112 675114 959168
rect 675170 959112 675175 959168
rect 672993 959110 675175 959112
rect 672993 959107 673059 959110
rect 675109 959107 675175 959110
rect 675753 958354 675819 958357
rect 676990 958354 676996 958356
rect 675753 958352 676996 958354
rect 675753 958296 675758 958352
rect 675814 958296 676996 958352
rect 675753 958294 676996 958296
rect 675753 958291 675819 958294
rect 676990 958292 676996 958294
rect 677060 958292 677066 958356
rect 40718 956524 40724 956588
rect 40788 956586 40794 956588
rect 41781 956586 41847 956589
rect 40788 956584 41847 956586
rect 40788 956528 41786 956584
rect 41842 956528 41847 956584
rect 40788 956526 41847 956528
rect 40788 956524 40794 956526
rect 41781 956523 41847 956526
rect 675753 956450 675819 956453
rect 676806 956450 676812 956452
rect 675753 956448 676812 956450
rect 675753 956392 675758 956448
rect 675814 956392 676812 956448
rect 675753 956390 676812 956392
rect 675753 956387 675819 956390
rect 676806 956388 676812 956390
rect 676876 956388 676882 956452
rect 40534 955436 40540 955500
rect 40604 955498 40610 955500
rect 41781 955498 41847 955501
rect 40604 955496 41847 955498
rect 40604 955440 41786 955496
rect 41842 955440 41847 955496
rect 40604 955438 41847 955440
rect 40604 955436 40610 955438
rect 41781 955435 41847 955438
rect 39297 952506 39363 952509
rect 41638 952506 41644 952508
rect 39297 952504 41644 952506
rect 39297 952448 39302 952504
rect 39358 952448 41644 952504
rect 39297 952446 41644 952448
rect 39297 952443 39363 952446
rect 41638 952444 41644 952446
rect 41708 952444 41714 952508
rect 37917 952234 37983 952237
rect 41454 952234 41460 952236
rect 37917 952232 41460 952234
rect 37917 952176 37922 952232
rect 37978 952176 41460 952232
rect 37917 952174 41460 952176
rect 37917 952171 37983 952174
rect 41454 952172 41460 952174
rect 41524 952172 41530 952236
rect 674097 952234 674163 952237
rect 675477 952234 675543 952237
rect 674097 952232 675543 952234
rect 674097 952176 674102 952232
rect 674158 952176 675482 952232
rect 675538 952176 675543 952232
rect 674097 952174 675543 952176
rect 674097 952171 674163 952174
rect 675477 952171 675543 952174
rect 40033 951690 40099 951693
rect 41270 951690 41276 951692
rect 40033 951688 41276 951690
rect 40033 951632 40038 951688
rect 40094 951632 41276 951688
rect 40033 951630 41276 951632
rect 40033 951627 40099 951630
rect 41270 951628 41276 951630
rect 41340 951628 41346 951692
rect 41505 951690 41571 951693
rect 42006 951690 42012 951692
rect 41505 951688 42012 951690
rect 41505 951632 41510 951688
rect 41566 951632 42012 951688
rect 41505 951630 42012 951632
rect 41505 951627 41571 951630
rect 42006 951628 42012 951630
rect 42076 951628 42082 951692
rect 676622 951492 676628 951556
rect 676692 951554 676698 951556
rect 677501 951554 677567 951557
rect 676692 951552 677567 951554
rect 676692 951496 677506 951552
rect 677562 951496 677567 951552
rect 676692 951494 677567 951496
rect 676692 951492 676698 951494
rect 677501 951491 677567 951494
rect 676070 949996 676076 950060
rect 676140 950058 676146 950060
rect 683297 950058 683363 950061
rect 676140 950056 683363 950058
rect 676140 950000 683302 950056
rect 683358 950000 683363 950056
rect 676140 949998 683363 950000
rect 676140 949996 676146 949998
rect 683297 949995 683363 949998
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 651557 949378 651623 949381
rect 650164 949376 651623 949378
rect 650164 949320 651562 949376
rect 651618 949320 651623 949376
rect 650164 949318 651623 949320
rect 651557 949315 651623 949318
rect 674925 948970 674991 948973
rect 675334 948970 675340 948972
rect 674925 948968 675340 948970
rect 674925 948912 674930 948968
rect 674986 948912 675340 948968
rect 674925 948910 675340 948912
rect 674925 948907 674991 948910
rect 675334 948908 675340 948910
rect 675404 948908 675410 948972
rect 43529 943530 43595 943533
rect 41492 943528 43595 943530
rect 41492 943472 43534 943528
rect 43590 943472 43595 943528
rect 41492 943470 43595 943472
rect 43529 943467 43595 943470
rect 44633 943122 44699 943125
rect 41492 943120 44699 943122
rect 41492 943064 44638 943120
rect 44694 943064 44699 943120
rect 41492 943062 44699 943064
rect 44633 943059 44699 943062
rect 47577 942714 47643 942717
rect 41492 942712 47643 942714
rect 41492 942656 47582 942712
rect 47638 942656 47643 942712
rect 41492 942654 47643 942656
rect 47577 942651 47643 942654
rect 43437 942306 43503 942309
rect 41492 942304 43503 942306
rect 41492 942248 43442 942304
rect 43498 942248 43503 942304
rect 41492 942246 43503 942248
rect 43437 942243 43503 942246
rect 41321 941898 41387 941901
rect 41308 941896 41387 941898
rect 41308 941840 41326 941896
rect 41382 941840 41387 941896
rect 41308 941838 41387 941840
rect 41321 941835 41387 941838
rect 674925 941898 674991 941901
rect 675845 941898 675911 941901
rect 674925 941896 675911 941898
rect 674925 941840 674930 941896
rect 674986 941840 675850 941896
rect 675906 941840 675911 941896
rect 674925 941838 675911 941840
rect 674925 941835 674991 941838
rect 675845 941835 675911 941838
rect 41324 941490 41890 941524
rect 41308 941464 41890 941490
rect 41308 941430 41384 941464
rect 41830 941354 41890 941464
rect 43621 941354 43687 941357
rect 41830 941352 43687 941354
rect 41830 941296 43626 941352
rect 43682 941296 43687 941352
rect 41830 941294 43687 941296
rect 43621 941291 43687 941294
rect 40953 941082 41019 941085
rect 40940 941080 41019 941082
rect 40940 941024 40958 941080
rect 41014 941024 41019 941080
rect 40940 941022 41019 941024
rect 40953 941019 41019 941022
rect 46197 940674 46263 940677
rect 41492 940672 46263 940674
rect 41492 940616 46202 940672
rect 46258 940616 46263 940672
rect 41492 940614 46263 940616
rect 46197 940611 46263 940614
rect 42057 940266 42123 940269
rect 41492 940264 42123 940266
rect 41492 940208 42062 940264
rect 42118 940208 42123 940264
rect 41492 940206 42123 940208
rect 42057 940203 42123 940206
rect 675477 939994 675543 939997
rect 675477 939992 676292 939994
rect 675477 939936 675482 939992
rect 675538 939936 676292 939992
rect 675477 939934 676292 939936
rect 675477 939931 675543 939934
rect 43437 939858 43503 939861
rect 41492 939856 43503 939858
rect 41492 939800 43442 939856
rect 43498 939800 43503 939856
rect 41492 939798 43503 939800
rect 43437 939795 43503 939798
rect 674925 939586 674991 939589
rect 674925 939584 676292 939586
rect 674925 939528 674930 939584
rect 674986 939528 676292 939584
rect 674925 939526 676292 939528
rect 674925 939523 674991 939526
rect 41137 939450 41203 939453
rect 41124 939448 41203 939450
rect 41124 939392 41142 939448
rect 41198 939392 41203 939448
rect 41124 939390 41203 939392
rect 41137 939387 41203 939390
rect 675293 939178 675359 939181
rect 675293 939176 676292 939178
rect 675293 939120 675298 939176
rect 675354 939120 676292 939176
rect 675293 939118 676292 939120
rect 675293 939115 675359 939118
rect 41822 939042 41828 939044
rect 41492 938982 41828 939042
rect 41822 938980 41828 938982
rect 41892 938980 41898 939044
rect 675477 938770 675543 938773
rect 675477 938768 676292 938770
rect 675477 938712 675482 938768
rect 675538 938712 676292 938768
rect 675477 938710 676292 938712
rect 675477 938707 675543 938710
rect 40910 938467 40970 938604
rect 35157 938464 35223 938467
rect 35157 938462 35266 938464
rect 35157 938406 35162 938462
rect 35218 938406 35266 938462
rect 35157 938401 35266 938406
rect 40910 938462 41019 938467
rect 40910 938406 40958 938462
rect 41014 938406 41019 938462
rect 40910 938404 41019 938406
rect 40953 938401 41019 938404
rect 35206 938196 35266 938401
rect 675477 938362 675543 938365
rect 675477 938360 676292 938362
rect 675477 938304 675482 938360
rect 675538 938304 676292 938360
rect 675477 938302 676292 938304
rect 675477 938299 675543 938302
rect 674925 937954 674991 937957
rect 674925 937952 676292 937954
rect 674925 937896 674930 937952
rect 674986 937896 676292 937952
rect 674925 937894 676292 937896
rect 674925 937891 674991 937894
rect 42241 937818 42307 937821
rect 41492 937816 42307 937818
rect 41492 937760 42246 937816
rect 42302 937760 42307 937816
rect 41492 937758 42307 937760
rect 42241 937755 42307 937758
rect 675293 937546 675359 937549
rect 675293 937544 676292 937546
rect 675293 937488 675298 937544
rect 675354 937488 676292 937544
rect 675293 937486 676292 937488
rect 675293 937483 675359 937486
rect 39297 937410 39363 937413
rect 39284 937408 39363 937410
rect 39284 937352 39302 937408
rect 39358 937352 39363 937408
rect 39284 937350 39363 937352
rect 39297 937347 39363 937350
rect 675477 937138 675543 937141
rect 675477 937136 676292 937138
rect 675477 937080 675482 937136
rect 675538 937080 676292 937136
rect 675477 937078 676292 937080
rect 675477 937075 675543 937078
rect 37917 937002 37983 937005
rect 62113 937002 62179 937005
rect 37917 937000 37996 937002
rect 37917 936944 37922 937000
rect 37978 936944 37996 937000
rect 37917 936942 37996 936944
rect 62113 937000 64492 937002
rect 62113 936944 62118 937000
rect 62174 936944 64492 937000
rect 62113 936942 64492 936944
rect 37917 936939 37983 936942
rect 62113 936939 62179 936942
rect 675661 936730 675727 936733
rect 675661 936728 676292 936730
rect 675661 936672 675666 936728
rect 675722 936672 676292 936728
rect 675661 936670 676292 936672
rect 675661 936667 675727 936670
rect 41822 936594 41828 936596
rect 41492 936534 41828 936594
rect 41822 936532 41828 936534
rect 41892 936532 41898 936596
rect 675477 936322 675543 936325
rect 675477 936320 676292 936322
rect 675477 936264 675482 936320
rect 675538 936264 676292 936320
rect 675477 936262 676292 936264
rect 675477 936259 675543 936262
rect 44817 936186 44883 936189
rect 651557 936186 651623 936189
rect 41492 936184 44883 936186
rect 41492 936128 44822 936184
rect 44878 936128 44883 936184
rect 41492 936126 44883 936128
rect 650164 936184 651623 936186
rect 650164 936128 651562 936184
rect 651618 936128 651623 936184
rect 650164 936126 651623 936128
rect 44817 936123 44883 936126
rect 651557 936123 651623 936126
rect 675293 935914 675359 935917
rect 675293 935912 676292 935914
rect 675293 935856 675298 935912
rect 675354 935856 676292 935912
rect 675293 935854 676292 935856
rect 675293 935851 675359 935854
rect 40033 935778 40099 935781
rect 40020 935776 40099 935778
rect 40020 935720 40038 935776
rect 40094 935720 40099 935776
rect 40020 935718 40099 935720
rect 40033 935715 40099 935718
rect 683297 935642 683363 935645
rect 683254 935640 683363 935642
rect 683254 935584 683302 935640
rect 683358 935584 683363 935640
rect 683254 935579 683363 935584
rect 683254 935476 683314 935579
rect 42793 935370 42859 935373
rect 41492 935368 42859 935370
rect 41492 935312 42798 935368
rect 42854 935312 42859 935368
rect 41492 935310 42859 935312
rect 42793 935307 42859 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 43069 934962 43135 934965
rect 41492 934960 43135 934962
rect 41492 934904 43074 934960
rect 43130 934904 43135 934960
rect 41492 934902 43135 934904
rect 43069 934899 43135 934902
rect 675845 934690 675911 934693
rect 675845 934688 676292 934690
rect 675845 934632 675850 934688
rect 675906 934632 676292 934688
rect 675845 934630 676292 934632
rect 675845 934627 675911 934630
rect 43253 934554 43319 934557
rect 41492 934552 43319 934554
rect 41492 934496 43258 934552
rect 43314 934496 43319 934552
rect 41492 934494 43319 934496
rect 43253 934491 43319 934494
rect 44449 934146 44515 934149
rect 41492 934144 44515 934146
rect 41492 934088 44454 934144
rect 44510 934088 44515 934144
rect 41492 934086 44515 934088
rect 44449 934083 44515 934086
rect 675109 934146 675175 934149
rect 676262 934146 676322 934252
rect 675109 934144 676322 934146
rect 675109 934088 675114 934144
rect 675170 934088 676322 934144
rect 675109 934086 676322 934088
rect 675109 934083 675175 934086
rect 675477 933874 675543 933877
rect 675477 933872 676292 933874
rect 675477 933816 675482 933872
rect 675538 933816 676292 933872
rect 675477 933814 676292 933816
rect 675477 933811 675543 933814
rect 44173 933738 44239 933741
rect 41492 933736 44239 933738
rect 41492 933680 44178 933736
rect 44234 933680 44239 933736
rect 41492 933678 44239 933680
rect 44173 933675 44239 933678
rect 674097 933466 674163 933469
rect 674097 933464 676292 933466
rect 674097 933408 674102 933464
rect 674158 933408 676292 933464
rect 674097 933406 676292 933408
rect 674097 933403 674163 933406
rect 43437 933330 43503 933333
rect 41492 933328 43503 933330
rect 41492 933272 43442 933328
rect 43498 933272 43503 933328
rect 41492 933270 43503 933272
rect 43437 933267 43503 933270
rect 675477 933058 675543 933061
rect 675477 933056 676292 933058
rect 675477 933000 675482 933056
rect 675538 933000 676292 933056
rect 675477 932998 676292 933000
rect 675477 932995 675543 932998
rect 42517 932922 42583 932925
rect 41492 932920 42583 932922
rect 27662 932484 27722 932892
rect 41492 932864 42522 932920
rect 42578 932864 42583 932920
rect 41492 932862 42583 932864
rect 42517 932859 42583 932862
rect 674649 932650 674715 932653
rect 674649 932648 676292 932650
rect 674649 932592 674654 932648
rect 674710 932592 676292 932648
rect 674649 932590 676292 932592
rect 674649 932587 674715 932590
rect 674281 932242 674347 932245
rect 674281 932240 676292 932242
rect 674281 932184 674286 932240
rect 674342 932184 676292 932240
rect 674281 932182 676292 932184
rect 674281 932179 674347 932182
rect 42793 932106 42859 932109
rect 41492 932104 42859 932106
rect 41492 932048 42798 932104
rect 42854 932048 42859 932104
rect 41492 932046 42859 932048
rect 42793 932043 42859 932046
rect 676806 931908 676812 931972
rect 676876 931908 676882 931972
rect 676814 931804 676874 931908
rect 674465 931426 674531 931429
rect 674465 931424 676292 931426
rect 674465 931368 674470 931424
rect 674526 931368 676292 931424
rect 674465 931366 676292 931368
rect 674465 931363 674531 931366
rect 677501 931154 677567 931157
rect 677501 931152 677610 931154
rect 677501 931096 677506 931152
rect 677562 931096 677610 931152
rect 677501 931091 677610 931096
rect 677550 930988 677610 931091
rect 676990 930684 676996 930748
rect 677060 930684 677066 930748
rect 676998 930580 677058 930684
rect 675477 930202 675543 930205
rect 675477 930200 676292 930202
rect 675477 930144 675482 930200
rect 675538 930144 676292 930200
rect 675477 930142 676292 930144
rect 675477 930139 675543 930142
rect 675477 929794 675543 929797
rect 675477 929792 676292 929794
rect 675477 929736 675482 929792
rect 675538 929736 676292 929792
rect 675477 929734 676292 929736
rect 675477 929731 675543 929734
rect 683113 929522 683179 929525
rect 683070 929520 683179 929522
rect 683070 929464 683118 929520
rect 683174 929464 683179 929520
rect 683070 929459 683179 929464
rect 683070 928948 683130 929459
rect 675477 928570 675543 928573
rect 675477 928568 676292 928570
rect 675477 928512 675482 928568
rect 675538 928512 676292 928568
rect 675477 928510 676292 928512
rect 675477 928507 675543 928510
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651557 922722 651623 922725
rect 650164 922720 651623 922722
rect 650164 922664 651562 922720
rect 651618 922664 651623 922720
rect 650164 922662 651623 922664
rect 651557 922659 651623 922662
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 651557 909530 651623 909533
rect 650164 909528 651623 909530
rect 650164 909472 651562 909528
rect 651618 909472 651623 909528
rect 650164 909470 651623 909472
rect 651557 909467 651623 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651557 896202 651623 896205
rect 650164 896200 651623 896202
rect 650164 896144 651562 896200
rect 651618 896144 651623 896200
rect 650164 896142 651623 896144
rect 651557 896139 651623 896142
rect 62113 884778 62179 884781
rect 62113 884776 64492 884778
rect 62113 884720 62118 884776
rect 62174 884720 64492 884776
rect 62113 884718 64492 884720
rect 62113 884715 62179 884718
rect 652385 882874 652451 882877
rect 650164 882872 652451 882874
rect 650164 882816 652390 882872
rect 652446 882816 652451 882872
rect 650164 882814 652451 882816
rect 652385 882811 652451 882814
rect 40677 881922 40743 881925
rect 42425 881922 42491 881925
rect 40677 881920 42491 881922
rect 40677 881864 40682 881920
rect 40738 881864 42430 881920
rect 42486 881864 42491 881920
rect 40677 881862 42491 881864
rect 40677 881859 40743 881862
rect 42425 881859 42491 881862
rect 675753 877162 675819 877165
rect 676070 877162 676076 877164
rect 675753 877160 676076 877162
rect 675753 877104 675758 877160
rect 675814 877104 676076 877160
rect 675753 877102 676076 877104
rect 675753 877099 675819 877102
rect 676070 877100 676076 877102
rect 676140 877100 676146 877164
rect 675293 876482 675359 876485
rect 676806 876482 676812 876484
rect 675293 876480 676812 876482
rect 675293 876424 675298 876480
rect 675354 876424 676812 876480
rect 675293 876422 676812 876424
rect 675293 876419 675359 876422
rect 676806 876420 676812 876422
rect 676876 876420 676882 876484
rect 675385 874036 675451 874037
rect 675334 874034 675340 874036
rect 675294 873974 675340 874034
rect 675404 874032 675451 874036
rect 675446 873976 675451 874032
rect 675334 873972 675340 873974
rect 675404 873972 675451 873976
rect 675385 873971 675451 873972
rect 672625 873626 672691 873629
rect 675385 873626 675451 873629
rect 672625 873624 675451 873626
rect 672625 873568 672630 873624
rect 672686 873568 675390 873624
rect 675446 873568 675451 873624
rect 672625 873566 675451 873568
rect 672625 873563 672691 873566
rect 675385 873563 675451 873566
rect 670417 872266 670483 872269
rect 675385 872266 675451 872269
rect 670417 872264 675451 872266
rect 670417 872208 670422 872264
rect 670478 872208 675390 872264
rect 675446 872208 675451 872264
rect 670417 872206 675451 872208
rect 670417 872203 670483 872206
rect 675385 872203 675451 872206
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 651557 869682 651623 869685
rect 650164 869680 651623 869682
rect 650164 869624 651562 869680
rect 651618 869624 651623 869680
rect 650164 869622 651623 869624
rect 651557 869619 651623 869622
rect 675661 869682 675727 869685
rect 675886 869682 675892 869684
rect 675661 869680 675892 869682
rect 675661 869624 675666 869680
rect 675722 869624 675892 869680
rect 675661 869622 675892 869624
rect 675661 869619 675727 869622
rect 675886 869620 675892 869622
rect 675956 869620 675962 869684
rect 674833 869546 674899 869549
rect 675334 869546 675340 869548
rect 674833 869544 675340 869546
rect 674833 869488 674838 869544
rect 674894 869488 675340 869544
rect 674833 869486 675340 869488
rect 674833 869483 674899 869486
rect 675334 869484 675340 869486
rect 675404 869484 675410 869548
rect 671797 868050 671863 868053
rect 675477 868050 675543 868053
rect 671797 868048 675543 868050
rect 671797 867992 671802 868048
rect 671858 867992 675482 868048
rect 675538 867992 675543 868048
rect 671797 867990 675543 867992
rect 671797 867987 671863 867990
rect 675477 867987 675543 867990
rect 62113 858666 62179 858669
rect 62113 858664 64492 858666
rect 62113 858608 62118 858664
rect 62174 858608 64492 858664
rect 62113 858606 64492 858608
rect 62113 858603 62179 858606
rect 651557 856354 651623 856357
rect 650164 856352 651623 856354
rect 650164 856296 651562 856352
rect 651618 856296 651623 856352
rect 650164 856294 651623 856296
rect 651557 856291 651623 856294
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 651557 843026 651623 843029
rect 650164 843024 651623 843026
rect 650164 842968 651562 843024
rect 651618 842968 651623 843024
rect 650164 842966 651623 842968
rect 651557 842963 651623 842966
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 651557 829834 651623 829837
rect 650164 829832 651623 829834
rect 650164 829776 651562 829832
rect 651618 829776 651623 829832
rect 650164 829774 651623 829776
rect 651557 829771 651623 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 39941 819090 40007 819093
rect 46197 819090 46263 819093
rect 39941 819088 46263 819090
rect 39941 819032 39946 819088
rect 40002 819032 46202 819088
rect 46258 819032 46263 819088
rect 39941 819030 46263 819032
rect 39941 819027 40007 819030
rect 46197 819027 46263 819030
rect 35617 818002 35683 818005
rect 35574 818000 35683 818002
rect 35574 817944 35622 818000
rect 35678 817944 35683 818000
rect 35574 817939 35683 817944
rect 40309 818002 40375 818005
rect 42057 818002 42123 818005
rect 40309 818000 42123 818002
rect 40309 817944 40314 818000
rect 40370 817944 42062 818000
rect 42118 817944 42123 818000
rect 40309 817942 42123 817944
rect 40309 817939 40375 817942
rect 42057 817939 42123 817942
rect 35574 817700 35634 817939
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 35249 816914 35315 816917
rect 35236 816912 35315 816914
rect 35236 816856 35254 816912
rect 35310 816856 35315 816912
rect 35236 816854 35315 816856
rect 35249 816851 35315 816854
rect 35433 816506 35499 816509
rect 651557 816506 651623 816509
rect 35420 816504 35499 816506
rect 35420 816448 35438 816504
rect 35494 816448 35499 816504
rect 35420 816446 35499 816448
rect 650164 816504 651623 816506
rect 650164 816448 651562 816504
rect 651618 816448 651623 816504
rect 650164 816446 651623 816448
rect 35433 816443 35499 816446
rect 651557 816443 651623 816446
rect 35801 816098 35867 816101
rect 35788 816096 35867 816098
rect 35788 816040 35806 816096
rect 35862 816040 35867 816096
rect 35788 816038 35867 816040
rect 35801 816035 35867 816038
rect 35617 815690 35683 815693
rect 35604 815688 35683 815690
rect 35604 815632 35622 815688
rect 35678 815632 35683 815688
rect 35604 815630 35683 815632
rect 35617 815627 35683 815630
rect 35433 815282 35499 815285
rect 35420 815280 35499 815282
rect 35420 815224 35438 815280
rect 35494 815224 35499 815280
rect 35420 815222 35499 815224
rect 35433 815219 35499 815222
rect 35617 814874 35683 814877
rect 35604 814872 35683 814874
rect 35604 814816 35622 814872
rect 35678 814816 35683 814872
rect 35604 814814 35683 814816
rect 35617 814811 35683 814814
rect 41873 814738 41939 814741
rect 42885 814738 42951 814741
rect 41873 814736 42951 814738
rect 41873 814680 41878 814736
rect 41934 814680 42890 814736
rect 42946 814680 42951 814736
rect 41873 814678 42951 814680
rect 41873 814675 41939 814678
rect 42885 814675 42951 814678
rect 35801 814466 35867 814469
rect 35788 814464 35867 814466
rect 35788 814408 35806 814464
rect 35862 814408 35867 814464
rect 35788 814406 35867 814408
rect 35801 814403 35867 814406
rect 41137 814058 41203 814061
rect 41124 814056 41203 814058
rect 41124 814000 41142 814056
rect 41198 814000 41203 814056
rect 41124 813998 41203 814000
rect 41137 813995 41203 813998
rect 43253 813650 43319 813653
rect 41492 813648 43319 813650
rect 41492 813592 43258 813648
rect 43314 813592 43319 813648
rect 41492 813590 43319 813592
rect 43253 813587 43319 813590
rect 42006 813242 42012 813244
rect 41492 813182 42012 813242
rect 42006 813180 42012 813182
rect 42076 813180 42082 813244
rect 41137 812834 41203 812837
rect 41124 812832 41203 812834
rect 41124 812776 41142 812832
rect 41198 812776 41203 812832
rect 41124 812774 41203 812776
rect 41137 812771 41203 812774
rect 41781 812834 41847 812837
rect 44449 812834 44515 812837
rect 41781 812832 44515 812834
rect 41781 812776 41786 812832
rect 41842 812776 44454 812832
rect 44510 812776 44515 812832
rect 41781 812774 44515 812776
rect 41781 812771 41847 812774
rect 44449 812771 44515 812774
rect 35157 812426 35223 812429
rect 35157 812424 35236 812426
rect 35157 812368 35162 812424
rect 35218 812368 35236 812424
rect 35157 812366 35236 812368
rect 35157 812363 35223 812366
rect 40953 812018 41019 812021
rect 40940 812016 41019 812018
rect 40940 811960 40958 812016
rect 41014 811960 41019 812016
rect 40940 811958 41019 811960
rect 40953 811955 41019 811958
rect 41321 811610 41387 811613
rect 41308 811608 41387 811610
rect 41308 811552 41326 811608
rect 41382 811552 41387 811608
rect 41308 811550 41387 811552
rect 41321 811547 41387 811550
rect 32397 811202 32463 811205
rect 32397 811200 32476 811202
rect 32397 811144 32402 811200
rect 32458 811144 32476 811200
rect 32397 811142 32476 811144
rect 32397 811139 32463 811142
rect 40542 810762 40602 810764
rect 40534 810698 40540 810762
rect 40604 810698 40610 810762
rect 41965 810386 42031 810389
rect 41492 810384 42031 810386
rect 41492 810328 41970 810384
rect 42026 810328 42031 810384
rect 41492 810326 42031 810328
rect 41965 810323 42031 810326
rect 31661 809978 31727 809981
rect 31661 809976 31740 809978
rect 31661 809920 31666 809976
rect 31722 809920 31740 809976
rect 31661 809918 31740 809920
rect 31661 809915 31727 809918
rect 33777 809570 33843 809573
rect 33764 809568 33843 809570
rect 33764 809512 33782 809568
rect 33838 809512 33843 809568
rect 33764 809510 33843 809512
rect 33777 809507 33843 809510
rect 36537 809162 36603 809165
rect 36524 809160 36603 809162
rect 36524 809104 36542 809160
rect 36598 809104 36603 809160
rect 36524 809102 36603 809104
rect 36537 809099 36603 809102
rect 43069 808754 43135 808757
rect 41492 808752 43135 808754
rect 41492 808696 43074 808752
rect 43130 808696 43135 808752
rect 41492 808694 43135 808696
rect 43069 808691 43135 808694
rect 42006 808346 42012 808348
rect 41492 808286 42012 808346
rect 42006 808284 42012 808286
rect 42076 808284 42082 808348
rect 44633 807938 44699 807941
rect 41492 807936 44699 807938
rect 41492 807880 44638 807936
rect 44694 807880 44699 807936
rect 41492 807878 44699 807880
rect 44633 807875 44699 807878
rect 41462 807360 41522 807500
rect 41462 807300 41844 807360
rect 41784 807258 41844 807300
rect 43621 807258 43687 807261
rect 41784 807256 43687 807258
rect 41784 807200 43626 807256
rect 43682 807200 43687 807256
rect 41784 807198 43687 807200
rect 43621 807195 43687 807198
rect 41462 806714 41522 807092
rect 42057 806714 42123 806717
rect 41462 806712 42123 806714
rect 41462 806684 42062 806712
rect 41492 806656 42062 806684
rect 42118 806656 42123 806712
rect 41492 806654 42123 806656
rect 42057 806651 42123 806654
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 46197 806306 46263 806309
rect 41492 806304 46263 806306
rect 41492 806248 46202 806304
rect 46258 806248 46263 806304
rect 41492 806246 46263 806248
rect 46197 806243 46263 806246
rect 40718 805292 40724 805356
rect 40788 805354 40794 805356
rect 41781 805354 41847 805357
rect 40788 805352 41847 805354
rect 40788 805296 41786 805352
rect 41842 805296 41847 805352
rect 40788 805294 41847 805296
rect 40788 805292 40794 805294
rect 41781 805291 41847 805294
rect 40902 805020 40908 805084
rect 40972 805082 40978 805084
rect 42006 805082 42012 805084
rect 40972 805022 42012 805082
rect 40972 805020 40978 805022
rect 42006 805020 42012 805022
rect 42076 805020 42082 805084
rect 40953 804810 41019 804813
rect 41638 804810 41644 804812
rect 40953 804808 41644 804810
rect 40953 804752 40958 804808
rect 41014 804752 41644 804808
rect 40953 804750 41644 804752
rect 40953 804747 41019 804750
rect 41638 804748 41644 804750
rect 41708 804748 41714 804812
rect 35157 803858 35223 803861
rect 41822 803858 41828 803860
rect 35157 803856 41828 803858
rect 35157 803800 35162 803856
rect 35218 803800 41828 803856
rect 35157 803798 41828 803800
rect 35157 803795 35223 803798
rect 41822 803796 41828 803798
rect 41892 803796 41898 803860
rect 651557 803314 651623 803317
rect 650164 803312 651623 803314
rect 650164 803256 651562 803312
rect 651618 803256 651623 803312
rect 650164 803254 651623 803256
rect 651557 803251 651623 803254
rect 39757 801954 39823 801957
rect 42609 801954 42675 801957
rect 39757 801952 42675 801954
rect 39757 801896 39762 801952
rect 39818 801896 42614 801952
rect 42670 801896 42675 801952
rect 39757 801894 42675 801896
rect 39757 801891 39823 801894
rect 42609 801891 42675 801894
rect 42333 801140 42399 801141
rect 42333 801136 42380 801140
rect 42444 801138 42450 801140
rect 42333 801080 42338 801136
rect 42333 801076 42380 801080
rect 42444 801078 42490 801138
rect 42444 801076 42450 801078
rect 42333 801075 42399 801076
rect 39849 801002 39915 801005
rect 41086 801002 41092 801004
rect 39849 801000 41092 801002
rect 39849 800944 39854 801000
rect 39910 800944 41092 801000
rect 39849 800942 41092 800944
rect 39849 800939 39915 800942
rect 41086 800940 41092 800942
rect 41156 800940 41162 801004
rect 41229 800866 41295 800869
rect 42333 800866 42399 800869
rect 41229 800864 42399 800866
rect 41229 800808 41234 800864
rect 41290 800808 42338 800864
rect 42394 800808 42399 800864
rect 41229 800806 42399 800808
rect 41229 800803 41295 800806
rect 42333 800803 42399 800806
rect 40033 800730 40099 800733
rect 40350 800730 40356 800732
rect 40033 800728 40356 800730
rect 40033 800672 40038 800728
rect 40094 800672 40356 800728
rect 40033 800670 40356 800672
rect 40033 800667 40099 800670
rect 40350 800668 40356 800670
rect 40420 800668 40426 800732
rect 41781 800322 41847 800325
rect 41781 800320 41890 800322
rect 41781 800264 41786 800320
rect 41842 800264 41890 800320
rect 41781 800259 41890 800264
rect 41830 799917 41890 800259
rect 41781 799912 41890 799917
rect 41781 799856 41786 799912
rect 41842 799856 41890 799912
rect 41781 799854 41890 799856
rect 41781 799851 41847 799854
rect 42149 797330 42215 797333
rect 43621 797330 43687 797333
rect 42149 797328 43687 797330
rect 42149 797272 42154 797328
rect 42210 797272 43626 797328
rect 43682 797272 43687 797328
rect 42149 797270 43687 797272
rect 42149 797267 42215 797270
rect 43621 797267 43687 797270
rect 40350 796180 40356 796244
rect 40420 796242 40426 796244
rect 41781 796242 41847 796245
rect 40420 796240 41847 796242
rect 40420 796184 41786 796240
rect 41842 796184 41847 796240
rect 40420 796182 41847 796184
rect 40420 796180 40426 796182
rect 41781 796179 41847 796182
rect 42057 795018 42123 795021
rect 44633 795018 44699 795021
rect 42057 795016 44699 795018
rect 42057 794960 42062 795016
rect 42118 794960 44638 795016
rect 44694 794960 44699 795016
rect 42057 794958 44699 794960
rect 42057 794955 42123 794958
rect 44633 794955 44699 794958
rect 41086 794412 41092 794476
rect 41156 794474 41162 794476
rect 41781 794474 41847 794477
rect 41156 794472 41847 794474
rect 41156 794416 41786 794472
rect 41842 794416 41847 794472
rect 41156 794414 41847 794416
rect 41156 794412 41162 794414
rect 41781 794411 41847 794414
rect 62113 793658 62179 793661
rect 62113 793656 64492 793658
rect 62113 793600 62118 793656
rect 62174 793600 64492 793656
rect 62113 793598 64492 793600
rect 62113 793595 62179 793598
rect 40902 793460 40908 793524
rect 40972 793522 40978 793524
rect 41781 793522 41847 793525
rect 40972 793520 41847 793522
rect 40972 793464 41786 793520
rect 41842 793464 41847 793520
rect 40972 793462 41847 793464
rect 40972 793460 40978 793462
rect 41781 793459 41847 793462
rect 42149 792978 42215 792981
rect 42374 792978 42380 792980
rect 42149 792976 42380 792978
rect 42149 792920 42154 792976
rect 42210 792920 42380 792976
rect 42149 792918 42380 792920
rect 42149 792915 42215 792918
rect 42374 792916 42380 792918
rect 42444 792916 42450 792980
rect 40718 791964 40724 792028
rect 40788 792026 40794 792028
rect 42425 792026 42491 792029
rect 40788 792024 42491 792026
rect 40788 791968 42430 792024
rect 42486 791968 42491 792024
rect 40788 791966 42491 791968
rect 40788 791964 40794 791966
rect 42425 791963 42491 791966
rect 40534 790060 40540 790124
rect 40604 790122 40610 790124
rect 42609 790122 42675 790125
rect 40604 790120 42675 790122
rect 40604 790064 42614 790120
rect 42670 790064 42675 790120
rect 40604 790062 42675 790064
rect 40604 790060 40610 790062
rect 42609 790059 42675 790062
rect 651557 789986 651623 789989
rect 650164 789984 651623 789986
rect 650164 789928 651562 789984
rect 651618 789928 651623 789984
rect 650164 789926 651623 789928
rect 651557 789923 651623 789926
rect 41638 789108 41644 789172
rect 41708 789170 41714 789172
rect 42333 789170 42399 789173
rect 41708 789168 42399 789170
rect 41708 789112 42338 789168
rect 42394 789112 42399 789168
rect 41708 789110 42399 789112
rect 41708 789108 41714 789110
rect 42333 789107 42399 789110
rect 41822 788428 41828 788492
rect 41892 788490 41898 788492
rect 41892 788430 42626 788490
rect 41892 788428 41898 788430
rect 41454 788156 41460 788220
rect 41524 788218 41530 788220
rect 42241 788218 42307 788221
rect 41524 788216 42307 788218
rect 41524 788160 42246 788216
rect 42302 788160 42307 788216
rect 41524 788158 42307 788160
rect 41524 788156 41530 788158
rect 42241 788155 42307 788158
rect 42566 787949 42626 788430
rect 42517 787944 42626 787949
rect 42517 787888 42522 787944
rect 42578 787888 42626 787944
rect 42517 787886 42626 787888
rect 42517 787883 42583 787886
rect 674230 784212 674236 784276
rect 674300 784274 674306 784276
rect 675293 784274 675359 784277
rect 674300 784272 675359 784274
rect 674300 784216 675298 784272
rect 675354 784216 675359 784272
rect 674300 784214 675359 784216
rect 674300 784212 674306 784214
rect 675293 784211 675359 784214
rect 674598 783940 674604 784004
rect 674668 784002 674674 784004
rect 675109 784002 675175 784005
rect 674668 784000 675175 784002
rect 674668 783944 675114 784000
rect 675170 783944 675175 784000
rect 674668 783942 675175 783944
rect 674668 783940 674674 783942
rect 675109 783939 675175 783942
rect 62113 780466 62179 780469
rect 62113 780464 64492 780466
rect 62113 780408 62118 780464
rect 62174 780408 64492 780464
rect 62113 780406 64492 780408
rect 62113 780403 62179 780406
rect 651557 776658 651623 776661
rect 650164 776656 651623 776658
rect 650164 776600 651562 776656
rect 651618 776600 651623 776656
rect 650164 776598 651623 776600
rect 651557 776595 651623 776598
rect 39757 775298 39823 775301
rect 44817 775298 44883 775301
rect 39757 775296 44883 775298
rect 39757 775240 39762 775296
rect 39818 775240 44822 775296
rect 44878 775240 44883 775296
rect 39757 775238 44883 775240
rect 39757 775235 39823 775238
rect 44817 775235 44883 775238
rect 670049 775026 670115 775029
rect 675477 775026 675543 775029
rect 670049 775024 675543 775026
rect 670049 774968 670054 775024
rect 670110 774968 675482 775024
rect 675538 774968 675543 775024
rect 670049 774966 675543 774968
rect 670049 774963 670115 774966
rect 675477 774963 675543 774966
rect 35758 774349 35818 774452
rect 35758 774344 35867 774349
rect 35758 774288 35806 774344
rect 35862 774288 35867 774344
rect 35758 774286 35867 774288
rect 35801 774283 35867 774286
rect 35758 773941 35818 774044
rect 35758 773936 35867 773941
rect 35758 773880 35806 773936
rect 35862 773880 35867 773936
rect 35758 773878 35867 773880
rect 35801 773875 35867 773878
rect 668577 773802 668643 773805
rect 675477 773802 675543 773805
rect 668577 773800 675543 773802
rect 668577 773744 668582 773800
rect 668638 773744 675482 773800
rect 675538 773744 675543 773800
rect 668577 773742 675543 773744
rect 668577 773739 668643 773742
rect 675477 773739 675543 773742
rect 35390 773533 35450 773636
rect 35341 773528 35450 773533
rect 35341 773472 35346 773528
rect 35402 773472 35450 773528
rect 35341 773470 35450 773472
rect 35341 773467 35407 773470
rect 35758 773125 35818 773228
rect 35525 773122 35591 773125
rect 35525 773120 35634 773122
rect 35525 773064 35530 773120
rect 35586 773064 35634 773120
rect 35525 773059 35634 773064
rect 35758 773120 35867 773125
rect 35758 773064 35806 773120
rect 35862 773064 35867 773120
rect 35758 773062 35867 773064
rect 35801 773059 35867 773062
rect 40861 773122 40927 773125
rect 43069 773122 43135 773125
rect 40861 773120 43135 773122
rect 40861 773064 40866 773120
rect 40922 773064 43074 773120
rect 43130 773064 43135 773120
rect 40861 773062 43135 773064
rect 40861 773059 40927 773062
rect 43069 773059 43135 773062
rect 35574 772820 35634 773059
rect 676070 772652 676076 772716
rect 676140 772714 676146 772716
rect 679617 772714 679683 772717
rect 676140 772712 679683 772714
rect 676140 772656 679622 772712
rect 679678 772656 679683 772712
rect 676140 772654 679683 772656
rect 676140 772652 676146 772654
rect 679617 772651 679683 772654
rect 674649 772442 674715 772445
rect 676029 772442 676095 772445
rect 674649 772440 676095 772442
rect 35390 772309 35450 772412
rect 674649 772384 674654 772440
rect 674710 772384 676034 772440
rect 676090 772384 676095 772440
rect 674649 772382 676095 772384
rect 674649 772379 674715 772382
rect 676029 772379 676095 772382
rect 35341 772304 35450 772309
rect 35341 772248 35346 772304
rect 35402 772248 35450 772304
rect 35341 772246 35450 772248
rect 35341 772243 35407 772246
rect 674649 772170 674715 772173
rect 675845 772170 675911 772173
rect 674649 772168 675911 772170
rect 674649 772112 674654 772168
rect 674710 772112 675850 772168
rect 675906 772112 675911 772168
rect 674649 772110 675911 772112
rect 674649 772107 674715 772110
rect 675845 772107 675911 772110
rect 35574 771901 35634 772004
rect 35525 771896 35634 771901
rect 35801 771898 35867 771901
rect 35525 771840 35530 771896
rect 35586 771840 35634 771896
rect 35525 771838 35634 771840
rect 35758 771896 35867 771898
rect 35758 771840 35806 771896
rect 35862 771840 35867 771896
rect 35525 771835 35591 771838
rect 35758 771835 35867 771840
rect 35758 771596 35818 771835
rect 35758 771085 35818 771188
rect 35758 771080 35867 771085
rect 35758 771024 35806 771080
rect 35862 771024 35867 771080
rect 35758 771022 35867 771024
rect 35801 771019 35867 771022
rect 35574 770677 35634 770780
rect 35574 770672 35683 770677
rect 35574 770616 35622 770672
rect 35678 770616 35683 770672
rect 35574 770614 35683 770616
rect 35617 770611 35683 770614
rect 39849 770674 39915 770677
rect 42885 770674 42951 770677
rect 39849 770672 42951 770674
rect 39849 770616 39854 770672
rect 39910 770616 42890 770672
rect 42946 770616 42951 770672
rect 39849 770614 42951 770616
rect 39849 770611 39915 770614
rect 42885 770611 42951 770614
rect 675109 770674 675175 770677
rect 675845 770674 675911 770677
rect 675109 770672 675911 770674
rect 675109 770616 675114 770672
rect 675170 770616 675850 770672
rect 675906 770616 675911 770672
rect 675109 770614 675911 770616
rect 675109 770611 675175 770614
rect 675845 770611 675911 770614
rect 35758 770269 35818 770372
rect 35758 770264 35867 770269
rect 35758 770208 35806 770264
rect 35862 770208 35867 770264
rect 35758 770206 35867 770208
rect 35801 770203 35867 770206
rect 39849 770266 39915 770269
rect 44265 770266 44331 770269
rect 39849 770264 44331 770266
rect 39849 770208 39854 770264
rect 39910 770208 44270 770264
rect 44326 770208 44331 770264
rect 39849 770206 44331 770208
rect 39849 770203 39915 770206
rect 44265 770203 44331 770206
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35574 769453 35634 769556
rect 35574 769448 35683 769453
rect 35574 769392 35622 769448
rect 35678 769392 35683 769448
rect 35574 769390 35683 769392
rect 35617 769387 35683 769390
rect 35758 769045 35818 769148
rect 35758 769040 35867 769045
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35758 768982 35867 768984
rect 35801 768979 35867 768982
rect 42517 768770 42583 768773
rect 41492 768768 42583 768770
rect 41492 768712 42522 768768
rect 42578 768712 42583 768768
rect 41492 768710 42583 768712
rect 42517 768707 42583 768710
rect 675886 768708 675892 768772
rect 675956 768770 675962 768772
rect 682377 768770 682443 768773
rect 675956 768768 682443 768770
rect 675956 768712 682382 768768
rect 682438 768712 682443 768768
rect 675956 768710 682443 768712
rect 675956 768708 675962 768710
rect 682377 768707 682443 768710
rect 35758 768229 35818 768332
rect 35758 768224 35867 768229
rect 35758 768168 35806 768224
rect 35862 768168 35867 768224
rect 35758 768166 35867 768168
rect 35801 768163 35867 768166
rect 35574 767821 35634 767924
rect 35574 767816 35683 767821
rect 35574 767760 35622 767816
rect 35678 767760 35683 767816
rect 35574 767758 35683 767760
rect 35617 767755 35683 767758
rect 32446 767413 32506 767516
rect 32397 767408 32506 767413
rect 32397 767352 32402 767408
rect 32458 767352 32506 767408
rect 32397 767350 32506 767352
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 32397 767347 32463 767350
rect 62113 767347 62179 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 35758 766597 35818 766700
rect 35758 766592 35867 766597
rect 35758 766536 35806 766592
rect 35862 766536 35867 766592
rect 35758 766534 35867 766536
rect 35801 766531 35867 766534
rect 674925 766594 674991 766597
rect 675702 766594 675708 766596
rect 674925 766592 675708 766594
rect 674925 766536 674930 766592
rect 674986 766536 675708 766592
rect 674925 766534 675708 766536
rect 674925 766531 674991 766534
rect 675702 766532 675708 766534
rect 675772 766532 675778 766596
rect 35758 766189 35818 766292
rect 35758 766184 35867 766189
rect 35758 766128 35806 766184
rect 35862 766128 35867 766184
rect 35758 766126 35867 766128
rect 35801 766123 35867 766126
rect 40910 765780 40970 765884
rect 40902 765716 40908 765780
rect 40972 765716 40978 765780
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40726 764964 40786 765068
rect 40718 764900 40724 764964
rect 40788 764900 40794 764964
rect 35758 764557 35818 764660
rect 35758 764552 35867 764557
rect 35758 764496 35806 764552
rect 35862 764496 35867 764552
rect 35758 764494 35867 764496
rect 35801 764491 35867 764494
rect 39757 764554 39823 764557
rect 43253 764554 43319 764557
rect 39757 764552 43319 764554
rect 39757 764496 39762 764552
rect 39818 764496 43258 764552
rect 43314 764496 43319 764552
rect 39757 764494 43319 764496
rect 39757 764491 39823 764494
rect 43253 764491 43319 764494
rect 35574 764149 35634 764252
rect 35574 764144 35683 764149
rect 35574 764088 35622 764144
rect 35678 764088 35683 764144
rect 35574 764086 35683 764088
rect 35617 764083 35683 764086
rect 35758 763333 35818 763844
rect 39113 763738 39179 763741
rect 45001 763738 45067 763741
rect 39113 763736 45067 763738
rect 39113 763680 39118 763736
rect 39174 763680 45006 763736
rect 45062 763680 45067 763736
rect 39113 763678 45067 763680
rect 39113 763675 39179 763678
rect 45001 763675 45067 763678
rect 35758 763328 35867 763333
rect 35758 763272 35806 763328
rect 35862 763272 35867 763328
rect 35758 763270 35867 763272
rect 35801 763267 35867 763270
rect 41689 763330 41755 763333
rect 47577 763330 47643 763333
rect 651557 763330 651623 763333
rect 41689 763328 47643 763330
rect 41689 763272 41694 763328
rect 41750 763272 47582 763328
rect 47638 763272 47643 763328
rect 41689 763270 47643 763272
rect 650164 763328 651623 763330
rect 650164 763272 651562 763328
rect 651618 763272 651623 763328
rect 650164 763270 651623 763272
rect 41689 763267 41755 763270
rect 47577 763267 47643 763270
rect 651557 763267 651623 763270
rect 35758 762925 35818 763028
rect 35758 762920 35867 762925
rect 35758 762864 35806 762920
rect 35862 762864 35867 762920
rect 35758 762862 35867 762864
rect 35801 762859 35867 762862
rect 675477 761562 675543 761565
rect 675477 761560 676292 761562
rect 675477 761504 675482 761560
rect 675538 761504 676292 761560
rect 675477 761502 676292 761504
rect 675477 761499 675543 761502
rect 675293 761154 675359 761157
rect 675293 761152 676292 761154
rect 675293 761096 675298 761152
rect 675354 761096 676292 761152
rect 675293 761094 676292 761096
rect 675293 761091 675359 761094
rect 675477 760746 675543 760749
rect 675477 760744 676292 760746
rect 675477 760688 675482 760744
rect 675538 760688 676292 760744
rect 675477 760686 676292 760688
rect 675477 760683 675543 760686
rect 675293 760338 675359 760341
rect 675293 760336 676292 760338
rect 675293 760280 675298 760336
rect 675354 760280 676292 760336
rect 675293 760278 676292 760280
rect 675293 760275 675359 760278
rect 675477 759930 675543 759933
rect 675477 759928 676292 759930
rect 675477 759872 675482 759928
rect 675538 759872 676292 759928
rect 675477 759870 676292 759872
rect 675477 759867 675543 759870
rect 32397 759658 32463 759661
rect 41638 759658 41644 759660
rect 32397 759656 41644 759658
rect 32397 759600 32402 759656
rect 32458 759600 41644 759656
rect 32397 759598 41644 759600
rect 32397 759595 32463 759598
rect 41638 759596 41644 759598
rect 41708 759596 41714 759660
rect 675477 759522 675543 759525
rect 675477 759520 676292 759522
rect 675477 759464 675482 759520
rect 675538 759464 676292 759520
rect 675477 759462 676292 759464
rect 675477 759459 675543 759462
rect 675477 759114 675543 759117
rect 675477 759112 676292 759114
rect 675477 759056 675482 759112
rect 675538 759056 676292 759112
rect 675477 759054 676292 759056
rect 675477 759051 675543 759054
rect 675477 758706 675543 758709
rect 675477 758704 676292 758706
rect 675477 758648 675482 758704
rect 675538 758648 676292 758704
rect 675477 758646 676292 758648
rect 675477 758643 675543 758646
rect 42241 758436 42307 758437
rect 42190 758434 42196 758436
rect 42150 758374 42196 758434
rect 42260 758432 42307 758436
rect 42302 758376 42307 758432
rect 42190 758372 42196 758374
rect 42260 758372 42307 758376
rect 42241 758371 42307 758372
rect 675477 758298 675543 758301
rect 675477 758296 676292 758298
rect 675477 758240 675482 758296
rect 675538 758240 676292 758296
rect 675477 758238 676292 758240
rect 675477 758235 675543 758238
rect 40217 758162 40283 758165
rect 44817 758162 44883 758165
rect 40217 758160 44883 758162
rect 40217 758104 40222 758160
rect 40278 758104 44822 758160
rect 44878 758104 44883 758160
rect 40217 758102 44883 758104
rect 40217 758099 40283 758102
rect 44817 758099 44883 758102
rect 41965 757890 42031 757893
rect 42425 757890 42491 757893
rect 41965 757888 42491 757890
rect 41965 757832 41970 757888
rect 42026 757832 42430 757888
rect 42486 757832 42491 757888
rect 41965 757830 42491 757832
rect 41965 757827 42031 757830
rect 42425 757827 42491 757830
rect 675477 757890 675543 757893
rect 675477 757888 676292 757890
rect 675477 757832 675482 757888
rect 675538 757832 676292 757888
rect 675477 757830 676292 757832
rect 675477 757827 675543 757830
rect 39297 757754 39363 757757
rect 41822 757754 41828 757756
rect 39297 757752 41828 757754
rect 39297 757696 39302 757752
rect 39358 757696 41828 757752
rect 39297 757694 41828 757696
rect 39297 757691 39363 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 39941 757482 40007 757485
rect 42241 757482 42307 757485
rect 39941 757480 42307 757482
rect 39941 757424 39946 757480
rect 40002 757424 42246 757480
rect 42302 757424 42307 757480
rect 39941 757422 42307 757424
rect 39941 757419 40007 757422
rect 42241 757419 42307 757422
rect 675477 757482 675543 757485
rect 675477 757480 676292 757482
rect 675477 757424 675482 757480
rect 675538 757424 676292 757480
rect 675477 757422 676292 757424
rect 675477 757419 675543 757422
rect 41781 757074 41847 757077
rect 42006 757074 42012 757076
rect 41781 757072 42012 757074
rect 41781 757016 41786 757072
rect 41842 757016 42012 757072
rect 41781 757014 42012 757016
rect 41781 757011 41847 757014
rect 42006 757012 42012 757014
rect 42076 757012 42082 757076
rect 675886 757012 675892 757076
rect 675956 757074 675962 757076
rect 675956 757014 676292 757074
rect 675956 757012 675962 757014
rect 684125 756666 684191 756669
rect 684125 756664 684204 756666
rect 684125 756608 684130 756664
rect 684186 756608 684204 756664
rect 684125 756606 684204 756608
rect 684125 756603 684191 756606
rect 679617 756258 679683 756261
rect 679604 756256 679683 756258
rect 679604 756200 679622 756256
rect 679678 756200 679683 756256
rect 679604 756198 679683 756200
rect 679617 756195 679683 756198
rect 675845 755850 675911 755853
rect 675845 755848 676292 755850
rect 675845 755792 675850 755848
rect 675906 755792 676292 755848
rect 675845 755790 676292 755792
rect 675845 755787 675911 755790
rect 41965 755444 42031 755445
rect 41965 755440 42012 755444
rect 42076 755442 42082 755444
rect 682377 755442 682443 755445
rect 41965 755384 41970 755440
rect 41965 755380 42012 755384
rect 42076 755382 42122 755442
rect 682364 755440 682443 755442
rect 682364 755384 682382 755440
rect 682438 755384 682443 755440
rect 682364 755382 682443 755384
rect 42076 755380 42082 755382
rect 41965 755379 42031 755380
rect 682377 755379 682443 755382
rect 675477 755034 675543 755037
rect 675477 755032 676292 755034
rect 675477 754976 675482 755032
rect 675538 754976 676292 755032
rect 675477 754974 676292 754976
rect 675477 754971 675543 754974
rect 42149 754900 42215 754901
rect 42149 754898 42196 754900
rect 42104 754896 42196 754898
rect 42104 754840 42154 754896
rect 42104 754838 42196 754840
rect 42149 754836 42196 754838
rect 42260 754836 42266 754900
rect 42149 754835 42215 754836
rect 675477 754626 675543 754629
rect 675477 754624 676292 754626
rect 675477 754568 675482 754624
rect 675538 754568 676292 754624
rect 675477 754566 676292 754568
rect 675477 754563 675543 754566
rect 62113 754354 62179 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 62113 754291 62179 754294
rect 675477 754218 675543 754221
rect 675477 754216 676292 754218
rect 675477 754160 675482 754216
rect 675538 754160 676292 754216
rect 675477 754158 676292 754160
rect 675477 754155 675543 754158
rect 42057 754082 42123 754085
rect 43437 754082 43503 754085
rect 42057 754080 43503 754082
rect 42057 754024 42062 754080
rect 42118 754024 43442 754080
rect 43498 754024 43503 754080
rect 42057 754022 43503 754024
rect 42057 754019 42123 754022
rect 43437 754019 43503 754022
rect 675109 753810 675175 753813
rect 675109 753808 676292 753810
rect 675109 753752 675114 753808
rect 675170 753752 676292 753808
rect 675109 753750 676292 753752
rect 675109 753747 675175 753750
rect 675477 753402 675543 753405
rect 675477 753400 676292 753402
rect 675477 753344 675482 753400
rect 675538 753344 676292 753400
rect 675477 753342 676292 753344
rect 675477 753339 675543 753342
rect 669221 752994 669287 752997
rect 675845 752994 675911 752997
rect 683297 752994 683363 752997
rect 669221 752992 675911 752994
rect 669221 752936 669226 752992
rect 669282 752936 675850 752992
rect 675906 752936 675911 752992
rect 669221 752934 675911 752936
rect 683284 752992 683363 752994
rect 683284 752936 683302 752992
rect 683358 752936 683363 752992
rect 683284 752934 683363 752936
rect 669221 752931 669287 752934
rect 675845 752931 675911 752934
rect 683297 752931 683363 752934
rect 670417 752722 670483 752725
rect 670417 752720 676230 752722
rect 670417 752664 670422 752720
rect 670478 752664 676230 752720
rect 670417 752662 676230 752664
rect 670417 752659 670483 752662
rect 676170 752586 676230 752662
rect 676170 752526 676292 752586
rect 674925 752450 674991 752453
rect 675886 752450 675892 752452
rect 674925 752448 675892 752450
rect 674925 752392 674930 752448
rect 674986 752392 675892 752448
rect 674925 752390 675892 752392
rect 674925 752387 674991 752390
rect 675886 752388 675892 752390
rect 675956 752388 675962 752452
rect 40718 752116 40724 752180
rect 40788 752178 40794 752180
rect 42241 752178 42307 752181
rect 40788 752176 42307 752178
rect 40788 752120 42246 752176
rect 42302 752120 42307 752176
rect 40788 752118 42307 752120
rect 40788 752116 40794 752118
rect 42241 752115 42307 752118
rect 675477 752178 675543 752181
rect 675477 752176 676292 752178
rect 675477 752120 675482 752176
rect 675538 752120 676292 752176
rect 675477 752118 676292 752120
rect 675477 752115 675543 752118
rect 42057 751770 42123 751773
rect 43437 751770 43503 751773
rect 42057 751768 43503 751770
rect 42057 751712 42062 751768
rect 42118 751712 43442 751768
rect 43498 751712 43503 751768
rect 42057 751710 43503 751712
rect 42057 751707 42123 751710
rect 43437 751707 43503 751710
rect 675477 751770 675543 751773
rect 675477 751768 676292 751770
rect 675477 751712 675482 751768
rect 675538 751712 676292 751768
rect 675477 751710 676292 751712
rect 675477 751707 675543 751710
rect 672349 751362 672415 751365
rect 672349 751360 676292 751362
rect 672349 751304 672354 751360
rect 672410 751304 676292 751360
rect 672349 751302 676292 751304
rect 672349 751299 672415 751302
rect 40902 751028 40908 751092
rect 40972 751090 40978 751092
rect 41781 751090 41847 751093
rect 40972 751088 41847 751090
rect 40972 751032 41786 751088
rect 41842 751032 41847 751088
rect 40972 751030 41847 751032
rect 40972 751028 40978 751030
rect 41781 751027 41847 751030
rect 683070 750753 683130 750924
rect 683070 750748 683179 750753
rect 683070 750692 683118 750748
rect 683174 750692 683179 750748
rect 683070 750687 683179 750692
rect 683070 750516 683130 750687
rect 651557 750138 651623 750141
rect 650164 750136 651623 750138
rect 650164 750080 651562 750136
rect 651618 750080 651623 750136
rect 650164 750078 651623 750080
rect 651557 750075 651623 750078
rect 675477 750138 675543 750141
rect 675477 750136 676292 750138
rect 675477 750080 675482 750136
rect 675538 750080 676292 750136
rect 675477 750078 676292 750080
rect 675477 750075 675543 750078
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 42241 749458 42307 749461
rect 40604 749456 42307 749458
rect 40604 749400 42246 749456
rect 42302 749400 42307 749456
rect 40604 749398 42307 749400
rect 40604 749396 40610 749398
rect 42241 749395 42307 749398
rect 41454 746540 41460 746604
rect 41524 746602 41530 746604
rect 42241 746602 42307 746605
rect 41524 746600 42307 746602
rect 41524 746544 42246 746600
rect 42302 746544 42307 746600
rect 41524 746542 42307 746544
rect 41524 746540 41530 746542
rect 42241 746539 42307 746542
rect 41638 746268 41644 746332
rect 41708 746330 41714 746332
rect 42425 746330 42491 746333
rect 41708 746328 42491 746330
rect 41708 746272 42430 746328
rect 42486 746272 42491 746328
rect 41708 746270 42491 746272
rect 41708 746268 41714 746270
rect 42425 746267 42491 746270
rect 42057 746058 42123 746061
rect 42609 746058 42675 746061
rect 42057 746056 42675 746058
rect 42057 746000 42062 746056
rect 42118 746000 42614 746056
rect 42670 746000 42675 746056
rect 42057 745998 42675 746000
rect 42057 745995 42123 745998
rect 42609 745995 42675 745998
rect 42057 745514 42123 745517
rect 42701 745514 42767 745517
rect 42057 745512 42767 745514
rect 42057 745456 42062 745512
rect 42118 745456 42706 745512
rect 42762 745456 42767 745512
rect 42057 745454 42767 745456
rect 42057 745451 42123 745454
rect 42701 745451 42767 745454
rect 41822 745044 41828 745108
rect 41892 745106 41898 745108
rect 42609 745106 42675 745109
rect 41892 745104 42675 745106
rect 41892 745048 42614 745104
rect 42670 745048 42675 745104
rect 41892 745046 42675 745048
rect 41892 745044 41898 745046
rect 42609 745043 42675 745046
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 674414 738108 674420 738172
rect 674484 738170 674490 738172
rect 675109 738170 675175 738173
rect 674484 738168 675175 738170
rect 674484 738112 675114 738168
rect 675170 738112 675175 738168
rect 674484 738110 675175 738112
rect 674484 738108 674490 738110
rect 675109 738107 675175 738110
rect 651557 736810 651623 736813
rect 650164 736808 651623 736810
rect 650164 736752 651562 736808
rect 651618 736752 651623 736808
rect 650164 736750 651623 736752
rect 651557 736747 651623 736750
rect 672533 734226 672599 734229
rect 675477 734226 675543 734229
rect 672533 734224 675543 734226
rect 672533 734168 672538 734224
rect 672594 734168 675482 734224
rect 675538 734168 675543 734224
rect 672533 734166 675543 734168
rect 672533 734163 672599 734166
rect 675477 734163 675543 734166
rect 671705 733682 671771 733685
rect 675477 733682 675543 733685
rect 671705 733680 675543 733682
rect 671705 733624 671710 733680
rect 671766 733624 675482 733680
rect 675538 733624 675543 733680
rect 671705 733622 675543 733624
rect 671705 733619 671771 733622
rect 675477 733619 675543 733622
rect 675109 733002 675175 733005
rect 677174 733002 677180 733004
rect 675109 733000 677180 733002
rect 675109 732944 675114 733000
rect 675170 732944 677180 733000
rect 675109 732942 677180 732944
rect 675109 732939 675175 732942
rect 677174 732940 677180 732942
rect 677244 732940 677250 733004
rect 673453 732730 673519 732733
rect 675477 732730 675543 732733
rect 673453 732728 675543 732730
rect 673453 732672 673458 732728
rect 673514 732672 675482 732728
rect 675538 732672 675543 732728
rect 673453 732670 675543 732672
rect 673453 732667 673519 732670
rect 675477 732667 675543 732670
rect 47761 731370 47827 731373
rect 41492 731368 47827 731370
rect 41492 731312 47766 731368
rect 47822 731312 47827 731368
rect 41492 731310 47827 731312
rect 47761 731307 47827 731310
rect 43253 730962 43319 730965
rect 41492 730960 43319 730962
rect 41492 730904 43258 730960
rect 43314 730904 43319 730960
rect 41492 730902 43319 730904
rect 43253 730899 43319 730902
rect 43437 730554 43503 730557
rect 41492 730552 43503 730554
rect 41492 730496 43442 730552
rect 43498 730496 43503 730552
rect 41492 730494 43503 730496
rect 43437 730491 43503 730494
rect 43069 730146 43135 730149
rect 41492 730144 43135 730146
rect 41492 730088 43074 730144
rect 43130 730088 43135 730144
rect 41492 730086 43135 730088
rect 43069 730083 43135 730086
rect 669037 730146 669103 730149
rect 675109 730146 675175 730149
rect 669037 730144 675175 730146
rect 669037 730088 669042 730144
rect 669098 730088 675114 730144
rect 675170 730088 675175 730144
rect 669037 730086 675175 730088
rect 669037 730083 669103 730086
rect 675109 730083 675175 730086
rect 44449 729738 44515 729741
rect 41492 729736 44515 729738
rect 41492 729680 44454 729736
rect 44510 729680 44515 729736
rect 41492 729678 44515 729680
rect 44449 729675 44515 729678
rect 42885 729330 42951 729333
rect 41492 729328 42951 729330
rect 41492 729272 42890 729328
rect 42946 729272 42951 729328
rect 41492 729270 42951 729272
rect 42885 729267 42951 729270
rect 41278 728687 41338 728892
rect 40861 728684 40927 728687
rect 40861 728682 40970 728684
rect 40861 728626 40866 728682
rect 40922 728626 40970 728682
rect 40861 728621 40970 728626
rect 41278 728682 41387 728687
rect 41278 728626 41326 728682
rect 41382 728626 41387 728682
rect 41278 728624 41387 728626
rect 41321 728621 41387 728624
rect 40910 728484 40970 728621
rect 62113 728242 62179 728245
rect 62113 728240 64492 728242
rect 62113 728184 62118 728240
rect 62174 728184 64492 728240
rect 62113 728182 64492 728184
rect 62113 728179 62179 728182
rect 42885 728106 42951 728109
rect 41492 728104 42951 728106
rect 41492 728048 42890 728104
rect 42946 728048 42951 728104
rect 41492 728046 42951 728048
rect 42885 728043 42951 728046
rect 674649 728106 674715 728109
rect 675845 728106 675911 728109
rect 674649 728104 675911 728106
rect 674649 728048 674654 728104
rect 674710 728048 675850 728104
rect 675906 728048 675911 728104
rect 674649 728046 675911 728048
rect 674649 728043 674715 728046
rect 675845 728043 675911 728046
rect 676254 728044 676260 728108
rect 676324 728106 676330 728108
rect 677501 728106 677567 728109
rect 676324 728104 677567 728106
rect 676324 728048 677506 728104
rect 677562 728048 677567 728104
rect 676324 728046 677567 728048
rect 676324 728044 676330 728046
rect 677501 728043 677567 728046
rect 674230 727772 674236 727836
rect 674300 727834 674306 727836
rect 683389 727834 683455 727837
rect 674300 727832 683455 727834
rect 674300 727776 683394 727832
rect 683450 727776 683455 727832
rect 674300 727774 683455 727776
rect 674300 727772 674306 727774
rect 683389 727771 683455 727774
rect 44633 727698 44699 727701
rect 41492 727696 44699 727698
rect 41492 727640 44638 727696
rect 44694 727640 44699 727696
rect 41492 727638 44699 727640
rect 44633 727635 44699 727638
rect 674189 727562 674255 727565
rect 676029 727562 676095 727565
rect 674189 727560 676095 727562
rect 674189 727504 674194 727560
rect 674250 727504 676034 727560
rect 676090 727504 676095 727560
rect 674189 727502 676095 727504
rect 674189 727499 674255 727502
rect 676029 727499 676095 727502
rect 41045 727460 41111 727463
rect 41045 727458 41154 727460
rect 41045 727402 41050 727458
rect 41106 727402 41154 727458
rect 41045 727397 41154 727402
rect 41094 727260 41154 727397
rect 41321 726882 41387 726885
rect 41308 726880 41387 726882
rect 41308 726824 41326 726880
rect 41382 726824 41387 726880
rect 41308 726822 41387 726824
rect 41321 726819 41387 726822
rect 42517 726474 42583 726477
rect 41492 726472 42583 726474
rect 41492 726416 42522 726472
rect 42578 726416 42583 726472
rect 41492 726414 42583 726416
rect 42517 726411 42583 726414
rect 40953 726236 41019 726239
rect 40910 726234 41019 726236
rect 40910 726178 40958 726234
rect 41014 726178 41019 726234
rect 40910 726173 41019 726178
rect 40910 726036 40970 726173
rect 41781 725796 41847 725797
rect 41781 725794 41828 725796
rect 41736 725792 41828 725794
rect 41736 725736 41786 725792
rect 41736 725734 41828 725736
rect 41781 725732 41828 725734
rect 41892 725732 41898 725796
rect 41781 725731 41847 725732
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 37917 725250 37983 725253
rect 37917 725248 37996 725250
rect 37917 725192 37922 725248
rect 37978 725192 37996 725248
rect 37917 725190 37996 725192
rect 37917 725187 37983 725190
rect 35157 724842 35223 724845
rect 35157 724840 35236 724842
rect 35157 724784 35162 724840
rect 35218 724784 35236 724840
rect 35157 724782 35236 724784
rect 35157 724779 35223 724782
rect 33041 724434 33107 724437
rect 33028 724432 33107 724434
rect 33028 724376 33046 724432
rect 33102 724376 33107 724432
rect 33028 724374 33107 724376
rect 33041 724371 33107 724374
rect 33734 723791 33794 723996
rect 33734 723786 33843 723791
rect 33734 723730 33782 723786
rect 33838 723730 33843 723786
rect 33734 723728 33843 723730
rect 33777 723725 33843 723728
rect 43253 723618 43319 723621
rect 41492 723616 43319 723618
rect 41492 723560 43258 723616
rect 43314 723560 43319 723616
rect 41492 723558 43319 723560
rect 43253 723555 43319 723558
rect 651557 723482 651623 723485
rect 650164 723480 651623 723482
rect 650164 723424 651562 723480
rect 651618 723424 651623 723480
rect 650164 723422 651623 723424
rect 651557 723419 651623 723422
rect 40677 723210 40743 723213
rect 40677 723208 40756 723210
rect 40677 723152 40682 723208
rect 40738 723152 40756 723208
rect 40677 723150 40756 723152
rect 40677 723147 40743 723150
rect 44173 722802 44239 722805
rect 41492 722800 44239 722802
rect 41492 722744 44178 722800
rect 44234 722744 44239 722800
rect 41492 722742 44239 722744
rect 44173 722739 44239 722742
rect 41781 722394 41847 722397
rect 41492 722392 41847 722394
rect 41492 722336 41786 722392
rect 41842 722336 41847 722392
rect 41492 722334 41847 722336
rect 41781 722331 41847 722334
rect 40726 721772 40786 721956
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 40902 721708 40908 721772
rect 40972 721708 40978 721772
rect 41137 721770 41203 721773
rect 41638 721770 41644 721772
rect 41137 721768 41644 721770
rect 41137 721712 41142 721768
rect 41198 721712 41644 721768
rect 41137 721710 41644 721712
rect 40910 721548 40970 721708
rect 41137 721707 41203 721710
rect 41638 721708 41644 721710
rect 41708 721708 41714 721772
rect 674833 721578 674899 721581
rect 676070 721578 676076 721580
rect 674833 721576 676076 721578
rect 674833 721520 674838 721576
rect 674894 721520 676076 721576
rect 674833 721518 676076 721520
rect 674833 721515 674899 721518
rect 676070 721516 676076 721518
rect 676140 721516 676146 721580
rect 46381 721170 46447 721173
rect 41492 721168 46447 721170
rect 41492 721112 46386 721168
rect 46442 721112 46447 721168
rect 41492 721110 46447 721112
rect 46381 721107 46447 721110
rect 31710 720357 31770 720732
rect 31710 720352 31819 720357
rect 31710 720324 31758 720352
rect 31740 720296 31758 720324
rect 31814 720296 31819 720352
rect 31740 720294 31819 720296
rect 31753 720291 31819 720294
rect 42333 719946 42399 719949
rect 41492 719944 42399 719946
rect 41492 719888 42338 719944
rect 42394 719888 42399 719944
rect 41492 719886 42399 719888
rect 42333 719883 42399 719886
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41781 718586 41847 718589
rect 40604 718584 41847 718586
rect 40604 718528 41786 718584
rect 41842 718528 41847 718584
rect 40604 718526 41847 718528
rect 40604 718524 40610 718526
rect 41781 718523 41847 718526
rect 41321 718314 41387 718317
rect 42333 718314 42399 718317
rect 41321 718312 42399 718314
rect 41321 718256 41326 718312
rect 41382 718256 42338 718312
rect 42394 718256 42399 718312
rect 41321 718254 42399 718256
rect 41321 718251 41387 718254
rect 42333 718251 42399 718254
rect 33041 716818 33107 716821
rect 41822 716818 41828 716820
rect 33041 716816 41828 716818
rect 33041 716760 33046 716816
rect 33102 716760 41828 716816
rect 33041 716758 41828 716760
rect 33041 716755 33107 716758
rect 41822 716756 41828 716758
rect 41892 716756 41898 716820
rect 675477 716546 675543 716549
rect 675477 716544 676292 716546
rect 675477 716488 675482 716544
rect 675538 716488 676292 716544
rect 675477 716486 676292 716488
rect 675477 716483 675543 716486
rect 675293 716138 675359 716141
rect 675293 716136 676292 716138
rect 675293 716080 675298 716136
rect 675354 716080 676292 716136
rect 675293 716078 676292 716080
rect 675293 716075 675359 716078
rect 675477 715730 675543 715733
rect 675477 715728 676292 715730
rect 675477 715672 675482 715728
rect 675538 715672 676292 715728
rect 675477 715670 676292 715672
rect 675477 715667 675543 715670
rect 62113 715322 62179 715325
rect 675109 715322 675175 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 675109 715320 676292 715322
rect 675109 715264 675114 715320
rect 675170 715264 676292 715320
rect 675109 715262 676292 715264
rect 62113 715259 62179 715262
rect 675109 715259 675175 715262
rect 42517 715186 42583 715189
rect 42517 715184 42626 715186
rect 42517 715128 42522 715184
rect 42578 715128 42626 715184
rect 42517 715123 42626 715128
rect 40309 714914 40375 714917
rect 42333 714914 42399 714917
rect 40309 714912 42399 714914
rect 40309 714856 40314 714912
rect 40370 714856 42338 714912
rect 42394 714856 42399 714912
rect 40309 714854 42399 714856
rect 40309 714851 40375 714854
rect 42333 714851 42399 714854
rect 42566 714780 42626 715123
rect 675477 714914 675543 714917
rect 675477 714912 676292 714914
rect 675477 714856 675482 714912
rect 675538 714856 676292 714912
rect 675477 714854 676292 714856
rect 675477 714851 675543 714854
rect 42558 714716 42564 714780
rect 42628 714716 42634 714780
rect 675477 714506 675543 714509
rect 675477 714504 676292 714506
rect 675477 714448 675482 714504
rect 675538 714448 676292 714504
rect 675477 714446 676292 714448
rect 675477 714443 675543 714446
rect 40677 714234 40743 714237
rect 41086 714234 41092 714236
rect 40677 714232 41092 714234
rect 40677 714176 40682 714232
rect 40738 714176 41092 714232
rect 40677 714174 41092 714176
rect 40677 714171 40743 714174
rect 41086 714172 41092 714174
rect 41156 714172 41162 714236
rect 675477 714098 675543 714101
rect 675477 714096 676292 714098
rect 675477 714040 675482 714096
rect 675538 714040 676292 714096
rect 675477 714038 676292 714040
rect 675477 714035 675543 714038
rect 41781 713962 41847 713965
rect 41781 713960 41890 713962
rect 41781 713904 41786 713960
rect 41842 713904 41890 713960
rect 41781 713899 41890 713904
rect 41830 713557 41890 713899
rect 675477 713690 675543 713693
rect 675477 713688 676292 713690
rect 675477 713632 675482 713688
rect 675538 713632 676292 713688
rect 675477 713630 676292 713632
rect 675477 713627 675543 713630
rect 41781 713552 41890 713557
rect 41781 713496 41786 713552
rect 41842 713496 41890 713552
rect 41781 713494 41890 713496
rect 41781 713491 41847 713494
rect 676765 713492 676831 713493
rect 676765 713488 676812 713492
rect 676876 713490 676882 713492
rect 676765 713432 676770 713488
rect 676765 713428 676812 713432
rect 676876 713430 676922 713490
rect 676876 713428 676882 713430
rect 676765 713427 676831 713428
rect 675477 713282 675543 713285
rect 675477 713280 676292 713282
rect 675477 713224 675482 713280
rect 675538 713224 676292 713280
rect 675477 713222 676292 713224
rect 675477 713219 675543 713222
rect 675477 712874 675543 712877
rect 675477 712872 676292 712874
rect 675477 712816 675482 712872
rect 675538 712816 676292 712872
rect 675477 712814 676292 712816
rect 675477 712811 675543 712814
rect 675477 712466 675543 712469
rect 675477 712464 676292 712466
rect 675477 712408 675482 712464
rect 675538 712408 676292 712464
rect 675477 712406 676292 712408
rect 675477 712403 675543 712406
rect 676029 712058 676095 712061
rect 676029 712056 676292 712058
rect 676029 712000 676034 712056
rect 676090 712000 676292 712056
rect 676029 711998 676292 712000
rect 676029 711995 676095 711998
rect 42149 711650 42215 711653
rect 42558 711650 42564 711652
rect 42149 711648 42564 711650
rect 42149 711592 42154 711648
rect 42210 711592 42564 711648
rect 42149 711590 42564 711592
rect 42149 711587 42215 711590
rect 42558 711588 42564 711590
rect 42628 711588 42634 711652
rect 676029 711650 676095 711653
rect 676029 711648 676292 711650
rect 676029 711592 676034 711648
rect 676090 711592 676292 711648
rect 676029 711590 676292 711592
rect 676029 711587 676095 711590
rect 675477 711242 675543 711245
rect 675477 711240 676292 711242
rect 675477 711184 675482 711240
rect 675538 711184 676292 711240
rect 675477 711182 676292 711184
rect 675477 711179 675543 711182
rect 684217 710834 684283 710837
rect 684204 710832 684283 710834
rect 684204 710776 684222 710832
rect 684278 710776 684283 710832
rect 684204 710774 684283 710776
rect 684217 710771 684283 710774
rect 670049 710698 670115 710701
rect 675845 710698 675911 710701
rect 670049 710696 675911 710698
rect 670049 710640 670054 710696
rect 670110 710640 675850 710696
rect 675906 710640 675911 710696
rect 670049 710638 675911 710640
rect 670049 710635 670115 710638
rect 675845 710635 675911 710638
rect 675293 710426 675359 710429
rect 675293 710424 676292 710426
rect 675293 710368 675298 710424
rect 675354 710368 676292 710424
rect 675293 710366 676292 710368
rect 675293 710363 675359 710366
rect 651557 710290 651623 710293
rect 650164 710288 651623 710290
rect 650164 710232 651562 710288
rect 651618 710232 651623 710288
rect 650164 710230 651623 710232
rect 651557 710227 651623 710230
rect 675477 710018 675543 710021
rect 675477 710016 676292 710018
rect 675477 709960 675482 710016
rect 675538 709960 676292 710016
rect 675477 709958 676292 709960
rect 675477 709955 675543 709958
rect 41086 709820 41092 709884
rect 41156 709882 41162 709884
rect 41781 709882 41847 709885
rect 41156 709880 41847 709882
rect 41156 709824 41786 709880
rect 41842 709824 41847 709880
rect 41156 709822 41847 709824
rect 41156 709820 41162 709822
rect 41781 709819 41847 709822
rect 675477 709610 675543 709613
rect 675477 709608 676292 709610
rect 675477 709552 675482 709608
rect 675538 709552 676292 709608
rect 675477 709550 676292 709552
rect 675477 709547 675543 709550
rect 683389 709202 683455 709205
rect 683389 709200 683468 709202
rect 683389 709144 683394 709200
rect 683450 709144 683468 709200
rect 683389 709142 683468 709144
rect 683389 709139 683455 709142
rect 674598 708732 674604 708796
rect 674668 708794 674674 708796
rect 674668 708734 676292 708794
rect 674668 708732 674674 708734
rect 40902 708460 40908 708524
rect 40972 708522 40978 708524
rect 41781 708522 41847 708525
rect 40972 708520 41847 708522
rect 40972 708464 41786 708520
rect 41842 708464 41847 708520
rect 40972 708462 41847 708464
rect 40972 708460 40978 708462
rect 41781 708459 41847 708462
rect 683205 708386 683271 708389
rect 683205 708384 683284 708386
rect 683205 708328 683210 708384
rect 683266 708328 683284 708384
rect 683205 708326 683284 708328
rect 683205 708323 683271 708326
rect 675477 707978 675543 707981
rect 675477 707976 676292 707978
rect 675477 707920 675482 707976
rect 675538 707920 676292 707976
rect 675477 707918 676292 707920
rect 675477 707915 675543 707918
rect 675477 707570 675543 707573
rect 675477 707568 676292 707570
rect 675477 707512 675482 707568
rect 675538 707512 676292 707568
rect 675477 707510 676292 707512
rect 675477 707507 675543 707510
rect 40718 707372 40724 707436
rect 40788 707434 40794 707436
rect 40788 707374 41890 707434
rect 40788 707372 40794 707374
rect 41830 707165 41890 707374
rect 41830 707160 41939 707165
rect 41830 707104 41878 707160
rect 41934 707104 41939 707160
rect 41830 707102 41939 707104
rect 41873 707099 41939 707102
rect 675477 707162 675543 707165
rect 675477 707160 676292 707162
rect 675477 707104 675482 707160
rect 675538 707104 676292 707160
rect 675477 707102 676292 707104
rect 675477 707099 675543 707102
rect 675477 706754 675543 706757
rect 675477 706752 676292 706754
rect 675477 706696 675482 706752
rect 675538 706696 676292 706752
rect 675477 706694 676292 706696
rect 675477 706691 675543 706694
rect 673310 706284 673316 706348
rect 673380 706346 673386 706348
rect 673380 706286 676292 706346
rect 673380 706284 673386 706286
rect 40534 706148 40540 706212
rect 40604 706210 40610 706212
rect 42241 706210 42307 706213
rect 40604 706208 42307 706210
rect 40604 706152 42246 706208
rect 42302 706152 42307 706208
rect 40604 706150 42307 706152
rect 40604 706148 40610 706150
rect 42241 706147 42307 706150
rect 677182 705530 677242 705908
rect 683113 705530 683179 705533
rect 677182 705528 683179 705530
rect 677182 705500 683118 705528
rect 677212 705472 683118 705500
rect 683174 705472 683179 705528
rect 677212 705470 683179 705472
rect 683113 705467 683179 705470
rect 675477 705122 675543 705125
rect 675477 705120 676292 705122
rect 675477 705064 675482 705120
rect 675538 705064 676292 705120
rect 675477 705062 676292 705064
rect 675477 705059 675543 705062
rect 41454 703700 41460 703764
rect 41524 703762 41530 703764
rect 42241 703762 42307 703765
rect 41524 703760 42307 703762
rect 41524 703704 42246 703760
rect 42302 703704 42307 703760
rect 41524 703702 42307 703704
rect 41524 703700 41530 703702
rect 42241 703699 42307 703702
rect 42057 703490 42123 703493
rect 43161 703490 43227 703493
rect 42057 703488 43227 703490
rect 42057 703432 42062 703488
rect 42118 703432 43166 703488
rect 43222 703432 43227 703488
rect 42057 703430 43227 703432
rect 42057 703427 42123 703430
rect 43161 703427 43227 703430
rect 42057 703082 42123 703085
rect 42701 703082 42767 703085
rect 42057 703080 42767 703082
rect 42057 703024 42062 703080
rect 42118 703024 42706 703080
rect 42762 703024 42767 703080
rect 42057 703022 42767 703024
rect 42057 703019 42123 703022
rect 42701 703019 42767 703022
rect 41638 702340 41644 702404
rect 41708 702402 41714 702404
rect 42609 702402 42675 702405
rect 41708 702400 42675 702402
rect 41708 702344 42614 702400
rect 42670 702344 42675 702400
rect 41708 702342 42675 702344
rect 41708 702340 41714 702342
rect 42609 702339 42675 702342
rect 62113 702266 62179 702269
rect 62113 702264 64492 702266
rect 62113 702208 62118 702264
rect 62174 702208 64492 702264
rect 62113 702206 64492 702208
rect 62113 702203 62179 702206
rect 41822 701796 41828 701860
rect 41892 701858 41898 701860
rect 42425 701858 42491 701861
rect 41892 701856 42491 701858
rect 41892 701800 42430 701856
rect 42486 701800 42491 701856
rect 41892 701798 42491 701800
rect 41892 701796 41898 701798
rect 42425 701795 42491 701798
rect 674598 698532 674604 698596
rect 674668 698594 674674 698596
rect 675385 698594 675451 698597
rect 674668 698592 675451 698594
rect 674668 698536 675390 698592
rect 675446 698536 675451 698592
rect 674668 698534 675451 698536
rect 674668 698532 674674 698534
rect 675385 698531 675451 698534
rect 651557 696962 651623 696965
rect 650164 696960 651623 696962
rect 650164 696904 651562 696960
rect 651618 696904 651623 696960
rect 650164 696902 651623 696904
rect 651557 696899 651623 696902
rect 675385 696828 675451 696829
rect 675334 696826 675340 696828
rect 675294 696766 675340 696826
rect 675404 696824 675451 696828
rect 675446 696768 675451 696824
rect 675334 696764 675340 696766
rect 675404 696764 675451 696768
rect 675385 696763 675451 696764
rect 675661 694378 675727 694381
rect 675661 694376 675954 694378
rect 675661 694320 675666 694376
rect 675722 694320 675954 694376
rect 675661 694318 675954 694320
rect 675661 694315 675727 694318
rect 675894 694106 675954 694318
rect 676806 694106 676812 694108
rect 675894 694046 676812 694106
rect 676806 694044 676812 694046
rect 676876 694044 676882 694108
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 672717 688666 672783 688669
rect 675477 688666 675543 688669
rect 672717 688664 675543 688666
rect 672717 688608 672722 688664
rect 672778 688608 675482 688664
rect 675538 688608 675543 688664
rect 672717 688606 675543 688608
rect 672717 688603 672783 688606
rect 675477 688603 675543 688606
rect 40953 688394 41019 688397
rect 40910 688392 41019 688394
rect 40910 688336 40958 688392
rect 41014 688336 41019 688392
rect 40910 688331 41019 688336
rect 40910 688092 40970 688331
rect 43253 687714 43319 687717
rect 41492 687712 43319 687714
rect 41492 687656 43258 687712
rect 43314 687656 43319 687712
rect 41492 687654 43319 687656
rect 43253 687651 43319 687654
rect 43437 687306 43503 687309
rect 41492 687304 43503 687306
rect 41492 687248 43442 687304
rect 43498 687248 43503 687304
rect 41492 687246 43503 687248
rect 43437 687243 43503 687246
rect 41137 686898 41203 686901
rect 41124 686896 41203 686898
rect 41124 686840 41142 686896
rect 41198 686840 41203 686896
rect 41124 686838 41203 686840
rect 41137 686835 41203 686838
rect 44265 686490 44331 686493
rect 41492 686488 44331 686490
rect 41492 686432 44270 686488
rect 44326 686432 44331 686488
rect 41492 686430 44331 686432
rect 44265 686427 44331 686430
rect 41278 685915 41338 686052
rect 40861 685912 40927 685915
rect 40861 685910 40970 685912
rect 40861 685854 40866 685910
rect 40922 685854 40970 685910
rect 40861 685849 40970 685854
rect 41278 685910 41387 685915
rect 41278 685854 41326 685910
rect 41382 685854 41387 685910
rect 41278 685852 41387 685854
rect 41321 685849 41387 685852
rect 40910 685644 40970 685849
rect 41137 685266 41203 685269
rect 41124 685264 41203 685266
rect 41124 685208 41142 685264
rect 41198 685208 41203 685264
rect 41124 685206 41203 685208
rect 41137 685203 41203 685206
rect 675017 685266 675083 685269
rect 675334 685266 675340 685268
rect 675017 685264 675340 685266
rect 675017 685208 675022 685264
rect 675078 685208 675340 685264
rect 675017 685206 675340 685208
rect 675017 685203 675083 685206
rect 675334 685204 675340 685206
rect 675404 685204 675410 685268
rect 667841 684994 667907 684997
rect 675477 684994 675543 684997
rect 667841 684992 675543 684994
rect 667841 684936 667846 684992
rect 667902 684936 675482 684992
rect 675538 684936 675543 684992
rect 667841 684934 675543 684936
rect 667841 684931 667907 684934
rect 675477 684931 675543 684934
rect 42701 684858 42767 684861
rect 41492 684856 42767 684858
rect 41492 684800 42706 684856
rect 42762 684800 42767 684856
rect 41492 684798 42767 684800
rect 42701 684795 42767 684798
rect 43069 684450 43135 684453
rect 41492 684448 43135 684450
rect 41492 684392 43074 684448
rect 43130 684392 43135 684448
rect 41492 684390 43135 684392
rect 43069 684387 43135 684390
rect 43253 684042 43319 684045
rect 41492 684040 43319 684042
rect 41492 683984 43258 684040
rect 43314 683984 43319 684040
rect 41492 683982 43319 683984
rect 43253 683979 43319 683982
rect 40953 683634 41019 683637
rect 651557 683634 651623 683637
rect 40940 683632 41019 683634
rect 40940 683576 40958 683632
rect 41014 683576 41019 683632
rect 40940 683574 41019 683576
rect 650164 683632 651623 683634
rect 650164 683576 651562 683632
rect 651618 683576 651623 683632
rect 650164 683574 651623 683576
rect 40953 683571 41019 683574
rect 651557 683571 651623 683574
rect 41321 683226 41387 683229
rect 41308 683224 41387 683226
rect 41308 683168 41326 683224
rect 41382 683168 41387 683224
rect 41308 683166 41387 683168
rect 41321 683163 41387 683166
rect 674005 683090 674071 683093
rect 675845 683090 675911 683093
rect 674005 683088 675911 683090
rect 674005 683032 674010 683088
rect 674066 683032 675850 683088
rect 675906 683032 675911 683088
rect 674005 683030 675911 683032
rect 674005 683027 674071 683030
rect 675845 683027 675911 683030
rect 40769 682818 40835 682821
rect 40756 682816 40835 682818
rect 40756 682760 40774 682816
rect 40830 682760 40835 682816
rect 40756 682758 40835 682760
rect 40769 682755 40835 682758
rect 40585 682410 40651 682413
rect 40572 682408 40651 682410
rect 40572 682352 40590 682408
rect 40646 682352 40651 682408
rect 40572 682350 40651 682352
rect 40585 682347 40651 682350
rect 41781 682412 41847 682413
rect 41781 682408 41828 682412
rect 41892 682410 41898 682412
rect 41781 682352 41786 682408
rect 41781 682348 41828 682352
rect 41892 682350 41938 682410
rect 41892 682348 41898 682350
rect 41781 682347 41847 682348
rect 37917 682002 37983 682005
rect 37917 682000 37996 682002
rect 37917 681944 37922 682000
rect 37978 681944 37996 682000
rect 37917 681942 37996 681944
rect 37917 681939 37983 681942
rect 36537 681594 36603 681597
rect 36524 681592 36603 681594
rect 36524 681536 36542 681592
rect 36598 681536 36603 681592
rect 36524 681534 36603 681536
rect 36537 681531 36603 681534
rect 32397 681186 32463 681189
rect 32397 681184 32476 681186
rect 32397 681128 32402 681184
rect 32458 681128 32476 681184
rect 32397 681126 32476 681128
rect 32397 681123 32463 681126
rect 33777 680778 33843 680781
rect 33764 680776 33843 680778
rect 33764 680720 33782 680776
rect 33838 680720 33843 680776
rect 33764 680718 33843 680720
rect 33777 680715 33843 680718
rect 43437 680370 43503 680373
rect 41492 680368 43503 680370
rect 41492 680312 43442 680368
rect 43498 680312 43503 680368
rect 41492 680310 43503 680312
rect 43437 680307 43503 680310
rect 45185 679962 45251 679965
rect 41492 679960 45251 679962
rect 41492 679904 45190 679960
rect 45246 679904 45251 679960
rect 41492 679902 45251 679904
rect 45185 679899 45251 679902
rect 44633 679554 44699 679557
rect 41492 679552 44699 679554
rect 41492 679496 44638 679552
rect 44694 679496 44699 679552
rect 41492 679494 44699 679496
rect 44633 679491 44699 679494
rect 40542 678992 40602 679116
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678928 40794 678992
rect 40726 678708 40786 678928
rect 41781 678876 41847 678877
rect 41781 678872 41828 678876
rect 41892 678874 41898 678876
rect 41781 678816 41786 678872
rect 41781 678812 41828 678816
rect 41892 678814 41938 678874
rect 41892 678812 41898 678814
rect 41781 678811 41847 678812
rect 43253 678330 43319 678333
rect 41492 678328 43319 678330
rect 41492 678272 43258 678328
rect 43314 678272 43319 678328
rect 41492 678270 43319 678272
rect 43253 678267 43319 678270
rect 676070 678268 676076 678332
rect 676140 678330 676146 678332
rect 678237 678330 678303 678333
rect 676140 678328 678303 678330
rect 676140 678272 678242 678328
rect 678298 678272 678303 678328
rect 676140 678270 678303 678272
rect 676140 678268 676146 678270
rect 678237 678267 678303 678270
rect 45001 677922 45067 677925
rect 41492 677920 45067 677922
rect 41492 677864 45006 677920
rect 45062 677864 45067 677920
rect 41492 677862 45067 677864
rect 45001 677859 45067 677862
rect 41094 677109 41154 677484
rect 41094 677104 41203 677109
rect 41094 677076 41142 677104
rect 41124 677048 41142 677076
rect 41198 677048 41203 677104
rect 41124 677046 41203 677048
rect 41137 677043 41203 677046
rect 43989 676698 44055 676701
rect 41492 676696 44055 676698
rect 41492 676640 43994 676696
rect 44050 676640 44055 676696
rect 41492 676638 44055 676640
rect 43989 676635 44055 676638
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 674414 674052 674420 674116
rect 674484 674114 674490 674116
rect 683205 674114 683271 674117
rect 674484 674112 683271 674114
rect 674484 674056 683210 674112
rect 683266 674056 683271 674112
rect 674484 674054 683271 674056
rect 674484 674052 674490 674054
rect 683205 674051 683271 674054
rect 32397 672754 32463 672757
rect 41822 672754 41828 672756
rect 32397 672752 41828 672754
rect 32397 672696 32402 672752
rect 32458 672696 41828 672752
rect 32397 672694 41828 672696
rect 32397 672691 32463 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 41137 672484 41203 672485
rect 41086 672420 41092 672484
rect 41156 672482 41203 672484
rect 41156 672480 41248 672482
rect 41198 672424 41248 672480
rect 41156 672422 41248 672424
rect 41156 672420 41203 672422
rect 41137 672419 41203 672420
rect 42241 672212 42307 672213
rect 42190 672148 42196 672212
rect 42260 672210 42307 672212
rect 42260 672208 42352 672210
rect 42302 672152 42352 672208
rect 42260 672150 42352 672152
rect 42260 672148 42307 672150
rect 42241 672147 42307 672148
rect 39481 671530 39547 671533
rect 42701 671530 42767 671533
rect 39481 671528 42767 671530
rect 39481 671472 39486 671528
rect 39542 671472 42706 671528
rect 42762 671472 42767 671528
rect 39481 671470 42767 671472
rect 39481 671467 39547 671470
rect 42701 671467 42767 671470
rect 675293 671394 675359 671397
rect 675293 671392 676292 671394
rect 675293 671336 675298 671392
rect 675354 671336 676292 671392
rect 675293 671334 676292 671336
rect 675293 671331 675359 671334
rect 40033 671258 40099 671261
rect 42701 671258 42767 671261
rect 40033 671256 42767 671258
rect 40033 671200 40038 671256
rect 40094 671200 42706 671256
rect 42762 671200 42767 671256
rect 40033 671198 42767 671200
rect 40033 671195 40099 671198
rect 42701 671195 42767 671198
rect 675477 670986 675543 670989
rect 675477 670984 676292 670986
rect 675477 670928 675482 670984
rect 675538 670928 676292 670984
rect 675477 670926 676292 670928
rect 675477 670923 675543 670926
rect 675661 670578 675727 670581
rect 675661 670576 676292 670578
rect 675661 670520 675666 670576
rect 675722 670520 676292 670576
rect 675661 670518 676292 670520
rect 675661 670515 675727 670518
rect 651557 670442 651623 670445
rect 650164 670440 651623 670442
rect 650164 670384 651562 670440
rect 651618 670384 651623 670440
rect 650164 670382 651623 670384
rect 651557 670379 651623 670382
rect 675293 670170 675359 670173
rect 675293 670168 676292 670170
rect 675293 670112 675298 670168
rect 675354 670112 676292 670168
rect 675293 670110 676292 670112
rect 675293 670107 675359 670110
rect 675477 669762 675543 669765
rect 675477 669760 676292 669762
rect 675477 669704 675482 669760
rect 675538 669704 676292 669760
rect 675477 669702 676292 669704
rect 675477 669699 675543 669702
rect 674833 669354 674899 669357
rect 674833 669352 676292 669354
rect 674833 669296 674838 669352
rect 674894 669296 676292 669352
rect 674833 669294 676292 669296
rect 674833 669291 674899 669294
rect 41086 669020 41092 669084
rect 41156 669082 41162 669084
rect 41781 669082 41847 669085
rect 41156 669080 41847 669082
rect 41156 669024 41786 669080
rect 41842 669024 41847 669080
rect 41156 669022 41847 669024
rect 41156 669020 41162 669022
rect 41781 669019 41847 669022
rect 675293 668946 675359 668949
rect 675293 668944 676292 668946
rect 675293 668888 675298 668944
rect 675354 668888 676292 668944
rect 675293 668886 676292 668888
rect 675293 668883 675359 668886
rect 675477 668538 675543 668541
rect 675477 668536 676292 668538
rect 675477 668480 675482 668536
rect 675538 668480 676292 668536
rect 675477 668478 676292 668480
rect 675477 668475 675543 668478
rect 675477 668130 675543 668133
rect 675477 668128 676292 668130
rect 675477 668072 675482 668128
rect 675538 668072 676292 668128
rect 675477 668070 676292 668072
rect 675477 668067 675543 668070
rect 42057 667722 42123 667725
rect 43621 667722 43687 667725
rect 42057 667720 43687 667722
rect 42057 667664 42062 667720
rect 42118 667664 43626 667720
rect 43682 667664 43687 667720
rect 42057 667662 43687 667664
rect 42057 667659 42123 667662
rect 43621 667659 43687 667662
rect 675477 667722 675543 667725
rect 675477 667720 676292 667722
rect 675477 667664 675482 667720
rect 675538 667664 676292 667720
rect 675477 667662 676292 667664
rect 675477 667659 675543 667662
rect 42190 667388 42196 667452
rect 42260 667450 42266 667452
rect 42425 667450 42491 667453
rect 42260 667448 42491 667450
rect 42260 667392 42430 667448
rect 42486 667392 42491 667448
rect 42260 667390 42491 667392
rect 42260 667388 42266 667390
rect 42425 667387 42491 667390
rect 675477 667314 675543 667317
rect 675477 667312 676292 667314
rect 675477 667256 675482 667312
rect 675538 667256 676292 667312
rect 675477 667254 676292 667256
rect 675477 667251 675543 667254
rect 678237 667042 678303 667045
rect 678237 667040 678346 667042
rect 678237 666984 678242 667040
rect 678298 666984 678346 667040
rect 678237 666979 678346 666984
rect 678286 666876 678346 666979
rect 675293 666498 675359 666501
rect 675293 666496 676292 666498
rect 675293 666440 675298 666496
rect 675354 666440 676292 666496
rect 675293 666438 676292 666440
rect 675293 666435 675359 666438
rect 675477 666090 675543 666093
rect 675477 666088 676292 666090
rect 675477 666032 675482 666088
rect 675538 666032 676292 666088
rect 675477 666030 676292 666032
rect 675477 666027 675543 666030
rect 675477 665682 675543 665685
rect 675477 665680 676292 665682
rect 675477 665624 675482 665680
rect 675538 665624 676292 665680
rect 675477 665622 676292 665624
rect 675477 665619 675543 665622
rect 676990 665348 676996 665412
rect 677060 665348 677066 665412
rect 676998 665244 677058 665348
rect 42057 665138 42123 665141
rect 43253 665138 43319 665141
rect 42057 665136 43319 665138
rect 42057 665080 42062 665136
rect 42118 665080 43258 665136
rect 43314 665080 43319 665136
rect 42057 665078 43319 665080
rect 42057 665075 42123 665078
rect 43253 665075 43319 665078
rect 675477 664866 675543 664869
rect 675477 664864 676292 664866
rect 675477 664808 675482 664864
rect 675538 664808 676292 664864
rect 675477 664806 676292 664808
rect 675477 664803 675543 664806
rect 675477 664458 675543 664461
rect 675477 664456 676292 664458
rect 675477 664400 675482 664456
rect 675538 664400 676292 664456
rect 675477 664398 676292 664400
rect 675477 664395 675543 664398
rect 40718 664124 40724 664188
rect 40788 664186 40794 664188
rect 41781 664186 41847 664189
rect 40788 664184 41847 664186
rect 40788 664128 41786 664184
rect 41842 664128 41847 664184
rect 40788 664126 41847 664128
rect 40788 664124 40794 664126
rect 41781 664123 41847 664126
rect 674465 664050 674531 664053
rect 674465 664048 676292 664050
rect 674465 663992 674470 664048
rect 674526 663992 676292 664048
rect 674465 663990 676292 663992
rect 674465 663987 674531 663990
rect 683389 663778 683455 663781
rect 683389 663776 683498 663778
rect 683389 663720 683394 663776
rect 683450 663720 683498 663776
rect 683389 663715 683498 663720
rect 683438 663612 683498 663715
rect 669037 663506 669103 663509
rect 675845 663506 675911 663509
rect 669037 663504 675911 663506
rect 669037 663448 669042 663504
rect 669098 663448 675850 663504
rect 675906 663448 675911 663504
rect 669037 663446 675911 663448
rect 669037 663443 669103 663446
rect 675845 663443 675911 663446
rect 675477 663234 675543 663237
rect 675477 663232 676292 663234
rect 675477 663176 675482 663232
rect 675538 663176 676292 663232
rect 675477 663174 676292 663176
rect 675477 663171 675543 663174
rect 62113 663098 62179 663101
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 62113 663035 62179 663038
rect 40534 662764 40540 662828
rect 40604 662826 40610 662828
rect 42149 662826 42215 662829
rect 40604 662824 42215 662826
rect 40604 662768 42154 662824
rect 42210 662768 42215 662824
rect 40604 662766 42215 662768
rect 40604 662764 40610 662766
rect 42149 662763 42215 662766
rect 675477 662826 675543 662829
rect 675477 662824 676292 662826
rect 675477 662768 675482 662824
rect 675538 662768 676292 662824
rect 675477 662766 676292 662768
rect 675477 662763 675543 662766
rect 683205 662554 683271 662557
rect 683205 662552 683314 662554
rect 683205 662496 683210 662552
rect 683266 662496 683314 662552
rect 683205 662491 683314 662496
rect 683254 662388 683314 662491
rect 675477 662010 675543 662013
rect 675477 662008 676292 662010
rect 675477 661952 675482 662008
rect 675538 661952 676292 662008
rect 675477 661950 676292 661952
rect 675477 661947 675543 661950
rect 675477 661602 675543 661605
rect 675477 661600 676292 661602
rect 675477 661544 675482 661600
rect 675538 661544 676292 661600
rect 675477 661542 676292 661544
rect 675477 661539 675543 661542
rect 675477 661194 675543 661197
rect 675477 661192 676292 661194
rect 675477 661136 675482 661192
rect 675538 661136 676292 661192
rect 675477 661134 676292 661136
rect 675477 661131 675543 661134
rect 41454 660316 41460 660380
rect 41524 660378 41530 660380
rect 42609 660378 42675 660381
rect 41524 660376 42675 660378
rect 41524 660320 42614 660376
rect 42670 660320 42675 660376
rect 41524 660318 42675 660320
rect 41524 660316 41530 660318
rect 42609 660315 42675 660318
rect 683070 660109 683130 660756
rect 683070 660104 683179 660109
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660046 683179 660048
rect 683113 660043 683179 660046
rect 675477 659970 675543 659973
rect 675477 659968 676292 659970
rect 675477 659912 675482 659968
rect 675538 659912 676292 659968
rect 675477 659910 676292 659912
rect 675477 659907 675543 659910
rect 41638 658820 41644 658884
rect 41708 658882 41714 658884
rect 42425 658882 42491 658885
rect 41708 658880 42491 658882
rect 41708 658824 42430 658880
rect 42486 658824 42491 658880
rect 41708 658822 42491 658824
rect 41708 658820 41714 658822
rect 42425 658819 42491 658822
rect 41822 658548 41828 658612
rect 41892 658610 41898 658612
rect 42241 658610 42307 658613
rect 41892 658608 42307 658610
rect 41892 658552 42246 658608
rect 42302 658552 42307 658608
rect 41892 658550 42307 658552
rect 41892 658548 41898 658550
rect 42241 658547 42307 658550
rect 651557 657114 651623 657117
rect 650164 657112 651623 657114
rect 650164 657056 651562 657112
rect 651618 657056 651623 657112
rect 650164 657054 651623 657056
rect 651557 657051 651623 657054
rect 675569 652900 675635 652901
rect 675518 652898 675524 652900
rect 675478 652838 675524 652898
rect 675588 652896 675635 652900
rect 675630 652840 675635 652896
rect 675518 652836 675524 652838
rect 675588 652836 675635 652840
rect 675569 652835 675635 652836
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 674833 649226 674899 649229
rect 675477 649226 675543 649229
rect 674833 649224 675543 649226
rect 674833 649168 674838 649224
rect 674894 649168 675482 649224
rect 675538 649168 675543 649224
rect 674833 649166 675543 649168
rect 674833 649163 674899 649166
rect 675477 649163 675543 649166
rect 674414 648620 674420 648684
rect 674484 648682 674490 648684
rect 675569 648682 675635 648685
rect 674484 648680 675635 648682
rect 674484 648624 675574 648680
rect 675630 648624 675635 648680
rect 674484 648622 675635 648624
rect 674484 648620 674490 648622
rect 675569 648619 675635 648622
rect 39389 646098 39455 646101
rect 47761 646098 47827 646101
rect 39389 646096 47827 646098
rect 39389 646040 39394 646096
rect 39450 646040 47766 646096
rect 47822 646040 47827 646096
rect 39389 646038 47827 646040
rect 39389 646035 39455 646038
rect 47761 646035 47827 646038
rect 675293 645828 675359 645829
rect 675293 645824 675340 645828
rect 675404 645826 675410 645828
rect 675293 645768 675298 645824
rect 675293 645764 675340 645768
rect 675404 645766 675450 645826
rect 675404 645764 675410 645766
rect 675293 645763 675359 645764
rect 672533 645418 672599 645421
rect 675477 645418 675543 645421
rect 672533 645416 675543 645418
rect 672533 645360 672538 645416
rect 672594 645360 675482 645416
rect 675538 645360 675543 645416
rect 672533 645358 675543 645360
rect 672533 645355 672599 645358
rect 675477 645355 675543 645358
rect 35574 644741 35634 644912
rect 35525 644736 35634 644741
rect 35801 644738 35867 644741
rect 35525 644680 35530 644736
rect 35586 644680 35634 644736
rect 35525 644678 35634 644680
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35525 644675 35591 644678
rect 35758 644675 35867 644680
rect 39757 644738 39823 644741
rect 43805 644738 43871 644741
rect 39757 644736 43871 644738
rect 39757 644680 39762 644736
rect 39818 644680 43810 644736
rect 43866 644680 43871 644736
rect 39757 644678 43871 644680
rect 39757 644675 39823 644678
rect 43805 644675 43871 644678
rect 674465 644738 674531 644741
rect 675385 644738 675451 644741
rect 674465 644736 675451 644738
rect 674465 644680 674470 644736
rect 674526 644680 675390 644736
rect 675446 644680 675451 644736
rect 674465 644678 675451 644680
rect 674465 644675 674531 644678
rect 675385 644675 675451 644678
rect 35758 644504 35818 644675
rect 674097 644330 674163 644333
rect 675385 644330 675451 644333
rect 674097 644328 675451 644330
rect 674097 644272 674102 644328
rect 674158 644272 675390 644328
rect 675446 644272 675451 644328
rect 674097 644270 675451 644272
rect 674097 644267 674163 644270
rect 675385 644267 675451 644270
rect 35390 643925 35450 644096
rect 35341 643920 35450 643925
rect 35341 643864 35346 643920
rect 35402 643864 35450 643920
rect 35341 643862 35450 643864
rect 39849 643922 39915 643925
rect 43069 643922 43135 643925
rect 39849 643920 43135 643922
rect 39849 643864 39854 643920
rect 39910 643864 43074 643920
rect 43130 643864 43135 643920
rect 39849 643862 43135 643864
rect 35341 643859 35407 643862
rect 39849 643859 39915 643862
rect 43069 643859 43135 643862
rect 651557 643786 651623 643789
rect 650164 643784 651623 643786
rect 650164 643728 651562 643784
rect 651618 643728 651623 643784
rect 650164 643726 651623 643728
rect 651557 643723 651623 643726
rect 35574 643517 35634 643688
rect 35525 643512 35634 643517
rect 35801 643514 35867 643517
rect 35525 643456 35530 643512
rect 35586 643456 35634 643512
rect 35525 643454 35634 643456
rect 35758 643512 35867 643514
rect 35758 643456 35806 643512
rect 35862 643456 35867 643512
rect 35525 643451 35591 643454
rect 35758 643451 35867 643456
rect 39665 643514 39731 643517
rect 44633 643514 44699 643517
rect 39665 643512 44699 643514
rect 39665 643456 39670 643512
rect 39726 643456 44638 643512
rect 44694 643456 44699 643512
rect 39665 643454 44699 643456
rect 39665 643451 39731 643454
rect 44633 643451 44699 643454
rect 671705 643514 671771 643517
rect 675477 643514 675543 643517
rect 671705 643512 675543 643514
rect 671705 643456 671710 643512
rect 671766 643456 675482 643512
rect 675538 643456 675543 643512
rect 671705 643454 675543 643456
rect 671705 643451 671771 643454
rect 675477 643451 675543 643454
rect 35758 643280 35818 643451
rect 39573 643106 39639 643109
rect 44265 643106 44331 643109
rect 39573 643104 44331 643106
rect 39573 643048 39578 643104
rect 39634 643048 44270 643104
rect 44326 643048 44331 643104
rect 39573 643046 44331 643048
rect 39573 643043 39639 643046
rect 44265 643043 44331 643046
rect 674833 643106 674899 643109
rect 675477 643106 675543 643109
rect 674833 643104 675543 643106
rect 674833 643048 674838 643104
rect 674894 643048 675482 643104
rect 675538 643048 675543 643104
rect 674833 643046 675543 643048
rect 674833 643043 674899 643046
rect 675477 643043 675543 643046
rect 35390 642701 35450 642872
rect 35390 642696 35499 642701
rect 35390 642640 35438 642696
rect 35494 642640 35499 642696
rect 35390 642638 35499 642640
rect 35433 642635 35499 642638
rect 35574 642293 35634 642464
rect 35574 642288 35683 642293
rect 35574 642232 35622 642288
rect 35678 642232 35683 642288
rect 35574 642230 35683 642232
rect 35617 642227 35683 642230
rect 38929 642290 38995 642293
rect 42885 642290 42951 642293
rect 38929 642288 42951 642290
rect 38929 642232 38934 642288
rect 38990 642232 42890 642288
rect 42946 642232 42951 642288
rect 38929 642230 42951 642232
rect 38929 642227 38995 642230
rect 42885 642227 42951 642230
rect 35758 641885 35818 642056
rect 35758 641880 35867 641885
rect 35758 641824 35806 641880
rect 35862 641824 35867 641880
rect 35758 641822 35867 641824
rect 35801 641819 35867 641822
rect 35758 641477 35818 641648
rect 35758 641472 35867 641477
rect 35758 641416 35806 641472
rect 35862 641416 35867 641472
rect 35758 641414 35867 641416
rect 35801 641411 35867 641414
rect 35574 641069 35634 641240
rect 35574 641064 35683 641069
rect 35574 641008 35622 641064
rect 35678 641008 35683 641064
rect 35574 641006 35683 641008
rect 35617 641003 35683 641006
rect 35758 640661 35818 640832
rect 35758 640656 35867 640661
rect 35758 640600 35806 640656
rect 35862 640600 35867 640656
rect 35758 640598 35867 640600
rect 35801 640595 35867 640598
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 674005 640522 674071 640525
rect 675477 640522 675543 640525
rect 674005 640520 675543 640522
rect 674005 640464 674010 640520
rect 674066 640464 675482 640520
rect 675538 640464 675543 640520
rect 674005 640462 675543 640464
rect 674005 640459 674071 640462
rect 675477 640459 675543 640462
rect 39665 640250 39731 640253
rect 43253 640250 43319 640253
rect 39665 640248 43319 640250
rect 39665 640192 39670 640248
rect 39726 640192 43258 640248
rect 43314 640192 43319 640248
rect 39665 640190 43319 640192
rect 39665 640187 39731 640190
rect 43253 640187 43319 640190
rect 35390 639845 35450 640016
rect 35341 639840 35450 639845
rect 35341 639784 35346 639840
rect 35402 639784 35450 639840
rect 35341 639782 35450 639784
rect 35341 639779 35407 639782
rect 35574 639437 35634 639608
rect 35525 639432 35634 639437
rect 35801 639434 35867 639437
rect 35525 639376 35530 639432
rect 35586 639376 35634 639432
rect 35525 639374 35634 639376
rect 35758 639432 35867 639434
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35525 639371 35591 639374
rect 35758 639371 35867 639376
rect 674833 639434 674899 639437
rect 675385 639434 675451 639437
rect 674833 639432 675451 639434
rect 674833 639376 674838 639432
rect 674894 639376 675390 639432
rect 675446 639376 675451 639432
rect 674833 639374 675451 639376
rect 674833 639371 674899 639374
rect 675385 639371 675451 639374
rect 35758 639200 35818 639371
rect 33734 638621 33794 638792
rect 33734 638616 33843 638621
rect 33734 638560 33782 638616
rect 33838 638560 33843 638616
rect 33734 638558 33843 638560
rect 33777 638555 33843 638558
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 41505 638210 41571 638213
rect 44357 638210 44423 638213
rect 41505 638208 44423 638210
rect 41505 638152 41510 638208
rect 41566 638152 44362 638208
rect 44418 638152 44423 638208
rect 41505 638150 44423 638152
rect 32397 638147 32463 638150
rect 41505 638147 41571 638150
rect 44357 638147 44423 638150
rect 675201 638210 675267 638213
rect 675753 638210 675819 638213
rect 675201 638208 675819 638210
rect 675201 638152 675206 638208
rect 675262 638152 675758 638208
rect 675814 638152 675819 638208
rect 675201 638150 675819 638152
rect 675201 638147 675267 638150
rect 675753 638147 675819 638150
rect 35758 637805 35818 637976
rect 35525 637802 35591 637805
rect 35525 637800 35634 637802
rect 35525 637744 35530 637800
rect 35586 637744 35634 637800
rect 35525 637739 35634 637744
rect 35758 637800 35867 637805
rect 35758 637744 35806 637800
rect 35862 637744 35867 637800
rect 35758 637742 35867 637744
rect 35801 637739 35867 637742
rect 40953 637802 41019 637805
rect 43621 637802 43687 637805
rect 675293 637804 675359 637805
rect 675293 637802 675340 637804
rect 40953 637800 43687 637802
rect 40953 637744 40958 637800
rect 41014 637744 43626 637800
rect 43682 637744 43687 637800
rect 40953 637742 43687 637744
rect 675248 637800 675340 637802
rect 675248 637744 675298 637800
rect 675248 637742 675340 637744
rect 40953 637739 41019 637742
rect 43621 637739 43687 637742
rect 675293 637740 675340 637742
rect 675404 637740 675410 637804
rect 675293 637739 675359 637740
rect 35574 637568 35634 637739
rect 675569 637668 675635 637669
rect 675518 637666 675524 637668
rect 675478 637606 675524 637666
rect 675588 637664 675635 637668
rect 675630 637608 675635 637664
rect 675518 637604 675524 637606
rect 675588 637604 675635 637608
rect 675569 637603 675635 637604
rect 40033 637394 40099 637397
rect 41638 637394 41644 637396
rect 40033 637392 41644 637394
rect 40033 637336 40038 637392
rect 40094 637336 41644 637392
rect 40033 637334 41644 637336
rect 40033 637331 40099 637334
rect 41638 637332 41644 637334
rect 41708 637332 41714 637396
rect 675017 637394 675083 637397
rect 676029 637394 676095 637397
rect 675017 637392 676095 637394
rect 675017 637336 675022 637392
rect 675078 637336 676034 637392
rect 676090 637336 676095 637392
rect 675017 637334 676095 637336
rect 675017 637331 675083 637334
rect 676029 637331 676095 637334
rect 40542 636988 40602 637160
rect 62113 637122 62179 637125
rect 673637 637122 673703 637125
rect 676029 637122 676095 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 673637 637120 676095 637122
rect 673637 637064 673642 637120
rect 673698 637064 676034 637120
rect 676090 637064 676095 637120
rect 673637 637062 676095 637064
rect 62113 637059 62179 637062
rect 673637 637059 673703 637062
rect 676029 637059 676095 637062
rect 40534 636924 40540 636988
rect 40604 636924 40610 636988
rect 35758 636581 35818 636752
rect 35758 636576 35867 636581
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35758 636518 35867 636520
rect 35801 636515 35867 636518
rect 40910 636172 40970 636344
rect 40902 636108 40908 636172
rect 40972 636108 40978 636172
rect 40726 635764 40786 635936
rect 40718 635700 40724 635764
rect 40788 635700 40794 635764
rect 35574 635357 35634 635528
rect 35574 635352 35683 635357
rect 35574 635296 35622 635352
rect 35678 635296 35683 635352
rect 35574 635294 35683 635296
rect 35617 635291 35683 635294
rect 40217 635354 40283 635357
rect 41822 635354 41828 635356
rect 40217 635352 41828 635354
rect 40217 635296 40222 635352
rect 40278 635296 41828 635352
rect 40217 635294 41828 635296
rect 40217 635291 40283 635294
rect 41822 635292 41828 635294
rect 41892 635292 41898 635356
rect 35758 634949 35818 635120
rect 35758 634944 35867 634949
rect 35758 634888 35806 634944
rect 35862 634888 35867 634944
rect 35758 634886 35867 634888
rect 35801 634883 35867 634886
rect 39573 634946 39639 634949
rect 43805 634946 43871 634949
rect 39573 634944 43871 634946
rect 39573 634888 39578 634944
rect 39634 634888 43810 634944
rect 43866 634888 43871 634944
rect 39573 634886 43871 634888
rect 39573 634883 39639 634886
rect 43805 634883 43871 634886
rect 35758 634541 35818 634712
rect 35758 634536 35867 634541
rect 35758 634480 35806 634536
rect 35862 634480 35867 634536
rect 35758 634478 35867 634480
rect 35801 634475 35867 634478
rect 40677 634538 40743 634541
rect 43989 634538 44055 634541
rect 40677 634536 44055 634538
rect 40677 634480 40682 634536
rect 40738 634480 43994 634536
rect 44050 634480 44055 634536
rect 40677 634478 44055 634480
rect 40677 634475 40743 634478
rect 43989 634475 44055 634478
rect 41462 633858 41522 634304
rect 42333 633858 42399 633861
rect 41462 633856 42399 633858
rect 41462 633800 42338 633856
rect 42394 633800 42399 633856
rect 41462 633798 42399 633800
rect 42333 633795 42399 633798
rect 35801 633722 35867 633725
rect 35758 633720 35867 633722
rect 35758 633664 35806 633720
rect 35862 633664 35867 633720
rect 35758 633659 35867 633664
rect 35758 633488 35818 633659
rect 40493 632090 40559 632093
rect 45185 632090 45251 632093
rect 40493 632088 45251 632090
rect 40493 632032 40498 632088
rect 40554 632032 45190 632088
rect 45246 632032 45251 632088
rect 40493 632030 45251 632032
rect 40493 632027 40559 632030
rect 45185 632027 45251 632030
rect 675569 631410 675635 631413
rect 676070 631410 676076 631412
rect 675569 631408 676076 631410
rect 675569 631352 675574 631408
rect 675630 631352 676076 631408
rect 675569 631350 676076 631352
rect 675569 631347 675635 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 651557 630594 651623 630597
rect 650164 630592 651623 630594
rect 650164 630536 651562 630592
rect 651618 630536 651623 630592
rect 650164 630534 651623 630536
rect 651557 630531 651623 630534
rect 675477 626378 675543 626381
rect 675477 626376 676292 626378
rect 675477 626320 675482 626376
rect 675538 626320 676292 626376
rect 675477 626318 676292 626320
rect 675477 626315 675543 626318
rect 675109 625970 675175 625973
rect 675109 625968 676292 625970
rect 675109 625912 675114 625968
rect 675170 625912 676292 625968
rect 675109 625910 676292 625912
rect 675109 625907 675175 625910
rect 675477 625562 675543 625565
rect 675477 625560 676292 625562
rect 675477 625504 675482 625560
rect 675538 625504 676292 625560
rect 675477 625502 676292 625504
rect 675477 625499 675543 625502
rect 40902 625364 40908 625428
rect 40972 625426 40978 625428
rect 42333 625426 42399 625429
rect 40972 625424 42399 625426
rect 40972 625368 42338 625424
rect 42394 625368 42399 625424
rect 40972 625366 42399 625368
rect 40972 625364 40978 625366
rect 42333 625363 42399 625366
rect 672165 625154 672231 625157
rect 672942 625154 672948 625156
rect 672165 625152 672948 625154
rect 672165 625096 672170 625152
rect 672226 625096 672948 625152
rect 672165 625094 672948 625096
rect 672165 625091 672231 625094
rect 672942 625092 672948 625094
rect 673012 625092 673018 625156
rect 675477 625154 675543 625157
rect 675477 625152 676292 625154
rect 675477 625096 675482 625152
rect 675538 625096 676292 625152
rect 675477 625094 676292 625096
rect 675477 625091 675543 625094
rect 675477 624746 675543 624749
rect 675477 624744 676292 624746
rect 675477 624688 675482 624744
rect 675538 624688 676292 624744
rect 675477 624686 676292 624688
rect 675477 624683 675543 624686
rect 42149 624610 42215 624613
rect 42885 624610 42951 624613
rect 42149 624608 42951 624610
rect 42149 624552 42154 624608
rect 42210 624552 42890 624608
rect 42946 624552 42951 624608
rect 42149 624550 42951 624552
rect 42149 624547 42215 624550
rect 42885 624547 42951 624550
rect 675477 624338 675543 624341
rect 675477 624336 676292 624338
rect 675477 624280 675482 624336
rect 675538 624280 676292 624336
rect 675477 624278 676292 624280
rect 675477 624275 675543 624278
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 674833 623930 674899 623933
rect 674833 623928 676292 623930
rect 674833 623872 674838 623928
rect 674894 623872 676292 623928
rect 674833 623870 676292 623872
rect 674833 623867 674899 623870
rect 675477 623522 675543 623525
rect 675477 623520 676292 623522
rect 675477 623464 675482 623520
rect 675538 623464 676292 623520
rect 675477 623462 676292 623464
rect 675477 623459 675543 623462
rect 42149 623386 42215 623389
rect 43989 623386 44055 623389
rect 42149 623384 44055 623386
rect 42149 623328 42154 623384
rect 42210 623328 43994 623384
rect 44050 623328 44055 623384
rect 42149 623326 44055 623328
rect 42149 623323 42215 623326
rect 43989 623323 44055 623326
rect 675477 623114 675543 623117
rect 675477 623112 676292 623114
rect 675477 623056 675482 623112
rect 675538 623056 676292 623112
rect 675477 623054 676292 623056
rect 675477 623051 675543 623054
rect 675477 622706 675543 622709
rect 675477 622704 676292 622706
rect 675477 622648 675482 622704
rect 675538 622648 676292 622704
rect 675477 622646 676292 622648
rect 675477 622643 675543 622646
rect 675477 622298 675543 622301
rect 675477 622296 676292 622298
rect 675477 622240 675482 622296
rect 675538 622240 676292 622296
rect 675477 622238 676292 622240
rect 675477 622235 675543 622238
rect 682561 622026 682627 622029
rect 682518 622024 682627 622026
rect 682518 621968 682566 622024
rect 682622 621968 682627 622024
rect 682518 621963 682627 621968
rect 682518 621860 682578 621963
rect 682377 621618 682443 621621
rect 682334 621616 682443 621618
rect 682334 621560 682382 621616
rect 682438 621560 682443 621616
rect 682334 621555 682443 621560
rect 682334 621452 682394 621555
rect 674598 621012 674604 621076
rect 674668 621074 674674 621076
rect 674668 621014 676292 621074
rect 674668 621012 674674 621014
rect 42057 620938 42123 620941
rect 45185 620938 45251 620941
rect 42057 620936 45251 620938
rect 42057 620880 42062 620936
rect 42118 620880 45190 620936
rect 45246 620880 45251 620936
rect 42057 620878 45251 620880
rect 42057 620875 42123 620878
rect 45185 620875 45251 620878
rect 683297 620802 683363 620805
rect 683254 620800 683363 620802
rect 683254 620744 683302 620800
rect 683358 620744 683363 620800
rect 683254 620739 683363 620744
rect 683254 620636 683314 620739
rect 42057 620258 42123 620261
rect 42701 620258 42767 620261
rect 42057 620256 42767 620258
rect 42057 620200 42062 620256
rect 42118 620200 42706 620256
rect 42762 620200 42767 620256
rect 42057 620198 42767 620200
rect 42057 620195 42123 620198
rect 42701 620195 42767 620198
rect 675477 620258 675543 620261
rect 675477 620256 676292 620258
rect 675477 620200 675482 620256
rect 675538 620200 676292 620256
rect 675477 620198 676292 620200
rect 675477 620195 675543 620198
rect 40718 619788 40724 619852
rect 40788 619850 40794 619852
rect 42241 619850 42307 619853
rect 40788 619848 42307 619850
rect 40788 619792 42246 619848
rect 42302 619792 42307 619848
rect 40788 619790 42307 619792
rect 40788 619788 40794 619790
rect 42241 619787 42307 619790
rect 675017 619850 675083 619853
rect 675017 619848 676292 619850
rect 675017 619792 675022 619848
rect 675078 619792 676292 619848
rect 675017 619790 676292 619792
rect 675017 619787 675083 619790
rect 675477 619442 675543 619445
rect 675477 619440 676292 619442
rect 675477 619384 675482 619440
rect 675538 619384 676292 619440
rect 675477 619382 676292 619384
rect 675477 619379 675543 619382
rect 676806 619108 676812 619172
rect 676876 619108 676882 619172
rect 40534 618972 40540 619036
rect 40604 619034 40610 619036
rect 42425 619034 42491 619037
rect 40604 619032 42491 619034
rect 40604 618976 42430 619032
rect 42486 618976 42491 619032
rect 676814 619004 676874 619108
rect 40604 618974 42491 618976
rect 40604 618972 40610 618974
rect 42425 618971 42491 618974
rect 41822 618700 41828 618764
rect 41892 618762 41898 618764
rect 42701 618762 42767 618765
rect 41892 618760 42767 618762
rect 41892 618704 42706 618760
rect 42762 618704 42767 618760
rect 41892 618702 42767 618704
rect 41892 618700 41898 618702
rect 42701 618699 42767 618702
rect 673821 618626 673887 618629
rect 673821 618624 676292 618626
rect 673821 618568 673826 618624
rect 673882 618568 676292 618624
rect 673821 618566 676292 618568
rect 673821 618563 673887 618566
rect 675661 618218 675727 618221
rect 675661 618216 676292 618218
rect 675661 618160 675666 618216
rect 675722 618160 676292 618216
rect 675661 618158 676292 618160
rect 675661 618155 675727 618158
rect 674281 617810 674347 617813
rect 674281 617808 676292 617810
rect 674281 617752 674286 617808
rect 674342 617752 676292 617808
rect 674281 617750 676292 617752
rect 674281 617747 674347 617750
rect 674649 617402 674715 617405
rect 674649 617400 676292 617402
rect 674649 617344 674654 617400
rect 674710 617344 676292 617400
rect 674649 617342 676292 617344
rect 674649 617339 674715 617342
rect 651557 617266 651623 617269
rect 650164 617264 651623 617266
rect 650164 617208 651562 617264
rect 651618 617208 651623 617264
rect 650164 617206 651623 617208
rect 651557 617203 651623 617206
rect 675477 616994 675543 616997
rect 675477 616992 676292 616994
rect 675477 616936 675482 616992
rect 675538 616936 676292 616992
rect 675477 616934 676292 616936
rect 675477 616931 675543 616934
rect 675477 616586 675543 616589
rect 675477 616584 676292 616586
rect 675477 616528 675482 616584
rect 675538 616528 676292 616584
rect 675477 616526 676292 616528
rect 675477 616523 675543 616526
rect 675477 616178 675543 616181
rect 675477 616176 676292 616178
rect 675477 616120 675482 616176
rect 675538 616120 676292 616176
rect 675477 616118 676292 616120
rect 675477 616115 675543 616118
rect 41454 615980 41460 616044
rect 41524 616042 41530 616044
rect 42241 616042 42307 616045
rect 41524 616040 42307 616042
rect 41524 615984 42246 616040
rect 42302 615984 42307 616040
rect 41524 615982 42307 615984
rect 41524 615980 41530 615982
rect 42241 615979 42307 615982
rect 667841 615906 667907 615909
rect 675845 615906 675911 615909
rect 667841 615904 675911 615906
rect 667841 615848 667846 615904
rect 667902 615848 675850 615904
rect 675906 615848 675911 615904
rect 667841 615846 675911 615848
rect 667841 615843 667907 615846
rect 675845 615843 675911 615846
rect 683070 615501 683130 615740
rect 683070 615498 683179 615501
rect 683070 615496 683260 615498
rect 683070 615440 683118 615496
rect 683174 615440 683260 615496
rect 683070 615438 683260 615440
rect 683070 615435 683179 615438
rect 683070 615332 683130 615435
rect 675477 614954 675543 614957
rect 675477 614952 676292 614954
rect 675477 614896 675482 614952
rect 675538 614896 676292 614952
rect 675477 614894 676292 614896
rect 675477 614891 675543 614894
rect 41781 612780 41847 612781
rect 41781 612776 41828 612780
rect 41892 612778 41898 612780
rect 41781 612720 41786 612776
rect 41781 612716 41828 612720
rect 41892 612718 41938 612778
rect 41892 612716 41898 612718
rect 41781 612715 41847 612716
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 674230 607820 674236 607884
rect 674300 607882 674306 607884
rect 675385 607882 675451 607885
rect 674300 607880 675451 607882
rect 674300 607824 675390 607880
rect 675446 607824 675451 607880
rect 674300 607822 675451 607824
rect 674300 607820 674306 607822
rect 675385 607819 675451 607822
rect 675753 607338 675819 607341
rect 677174 607338 677180 607340
rect 675753 607336 677180 607338
rect 675753 607280 675758 607336
rect 675814 607280 677180 607336
rect 675753 607278 677180 607280
rect 675753 607275 675819 607278
rect 677174 607276 677180 607278
rect 677244 607276 677250 607340
rect 670141 607202 670207 607205
rect 670141 607200 670434 607202
rect 670141 607144 670146 607200
rect 670202 607144 670434 607200
rect 670141 607142 670434 607144
rect 670141 607139 670207 607142
rect 670374 606933 670434 607142
rect 670325 606928 670434 606933
rect 670325 606872 670330 606928
rect 670386 606872 670434 606928
rect 670325 606870 670434 606872
rect 670325 606867 670391 606870
rect 652569 603938 652635 603941
rect 650164 603936 652635 603938
rect 650164 603880 652574 603936
rect 652630 603880 652635 603936
rect 650164 603878 652635 603880
rect 652569 603875 652635 603878
rect 674598 602924 674604 602988
rect 674668 602986 674674 602988
rect 675293 602986 675359 602989
rect 674668 602984 675359 602986
rect 674668 602928 675298 602984
rect 675354 602928 675359 602984
rect 674668 602926 675359 602928
rect 674668 602924 674674 602926
rect 675293 602923 675359 602926
rect 35801 601762 35867 601765
rect 35788 601760 35867 601762
rect 35788 601704 35806 601760
rect 35862 601704 35867 601760
rect 35788 601702 35867 601704
rect 35801 601699 35867 601702
rect 47761 601354 47827 601357
rect 41492 601352 47827 601354
rect 41492 601296 47766 601352
rect 47822 601296 47827 601352
rect 41492 601294 47827 601296
rect 47761 601291 47827 601294
rect 674833 601218 674899 601221
rect 675385 601218 675451 601221
rect 674833 601216 675451 601218
rect 674833 601160 674838 601216
rect 674894 601160 675390 601216
rect 675446 601160 675451 601216
rect 674833 601158 675451 601160
rect 674833 601155 674899 601158
rect 675385 601155 675451 601158
rect 43805 600946 43871 600949
rect 41492 600944 43871 600946
rect 41492 600888 43810 600944
rect 43866 600888 43871 600944
rect 41492 600886 43871 600888
rect 43805 600883 43871 600886
rect 44541 600538 44607 600541
rect 41492 600536 44607 600538
rect 41492 600480 44546 600536
rect 44602 600480 44607 600536
rect 41492 600478 44607 600480
rect 44541 600475 44607 600478
rect 44357 600130 44423 600133
rect 41492 600128 44423 600130
rect 41492 600072 44362 600128
rect 44418 600072 44423 600128
rect 41492 600070 44423 600072
rect 44357 600067 44423 600070
rect 44173 599722 44239 599725
rect 41492 599720 44239 599722
rect 41492 599664 44178 599720
rect 44234 599664 44239 599720
rect 41492 599662 44239 599664
rect 44173 599659 44239 599662
rect 41321 599314 41387 599317
rect 41308 599312 41387 599314
rect 41308 599256 41326 599312
rect 41382 599256 41387 599312
rect 41308 599254 41387 599256
rect 41321 599251 41387 599254
rect 673913 599178 673979 599181
rect 675477 599178 675543 599181
rect 673913 599176 675543 599178
rect 673913 599120 673918 599176
rect 673974 599120 675482 599176
rect 675538 599120 675543 599176
rect 673913 599118 675543 599120
rect 673913 599115 673979 599118
rect 675477 599115 675543 599118
rect 40861 598906 40927 598909
rect 40861 598904 40940 598906
rect 40861 598848 40866 598904
rect 40922 598848 40940 598904
rect 40861 598846 40940 598848
rect 40861 598843 40927 598846
rect 42701 598498 42767 598501
rect 41492 598496 42767 598498
rect 41492 598440 42706 598496
rect 42762 598440 42767 598496
rect 41492 598438 42767 598440
rect 42701 598435 42767 598438
rect 672717 598498 672783 598501
rect 675477 598498 675543 598501
rect 672717 598496 675543 598498
rect 672717 598440 672722 598496
rect 672778 598440 675482 598496
rect 675538 598440 675543 598496
rect 672717 598438 675543 598440
rect 672717 598435 672783 598438
rect 675477 598435 675543 598438
rect 41094 597855 41154 598060
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 41045 597850 41154 597855
rect 41321 597852 41387 597855
rect 41045 597794 41050 597850
rect 41106 597794 41154 597850
rect 41045 597792 41154 597794
rect 41278 597850 41387 597852
rect 41278 597794 41326 597850
rect 41382 597794 41387 597850
rect 41045 597789 41111 597792
rect 41278 597789 41387 597794
rect 41278 597652 41338 597789
rect 674925 597684 674991 597685
rect 674925 597682 674972 597684
rect 674880 597680 674972 597682
rect 674880 597624 674930 597680
rect 674880 597622 674972 597624
rect 674925 597620 674972 597622
rect 675036 597620 675042 597684
rect 674925 597619 674991 597620
rect 673821 597410 673887 597413
rect 675477 597410 675543 597413
rect 673821 597408 675543 597410
rect 673821 597352 673826 597408
rect 673882 597352 675482 597408
rect 675538 597352 675543 597408
rect 673821 597350 675543 597352
rect 673821 597347 673887 597350
rect 675477 597347 675543 597350
rect 41137 597274 41203 597277
rect 41124 597272 41203 597274
rect 41124 597216 41142 597272
rect 41198 597216 41203 597272
rect 41124 597214 41203 597216
rect 41137 597211 41203 597214
rect 42241 596866 42307 596869
rect 41492 596864 42307 596866
rect 41492 596808 42246 596864
rect 42302 596808 42307 596864
rect 41492 596806 42307 596808
rect 42241 596803 42307 596806
rect 42190 596458 42196 596460
rect 41492 596398 42196 596458
rect 42190 596396 42196 596398
rect 42260 596396 42266 596460
rect 42057 596050 42123 596053
rect 41492 596048 42123 596050
rect 41492 595992 42062 596048
rect 42118 595992 42123 596048
rect 41492 595990 42123 595992
rect 42057 595987 42123 595990
rect 41689 595778 41755 595781
rect 42006 595778 42012 595780
rect 41689 595776 42012 595778
rect 41689 595720 41694 595776
rect 41750 595720 42012 595776
rect 41689 595718 42012 595720
rect 41689 595715 41755 595718
rect 42006 595716 42012 595718
rect 42076 595716 42082 595780
rect 33041 595642 33107 595645
rect 33028 595640 33107 595642
rect 33028 595584 33046 595640
rect 33102 595584 33107 595640
rect 33028 595582 33107 595584
rect 33041 595579 33107 595582
rect 35157 595234 35223 595237
rect 35157 595232 35236 595234
rect 35157 595176 35162 595232
rect 35218 595176 35236 595232
rect 35157 595174 35236 595176
rect 35157 595171 35223 595174
rect 34421 594826 34487 594829
rect 34421 594824 34500 594826
rect 34421 594768 34426 594824
rect 34482 594768 34500 594824
rect 34421 594766 34500 594768
rect 675477 594824 675543 594829
rect 675477 594768 675482 594824
rect 675538 594768 675543 594824
rect 34421 594763 34487 594766
rect 675477 594763 675543 594768
rect 675017 594554 675083 594557
rect 675480 594554 675540 594763
rect 675017 594552 675540 594554
rect 675017 594496 675022 594552
rect 675078 594496 675540 594552
rect 675017 594494 675540 594496
rect 675017 594491 675083 594494
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 41822 594010 41828 594012
rect 41492 593950 41828 594010
rect 41822 593948 41828 593950
rect 41892 593948 41898 594012
rect 36537 593602 36603 593605
rect 36524 593600 36603 593602
rect 36524 593544 36542 593600
rect 36598 593544 36603 593600
rect 36524 593542 36603 593544
rect 36537 593539 36603 593542
rect 42977 593194 43043 593197
rect 41492 593192 43043 593194
rect 41492 593136 42982 593192
rect 43038 593136 43043 593192
rect 41492 593134 43043 593136
rect 42977 593131 43043 593134
rect 41689 592922 41755 592925
rect 41646 592920 41755 592922
rect 41646 592864 41694 592920
rect 41750 592864 41755 592920
rect 41646 592859 41755 592864
rect 673453 592922 673519 592925
rect 675845 592922 675911 592925
rect 673453 592920 675911 592922
rect 673453 592864 673458 592920
rect 673514 592864 675850 592920
rect 675906 592864 675911 592920
rect 673453 592862 675911 592864
rect 673453 592859 673519 592862
rect 675845 592859 675911 592862
rect 41646 592820 41706 592859
rect 41462 592760 41706 592820
rect 41462 592756 41522 592760
rect 674966 592452 674972 592516
rect 675036 592514 675042 592516
rect 675845 592514 675911 592517
rect 675036 592512 675911 592514
rect 675036 592456 675850 592512
rect 675906 592456 675911 592512
rect 675036 592454 675911 592456
rect 675036 592452 675042 592454
rect 675845 592451 675911 592454
rect 41781 592378 41847 592381
rect 41492 592376 41847 592378
rect 41492 592320 41786 592376
rect 41842 592320 41847 592376
rect 41492 592318 41847 592320
rect 41781 592315 41847 592318
rect 674465 592242 674531 592245
rect 675845 592242 675911 592245
rect 674465 592240 675911 592242
rect 674465 592184 674470 592240
rect 674526 592184 675850 592240
rect 675906 592184 675911 592240
rect 674465 592182 675911 592184
rect 674465 592179 674531 592182
rect 675845 592179 675911 592182
rect 44633 591970 44699 591973
rect 41492 591968 44699 591970
rect 41492 591912 44638 591968
rect 44694 591912 44699 591968
rect 41492 591910 44699 591912
rect 44633 591907 44699 591910
rect 43253 591562 43319 591565
rect 41492 591560 43319 591562
rect 41492 591504 43258 591560
rect 43314 591504 43319 591560
rect 41492 591502 43319 591504
rect 43253 591499 43319 591502
rect 674189 591290 674255 591293
rect 675845 591290 675911 591293
rect 674189 591288 675911 591290
rect 674189 591232 674194 591288
rect 674250 591232 675850 591288
rect 675906 591232 675911 591288
rect 674189 591230 675911 591232
rect 674189 591227 674255 591230
rect 675845 591227 675911 591230
rect 39990 590749 40050 591124
rect 39941 590744 40050 590749
rect 651557 590746 651623 590749
rect 39941 590688 39946 590744
rect 40002 590716 40050 590744
rect 650164 590744 651623 590746
rect 40002 590688 40020 590716
rect 39941 590686 40020 590688
rect 650164 590688 651562 590744
rect 651618 590688 651623 590744
rect 650164 590686 651623 590688
rect 39941 590683 40007 590686
rect 651557 590683 651623 590686
rect 47761 590338 47827 590341
rect 41492 590336 47827 590338
rect 41492 590280 47766 590336
rect 47822 590280 47827 590336
rect 41492 590278 47827 590280
rect 47761 590275 47827 590278
rect 40769 589660 40835 589661
rect 40718 589658 40724 589660
rect 40678 589598 40724 589658
rect 40788 589656 40835 589660
rect 40830 589600 40835 589656
rect 40718 589596 40724 589598
rect 40788 589596 40835 589600
rect 40769 589595 40835 589596
rect 40902 589460 40908 589524
rect 40972 589522 40978 589524
rect 41781 589522 41847 589525
rect 40972 589520 41847 589522
rect 40972 589464 41786 589520
rect 41842 589464 41847 589520
rect 40972 589462 41847 589464
rect 40972 589460 40978 589462
rect 41781 589459 41847 589462
rect 676070 589188 676076 589252
rect 676140 589250 676146 589252
rect 682377 589250 682443 589253
rect 676140 589248 682443 589250
rect 676140 589192 682382 589248
rect 682438 589192 682443 589248
rect 676140 589190 682443 589192
rect 676140 589188 676146 589190
rect 682377 589187 682443 589190
rect 34421 587210 34487 587213
rect 41822 587210 41828 587212
rect 34421 587208 41828 587210
rect 34421 587152 34426 587208
rect 34482 587152 41828 587208
rect 34421 587150 41828 587152
rect 34421 587147 34487 587150
rect 41822 587148 41828 587150
rect 41892 587148 41898 587212
rect 39573 586666 39639 586669
rect 42190 586666 42196 586668
rect 39573 586664 42196 586666
rect 39573 586608 39578 586664
rect 39634 586608 42196 586664
rect 39573 586606 42196 586608
rect 39573 586603 39639 586606
rect 42190 586604 42196 586606
rect 42260 586604 42266 586668
rect 672349 586258 672415 586261
rect 672942 586258 672948 586260
rect 672349 586256 672948 586258
rect 672349 586200 672354 586256
rect 672410 586200 672948 586256
rect 672349 586198 672948 586200
rect 672349 586195 672415 586198
rect 672942 586196 672948 586198
rect 673012 586196 673018 586260
rect 675293 586258 675359 586261
rect 676070 586258 676076 586260
rect 675293 586256 676076 586258
rect 675293 586200 675298 586256
rect 675354 586200 676076 586256
rect 675293 586198 676076 586200
rect 675293 586195 675359 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 39573 585850 39639 585853
rect 41086 585850 41092 585852
rect 39573 585848 41092 585850
rect 39573 585792 39578 585848
rect 39634 585792 41092 585848
rect 39573 585790 41092 585792
rect 39573 585787 39639 585790
rect 41086 585788 41092 585790
rect 41156 585788 41162 585852
rect 39941 585578 40007 585581
rect 41270 585578 41276 585580
rect 39941 585576 41276 585578
rect 39941 585520 39946 585576
rect 40002 585520 41276 585576
rect 39941 585518 41276 585520
rect 39941 585515 40007 585518
rect 41270 585516 41276 585518
rect 41340 585516 41346 585580
rect 42425 585444 42491 585445
rect 42374 585380 42380 585444
rect 42444 585442 42491 585444
rect 42444 585440 42536 585442
rect 42486 585384 42536 585440
rect 42444 585382 42536 585384
rect 42444 585380 42491 585382
rect 42425 585379 42491 585380
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 40493 584762 40559 584765
rect 42057 584762 42123 584765
rect 40493 584760 42123 584762
rect 40493 584704 40498 584760
rect 40554 584704 42062 584760
rect 42118 584704 42123 584760
rect 40493 584702 42123 584704
rect 40493 584699 40559 584702
rect 42057 584699 42123 584702
rect 39665 584626 39731 584629
rect 40350 584626 40356 584628
rect 39665 584624 40356 584626
rect 39665 584568 39670 584624
rect 39726 584568 40356 584624
rect 39665 584566 40356 584568
rect 39665 584563 39731 584566
rect 40350 584564 40356 584566
rect 40420 584564 40426 584628
rect 41270 582524 41276 582588
rect 41340 582586 41346 582588
rect 41781 582586 41847 582589
rect 41340 582584 41847 582586
rect 41340 582528 41786 582584
rect 41842 582528 41847 582584
rect 41340 582526 41847 582528
rect 41340 582524 41346 582526
rect 41781 582523 41847 582526
rect 42425 581636 42491 581637
rect 42374 581572 42380 581636
rect 42444 581634 42491 581636
rect 42444 581632 42536 581634
rect 42486 581576 42536 581632
rect 42444 581574 42536 581576
rect 42444 581572 42491 581574
rect 42425 581571 42491 581572
rect 41086 581436 41092 581500
rect 41156 581498 41162 581500
rect 42241 581498 42307 581501
rect 41156 581496 42307 581498
rect 41156 581440 42246 581496
rect 42302 581440 42307 581496
rect 41156 581438 42307 581440
rect 41156 581436 41162 581438
rect 42241 581435 42307 581438
rect 42057 581226 42123 581229
rect 43437 581226 43503 581229
rect 42057 581224 43503 581226
rect 42057 581168 42062 581224
rect 42118 581168 43442 581224
rect 43498 581168 43503 581224
rect 42057 581166 43503 581168
rect 42057 581163 42123 581166
rect 43437 581163 43503 581166
rect 675477 581090 675543 581093
rect 675477 581088 676292 581090
rect 675477 581032 675482 581088
rect 675538 581032 676292 581088
rect 675477 581030 676292 581032
rect 675477 581027 675543 581030
rect 674925 580682 674991 580685
rect 674925 580680 676292 580682
rect 674925 580624 674930 580680
rect 674986 580624 676292 580680
rect 674925 580622 676292 580624
rect 674925 580619 674991 580622
rect 675293 580274 675359 580277
rect 675293 580272 676292 580274
rect 675293 580216 675298 580272
rect 675354 580216 676292 580272
rect 675293 580214 676292 580216
rect 675293 580211 675359 580214
rect 40902 580076 40908 580140
rect 40972 580138 40978 580140
rect 42241 580138 42307 580141
rect 40972 580136 42307 580138
rect 40972 580080 42246 580136
rect 42302 580080 42307 580136
rect 40972 580078 42307 580080
rect 40972 580076 40978 580078
rect 42241 580075 42307 580078
rect 40350 579804 40356 579868
rect 40420 579866 40426 579868
rect 42609 579866 42675 579869
rect 40420 579864 42675 579866
rect 40420 579808 42614 579864
rect 42670 579808 42675 579864
rect 40420 579806 42675 579808
rect 40420 579804 40426 579806
rect 42609 579803 42675 579806
rect 675477 579866 675543 579869
rect 675477 579864 676292 579866
rect 675477 579808 675482 579864
rect 675538 579808 676292 579864
rect 675477 579806 676292 579808
rect 675477 579803 675543 579806
rect 40718 579532 40724 579596
rect 40788 579594 40794 579596
rect 42374 579594 42380 579596
rect 40788 579534 42380 579594
rect 40788 579532 40794 579534
rect 42374 579532 42380 579534
rect 42444 579532 42450 579596
rect 674925 579458 674991 579461
rect 674925 579456 676292 579458
rect 674925 579400 674930 579456
rect 674986 579400 676292 579456
rect 674925 579398 676292 579400
rect 674925 579395 674991 579398
rect 675293 579050 675359 579053
rect 675293 579048 676292 579050
rect 675293 578992 675298 579048
rect 675354 578992 676292 579048
rect 675293 578990 676292 578992
rect 675293 578987 675359 578990
rect 42057 578914 42123 578917
rect 43161 578914 43227 578917
rect 42057 578912 43227 578914
rect 42057 578856 42062 578912
rect 42118 578856 43166 578912
rect 43222 578856 43227 578912
rect 42057 578854 43227 578856
rect 42057 578851 42123 578854
rect 43161 578851 43227 578854
rect 675477 578642 675543 578645
rect 675477 578640 676292 578642
rect 675477 578584 675482 578640
rect 675538 578584 676292 578640
rect 675477 578582 676292 578584
rect 675477 578579 675543 578582
rect 42149 578234 42215 578237
rect 42977 578234 43043 578237
rect 42149 578232 43043 578234
rect 42149 578176 42154 578232
rect 42210 578176 42982 578232
rect 43038 578176 43043 578232
rect 42149 578174 43043 578176
rect 42149 578171 42215 578174
rect 42977 578171 43043 578174
rect 675477 578234 675543 578237
rect 675477 578232 676292 578234
rect 675477 578176 675482 578232
rect 675538 578176 676292 578232
rect 675477 578174 676292 578176
rect 675477 578171 675543 578174
rect 675293 577826 675359 577829
rect 675293 577824 676292 577826
rect 675293 577768 675298 577824
rect 675354 577768 676292 577824
rect 675293 577766 676292 577768
rect 675293 577763 675359 577766
rect 651557 577418 651623 577421
rect 650164 577416 651623 577418
rect 650164 577360 651562 577416
rect 651618 577360 651623 577416
rect 650164 577358 651623 577360
rect 651557 577355 651623 577358
rect 675477 577418 675543 577421
rect 675477 577416 676292 577418
rect 675477 577360 675482 577416
rect 675538 577360 676292 577416
rect 675477 577358 676292 577360
rect 675477 577355 675543 577358
rect 42149 577012 42215 577013
rect 42149 577010 42196 577012
rect 42104 577008 42196 577010
rect 42104 576952 42154 577008
rect 42104 576950 42196 576952
rect 42149 576948 42196 576950
rect 42260 576948 42266 577012
rect 675477 577010 675543 577013
rect 675477 577008 676292 577010
rect 675477 576952 675482 577008
rect 675538 576952 676292 577008
rect 675477 576950 676292 576952
rect 42149 576947 42215 576948
rect 675477 576947 675543 576950
rect 675477 576602 675543 576605
rect 675477 576600 676292 576602
rect 675477 576544 675482 576600
rect 675538 576544 676292 576600
rect 675477 576542 676292 576544
rect 675477 576539 675543 576542
rect 683297 576466 683363 576469
rect 683254 576464 683363 576466
rect 683254 576408 683302 576464
rect 683358 576408 683363 576464
rect 683254 576403 683363 576408
rect 683254 576164 683314 576403
rect 682377 576058 682443 576061
rect 682334 576056 682443 576058
rect 682334 576000 682382 576056
rect 682438 576000 682443 576056
rect 682334 575995 682443 576000
rect 682334 575756 682394 575995
rect 40534 575588 40540 575652
rect 40604 575650 40610 575652
rect 42241 575650 42307 575653
rect 40604 575648 42307 575650
rect 40604 575592 42246 575648
rect 42302 575592 42307 575648
rect 40604 575590 42307 575592
rect 40604 575588 40610 575590
rect 42241 575587 42307 575590
rect 678237 575650 678303 575653
rect 678237 575648 678346 575650
rect 678237 575592 678242 575648
rect 678298 575592 678346 575648
rect 678237 575587 678346 575592
rect 678286 575348 678346 575587
rect 675477 574970 675543 574973
rect 675477 574968 676292 574970
rect 675477 574912 675482 574968
rect 675538 574912 676292 574968
rect 675477 574910 676292 574912
rect 675477 574907 675543 574910
rect 42057 574698 42123 574701
rect 42374 574698 42380 574700
rect 42057 574696 42380 574698
rect 42057 574640 42062 574696
rect 42118 574640 42380 574696
rect 42057 574638 42380 574640
rect 42057 574635 42123 574638
rect 42374 574636 42380 574638
rect 42444 574636 42450 574700
rect 675293 574562 675359 574565
rect 675293 574560 676292 574562
rect 675293 574504 675298 574560
rect 675354 574504 676292 574560
rect 675293 574502 676292 574504
rect 675293 574499 675359 574502
rect 675477 574154 675543 574157
rect 675477 574152 676292 574154
rect 675477 574096 675482 574152
rect 675538 574096 676292 574152
rect 675477 574094 676292 574096
rect 675477 574091 675543 574094
rect 675293 573746 675359 573749
rect 675293 573744 676292 573746
rect 675293 573688 675298 573744
rect 675354 573688 676292 573744
rect 675293 573686 676292 573688
rect 675293 573683 675359 573686
rect 674414 573276 674420 573340
rect 674484 573338 674490 573340
rect 674484 573278 676292 573338
rect 674484 573276 674490 573278
rect 675477 572930 675543 572933
rect 675477 572928 676292 572930
rect 675477 572872 675482 572928
rect 675538 572872 676292 572928
rect 675477 572870 676292 572872
rect 675477 572867 675543 572870
rect 41454 572732 41460 572796
rect 41524 572794 41530 572796
rect 42609 572794 42675 572797
rect 41524 572792 42675 572794
rect 41524 572736 42614 572792
rect 42670 572736 42675 572792
rect 41524 572734 42675 572736
rect 41524 572732 41530 572734
rect 42609 572731 42675 572734
rect 684125 572794 684191 572797
rect 684125 572792 684234 572794
rect 684125 572736 684130 572792
rect 684186 572736 684234 572792
rect 684125 572731 684234 572736
rect 684174 572492 684234 572731
rect 41638 572052 41644 572116
rect 41708 572114 41714 572116
rect 42517 572114 42583 572117
rect 41708 572112 42583 572114
rect 41708 572056 42522 572112
rect 42578 572056 42583 572112
rect 41708 572054 42583 572056
rect 41708 572052 41714 572054
rect 42517 572051 42583 572054
rect 669221 572114 669287 572117
rect 669221 572112 676292 572114
rect 669221 572056 669226 572112
rect 669282 572056 676292 572112
rect 669221 572054 676292 572056
rect 669221 572051 669287 572054
rect 683481 571978 683547 571981
rect 683438 571976 683547 571978
rect 683438 571920 683486 571976
rect 683542 571920 683547 571976
rect 683438 571915 683547 571920
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 683438 571676 683498 571915
rect 675293 571298 675359 571301
rect 675293 571296 676292 571298
rect 675293 571240 675298 571296
rect 675354 571240 676292 571296
rect 675293 571238 676292 571240
rect 675293 571235 675359 571238
rect 676262 570757 676322 570860
rect 676213 570752 676322 570757
rect 676213 570696 676218 570752
rect 676274 570696 676322 570752
rect 676213 570694 676322 570696
rect 676213 570691 676279 570694
rect 682886 570346 682946 570452
rect 683113 570346 683179 570349
rect 682886 570344 683179 570346
rect 682886 570288 683118 570344
rect 683174 570288 683179 570344
rect 682886 570286 683179 570288
rect 41781 570212 41847 570213
rect 41781 570208 41828 570212
rect 41892 570210 41898 570212
rect 41781 570152 41786 570208
rect 41781 570148 41828 570152
rect 41892 570150 41938 570210
rect 41892 570148 41898 570150
rect 41781 570147 41847 570148
rect 682886 570044 682946 570286
rect 683113 570283 683179 570286
rect 675477 569666 675543 569669
rect 675477 569664 676292 569666
rect 675477 569608 675482 569664
rect 675538 569608 676292 569664
rect 675477 569606 676292 569608
rect 675477 569603 675543 569606
rect 652385 564090 652451 564093
rect 650164 564088 652451 564090
rect 650164 564032 652390 564088
rect 652446 564032 652451 564088
rect 650164 564030 652451 564032
rect 652385 564027 652451 564030
rect 668761 563954 668827 563957
rect 675845 563954 675911 563957
rect 668761 563952 675911 563954
rect 668761 563896 668766 563952
rect 668822 563896 675850 563952
rect 675906 563896 675911 563952
rect 668761 563894 675911 563896
rect 668761 563891 668827 563894
rect 675845 563891 675911 563894
rect 675385 561916 675451 561917
rect 675334 561914 675340 561916
rect 675294 561854 675340 561914
rect 675404 561912 675451 561916
rect 675446 561856 675451 561912
rect 675334 561852 675340 561854
rect 675404 561852 675451 561856
rect 675385 561851 675451 561852
rect 675477 559468 675543 559469
rect 675477 559464 675524 559468
rect 675588 559466 675594 559468
rect 675477 559408 675482 559464
rect 675477 559404 675524 559408
rect 675588 559406 675634 559466
rect 675588 559404 675594 559406
rect 675477 559403 675543 559404
rect 675753 559058 675819 559061
rect 676806 559058 676812 559060
rect 675753 559056 676812 559058
rect 675753 559000 675758 559056
rect 675814 559000 676812 559056
rect 675753 558998 676812 559000
rect 675753 558995 675819 558998
rect 676806 558996 676812 558998
rect 676876 558996 676882 559060
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 43253 558514 43319 558517
rect 41492 558512 43319 558514
rect 41492 558456 43258 558512
rect 43314 558456 43319 558512
rect 41492 558454 43319 558456
rect 43253 558451 43319 558454
rect 43437 558106 43503 558109
rect 41492 558104 43503 558106
rect 41492 558048 43442 558104
rect 43498 558048 43503 558104
rect 41492 558046 43503 558048
rect 43437 558043 43503 558046
rect 43437 557698 43503 557701
rect 41492 557696 43503 557698
rect 41492 557640 43442 557696
rect 43498 557640 43503 557696
rect 41492 557638 43503 557640
rect 43437 557635 43503 557638
rect 44265 557290 44331 557293
rect 41492 557288 44331 557290
rect 41492 557232 44270 557288
rect 44326 557232 44331 557288
rect 41492 557230 44331 557232
rect 44265 557227 44331 557230
rect 44633 556882 44699 556885
rect 41492 556880 44699 556882
rect 41492 556824 44638 556880
rect 44694 556824 44699 556880
rect 41492 556822 44699 556824
rect 44633 556819 44699 556822
rect 44449 556474 44515 556477
rect 41492 556472 44515 556474
rect 41492 556416 44454 556472
rect 44510 556416 44515 556472
rect 41492 556414 44515 556416
rect 44449 556411 44515 556414
rect 40585 556066 40651 556069
rect 40572 556064 40651 556066
rect 40572 556008 40590 556064
rect 40646 556008 40651 556064
rect 40572 556006 40651 556008
rect 40585 556003 40651 556006
rect 40861 555658 40927 555661
rect 40861 555656 40940 555658
rect 40861 555600 40866 555656
rect 40922 555600 40940 555656
rect 40861 555598 40940 555600
rect 40861 555595 40927 555598
rect 42977 555250 43043 555253
rect 41492 555248 43043 555250
rect 41492 555192 42982 555248
rect 43038 555192 43043 555248
rect 41492 555190 43043 555192
rect 42977 555187 43043 555190
rect 43805 554842 43871 554845
rect 41492 554840 43871 554842
rect 41492 554784 43810 554840
rect 43866 554784 43871 554840
rect 41492 554782 43871 554784
rect 43805 554779 43871 554782
rect 43805 554434 43871 554437
rect 41492 554432 43871 554434
rect 41492 554376 43810 554432
rect 43866 554376 43871 554432
rect 41492 554374 43871 554376
rect 43805 554371 43871 554374
rect 42190 554026 42196 554028
rect 41492 553966 42196 554026
rect 42190 553964 42196 553966
rect 42260 553964 42266 554028
rect 39990 553413 40050 553588
rect 671981 553482 672047 553485
rect 675385 553482 675451 553485
rect 671981 553480 675451 553482
rect 671981 553424 671986 553480
rect 672042 553424 675390 553480
rect 675446 553424 675451 553480
rect 671981 553422 675451 553424
rect 671981 553419 672047 553422
rect 675385 553419 675451 553422
rect 39990 553408 40099 553413
rect 39990 553352 40038 553408
rect 40094 553352 40099 553408
rect 39990 553350 40099 553352
rect 40033 553347 40099 553350
rect 40861 553410 40927 553413
rect 40861 553408 40970 553410
rect 40861 553352 40866 553408
rect 40922 553352 40970 553408
rect 40861 553347 40970 553352
rect 40910 553180 40970 553347
rect 42374 552802 42380 552804
rect 41492 552742 42380 552802
rect 42374 552740 42380 552742
rect 42444 552740 42450 552804
rect 45369 552394 45435 552397
rect 41492 552392 45435 552394
rect 41492 552336 45374 552392
rect 45430 552336 45435 552392
rect 41492 552334 45435 552336
rect 45369 552331 45435 552334
rect 675753 552122 675819 552125
rect 676990 552122 676996 552124
rect 675753 552120 676996 552122
rect 675753 552064 675758 552120
rect 675814 552064 676996 552120
rect 675753 552062 676996 552064
rect 675753 552059 675819 552062
rect 676990 552060 676996 552062
rect 677060 552060 677066 552124
rect 34421 551986 34487 551989
rect 34421 551984 34500 551986
rect 34421 551928 34426 551984
rect 34482 551928 34500 551984
rect 34421 551926 34500 551928
rect 34421 551923 34487 551926
rect 43345 551578 43411 551581
rect 41492 551576 43411 551578
rect 41492 551520 43350 551576
rect 43406 551520 43411 551576
rect 41492 551518 43411 551520
rect 43345 551515 43411 551518
rect 45185 551170 45251 551173
rect 41492 551168 45251 551170
rect 41492 551112 45190 551168
rect 45246 551112 45251 551168
rect 41492 551110 45251 551112
rect 45185 551107 45251 551110
rect 651557 550898 651623 550901
rect 650164 550896 651623 550898
rect 650164 550840 651562 550896
rect 651618 550840 651623 550896
rect 650164 550838 651623 550840
rect 651557 550835 651623 550838
rect 41492 550702 41890 550762
rect 41830 550629 41890 550702
rect 41830 550624 41939 550629
rect 41830 550568 41878 550624
rect 41934 550568 41939 550624
rect 41830 550566 41939 550568
rect 41873 550563 41939 550566
rect 42006 550354 42012 550356
rect 41492 550294 42012 550354
rect 42006 550292 42012 550294
rect 42076 550292 42082 550356
rect 42149 549946 42215 549949
rect 41492 549944 42215 549946
rect 41492 549888 42154 549944
rect 42210 549888 42215 549944
rect 41492 549886 42215 549888
rect 42149 549883 42215 549886
rect 675477 549676 675543 549677
rect 675477 549674 675524 549676
rect 675432 549672 675524 549674
rect 675432 549616 675482 549672
rect 675432 549614 675524 549616
rect 675477 549612 675524 549614
rect 675588 549612 675594 549676
rect 675477 549611 675543 549612
rect 41965 549538 42031 549541
rect 41492 549536 42031 549538
rect 41492 549480 41970 549536
rect 42026 549480 42031 549536
rect 41492 549478 42031 549480
rect 41965 549475 42031 549478
rect 43989 549130 44055 549133
rect 41492 549128 44055 549130
rect 41492 549072 43994 549128
rect 44050 549072 44055 549128
rect 41492 549070 44055 549072
rect 43989 549067 44055 549070
rect 44173 548722 44239 548725
rect 41492 548720 44239 548722
rect 41492 548664 44178 548720
rect 44234 548664 44239 548720
rect 41492 548662 44239 548664
rect 44173 548659 44239 548662
rect 670233 548450 670299 548453
rect 675477 548450 675543 548453
rect 670233 548448 675543 548450
rect 670233 548392 670238 548448
rect 670294 548392 675482 548448
rect 675538 548392 675543 548448
rect 670233 548390 675543 548392
rect 670233 548387 670299 548390
rect 675477 548387 675543 548390
rect 41094 548147 41154 548284
rect 41094 548142 41203 548147
rect 41094 548086 41142 548142
rect 41198 548086 41203 548142
rect 41094 548084 41203 548086
rect 41137 548081 41203 548084
rect 28766 547498 28826 547890
rect 675334 547844 675340 547908
rect 675404 547906 675410 547908
rect 675753 547906 675819 547909
rect 675404 547904 675819 547906
rect 675404 547848 675758 547904
rect 675814 547848 675819 547904
rect 675404 547846 675819 547848
rect 675404 547844 675410 547846
rect 675753 547843 675819 547846
rect 41689 547770 41755 547773
rect 43437 547770 43503 547773
rect 41689 547768 43503 547770
rect 41689 547712 41694 547768
rect 41750 547712 43442 547768
rect 43498 547712 43503 547768
rect 41689 547710 43503 547712
rect 41689 547707 41755 547710
rect 43437 547707 43503 547710
rect 674925 547634 674991 547637
rect 675937 547634 676003 547637
rect 674925 547632 676003 547634
rect 674925 547576 674930 547632
rect 674986 547576 675942 547632
rect 675998 547576 676003 547632
rect 674925 547574 676003 547576
rect 674925 547571 674991 547574
rect 675937 547571 676003 547574
rect 677174 547572 677180 547636
rect 677244 547634 677250 547636
rect 677501 547634 677567 547637
rect 677244 547632 677567 547634
rect 677244 547576 677506 547632
rect 677562 547576 677567 547632
rect 677244 547574 677567 547576
rect 677244 547572 677250 547574
rect 677501 547571 677567 547574
rect 31753 547498 31819 547501
rect 28766 547496 31819 547498
rect 28766 547468 31758 547496
rect 28796 547440 31758 547468
rect 31814 547440 31819 547496
rect 28796 547438 31819 547440
rect 31753 547435 31819 547438
rect 674189 547362 674255 547365
rect 676121 547362 676187 547365
rect 674189 547360 676187 547362
rect 674189 547304 674194 547360
rect 674250 547304 676126 547360
rect 676182 547304 676187 547360
rect 674189 547302 676187 547304
rect 674189 547299 674255 547302
rect 676121 547299 676187 547302
rect 43437 547090 43503 547093
rect 41492 547088 43503 547090
rect 41492 547032 43442 547088
rect 43498 547032 43503 547088
rect 41492 547030 43503 547032
rect 43437 547027 43503 547030
rect 674230 547028 674236 547092
rect 674300 547090 674306 547092
rect 683389 547090 683455 547093
rect 674300 547088 683455 547090
rect 674300 547032 683394 547088
rect 683450 547032 683455 547088
rect 674300 547030 683455 547032
rect 674300 547028 674306 547030
rect 683389 547027 683455 547030
rect 676070 546756 676076 546820
rect 676140 546818 676146 546820
rect 679617 546818 679683 546821
rect 676140 546816 679683 546818
rect 676140 546760 679622 546816
rect 679678 546760 679683 546816
rect 676140 546758 679683 546760
rect 676140 546756 676146 546758
rect 679617 546755 679683 546758
rect 41638 546348 41644 546412
rect 41708 546410 41714 546412
rect 42374 546410 42380 546412
rect 41708 546350 42380 546410
rect 41708 546348 41714 546350
rect 42374 546348 42380 546350
rect 42444 546348 42450 546412
rect 40861 545866 40927 545869
rect 41822 545866 41828 545868
rect 40861 545864 41828 545866
rect 40861 545808 40866 545864
rect 40922 545808 41828 545864
rect 40861 545806 41828 545808
rect 40861 545803 40927 545806
rect 41822 545804 41828 545806
rect 41892 545804 41898 545868
rect 62113 545866 62179 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 62113 545803 62179 545806
rect 40718 545532 40724 545596
rect 40788 545594 40794 545596
rect 42149 545594 42215 545597
rect 40788 545592 42215 545594
rect 40788 545536 42154 545592
rect 42210 545536 42215 545592
rect 40788 545534 42215 545536
rect 40788 545532 40794 545534
rect 42149 545531 42215 545534
rect 40534 545260 40540 545324
rect 40604 545322 40610 545324
rect 41965 545322 42031 545325
rect 40604 545320 42031 545322
rect 40604 545264 41970 545320
rect 42026 545264 42031 545320
rect 40604 545262 42031 545264
rect 40604 545260 40610 545262
rect 41965 545259 42031 545262
rect 39757 542194 39823 542197
rect 42333 542194 42399 542197
rect 39757 542192 42399 542194
rect 39757 542136 39762 542192
rect 39818 542136 42338 542192
rect 42394 542136 42399 542192
rect 39757 542134 42399 542136
rect 39757 542131 39823 542134
rect 42333 542131 42399 542134
rect 39481 541922 39547 541925
rect 42057 541922 42123 541925
rect 39481 541920 42123 541922
rect 39481 541864 39486 541920
rect 39542 541864 42062 541920
rect 42118 541864 42123 541920
rect 39481 541862 42123 541864
rect 39481 541859 39547 541862
rect 42057 541859 42123 541862
rect 40902 538188 40908 538252
rect 40972 538250 40978 538252
rect 42333 538250 42399 538253
rect 40972 538248 42399 538250
rect 40972 538192 42338 538248
rect 42394 538192 42399 538248
rect 40972 538190 42399 538192
rect 40972 538188 40978 538190
rect 42333 538187 42399 538190
rect 42149 537978 42215 537981
rect 42701 537978 42767 537981
rect 42149 537976 42767 537978
rect 42149 537920 42154 537976
rect 42210 537920 42706 537976
rect 42762 537920 42767 537976
rect 42149 537918 42767 537920
rect 42149 537915 42215 537918
rect 42701 537915 42767 537918
rect 651557 537570 651623 537573
rect 650164 537568 651623 537570
rect 650164 537512 651562 537568
rect 651618 537512 651623 537568
rect 650164 537510 651623 537512
rect 651557 537507 651623 537510
rect 675477 536074 675543 536077
rect 676262 536074 676322 536112
rect 675477 536072 676322 536074
rect 675477 536016 675482 536072
rect 675538 536016 676322 536072
rect 675477 536014 676322 536016
rect 675477 536011 675543 536014
rect 675477 535530 675543 535533
rect 676262 535530 676322 535704
rect 675477 535528 676322 535530
rect 675477 535472 675482 535528
rect 675538 535472 676322 535528
rect 675477 535470 676322 535472
rect 675477 535467 675543 535470
rect 40718 535196 40724 535260
rect 40788 535258 40794 535260
rect 41781 535258 41847 535261
rect 40788 535256 41847 535258
rect 40788 535200 41786 535256
rect 41842 535200 41847 535256
rect 40788 535198 41847 535200
rect 40788 535196 40794 535198
rect 41781 535195 41847 535198
rect 674465 535122 674531 535125
rect 676262 535122 676322 535296
rect 674465 535120 676322 535122
rect 674465 535064 674470 535120
rect 674526 535064 676322 535120
rect 674465 535062 676322 535064
rect 674465 535059 674531 535062
rect 675477 534850 675543 534853
rect 676262 534850 676322 534888
rect 675477 534848 676322 534850
rect 675477 534792 675482 534848
rect 675538 534792 676322 534848
rect 675477 534790 676322 534792
rect 675477 534787 675543 534790
rect 675477 534306 675543 534309
rect 676262 534306 676322 534480
rect 675477 534304 676322 534306
rect 675477 534248 675482 534304
rect 675538 534248 676322 534304
rect 675477 534246 676322 534248
rect 675477 534243 675543 534246
rect 674925 534034 674991 534037
rect 676262 534034 676322 534090
rect 674925 534032 676322 534034
rect 674925 533976 674930 534032
rect 674986 533976 676322 534032
rect 674925 533974 676322 533976
rect 674925 533971 674991 533974
rect 674281 533626 674347 533629
rect 676262 533626 676322 533664
rect 674281 533624 676322 533626
rect 674281 533568 674286 533624
rect 674342 533568 676322 533624
rect 674281 533566 676322 533568
rect 674281 533563 674347 533566
rect 40534 533292 40540 533356
rect 40604 533354 40610 533356
rect 42241 533354 42307 533357
rect 40604 533352 42307 533354
rect 40604 533296 42246 533352
rect 42302 533296 42307 533352
rect 40604 533294 42307 533296
rect 40604 533292 40610 533294
rect 42241 533291 42307 533294
rect 675477 533354 675543 533357
rect 675477 533352 676322 533354
rect 675477 533296 675482 533352
rect 675538 533296 676322 533352
rect 675477 533294 676322 533296
rect 675477 533291 675543 533294
rect 676262 533256 676322 533294
rect 62757 532810 62823 532813
rect 675477 532810 675543 532813
rect 676262 532810 676322 532848
rect 62757 532808 64492 532810
rect 62757 532752 62762 532808
rect 62818 532752 64492 532808
rect 62757 532750 64492 532752
rect 675477 532808 676322 532810
rect 675477 532752 675482 532808
rect 675538 532752 676322 532808
rect 675477 532750 676322 532752
rect 62757 532747 62823 532750
rect 675477 532747 675543 532750
rect 675477 532538 675543 532541
rect 675477 532536 676322 532538
rect 675477 532480 675482 532536
rect 675538 532480 676322 532536
rect 675477 532478 676322 532480
rect 675477 532475 675543 532478
rect 676262 532440 676322 532478
rect 674465 531994 674531 531997
rect 676262 531994 676322 532032
rect 674465 531992 676322 531994
rect 674465 531936 674470 531992
rect 674526 531936 676322 531992
rect 674465 531934 676322 531936
rect 674465 531931 674531 531934
rect 675477 531586 675543 531589
rect 676262 531586 676322 531624
rect 675477 531584 676322 531586
rect 675477 531528 675482 531584
rect 675538 531528 676322 531584
rect 675477 531526 676322 531528
rect 675477 531523 675543 531526
rect 674925 531178 674991 531181
rect 676262 531178 676322 531216
rect 674925 531176 676322 531178
rect 674925 531120 674930 531176
rect 674986 531120 676322 531176
rect 674925 531118 676322 531120
rect 674925 531115 674991 531118
rect 683389 531042 683455 531045
rect 683389 531040 683498 531042
rect 683389 530984 683394 531040
rect 683450 530984 683498 531040
rect 683389 530979 683498 530984
rect 683438 530808 683498 530979
rect 679617 530634 679683 530637
rect 679574 530632 679683 530634
rect 679574 530576 679622 530632
rect 679678 530576 679683 530632
rect 679574 530571 679683 530576
rect 679574 530400 679634 530571
rect 41454 530164 41460 530228
rect 41524 530226 41530 530228
rect 42609 530226 42675 530229
rect 41524 530224 42675 530226
rect 41524 530168 42614 530224
rect 42670 530168 42675 530224
rect 41524 530166 42675 530168
rect 41524 530164 41530 530166
rect 42609 530163 42675 530166
rect 675477 530090 675543 530093
rect 675477 530088 676322 530090
rect 675477 530032 675482 530088
rect 675538 530032 676322 530088
rect 675477 530030 676322 530032
rect 675477 530027 675543 530030
rect 676262 529992 676322 530030
rect 41822 529756 41828 529820
rect 41892 529818 41898 529820
rect 42701 529818 42767 529821
rect 41892 529816 42767 529818
rect 41892 529760 42706 529816
rect 42762 529760 42767 529816
rect 41892 529758 42767 529760
rect 41892 529756 41898 529758
rect 42701 529755 42767 529758
rect 675477 529546 675543 529549
rect 676262 529546 676322 529584
rect 675477 529544 676322 529546
rect 675477 529488 675482 529544
rect 675538 529488 676322 529544
rect 675477 529486 676322 529488
rect 675477 529483 675543 529486
rect 41781 529412 41847 529413
rect 41781 529408 41828 529412
rect 41892 529410 41898 529412
rect 677501 529410 677567 529413
rect 41781 529352 41786 529408
rect 41781 529348 41828 529352
rect 41892 529350 41938 529410
rect 677501 529408 677610 529410
rect 677501 529352 677506 529408
rect 677562 529352 677610 529408
rect 41892 529348 41898 529350
rect 41781 529347 41847 529348
rect 677501 529347 677610 529352
rect 677550 529176 677610 529347
rect 683205 529002 683271 529005
rect 683205 529000 683314 529002
rect 683205 528944 683210 529000
rect 683266 528944 683314 529000
rect 683205 528939 683314 528944
rect 683254 528768 683314 528939
rect 675477 528458 675543 528461
rect 675477 528456 676322 528458
rect 675477 528400 675482 528456
rect 675538 528400 676322 528456
rect 675477 528398 676322 528400
rect 675477 528395 675543 528398
rect 676262 528360 676322 528398
rect 675477 528050 675543 528053
rect 675477 528048 676322 528050
rect 675477 527992 675482 528048
rect 675538 527992 676322 528048
rect 675477 527990 676322 527992
rect 675477 527987 675543 527990
rect 676262 527952 676322 527990
rect 674005 527642 674071 527645
rect 674005 527640 676322 527642
rect 674005 527584 674010 527640
rect 674066 527584 676322 527640
rect 674005 527582 676322 527584
rect 674005 527579 674071 527582
rect 676262 527544 676322 527582
rect 674598 527036 674604 527100
rect 674668 527098 674674 527100
rect 676262 527098 676322 527136
rect 674668 527038 676322 527098
rect 674668 527036 674674 527038
rect 675477 526826 675543 526829
rect 675477 526824 676322 526826
rect 675477 526768 675482 526824
rect 675538 526768 676322 526824
rect 675477 526766 676322 526768
rect 675477 526763 675543 526766
rect 676262 526728 676322 526766
rect 675477 526418 675543 526421
rect 675477 526416 676322 526418
rect 675477 526360 675482 526416
rect 675538 526360 676322 526416
rect 675477 526358 676322 526360
rect 675477 526355 675543 526358
rect 676262 526320 676322 526358
rect 675477 525874 675543 525877
rect 676262 525874 676322 525912
rect 675477 525872 676322 525874
rect 675477 525816 675482 525872
rect 675538 525816 676322 525872
rect 675477 525814 676322 525816
rect 675477 525811 675543 525814
rect 683113 525738 683179 525741
rect 683070 525736 683179 525738
rect 683070 525680 683118 525736
rect 683174 525680 683179 525736
rect 683070 525675 683179 525680
rect 683070 525096 683130 525675
rect 673862 524452 673868 524516
rect 673932 524514 673938 524516
rect 676262 524514 676322 524688
rect 673932 524454 676322 524514
rect 673932 524452 673938 524454
rect 651557 524242 651623 524245
rect 650164 524240 651623 524242
rect 650164 524184 651562 524240
rect 651618 524184 651623 524240
rect 650164 524182 651623 524184
rect 651557 524179 651623 524182
rect 40677 522746 40743 522749
rect 43253 522746 43319 522749
rect 40677 522744 43319 522746
rect 40677 522688 40682 522744
rect 40738 522688 43258 522744
rect 43314 522688 43319 522744
rect 40677 522686 43319 522688
rect 40677 522683 40743 522686
rect 43253 522683 43319 522686
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 651557 511050 651623 511053
rect 650164 511048 651623 511050
rect 650164 510992 651562 511048
rect 651618 510992 651623 511048
rect 650164 510990 651623 510992
rect 651557 510987 651623 510990
rect 675109 508874 675175 508877
rect 676029 508874 676095 508877
rect 675109 508872 676095 508874
rect 675109 508816 675114 508872
rect 675170 508816 676034 508872
rect 676090 508816 676095 508872
rect 675109 508814 676095 508816
rect 675109 508811 675175 508814
rect 676029 508811 676095 508814
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 675293 500306 675359 500309
rect 676029 500306 676095 500309
rect 675293 500304 676095 500306
rect 675293 500248 675298 500304
rect 675354 500248 676034 500304
rect 676090 500248 676095 500304
rect 675293 500246 676095 500248
rect 675293 500243 675359 500246
rect 676029 500243 676095 500246
rect 651557 497722 651623 497725
rect 650164 497720 651623 497722
rect 650164 497664 651562 497720
rect 651618 497664 651623 497720
rect 650164 497662 651623 497664
rect 651557 497659 651623 497662
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 675293 492146 675359 492149
rect 675293 492144 676292 492146
rect 675293 492088 675298 492144
rect 675354 492088 676292 492144
rect 675293 492086 676292 492088
rect 675293 492083 675359 492086
rect 675477 491738 675543 491741
rect 675477 491736 676292 491738
rect 675477 491680 675482 491736
rect 675538 491680 676292 491736
rect 675477 491678 676292 491680
rect 675477 491675 675543 491678
rect 675477 491330 675543 491333
rect 675477 491328 676292 491330
rect 675477 491272 675482 491328
rect 675538 491272 676292 491328
rect 675477 491270 676292 491272
rect 675477 491267 675543 491270
rect 675477 490922 675543 490925
rect 675477 490920 676292 490922
rect 675477 490864 675482 490920
rect 675538 490864 676292 490920
rect 675477 490862 676292 490864
rect 675477 490859 675543 490862
rect 676029 490514 676095 490517
rect 676029 490512 676292 490514
rect 676029 490456 676034 490512
rect 676090 490456 676292 490512
rect 676029 490454 676292 490456
rect 676029 490451 676095 490454
rect 674281 490106 674347 490109
rect 674281 490104 676292 490106
rect 674281 490048 674286 490104
rect 674342 490048 676292 490104
rect 674281 490046 676292 490048
rect 674281 490043 674347 490046
rect 676029 489698 676095 489701
rect 676029 489696 676292 489698
rect 676029 489640 676034 489696
rect 676090 489640 676292 489696
rect 676029 489638 676292 489640
rect 676029 489635 676095 489638
rect 675477 489290 675543 489293
rect 675477 489288 676292 489290
rect 675477 489232 675482 489288
rect 675538 489232 676292 489288
rect 675477 489230 676292 489232
rect 675477 489227 675543 489230
rect 675661 488882 675727 488885
rect 675661 488880 676292 488882
rect 675661 488824 675666 488880
rect 675722 488824 676292 488880
rect 675661 488822 676292 488824
rect 675661 488819 675727 488822
rect 674465 488474 674531 488477
rect 674465 488472 676292 488474
rect 674465 488416 674470 488472
rect 674526 488416 676292 488472
rect 674465 488414 676292 488416
rect 674465 488411 674531 488414
rect 676029 488066 676095 488069
rect 676029 488064 676292 488066
rect 676029 488008 676034 488064
rect 676090 488008 676292 488064
rect 676029 488006 676292 488008
rect 676029 488003 676095 488006
rect 675845 487658 675911 487661
rect 675845 487656 676292 487658
rect 675845 487600 675850 487656
rect 675906 487600 676292 487656
rect 675845 487598 676292 487600
rect 675845 487595 675911 487598
rect 679617 487250 679683 487253
rect 679604 487248 679683 487250
rect 679604 487192 679622 487248
rect 679678 487192 679683 487248
rect 679604 487190 679683 487192
rect 679617 487187 679683 487190
rect 675293 486842 675359 486845
rect 675293 486840 676292 486842
rect 675293 486784 675298 486840
rect 675354 486784 676292 486840
rect 675293 486782 676292 486784
rect 675293 486779 675359 486782
rect 679801 486434 679867 486437
rect 679788 486432 679867 486434
rect 679788 486376 679806 486432
rect 679862 486376 679867 486432
rect 679788 486374 679867 486376
rect 679801 486371 679867 486374
rect 675477 486026 675543 486029
rect 675477 486024 676292 486026
rect 675477 485968 675482 486024
rect 675538 485968 676292 486024
rect 675477 485966 676292 485968
rect 675477 485963 675543 485966
rect 675477 485618 675543 485621
rect 675477 485616 676292 485618
rect 675477 485560 675482 485616
rect 675538 485560 676292 485616
rect 675477 485558 676292 485560
rect 675477 485555 675543 485558
rect 675477 485210 675543 485213
rect 675477 485208 676292 485210
rect 675477 485152 675482 485208
rect 675538 485152 676292 485208
rect 675477 485150 676292 485152
rect 675477 485147 675543 485150
rect 675886 484740 675892 484804
rect 675956 484802 675962 484804
rect 675956 484742 676292 484802
rect 675956 484740 675962 484742
rect 651557 484530 651623 484533
rect 650164 484528 651623 484530
rect 650164 484472 651562 484528
rect 651618 484472 651623 484528
rect 650164 484470 651623 484472
rect 651557 484467 651623 484470
rect 674649 484394 674715 484397
rect 674649 484392 676292 484394
rect 674649 484336 674654 484392
rect 674710 484336 676292 484392
rect 674649 484334 676292 484336
rect 674649 484331 674715 484334
rect 675886 483924 675892 483988
rect 675956 483986 675962 483988
rect 675956 483926 676292 483986
rect 675956 483924 675962 483926
rect 675477 483578 675543 483581
rect 675477 483576 676292 483578
rect 675477 483520 675482 483576
rect 675538 483520 676292 483576
rect 675477 483518 676292 483520
rect 675477 483515 675543 483518
rect 675477 483170 675543 483173
rect 675477 483168 676292 483170
rect 675477 483112 675482 483168
rect 675538 483112 676292 483168
rect 675477 483110 676292 483112
rect 675477 483107 675543 483110
rect 675477 482762 675543 482765
rect 675477 482760 676292 482762
rect 675477 482704 675482 482760
rect 675538 482704 676292 482760
rect 675477 482702 676292 482704
rect 675477 482699 675543 482702
rect 675477 482354 675543 482357
rect 675477 482352 676292 482354
rect 675477 482296 675482 482352
rect 675538 482296 676292 482352
rect 675477 482294 676292 482296
rect 675477 482291 675543 482294
rect 675477 481946 675543 481949
rect 675477 481944 676292 481946
rect 675477 481888 675482 481944
rect 675538 481888 676292 481944
rect 675477 481886 676292 481888
rect 675477 481883 675543 481886
rect 674925 481538 674991 481541
rect 674925 481536 676292 481538
rect 674925 481480 674930 481536
rect 674986 481508 676292 481536
rect 674986 481480 676322 481508
rect 674925 481478 676322 481480
rect 674925 481475 674991 481478
rect 676262 481100 676322 481478
rect 675477 480722 675543 480725
rect 675477 480720 676292 480722
rect 675477 480664 675482 480720
rect 675538 480664 676292 480720
rect 675477 480662 676292 480664
rect 675477 480659 675543 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 672625 474874 672691 474877
rect 673310 474874 673316 474876
rect 672625 474872 673316 474874
rect 672625 474816 672630 474872
rect 672686 474816 673316 474872
rect 672625 474814 673316 474816
rect 672625 474811 672691 474814
rect 673310 474812 673316 474814
rect 673380 474812 673386 474876
rect 651557 471202 651623 471205
rect 650164 471200 651623 471202
rect 650164 471144 651562 471200
rect 651618 471144 651623 471200
rect 650164 471142 651623 471144
rect 651557 471139 651623 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 651557 457874 651623 457877
rect 650164 457872 651623 457874
rect 650164 457816 651562 457872
rect 651618 457816 651623 457872
rect 650164 457814 651623 457816
rect 651557 457811 651623 457814
rect 62113 454610 62179 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 62113 454547 62179 454550
rect 651557 444546 651623 444549
rect 650164 444544 651623 444546
rect 650164 444488 651562 444544
rect 651618 444488 651623 444544
rect 650164 444486 651623 444488
rect 651557 444483 651623 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 651557 431354 651623 431357
rect 650164 431352 651623 431354
rect 650164 431296 651562 431352
rect 651618 431296 651623 431352
rect 650164 431294 651623 431296
rect 651557 431291 651623 431294
rect 40677 431218 40743 431221
rect 40677 431216 40786 431218
rect 40677 431160 40682 431216
rect 40738 431160 40786 431216
rect 40677 431155 40786 431160
rect 40726 430916 40786 431155
rect 41321 430538 41387 430541
rect 41308 430536 41387 430538
rect 41308 430480 41326 430536
rect 41382 430480 41387 430536
rect 41308 430478 41387 430480
rect 41321 430475 41387 430478
rect 41137 430130 41203 430133
rect 41124 430128 41203 430130
rect 41124 430072 41142 430128
rect 41198 430072 41203 430128
rect 41124 430070 41203 430072
rect 41137 430067 41203 430070
rect 40910 429487 40970 429692
rect 40910 429482 41019 429487
rect 41321 429484 41387 429487
rect 40910 429426 40958 429482
rect 41014 429426 41019 429482
rect 40910 429424 41019 429426
rect 40953 429421 41019 429424
rect 41278 429482 41387 429484
rect 41278 429426 41326 429482
rect 41382 429426 41387 429482
rect 41278 429421 41387 429426
rect 41278 429284 41338 429421
rect 41137 428906 41203 428909
rect 41124 428904 41203 428906
rect 41124 428848 41142 428904
rect 41198 428848 41203 428904
rect 41124 428846 41203 428848
rect 41137 428843 41203 428846
rect 42701 428498 42767 428501
rect 41492 428496 42767 428498
rect 41492 428440 42706 428496
rect 42762 428440 42767 428496
rect 41492 428438 42767 428440
rect 42701 428435 42767 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 41278 427855 41338 428060
rect 41278 427850 41387 427855
rect 41278 427794 41326 427850
rect 41382 427794 41387 427850
rect 41278 427792 41387 427794
rect 41321 427789 41387 427792
rect 40953 427682 41019 427685
rect 40940 427680 41019 427682
rect 40940 427624 40958 427680
rect 41014 427624 41019 427680
rect 40940 427622 41019 427624
rect 40953 427619 41019 427622
rect 41137 427274 41203 427277
rect 41124 427272 41203 427274
rect 41124 427216 41142 427272
rect 41198 427216 41203 427272
rect 41124 427214 41203 427216
rect 41137 427211 41203 427214
rect 44541 426866 44607 426869
rect 41492 426864 44607 426866
rect 41492 426808 44546 426864
rect 44602 426808 44607 426864
rect 41492 426806 44607 426808
rect 44541 426803 44607 426806
rect 41822 426458 41828 426460
rect 41492 426398 41828 426458
rect 41822 426396 41828 426398
rect 41892 426396 41898 426460
rect 41321 426050 41387 426053
rect 41308 426048 41387 426050
rect 41308 425992 41326 426048
rect 41382 425992 41387 426048
rect 41308 425990 41387 425992
rect 41321 425987 41387 425990
rect 41822 425642 41828 425644
rect 41492 425582 41828 425642
rect 41822 425580 41828 425582
rect 41892 425580 41898 425644
rect 40769 425234 40835 425237
rect 40756 425232 40835 425234
rect 40756 425176 40774 425232
rect 40830 425176 40835 425232
rect 40756 425174 40835 425176
rect 40769 425171 40835 425174
rect 45553 424826 45619 424829
rect 41492 424824 45619 424826
rect 41492 424768 45558 424824
rect 45614 424768 45619 424824
rect 41492 424766 45619 424768
rect 45553 424763 45619 424766
rect 42609 424418 42675 424421
rect 41492 424416 42675 424418
rect 41492 424360 42614 424416
rect 42670 424360 42675 424416
rect 41492 424358 42675 424360
rect 42609 424355 42675 424358
rect 43989 424010 44055 424013
rect 41492 424008 44055 424010
rect 41492 423952 43994 424008
rect 44050 423952 44055 424008
rect 41492 423950 44055 423952
rect 43989 423947 44055 423950
rect 45185 423602 45251 423605
rect 41492 423600 45251 423602
rect 41492 423544 45190 423600
rect 45246 423544 45251 423600
rect 41492 423542 45251 423544
rect 45185 423539 45251 423542
rect 43805 423194 43871 423197
rect 41492 423192 43871 423194
rect 41492 423136 43810 423192
rect 43866 423136 43871 423192
rect 41492 423134 43871 423136
rect 43805 423131 43871 423134
rect 43437 422786 43503 422789
rect 41492 422784 43503 422786
rect 41492 422728 43442 422784
rect 43498 422728 43503 422784
rect 41492 422726 43503 422728
rect 43437 422723 43503 422726
rect 40726 422312 40786 422348
rect 40718 422248 40724 422312
rect 40788 422248 40794 422312
rect 42006 421970 42012 421972
rect 41492 421910 42012 421970
rect 42006 421908 42012 421910
rect 42076 421908 42082 421972
rect 43069 421562 43135 421565
rect 41492 421560 43135 421562
rect 41492 421504 43074 421560
rect 43130 421504 43135 421560
rect 41492 421502 43135 421504
rect 43069 421499 43135 421502
rect 41462 421290 42074 421324
rect 45369 421290 45435 421293
rect 41462 421288 45435 421290
rect 41462 421264 45374 421288
rect 41462 421124 41522 421264
rect 42014 421232 45374 421264
rect 45430 421232 45435 421288
rect 42014 421230 45435 421232
rect 45369 421227 45435 421230
rect 41781 421156 41847 421157
rect 41781 421152 41828 421156
rect 41892 421154 41898 421156
rect 41781 421096 41786 421152
rect 41781 421092 41828 421096
rect 41892 421094 41938 421154
rect 41892 421092 41898 421094
rect 41781 421091 41847 421092
rect 42425 420746 42491 420749
rect 41492 420744 42491 420746
rect 41492 420688 42430 420744
rect 42486 420688 42491 420744
rect 41492 420686 42491 420688
rect 42425 420683 42491 420686
rect 41462 419930 41522 420308
rect 41873 419930 41939 419933
rect 41462 419928 41939 419930
rect 41462 419900 41878 419928
rect 41492 419872 41878 419900
rect 41934 419872 41939 419928
rect 41492 419870 41939 419872
rect 41873 419867 41939 419870
rect 45737 419522 45803 419525
rect 41492 419520 45803 419522
rect 41492 419464 45742 419520
rect 45798 419464 45803 419520
rect 41492 419462 45803 419464
rect 45737 419459 45803 419462
rect 40534 418644 40540 418708
rect 40604 418706 40610 418708
rect 42006 418706 42012 418708
rect 40604 418646 42012 418706
rect 40604 418644 40610 418646
rect 42006 418644 42012 418646
rect 42076 418644 42082 418708
rect 651557 418026 651623 418029
rect 650164 418024 651623 418026
rect 650164 417968 651562 418024
rect 651618 417968 651623 418024
rect 650164 417966 651623 417968
rect 651557 417963 651623 417966
rect 62113 415442 62179 415445
rect 62113 415440 64492 415442
rect 62113 415384 62118 415440
rect 62174 415384 64492 415440
rect 62113 415382 64492 415384
rect 62113 415379 62179 415382
rect 42057 412994 42123 412997
rect 42609 412994 42675 412997
rect 42057 412992 42675 412994
rect 42057 412936 42062 412992
rect 42118 412936 42614 412992
rect 42670 412936 42675 412992
rect 42057 412934 42675 412936
rect 42057 412931 42123 412934
rect 42609 412931 42675 412934
rect 40718 407492 40724 407556
rect 40788 407554 40794 407556
rect 41781 407554 41847 407557
rect 40788 407552 41847 407554
rect 40788 407496 41786 407552
rect 41842 407496 41847 407552
rect 40788 407494 41847 407496
rect 40788 407492 40794 407494
rect 41781 407491 41847 407494
rect 651557 404698 651623 404701
rect 650164 404696 651623 404698
rect 650164 404640 651562 404696
rect 651618 404640 651623 404696
rect 650164 404638 651623 404640
rect 651557 404635 651623 404638
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 675477 403882 675543 403885
rect 675477 403880 676292 403882
rect 675477 403824 675482 403880
rect 675538 403824 676292 403880
rect 675477 403822 676292 403824
rect 675477 403819 675543 403822
rect 675293 403474 675359 403477
rect 675293 403472 676292 403474
rect 675293 403416 675298 403472
rect 675354 403416 676292 403472
rect 675293 403414 676292 403416
rect 675293 403411 675359 403414
rect 675477 403066 675543 403069
rect 675477 403064 676292 403066
rect 675477 403008 675482 403064
rect 675538 403008 676292 403064
rect 675477 403006 676292 403008
rect 675477 403003 675543 403006
rect 677409 402930 677475 402933
rect 677366 402928 677475 402930
rect 677366 402872 677414 402928
rect 677470 402872 677475 402928
rect 677366 402867 677475 402872
rect 677366 402628 677426 402867
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 674649 402250 674715 402253
rect 674649 402248 676292 402250
rect 674649 402192 674654 402248
rect 674710 402192 676292 402248
rect 674649 402190 676292 402192
rect 674649 402187 674715 402190
rect 677225 402114 677291 402117
rect 677182 402112 677291 402114
rect 677182 402056 677230 402112
rect 677286 402056 677291 402112
rect 677182 402051 677291 402056
rect 41781 401980 41847 401981
rect 41781 401976 41828 401980
rect 41892 401978 41898 401980
rect 41781 401920 41786 401976
rect 41781 401916 41828 401920
rect 41892 401918 41938 401978
rect 41892 401916 41898 401918
rect 41781 401915 41847 401916
rect 677182 401812 677242 402051
rect 674465 401434 674531 401437
rect 674465 401432 676292 401434
rect 674465 401376 674470 401432
rect 674526 401376 676292 401432
rect 674465 401374 676292 401376
rect 674465 401371 674531 401374
rect 675937 401026 676003 401029
rect 675937 401024 676292 401026
rect 675937 400968 675942 401024
rect 675998 400968 676292 401024
rect 675937 400966 676292 400968
rect 675937 400963 676003 400966
rect 675477 400618 675543 400621
rect 675477 400616 676292 400618
rect 675477 400560 675482 400616
rect 675538 400560 676292 400616
rect 675477 400558 676292 400560
rect 675477 400555 675543 400558
rect 675937 400210 676003 400213
rect 675937 400208 676292 400210
rect 675937 400152 675942 400208
rect 675998 400152 676292 400208
rect 675937 400150 676292 400152
rect 675937 400147 676003 400150
rect 41454 400012 41460 400076
rect 41524 400074 41530 400076
rect 41781 400074 41847 400077
rect 41524 400072 41847 400074
rect 41524 400016 41786 400072
rect 41842 400016 41847 400072
rect 41524 400014 41847 400016
rect 41524 400012 41530 400014
rect 41781 400011 41847 400014
rect 675477 399802 675543 399805
rect 675477 399800 676292 399802
rect 675477 399744 675482 399800
rect 675538 399744 676292 399800
rect 675477 399742 676292 399744
rect 675477 399739 675543 399742
rect 674925 399394 674991 399397
rect 674925 399392 676292 399394
rect 674925 399336 674930 399392
rect 674986 399336 676292 399392
rect 674925 399334 676292 399336
rect 674925 399331 674991 399334
rect 41873 398852 41939 398853
rect 41822 398850 41828 398852
rect 41782 398790 41828 398850
rect 41892 398848 41939 398852
rect 41934 398792 41939 398848
rect 41822 398788 41828 398790
rect 41892 398788 41939 398792
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 41873 398787 41939 398788
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 675109 398170 675175 398173
rect 675109 398168 676292 398170
rect 675109 398112 675114 398168
rect 675170 398112 676292 398168
rect 675109 398110 676292 398112
rect 675109 398107 675175 398110
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 675477 397354 675543 397357
rect 675477 397352 676292 397354
rect 675477 397296 675482 397352
rect 675538 397296 676292 397352
rect 675477 397294 676292 397296
rect 675477 397291 675543 397294
rect 676262 396812 676322 396916
rect 676254 396748 676260 396812
rect 676324 396748 676330 396812
rect 681230 396405 681290 396508
rect 681181 396400 681290 396405
rect 681181 396344 681186 396400
rect 681242 396344 681290 396400
rect 681181 396342 681290 396344
rect 681181 396339 681247 396342
rect 675477 396130 675543 396133
rect 675477 396128 676292 396130
rect 675477 396072 675482 396128
rect 675538 396072 676292 396128
rect 675477 396070 676292 396072
rect 675477 396067 675543 396070
rect 675477 395722 675543 395725
rect 675477 395720 676292 395722
rect 675477 395664 675482 395720
rect 675538 395664 676292 395720
rect 675477 395662 676292 395664
rect 675477 395659 675543 395662
rect 676630 395180 676690 395284
rect 676622 395116 676628 395180
rect 676692 395116 676698 395180
rect 676446 394772 676506 394876
rect 676438 394708 676444 394772
rect 676508 394708 676514 394772
rect 675477 394498 675543 394501
rect 675477 394496 676292 394498
rect 675477 394440 675482 394496
rect 675538 394440 676292 394496
rect 675477 394438 676292 394440
rect 675477 394435 675543 394438
rect 675477 394090 675543 394093
rect 675477 394088 676292 394090
rect 675477 394032 675482 394088
rect 675538 394032 676292 394088
rect 675477 394030 676292 394032
rect 675477 394027 675543 394030
rect 674281 393682 674347 393685
rect 674281 393680 676292 393682
rect 674281 393624 674286 393680
rect 674342 393624 676292 393680
rect 674281 393622 676292 393624
rect 674281 393619 674347 393622
rect 672349 393274 672415 393277
rect 672942 393274 672948 393276
rect 672349 393272 672948 393274
rect 672349 393216 672354 393272
rect 672410 393216 672948 393272
rect 672349 393214 672948 393216
rect 672349 393211 672415 393214
rect 672942 393212 672948 393214
rect 673012 393212 673018 393276
rect 683070 392733 683130 393244
rect 683070 392728 683179 392733
rect 683070 392672 683118 392728
rect 683174 392672 683179 392728
rect 683070 392670 683179 392672
rect 683113 392667 683179 392670
rect 675477 392458 675543 392461
rect 675477 392456 676292 392458
rect 675477 392400 675482 392456
rect 675538 392400 676292 392456
rect 675477 392398 676292 392400
rect 675477 392395 675543 392398
rect 651557 391506 651623 391509
rect 650164 391504 651623 391506
rect 650164 391448 651562 391504
rect 651618 391448 651623 391504
rect 650164 391446 651623 391448
rect 651557 391443 651623 391446
rect 62113 389330 62179 389333
rect 672809 389330 672875 389333
rect 675845 389330 675911 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 672809 389328 675911 389330
rect 672809 389272 672814 389328
rect 672870 389272 675850 389328
rect 675906 389272 675911 389328
rect 672809 389270 675911 389272
rect 62113 389267 62179 389270
rect 672809 389267 672875 389270
rect 675845 389267 675911 389270
rect 675886 388452 675892 388516
rect 675956 388514 675962 388516
rect 680997 388514 681063 388517
rect 675956 388512 681063 388514
rect 675956 388456 681002 388512
rect 681058 388456 681063 388512
rect 675956 388454 681063 388456
rect 675956 388452 675962 388454
rect 680997 388451 681063 388454
rect 35390 387565 35450 387668
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 681181 387698 681247 387701
rect 675772 387696 681247 387698
rect 675772 387640 681186 387696
rect 681242 387640 681247 387696
rect 675772 387638 681247 387640
rect 675772 387636 675778 387638
rect 681181 387635 681247 387638
rect 35390 387560 35499 387565
rect 35801 387562 35867 387565
rect 35390 387504 35438 387560
rect 35494 387504 35499 387560
rect 35390 387502 35499 387504
rect 35433 387499 35499 387502
rect 35758 387560 35867 387562
rect 35758 387504 35806 387560
rect 35862 387504 35867 387560
rect 35758 387499 35867 387504
rect 35758 387260 35818 387499
rect 39941 387154 40007 387157
rect 43253 387154 43319 387157
rect 39941 387152 43319 387154
rect 39941 387096 39946 387152
rect 40002 387096 43258 387152
rect 43314 387096 43319 387152
rect 39941 387094 43319 387096
rect 39941 387091 40007 387094
rect 43253 387091 43319 387094
rect 35758 386749 35818 386852
rect 35758 386744 35867 386749
rect 35758 386688 35806 386744
rect 35862 386688 35867 386744
rect 35758 386686 35867 386688
rect 35801 386683 35867 386686
rect 40125 386746 40191 386749
rect 43621 386746 43687 386749
rect 40125 386744 43687 386746
rect 40125 386688 40130 386744
rect 40186 386688 43626 386744
rect 43682 386688 43687 386744
rect 40125 386686 43687 386688
rect 40125 386683 40191 386686
rect 43621 386683 43687 386686
rect 35574 386341 35634 386444
rect 35574 386336 35683 386341
rect 35574 386280 35622 386336
rect 35678 386280 35683 386336
rect 35574 386278 35683 386280
rect 35617 386275 35683 386278
rect 35390 385933 35450 386036
rect 35341 385928 35450 385933
rect 35341 385872 35346 385928
rect 35402 385872 35450 385928
rect 35341 385870 35450 385872
rect 35341 385867 35407 385870
rect 35574 385525 35634 385628
rect 35525 385520 35634 385525
rect 35801 385522 35867 385525
rect 35525 385464 35530 385520
rect 35586 385464 35634 385520
rect 35525 385462 35634 385464
rect 35758 385520 35867 385522
rect 35758 385464 35806 385520
rect 35862 385464 35867 385520
rect 35525 385459 35591 385462
rect 35758 385459 35867 385464
rect 35758 385220 35818 385459
rect 39941 385114 40007 385117
rect 44357 385114 44423 385117
rect 39941 385112 44423 385114
rect 39941 385056 39946 385112
rect 40002 385056 44362 385112
rect 44418 385056 44423 385112
rect 39941 385054 44423 385056
rect 39941 385051 40007 385054
rect 44357 385051 44423 385054
rect 35574 384709 35634 384812
rect 35574 384704 35683 384709
rect 35574 384648 35622 384704
rect 35678 384648 35683 384704
rect 35574 384646 35683 384648
rect 35617 384643 35683 384646
rect 35758 384301 35818 384404
rect 35758 384296 35867 384301
rect 35758 384240 35806 384296
rect 35862 384240 35867 384296
rect 35758 384238 35867 384240
rect 35801 384235 35867 384238
rect 35758 383893 35818 383996
rect 35758 383888 35867 383893
rect 35758 383832 35806 383888
rect 35862 383832 35867 383888
rect 35758 383830 35867 383832
rect 35801 383827 35867 383830
rect 39757 383890 39823 383893
rect 42793 383890 42859 383893
rect 39757 383888 42859 383890
rect 39757 383832 39762 383888
rect 39818 383832 42798 383888
rect 42854 383832 42859 383888
rect 39757 383830 42859 383832
rect 39757 383827 39823 383830
rect 42793 383827 42859 383830
rect 675293 383618 675359 383621
rect 676254 383618 676260 383620
rect 675293 383616 676260 383618
rect 35206 383485 35266 383588
rect 675293 383560 675298 383616
rect 675354 383560 676260 383616
rect 675293 383558 676260 383560
rect 675293 383555 675359 383558
rect 676254 383556 676260 383558
rect 676324 383556 676330 383620
rect 35206 383480 35315 383485
rect 35206 383424 35254 383480
rect 35310 383424 35315 383480
rect 35206 383422 35315 383424
rect 35249 383419 35315 383422
rect 40125 383482 40191 383485
rect 44633 383482 44699 383485
rect 40125 383480 44699 383482
rect 40125 383424 40130 383480
rect 40186 383424 44638 383480
rect 44694 383424 44699 383480
rect 40125 383422 44699 383424
rect 40125 383419 40191 383422
rect 44633 383419 44699 383422
rect 35390 383077 35450 383180
rect 35390 383072 35499 383077
rect 35390 383016 35438 383072
rect 35494 383016 35499 383072
rect 35390 383014 35499 383016
rect 35433 383011 35499 383014
rect 35758 382669 35818 382772
rect 35758 382664 35867 382669
rect 35758 382608 35806 382664
rect 35862 382608 35867 382664
rect 35758 382606 35867 382608
rect 35801 382603 35867 382606
rect 35574 382261 35634 382364
rect 35574 382256 35683 382261
rect 35574 382200 35622 382256
rect 35678 382200 35683 382256
rect 35574 382198 35683 382200
rect 35617 382195 35683 382198
rect 40033 382258 40099 382261
rect 675753 382260 675819 382261
rect 41454 382258 41460 382260
rect 40033 382256 41460 382258
rect 40033 382200 40038 382256
rect 40094 382200 41460 382256
rect 40033 382198 41460 382200
rect 40033 382195 40099 382198
rect 41454 382196 41460 382198
rect 41524 382196 41530 382260
rect 675702 382258 675708 382260
rect 675662 382198 675708 382258
rect 675772 382256 675819 382260
rect 675814 382200 675819 382256
rect 675702 382196 675708 382198
rect 675772 382196 675819 382200
rect 675753 382195 675819 382196
rect 35574 381853 35634 381956
rect 35574 381848 35683 381853
rect 35574 381792 35622 381848
rect 35678 381792 35683 381848
rect 35574 381790 35683 381792
rect 35617 381787 35683 381790
rect 39021 381850 39087 381853
rect 43621 381850 43687 381853
rect 39021 381848 43687 381850
rect 39021 381792 39026 381848
rect 39082 381792 43626 381848
rect 43682 381792 43687 381848
rect 39021 381790 43687 381792
rect 39021 381787 39087 381790
rect 43621 381787 43687 381790
rect 32446 381445 32506 381548
rect 32397 381440 32506 381445
rect 32397 381384 32402 381440
rect 32458 381384 32506 381440
rect 32397 381382 32506 381384
rect 32397 381379 32463 381382
rect 35758 381037 35818 381140
rect 35758 381032 35867 381037
rect 35758 380976 35806 381032
rect 35862 380976 35867 381032
rect 35758 380974 35867 380976
rect 35801 380971 35867 380974
rect 41413 381034 41479 381037
rect 44173 381034 44239 381037
rect 41413 381032 44239 381034
rect 41413 380976 41418 381032
rect 41474 380976 44178 381032
rect 44234 380976 44239 381032
rect 41413 380974 44239 380976
rect 41413 380971 41479 380974
rect 44173 380971 44239 380974
rect 35574 380629 35634 380732
rect 35574 380624 35683 380629
rect 35574 380568 35622 380624
rect 35678 380568 35683 380624
rect 35574 380566 35683 380568
rect 35617 380563 35683 380566
rect 675753 380626 675819 380629
rect 676438 380626 676444 380628
rect 675753 380624 676444 380626
rect 675753 380568 675758 380624
rect 675814 380568 676444 380624
rect 675753 380566 676444 380568
rect 675753 380563 675819 380566
rect 676438 380564 676444 380566
rect 676508 380564 676514 380628
rect 35758 380221 35818 380324
rect 35758 380216 35867 380221
rect 35758 380160 35806 380216
rect 35862 380160 35867 380216
rect 35758 380158 35867 380160
rect 35801 380155 35867 380158
rect 40033 380218 40099 380221
rect 41638 380218 41644 380220
rect 40033 380216 41644 380218
rect 40033 380160 40038 380216
rect 40094 380160 41644 380216
rect 40033 380158 41644 380160
rect 40033 380155 40099 380158
rect 41638 380156 41644 380158
rect 41708 380156 41714 380220
rect 35758 379813 35818 379916
rect 35758 379808 35867 379813
rect 35758 379752 35806 379808
rect 35862 379752 35867 379808
rect 35758 379750 35867 379752
rect 35801 379747 35867 379750
rect 40910 379404 40970 379508
rect 40902 379340 40908 379404
rect 40972 379340 40978 379404
rect 35758 378997 35818 379100
rect 35758 378992 35867 378997
rect 35758 378936 35806 378992
rect 35862 378936 35867 378992
rect 35758 378934 35867 378936
rect 35801 378931 35867 378934
rect 40217 378994 40283 378997
rect 41822 378994 41828 378996
rect 40217 378992 41828 378994
rect 40217 378936 40222 378992
rect 40278 378936 41828 378992
rect 40217 378934 41828 378936
rect 40217 378931 40283 378934
rect 41822 378932 41828 378934
rect 41892 378932 41898 378996
rect 40542 378588 40602 378692
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 41505 378586 41571 378589
rect 44357 378586 44423 378589
rect 41505 378584 44423 378586
rect 41505 378528 41510 378584
rect 41566 378528 44362 378584
rect 44418 378528 44423 378584
rect 41505 378526 44423 378528
rect 41505 378523 41571 378526
rect 44357 378523 44423 378526
rect 675661 378586 675727 378589
rect 675886 378586 675892 378588
rect 675661 378584 675892 378586
rect 675661 378528 675666 378584
rect 675722 378528 675892 378584
rect 675661 378526 675892 378528
rect 675661 378523 675727 378526
rect 675886 378524 675892 378526
rect 675956 378524 675962 378588
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 41229 378178 41295 378181
rect 43805 378178 43871 378181
rect 651557 378178 651623 378181
rect 41229 378176 43871 378178
rect 41229 378120 41234 378176
rect 41290 378120 43810 378176
rect 43866 378120 43871 378176
rect 41229 378118 43871 378120
rect 650164 378176 651623 378178
rect 650164 378120 651562 378176
rect 651618 378120 651623 378176
rect 650164 378118 651623 378120
rect 41229 378115 41295 378118
rect 43805 378115 43871 378118
rect 651557 378115 651623 378118
rect 35574 377773 35634 377876
rect 35574 377768 35683 377773
rect 35574 377712 35622 377768
rect 35678 377712 35683 377768
rect 35574 377710 35683 377712
rect 35617 377707 35683 377710
rect 39941 377770 40007 377773
rect 42977 377770 43043 377773
rect 39941 377768 43043 377770
rect 39941 377712 39946 377768
rect 40002 377712 42982 377768
rect 43038 377712 43043 377768
rect 39941 377710 43043 377712
rect 39941 377707 40007 377710
rect 42977 377707 43043 377710
rect 671153 377770 671219 377773
rect 674782 377770 674788 377772
rect 671153 377768 674788 377770
rect 671153 377712 671158 377768
rect 671214 377712 674788 377768
rect 671153 377710 674788 377712
rect 671153 377707 671219 377710
rect 674782 377708 674788 377710
rect 674852 377708 674858 377772
rect 35758 377365 35818 377468
rect 35758 377360 35867 377365
rect 35758 377304 35806 377360
rect 35862 377304 35867 377360
rect 35758 377302 35867 377304
rect 35801 377299 35867 377302
rect 39573 377362 39639 377365
rect 43253 377362 43319 377365
rect 39573 377360 43319 377362
rect 39573 377304 39578 377360
rect 39634 377304 43258 377360
rect 43314 377304 43319 377360
rect 39573 377302 43319 377304
rect 39573 377299 39639 377302
rect 43253 377299 43319 377302
rect 675753 377362 675819 377365
rect 676622 377362 676628 377364
rect 675753 377360 676628 377362
rect 675753 377304 675758 377360
rect 675814 377304 676628 377360
rect 675753 377302 676628 377304
rect 675753 377299 675819 377302
rect 676622 377300 676628 377302
rect 676692 377300 676698 377364
rect 28766 376549 28826 377060
rect 41689 376954 41755 376957
rect 45185 376954 45251 376957
rect 41689 376952 45251 376954
rect 41689 376896 41694 376952
rect 41750 376896 45190 376952
rect 45246 376896 45251 376952
rect 41689 376894 45251 376896
rect 41689 376891 41755 376894
rect 45185 376891 45251 376894
rect 673913 376818 673979 376821
rect 674925 376818 674991 376821
rect 673913 376816 674991 376818
rect 673913 376760 673918 376816
rect 673974 376760 674930 376816
rect 674986 376760 674991 376816
rect 673913 376758 674991 376760
rect 673913 376755 673979 376758
rect 674925 376755 674991 376758
rect 28766 376544 28875 376549
rect 28766 376488 28814 376544
rect 28870 376488 28875 376544
rect 28766 376486 28875 376488
rect 28809 376483 28875 376486
rect 62113 376274 62179 376277
rect 62113 376272 64492 376274
rect 35758 376141 35818 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 62113 376211 62179 376214
rect 35758 376136 35867 376141
rect 35758 376080 35806 376136
rect 35862 376080 35867 376136
rect 35758 376078 35867 376080
rect 35801 376075 35867 376078
rect 675293 375050 675359 375053
rect 676070 375050 676076 375052
rect 675293 375048 676076 375050
rect 675293 374992 675298 375048
rect 675354 374992 676076 375048
rect 675293 374990 676076 374992
rect 675293 374987 675359 374990
rect 676070 374988 676076 374990
rect 676140 374988 676146 375052
rect 674782 372540 674788 372604
rect 674852 372602 674858 372604
rect 675109 372602 675175 372605
rect 674852 372600 675175 372602
rect 674852 372544 675114 372600
rect 675170 372544 675175 372600
rect 674852 372542 675175 372544
rect 674852 372540 674858 372542
rect 675109 372539 675175 372542
rect 42057 369746 42123 369749
rect 44173 369746 44239 369749
rect 42057 369744 44239 369746
rect 42057 369688 42062 369744
rect 42118 369688 44178 369744
rect 44234 369688 44239 369744
rect 42057 369686 44239 369688
rect 42057 369683 42123 369686
rect 44173 369683 44239 369686
rect 40902 365604 40908 365668
rect 40972 365666 40978 365668
rect 41781 365666 41847 365669
rect 40972 365664 41847 365666
rect 40972 365608 41786 365664
rect 41842 365608 41847 365664
rect 40972 365606 41847 365608
rect 40972 365604 40978 365606
rect 41781 365603 41847 365606
rect 651557 364850 651623 364853
rect 650164 364848 651623 364850
rect 650164 364792 651562 364848
rect 651618 364792 651623 364848
rect 650164 364790 651623 364792
rect 651557 364787 651623 364790
rect 40718 363700 40724 363764
rect 40788 363762 40794 363764
rect 41781 363762 41847 363765
rect 40788 363760 41847 363762
rect 40788 363704 41786 363760
rect 41842 363704 41847 363760
rect 40788 363702 41847 363704
rect 40788 363700 40794 363702
rect 41781 363699 41847 363702
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 40534 360572 40540 360636
rect 40604 360634 40610 360636
rect 41781 360634 41847 360637
rect 40604 360632 41847 360634
rect 40604 360576 41786 360632
rect 41842 360576 41847 360632
rect 40604 360574 41847 360576
rect 40604 360572 40610 360574
rect 41781 360571 41847 360574
rect 41873 358732 41939 358733
rect 41822 358730 41828 358732
rect 41782 358670 41828 358730
rect 41892 358728 41939 358732
rect 41934 358672 41939 358728
rect 41822 358668 41828 358670
rect 41892 358668 41939 358672
rect 41873 358667 41939 358668
rect 675293 358730 675359 358733
rect 675293 358728 676292 358730
rect 675293 358672 675298 358728
rect 675354 358672 676292 358728
rect 675293 358670 676292 358672
rect 675293 358667 675359 358670
rect 675109 358322 675175 358325
rect 675109 358320 676292 358322
rect 675109 358264 675114 358320
rect 675170 358264 676292 358320
rect 675109 358262 676292 358264
rect 675109 358259 675175 358262
rect 675477 357914 675543 357917
rect 675477 357912 676292 357914
rect 675477 357856 675482 357912
rect 675538 357856 676292 357912
rect 675477 357854 676292 357856
rect 675477 357851 675543 357854
rect 674649 357506 674715 357509
rect 674649 357504 676292 357506
rect 674649 357448 674654 357504
rect 674710 357448 676292 357504
rect 674649 357446 676292 357448
rect 674649 357443 674715 357446
rect 675477 357098 675543 357101
rect 675477 357096 676292 357098
rect 675477 357040 675482 357096
rect 675538 357040 676292 357096
rect 675477 357038 676292 357040
rect 675477 357035 675543 357038
rect 41454 356900 41460 356964
rect 41524 356962 41530 356964
rect 41781 356962 41847 356965
rect 41524 356960 41847 356962
rect 41524 356904 41786 356960
rect 41842 356904 41847 356960
rect 41524 356902 41847 356904
rect 41524 356900 41530 356902
rect 41781 356899 41847 356902
rect 674465 356690 674531 356693
rect 674465 356688 676292 356690
rect 674465 356632 674470 356688
rect 674526 356632 676292 356688
rect 674465 356630 676292 356632
rect 674465 356627 674531 356630
rect 674649 356282 674715 356285
rect 674649 356280 676292 356282
rect 674649 356224 674654 356280
rect 674710 356224 676292 356280
rect 674649 356222 676292 356224
rect 674649 356219 674715 356222
rect 675477 355874 675543 355877
rect 675477 355872 676292 355874
rect 675477 355816 675482 355872
rect 675538 355816 676292 355872
rect 675477 355814 676292 355816
rect 675477 355811 675543 355814
rect 41965 355740 42031 355741
rect 41965 355736 42012 355740
rect 42076 355738 42082 355740
rect 41965 355680 41970 355736
rect 41965 355676 42012 355680
rect 42076 355678 42122 355738
rect 42076 355676 42082 355678
rect 41965 355675 42031 355676
rect 675477 355466 675543 355469
rect 675477 355464 676292 355466
rect 675477 355408 675482 355464
rect 675538 355408 676292 355464
rect 675477 355406 676292 355408
rect 675477 355403 675543 355406
rect 675477 355058 675543 355061
rect 675477 355056 676292 355058
rect 675477 355000 675482 355056
rect 675538 355000 676292 355056
rect 675477 354998 676292 355000
rect 675477 354995 675543 354998
rect 675477 354650 675543 354653
rect 675477 354648 676292 354650
rect 675477 354592 675482 354648
rect 675538 354592 676292 354648
rect 675477 354590 676292 354592
rect 675477 354587 675543 354590
rect 675334 354180 675340 354244
rect 675404 354242 675410 354244
rect 675404 354182 676292 354242
rect 675404 354180 675410 354182
rect 675477 353834 675543 353837
rect 675477 353832 676292 353834
rect 675477 353776 675482 353832
rect 675538 353776 676292 353832
rect 675477 353774 676292 353776
rect 675477 353771 675543 353774
rect 675477 353426 675543 353429
rect 675477 353424 676292 353426
rect 675477 353368 675482 353424
rect 675538 353368 676292 353424
rect 675477 353366 676292 353368
rect 675477 353363 675543 353366
rect 675518 352956 675524 353020
rect 675588 353018 675594 353020
rect 675588 352958 676292 353018
rect 675588 352956 675594 352958
rect 675477 352610 675543 352613
rect 675477 352608 676292 352610
rect 675477 352552 675482 352608
rect 675538 352552 676292 352608
rect 675477 352550 676292 352552
rect 675477 352547 675543 352550
rect 675702 352140 675708 352204
rect 675772 352202 675778 352204
rect 675772 352142 676292 352202
rect 675772 352140 675778 352142
rect 675886 351868 675892 351932
rect 675956 351930 675962 351932
rect 675956 351870 676230 351930
rect 675956 351868 675962 351870
rect 676170 351794 676230 351870
rect 676170 351734 676292 351794
rect 652017 351658 652083 351661
rect 650164 351656 652083 351658
rect 650164 351600 652022 351656
rect 652078 351600 652083 351656
rect 650164 351598 652083 351600
rect 652017 351595 652083 351598
rect 674465 351386 674531 351389
rect 674465 351384 676292 351386
rect 674465 351328 674470 351384
rect 674526 351328 676292 351384
rect 674465 351326 676292 351328
rect 674465 351323 674531 351326
rect 676029 350978 676095 350981
rect 676029 350976 676292 350978
rect 676029 350920 676034 350976
rect 676090 350920 676292 350976
rect 676029 350918 676292 350920
rect 676029 350915 676095 350918
rect 675845 350570 675911 350573
rect 675845 350568 676292 350570
rect 675845 350512 675850 350568
rect 675906 350512 676292 350568
rect 675845 350510 676292 350512
rect 675845 350507 675911 350510
rect 62113 350298 62179 350301
rect 62113 350296 64492 350298
rect 62113 350240 62118 350296
rect 62174 350240 64492 350296
rect 62113 350238 64492 350240
rect 62113 350235 62179 350238
rect 675477 350162 675543 350165
rect 675477 350160 676292 350162
rect 675477 350104 675482 350160
rect 675538 350104 676292 350160
rect 675477 350102 676292 350104
rect 675477 350099 675543 350102
rect 675477 349754 675543 349757
rect 675477 349752 676292 349754
rect 675477 349696 675482 349752
rect 675538 349696 676292 349752
rect 675477 349694 676292 349696
rect 675477 349691 675543 349694
rect 675477 349346 675543 349349
rect 675477 349344 676292 349346
rect 675477 349288 675482 349344
rect 675538 349288 676292 349344
rect 675477 349286 676292 349288
rect 675477 349283 675543 349286
rect 675477 348938 675543 348941
rect 675477 348936 676292 348938
rect 675477 348880 675482 348936
rect 675538 348880 676292 348936
rect 675477 348878 676292 348880
rect 675477 348875 675543 348878
rect 675477 348530 675543 348533
rect 675477 348528 676292 348530
rect 675477 348472 675482 348528
rect 675538 348472 676292 348528
rect 675477 348470 676292 348472
rect 675477 348467 675543 348470
rect 683070 347717 683130 348092
rect 683070 347712 683179 347717
rect 683070 347684 683118 347712
rect 683100 347656 683118 347684
rect 683174 347656 683179 347712
rect 683100 347654 683179 347656
rect 683113 347651 683179 347654
rect 675477 347306 675543 347309
rect 675477 347304 676292 347306
rect 675477 347248 675482 347304
rect 675538 347248 676292 347304
rect 675477 347246 676292 347248
rect 675477 347243 675543 347246
rect 676029 346626 676095 346629
rect 676438 346626 676444 346628
rect 676029 346624 676444 346626
rect 676029 346568 676034 346624
rect 676090 346568 676444 346624
rect 676029 346566 676444 346568
rect 676029 346563 676095 346566
rect 676438 346564 676444 346566
rect 676508 346564 676514 346628
rect 676581 346492 676647 346493
rect 676581 346488 676628 346492
rect 676692 346490 676698 346492
rect 676581 346432 676586 346488
rect 676581 346428 676628 346432
rect 676692 346430 676738 346490
rect 676692 346428 676698 346430
rect 676581 346427 676647 346428
rect 39205 345946 39271 345949
rect 46565 345946 46631 345949
rect 39205 345944 46631 345946
rect 39205 345888 39210 345944
rect 39266 345888 46570 345944
rect 46626 345888 46631 345944
rect 39205 345886 46631 345888
rect 39205 345883 39271 345886
rect 46565 345883 46631 345886
rect 35758 344317 35818 344556
rect 35758 344312 35867 344317
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35758 344254 35867 344256
rect 35801 344251 35867 344254
rect 35574 343909 35634 344148
rect 35574 343904 35683 343909
rect 35574 343848 35622 343904
rect 35678 343848 35683 343904
rect 35574 343846 35683 343848
rect 35617 343843 35683 343846
rect 35758 343501 35818 343740
rect 35758 343496 35867 343501
rect 35758 343440 35806 343496
rect 35862 343440 35867 343496
rect 35758 343438 35867 343440
rect 35801 343435 35867 343438
rect 35574 343093 35634 343332
rect 35574 343088 35683 343093
rect 35574 343032 35622 343088
rect 35678 343032 35683 343088
rect 35574 343030 35683 343032
rect 35617 343027 35683 343030
rect 40033 343090 40099 343093
rect 45369 343090 45435 343093
rect 40033 343088 45435 343090
rect 40033 343032 40038 343088
rect 40094 343032 45374 343088
rect 45430 343032 45435 343088
rect 40033 343030 45435 343032
rect 40033 343027 40099 343030
rect 45369 343027 45435 343030
rect 35758 342685 35818 342924
rect 35758 342680 35867 342685
rect 35758 342624 35806 342680
rect 35862 342624 35867 342680
rect 35758 342622 35867 342624
rect 35801 342619 35867 342622
rect 40309 342682 40375 342685
rect 43253 342682 43319 342685
rect 40309 342680 43319 342682
rect 40309 342624 40314 342680
rect 40370 342624 43258 342680
rect 43314 342624 43319 342680
rect 40309 342622 43319 342624
rect 40309 342619 40375 342622
rect 43253 342619 43319 342622
rect 35574 342277 35634 342516
rect 35574 342272 35683 342277
rect 35574 342216 35622 342272
rect 35678 342216 35683 342272
rect 35574 342214 35683 342216
rect 35617 342211 35683 342214
rect 670233 342274 670299 342277
rect 675845 342274 675911 342277
rect 670233 342272 675911 342274
rect 670233 342216 670238 342272
rect 670294 342216 675850 342272
rect 675906 342216 675911 342272
rect 670233 342214 675911 342216
rect 670233 342211 670299 342214
rect 675845 342211 675911 342214
rect 35758 341869 35818 342108
rect 35758 341864 35867 341869
rect 35758 341808 35806 341864
rect 35862 341808 35867 341864
rect 35758 341806 35867 341808
rect 35801 341803 35867 341806
rect 35390 341461 35450 341700
rect 35341 341456 35450 341461
rect 35617 341458 35683 341461
rect 35341 341400 35346 341456
rect 35402 341400 35450 341456
rect 35341 341398 35450 341400
rect 35574 341456 35683 341458
rect 35574 341400 35622 341456
rect 35678 341400 35683 341456
rect 35341 341395 35407 341398
rect 35574 341395 35683 341400
rect 35574 341292 35634 341395
rect 35801 341050 35867 341053
rect 35758 341048 35867 341050
rect 35758 340992 35806 341048
rect 35862 340992 35867 341048
rect 35758 340987 35867 340992
rect 35758 340884 35818 340987
rect 35758 340237 35818 340476
rect 35758 340232 35867 340237
rect 35758 340176 35806 340232
rect 35862 340176 35867 340232
rect 35758 340174 35867 340176
rect 35801 340171 35867 340174
rect 675753 340234 675819 340237
rect 676254 340234 676260 340236
rect 675753 340232 676260 340234
rect 675753 340176 675758 340232
rect 675814 340176 676260 340232
rect 675753 340174 676260 340176
rect 675753 340171 675819 340174
rect 676254 340172 676260 340174
rect 676324 340172 676330 340236
rect 41462 339828 41522 340068
rect 41454 339764 41460 339828
rect 41524 339764 41530 339828
rect 41278 339554 41338 339660
rect 41822 339554 41828 339556
rect 41278 339494 41828 339554
rect 41822 339492 41828 339494
rect 41892 339492 41898 339556
rect 35574 339013 35634 339252
rect 35574 339008 35683 339013
rect 35574 338952 35622 339008
rect 35678 338952 35683 339008
rect 35574 338950 35683 338952
rect 35617 338947 35683 338950
rect 41413 339010 41479 339013
rect 44265 339010 44331 339013
rect 675385 339012 675451 339013
rect 675334 339010 675340 339012
rect 41413 339008 44331 339010
rect 41413 338952 41418 339008
rect 41474 338952 44270 339008
rect 44326 338952 44331 339008
rect 41413 338950 44331 338952
rect 675294 338950 675340 339010
rect 675404 339008 675451 339012
rect 675446 338952 675451 339008
rect 41413 338947 41479 338950
rect 44265 338947 44331 338950
rect 675334 338948 675340 338950
rect 675404 338948 675451 338952
rect 675385 338947 675451 338948
rect 35801 338602 35867 338605
rect 35758 338600 35867 338602
rect 35758 338544 35806 338600
rect 35862 338544 35867 338600
rect 35758 338539 35867 338544
rect 41462 338602 41522 338844
rect 41781 338738 41847 338741
rect 45553 338738 45619 338741
rect 41781 338736 45619 338738
rect 41781 338680 41786 338736
rect 41842 338680 45558 338736
rect 45614 338680 45619 338736
rect 41781 338678 45619 338680
rect 41781 338675 41847 338678
rect 45553 338675 45619 338678
rect 41638 338602 41644 338604
rect 41462 338542 41644 338602
rect 41638 338540 41644 338542
rect 41708 338540 41714 338604
rect 35758 338436 35818 338539
rect 652201 338330 652267 338333
rect 650164 338328 652267 338330
rect 650164 338272 652206 338328
rect 652262 338272 652267 338328
rect 650164 338270 652267 338272
rect 652201 338267 652267 338270
rect 41689 338194 41755 338197
rect 45369 338194 45435 338197
rect 41689 338192 45435 338194
rect 41689 338136 41694 338192
rect 41750 338136 45374 338192
rect 45430 338136 45435 338192
rect 41689 338134 45435 338136
rect 41689 338131 41755 338134
rect 45369 338131 45435 338134
rect 35758 337789 35818 338028
rect 35758 337784 35867 337789
rect 35758 337728 35806 337784
rect 35862 337728 35867 337784
rect 35758 337726 35867 337728
rect 35801 337723 35867 337726
rect 675661 337786 675727 337789
rect 675886 337786 675892 337788
rect 675661 337784 675892 337786
rect 675661 337728 675666 337784
rect 675722 337728 675892 337784
rect 675661 337726 675892 337728
rect 675661 337723 675727 337726
rect 675886 337724 675892 337726
rect 675956 337724 675962 337788
rect 40542 337380 40602 337620
rect 40534 337316 40540 337380
rect 40604 337316 40610 337380
rect 62113 337242 62179 337245
rect 62113 337240 64492 337242
rect 35574 336973 35634 337212
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 62113 337179 62179 337182
rect 35525 336968 35634 336973
rect 35801 336970 35867 336973
rect 35525 336912 35530 336968
rect 35586 336912 35634 336968
rect 35525 336910 35634 336912
rect 35758 336968 35867 336970
rect 35758 336912 35806 336968
rect 35862 336912 35867 336968
rect 35525 336907 35591 336910
rect 35758 336907 35867 336912
rect 35758 336804 35818 336907
rect 40726 336156 40786 336396
rect 40718 336092 40724 336156
rect 40788 336092 40794 336156
rect 35574 335749 35634 335988
rect 35574 335744 35683 335749
rect 35574 335688 35622 335744
rect 35678 335688 35683 335744
rect 35574 335686 35683 335688
rect 35617 335683 35683 335686
rect 40309 335746 40375 335749
rect 43805 335746 43871 335749
rect 40309 335744 43871 335746
rect 40309 335688 40314 335744
rect 40370 335688 43810 335744
rect 43866 335688 43871 335744
rect 40309 335686 43871 335688
rect 40309 335683 40375 335686
rect 43805 335683 43871 335686
rect 35801 335610 35867 335613
rect 35788 335608 35867 335610
rect 35788 335552 35806 335608
rect 35862 335552 35867 335608
rect 35788 335550 35867 335552
rect 35801 335547 35867 335550
rect 675293 335338 675359 335341
rect 676438 335338 676444 335340
rect 675293 335336 676444 335338
rect 675293 335280 675298 335336
rect 675354 335280 676444 335336
rect 675293 335278 676444 335280
rect 675293 335275 675359 335278
rect 676438 335276 676444 335278
rect 676508 335276 676514 335340
rect 35574 334933 35634 335172
rect 35574 334928 35683 334933
rect 35574 334872 35622 334928
rect 35678 334872 35683 334928
rect 35574 334870 35683 334872
rect 35617 334867 35683 334870
rect 40217 334930 40283 334933
rect 43989 334930 44055 334933
rect 40217 334928 44055 334930
rect 40217 334872 40222 334928
rect 40278 334872 43994 334928
rect 44050 334872 44055 334928
rect 40217 334870 44055 334872
rect 40217 334867 40283 334870
rect 43989 334867 44055 334870
rect 35390 334525 35450 334764
rect 35390 334520 35499 334525
rect 35801 334522 35867 334525
rect 35390 334464 35438 334520
rect 35494 334464 35499 334520
rect 35390 334462 35499 334464
rect 35433 334459 35499 334462
rect 35758 334520 35867 334522
rect 35758 334464 35806 334520
rect 35862 334464 35867 334520
rect 35758 334459 35867 334464
rect 35758 334356 35818 334459
rect 35758 333301 35818 333948
rect 40309 333706 40375 333709
rect 46013 333706 46079 333709
rect 40309 333704 46079 333706
rect 40309 333648 40314 333704
rect 40370 333648 46018 333704
rect 46074 333648 46079 333704
rect 40309 333646 46079 333648
rect 40309 333643 40375 333646
rect 46013 333643 46079 333646
rect 35758 333296 35867 333301
rect 35758 333240 35806 333296
rect 35862 333240 35867 333296
rect 35758 333238 35867 333240
rect 35801 333235 35867 333238
rect 35758 332893 35818 333132
rect 35758 332888 35867 332893
rect 35758 332832 35806 332888
rect 35862 332832 35867 332888
rect 35758 332830 35867 332832
rect 35801 332827 35867 332830
rect 39849 332890 39915 332893
rect 45829 332890 45895 332893
rect 39849 332888 45895 332890
rect 39849 332832 39854 332888
rect 39910 332832 45834 332888
rect 45890 332832 45895 332888
rect 39849 332830 45895 332832
rect 39849 332827 39915 332830
rect 45829 332827 45895 332830
rect 40861 332482 40927 332485
rect 43069 332482 43135 332485
rect 40861 332480 43135 332482
rect 40861 332424 40866 332480
rect 40922 332424 43074 332480
rect 43130 332424 43135 332480
rect 40861 332422 43135 332424
rect 40861 332419 40927 332422
rect 43069 332419 43135 332422
rect 40125 331258 40191 331261
rect 46749 331258 46815 331261
rect 676622 331258 676628 331260
rect 40125 331256 46815 331258
rect 40125 331200 40130 331256
rect 40186 331200 46754 331256
rect 46810 331200 46815 331256
rect 40125 331198 46815 331200
rect 40125 331195 40191 331198
rect 46749 331195 46815 331198
rect 675342 331198 676628 331258
rect 675342 331125 675402 331198
rect 676622 331196 676628 331198
rect 676692 331196 676698 331260
rect 675293 331120 675402 331125
rect 675293 331064 675298 331120
rect 675354 331064 675402 331120
rect 675293 331062 675402 331064
rect 675293 331059 675359 331062
rect 39297 330714 39363 330717
rect 44633 330714 44699 330717
rect 39297 330712 44699 330714
rect 39297 330656 39302 330712
rect 39358 330656 44638 330712
rect 44694 330656 44699 330712
rect 39297 330654 44699 330656
rect 39297 330651 39363 330654
rect 44633 330651 44699 330654
rect 675753 326906 675819 326909
rect 676070 326906 676076 326908
rect 675753 326904 676076 326906
rect 675753 326848 675758 326904
rect 675814 326848 676076 326904
rect 675753 326846 676076 326848
rect 675753 326843 675819 326846
rect 676070 326844 676076 326846
rect 676140 326844 676146 326908
rect 651557 325002 651623 325005
rect 650164 325000 651623 325002
rect 650164 324944 651562 325000
rect 651618 324944 651623 325000
rect 650164 324942 651623 324944
rect 651557 324939 651623 324942
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 62757 324186 62823 324189
rect 62757 324184 64492 324186
rect 62757 324128 62762 324184
rect 62818 324128 64492 324184
rect 62757 324126 64492 324128
rect 62757 324123 62823 324126
rect 40718 322764 40724 322828
rect 40788 322826 40794 322828
rect 41781 322826 41847 322829
rect 40788 322824 41847 322826
rect 40788 322768 41786 322824
rect 41842 322768 41847 322824
rect 40788 322766 41847 322768
rect 40788 322764 40794 322766
rect 41781 322763 41847 322766
rect 41781 315620 41847 315621
rect 41781 315616 41828 315620
rect 41892 315618 41898 315620
rect 41781 315560 41786 315616
rect 41781 315556 41828 315560
rect 41892 315558 41938 315618
rect 41892 315556 41898 315558
rect 41781 315555 41847 315556
rect 41454 313652 41460 313716
rect 41524 313714 41530 313716
rect 41781 313714 41847 313717
rect 41524 313712 41847 313714
rect 41524 313656 41786 313712
rect 41842 313656 41847 313712
rect 41524 313654 41847 313656
rect 41524 313652 41530 313654
rect 41781 313651 41847 313654
rect 675477 313714 675543 313717
rect 675477 313712 676292 313714
rect 675477 313656 675482 313712
rect 675538 313656 676292 313712
rect 675477 313654 676292 313656
rect 675477 313651 675543 313654
rect 675477 313306 675543 313309
rect 675477 313304 676292 313306
rect 675477 313248 675482 313304
rect 675538 313248 676292 313304
rect 675477 313246 676292 313248
rect 675477 313243 675543 313246
rect 40534 312972 40540 313036
rect 40604 313034 40610 313036
rect 41781 313034 41847 313037
rect 40604 313032 41847 313034
rect 40604 312976 41786 313032
rect 41842 312976 41847 313032
rect 40604 312974 41847 312976
rect 40604 312972 40610 312974
rect 41781 312971 41847 312974
rect 675293 312898 675359 312901
rect 675293 312896 676292 312898
rect 675293 312840 675298 312896
rect 675354 312840 676292 312896
rect 675293 312838 676292 312840
rect 675293 312835 675359 312838
rect 675477 312490 675543 312493
rect 675477 312488 676292 312490
rect 675477 312432 675482 312488
rect 675538 312432 676292 312488
rect 675477 312430 676292 312432
rect 675477 312427 675543 312430
rect 675477 312082 675543 312085
rect 675477 312080 676292 312082
rect 675477 312024 675482 312080
rect 675538 312024 676292 312080
rect 675477 312022 676292 312024
rect 675477 312019 675543 312022
rect 651557 311810 651623 311813
rect 650164 311808 651623 311810
rect 650164 311752 651562 311808
rect 651618 311752 651623 311808
rect 650164 311750 651623 311752
rect 651557 311747 651623 311750
rect 674649 311674 674715 311677
rect 674649 311672 676292 311674
rect 674649 311616 674654 311672
rect 674710 311616 676292 311672
rect 674649 311614 676292 311616
rect 674649 311611 674715 311614
rect 675477 311266 675543 311269
rect 675477 311264 676292 311266
rect 675477 311208 675482 311264
rect 675538 311208 676292 311264
rect 675477 311206 676292 311208
rect 675477 311203 675543 311206
rect 62757 311130 62823 311133
rect 62757 311128 64492 311130
rect 62757 311072 62762 311128
rect 62818 311072 64492 311128
rect 62757 311070 64492 311072
rect 62757 311067 62823 311070
rect 672717 310858 672783 310861
rect 672717 310856 676292 310858
rect 672717 310800 672722 310856
rect 672778 310800 676292 310856
rect 672717 310798 676292 310800
rect 672717 310795 672783 310798
rect 675477 310450 675543 310453
rect 675477 310448 676292 310450
rect 675477 310392 675482 310448
rect 675538 310392 676292 310448
rect 675477 310390 676292 310392
rect 675477 310387 675543 310390
rect 675477 310042 675543 310045
rect 675477 310040 676292 310042
rect 675477 309984 675482 310040
rect 675538 309984 676292 310040
rect 675477 309982 676292 309984
rect 675477 309979 675543 309982
rect 675477 309634 675543 309637
rect 675477 309632 676292 309634
rect 675477 309576 675482 309632
rect 675538 309576 676292 309632
rect 675477 309574 676292 309576
rect 675477 309571 675543 309574
rect 675201 309226 675267 309229
rect 675201 309224 676292 309226
rect 675201 309168 675206 309224
rect 675262 309168 676292 309224
rect 675201 309166 676292 309168
rect 675201 309163 675267 309166
rect 675518 308756 675524 308820
rect 675588 308818 675594 308820
rect 675588 308758 676292 308818
rect 675588 308756 675594 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675017 308002 675083 308005
rect 675017 308000 676292 308002
rect 675017 307944 675022 308000
rect 675078 307944 676292 308000
rect 675017 307942 676292 307944
rect 675017 307939 675083 307942
rect 674833 307594 674899 307597
rect 674833 307592 676292 307594
rect 674833 307536 674838 307592
rect 674894 307536 676292 307592
rect 674833 307534 676292 307536
rect 674833 307531 674899 307534
rect 678237 307186 678303 307189
rect 678237 307184 678316 307186
rect 678237 307128 678242 307184
rect 678298 307128 678316 307184
rect 678237 307126 678316 307128
rect 678237 307123 678303 307126
rect 680997 306778 681063 306781
rect 680997 306776 681076 306778
rect 680997 306720 681002 306776
rect 681058 306720 681076 306776
rect 680997 306718 681076 306720
rect 680997 306715 681063 306718
rect 674465 306370 674531 306373
rect 674465 306368 676292 306370
rect 674465 306312 674470 306368
rect 674526 306312 676292 306368
rect 674465 306310 676292 306312
rect 674465 306307 674531 306310
rect 675702 305900 675708 305964
rect 675772 305962 675778 305964
rect 675772 305902 676292 305962
rect 675772 305900 675778 305902
rect 675477 305554 675543 305557
rect 675477 305552 676292 305554
rect 675477 305496 675482 305552
rect 675538 305496 676292 305552
rect 675477 305494 676292 305496
rect 675477 305491 675543 305494
rect 675845 305146 675911 305149
rect 675845 305144 676292 305146
rect 675845 305088 675850 305144
rect 675906 305088 676292 305144
rect 675845 305086 676292 305088
rect 675845 305083 675911 305086
rect 676029 304738 676095 304741
rect 676029 304736 676292 304738
rect 676029 304680 676034 304736
rect 676090 304680 676292 304736
rect 676029 304678 676292 304680
rect 676029 304675 676095 304678
rect 674649 304330 674715 304333
rect 674649 304328 676292 304330
rect 674649 304272 674654 304328
rect 674710 304272 676292 304328
rect 674649 304270 676292 304272
rect 674649 304267 674715 304270
rect 675477 303922 675543 303925
rect 675477 303920 676292 303922
rect 675477 303864 675482 303920
rect 675538 303864 676292 303920
rect 675477 303862 676292 303864
rect 675477 303859 675543 303862
rect 675477 303514 675543 303517
rect 675477 303512 676292 303514
rect 675477 303456 675482 303512
rect 675538 303456 676292 303512
rect 675477 303454 676292 303456
rect 675477 303451 675543 303454
rect 676029 302972 676095 302973
rect 676029 302970 676076 302972
rect 675984 302968 676076 302970
rect 675984 302912 676034 302968
rect 675984 302910 676076 302912
rect 676029 302908 676076 302910
rect 676140 302908 676146 302972
rect 676029 302907 676095 302908
rect 677182 302698 677242 303076
rect 683113 302698 683179 302701
rect 677182 302696 683179 302698
rect 677182 302668 683118 302696
rect 677212 302640 683118 302668
rect 683174 302640 683179 302696
rect 677212 302638 683179 302640
rect 683113 302635 683179 302638
rect 675477 302290 675543 302293
rect 675477 302288 676292 302290
rect 675477 302232 675482 302288
rect 675538 302232 676292 302288
rect 675477 302230 676292 302232
rect 675477 302227 675543 302230
rect 675845 301610 675911 301613
rect 676622 301610 676628 301612
rect 675845 301608 676628 301610
rect 675845 301552 675850 301608
rect 675906 301552 676628 301608
rect 675845 301550 676628 301552
rect 675845 301547 675911 301550
rect 676622 301548 676628 301550
rect 676692 301548 676698 301612
rect 43069 301338 43135 301341
rect 41492 301336 43135 301338
rect 41492 301280 43074 301336
rect 43130 301280 43135 301336
rect 41492 301278 43135 301280
rect 43069 301275 43135 301278
rect 43621 300930 43687 300933
rect 41492 300928 43687 300930
rect 41492 300872 43626 300928
rect 43682 300872 43687 300928
rect 41492 300870 43687 300872
rect 43621 300867 43687 300870
rect 40953 300522 41019 300525
rect 40940 300520 41019 300522
rect 40940 300464 40958 300520
rect 41014 300464 41019 300520
rect 40940 300462 41019 300464
rect 40953 300459 41019 300462
rect 41137 300114 41203 300117
rect 41124 300112 41203 300114
rect 41124 300056 41142 300112
rect 41198 300056 41203 300112
rect 41124 300054 41203 300056
rect 41137 300051 41203 300054
rect 43069 299706 43135 299709
rect 41492 299704 43135 299706
rect 41492 299648 43074 299704
rect 43130 299648 43135 299704
rect 41492 299646 43135 299648
rect 43069 299643 43135 299646
rect 675886 299372 675892 299436
rect 675956 299434 675962 299436
rect 680353 299434 680419 299437
rect 675956 299432 680419 299434
rect 675956 299376 680358 299432
rect 680414 299376 680419 299432
rect 675956 299374 680419 299376
rect 675956 299372 675962 299374
rect 680353 299371 680419 299374
rect 41137 299298 41203 299301
rect 41124 299296 41203 299298
rect 41124 299240 41142 299296
rect 41198 299240 41203 299296
rect 41124 299238 41203 299240
rect 41137 299235 41203 299238
rect 42701 298890 42767 298893
rect 41492 298888 42767 298890
rect 41492 298832 42706 298888
rect 42762 298832 42767 298888
rect 41492 298830 42767 298832
rect 42701 298827 42767 298830
rect 40953 298482 41019 298485
rect 652201 298482 652267 298485
rect 40940 298480 41019 298482
rect 40940 298424 40958 298480
rect 41014 298424 41019 298480
rect 40940 298422 41019 298424
rect 650164 298480 652267 298482
rect 650164 298424 652206 298480
rect 652262 298424 652267 298480
rect 650164 298422 652267 298424
rect 40953 298419 41019 298422
rect 652201 298419 652267 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 40953 298074 41019 298077
rect 40940 298072 41019 298074
rect 40940 298016 40958 298072
rect 41014 298016 41019 298072
rect 40940 298014 41019 298016
rect 40953 298011 41019 298014
rect 41137 297666 41203 297669
rect 41124 297664 41203 297666
rect 41124 297608 41142 297664
rect 41198 297608 41203 297664
rect 41124 297606 41203 297608
rect 41137 297603 41203 297606
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 678237 297394 678303 297397
rect 675772 297392 678303 297394
rect 675772 297336 678242 297392
rect 678298 297336 678303 297392
rect 675772 297334 678303 297336
rect 675772 297332 675778 297334
rect 678237 297331 678303 297334
rect 44357 297258 44423 297261
rect 41492 297256 44423 297258
rect 41492 297200 44362 297256
rect 44418 297200 44423 297256
rect 41492 297198 44423 297200
rect 44357 297195 44423 297198
rect 41822 296850 41828 296852
rect 41492 296790 41828 296850
rect 41822 296788 41828 296790
rect 41892 296788 41898 296852
rect 42006 296442 42012 296444
rect 41492 296382 42012 296442
rect 42006 296380 42012 296382
rect 42076 296380 42082 296444
rect 45553 296034 45619 296037
rect 41492 296032 45619 296034
rect 41492 295976 45558 296032
rect 45614 295976 45619 296032
rect 41492 295974 45619 295976
rect 45553 295971 45619 295974
rect 40769 295626 40835 295629
rect 40756 295624 40835 295626
rect 40756 295568 40774 295624
rect 40830 295568 40835 295624
rect 40756 295566 40835 295568
rect 40769 295563 40835 295566
rect 41781 295218 41847 295221
rect 41492 295216 41847 295218
rect 41492 295160 41786 295216
rect 41842 295160 41847 295216
rect 41492 295158 41847 295160
rect 41781 295155 41847 295158
rect 37917 294810 37983 294813
rect 37917 294808 37996 294810
rect 37917 294752 37922 294808
rect 37978 294752 37996 294808
rect 37917 294750 37996 294752
rect 37917 294747 37983 294750
rect 41781 294538 41847 294541
rect 47025 294538 47091 294541
rect 41781 294536 47091 294538
rect 41781 294480 41786 294536
rect 41842 294480 47030 294536
rect 47086 294480 47091 294536
rect 41781 294478 47091 294480
rect 41781 294475 41847 294478
rect 47025 294475 47091 294478
rect 41321 294402 41387 294405
rect 41308 294400 41387 294402
rect 41308 294344 41326 294400
rect 41382 294344 41387 294400
rect 41308 294342 41387 294344
rect 41321 294339 41387 294342
rect 45369 293994 45435 293997
rect 41492 293992 45435 293994
rect 41492 293936 45374 293992
rect 45430 293936 45435 293992
rect 41492 293934 45435 293936
rect 45369 293931 45435 293934
rect 41781 293586 41847 293589
rect 41492 293584 41847 293586
rect 41492 293528 41786 293584
rect 41842 293528 41847 293584
rect 41492 293526 41847 293528
rect 41781 293523 41847 293526
rect 42977 293178 43043 293181
rect 41492 293176 43043 293178
rect 41492 293120 42982 293176
rect 43038 293120 43043 293176
rect 41492 293118 43043 293120
rect 42977 293115 43043 293118
rect 40493 292592 40559 292593
rect 40726 292592 40786 292740
rect 40493 292590 40540 292592
rect 40448 292588 40540 292590
rect 40448 292532 40498 292588
rect 40448 292530 40540 292532
rect 40493 292528 40540 292530
rect 40604 292528 40610 292592
rect 40718 292528 40724 292592
rect 40788 292528 40794 292592
rect 40902 292528 40908 292592
rect 40972 292528 40978 292592
rect 40493 292527 40559 292528
rect 40910 292332 40970 292528
rect 41781 292092 41847 292093
rect 41781 292088 41828 292092
rect 41892 292090 41898 292092
rect 41781 292032 41786 292088
rect 41781 292028 41828 292032
rect 41892 292030 41938 292090
rect 41892 292028 41898 292030
rect 41781 292027 41847 292028
rect 41137 291954 41203 291957
rect 41124 291952 41203 291954
rect 41124 291896 41142 291952
rect 41198 291896 41203 291952
rect 41124 291894 41203 291896
rect 41137 291891 41203 291894
rect 44173 291546 44239 291549
rect 41492 291544 44239 291546
rect 41492 291488 44178 291544
rect 44234 291488 44239 291544
rect 41492 291486 44239 291488
rect 44173 291483 44239 291486
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 40953 291138 41019 291141
rect 40940 291136 41019 291138
rect 40940 291080 40958 291136
rect 41014 291080 41019 291136
rect 40940 291078 41019 291080
rect 40953 291075 41019 291078
rect 675753 291002 675819 291005
rect 676254 291002 676260 291004
rect 675753 291000 676260 291002
rect 675753 290944 675758 291000
rect 675814 290944 676260 291000
rect 675753 290942 676260 290944
rect 675753 290939 675819 290942
rect 676254 290940 676260 290942
rect 676324 290940 676330 291004
rect 43621 290730 43687 290733
rect 41492 290728 43687 290730
rect 41492 290672 43626 290728
rect 43682 290672 43687 290728
rect 41492 290670 43687 290672
rect 43621 290667 43687 290670
rect 41137 290322 41203 290325
rect 41124 290320 41203 290322
rect 41124 290264 41142 290320
rect 41198 290264 41203 290320
rect 41124 290262 41203 290264
rect 41137 290259 41203 290262
rect 41278 289830 41338 289884
rect 41278 289770 42074 289830
rect 42014 289645 42074 289770
rect 41965 289640 42074 289645
rect 41965 289584 41970 289640
rect 42026 289584 42074 289640
rect 41965 289582 42074 289584
rect 41965 289579 42031 289582
rect 675753 287058 675819 287061
rect 676622 287058 676628 287060
rect 675753 287056 676628 287058
rect 675753 287000 675758 287056
rect 675814 287000 676628 287056
rect 675753 286998 676628 287000
rect 675753 286995 675819 286998
rect 676622 286996 676628 286998
rect 676692 286996 676698 287060
rect 673085 286514 673151 286517
rect 675385 286514 675451 286517
rect 673085 286512 675451 286514
rect 673085 286456 673090 286512
rect 673146 286456 675390 286512
rect 675446 286456 675451 286512
rect 673085 286454 675451 286456
rect 673085 286451 673151 286454
rect 675385 286451 675451 286454
rect 673269 285562 673335 285565
rect 675109 285562 675175 285565
rect 673269 285560 675175 285562
rect 673269 285504 673274 285560
rect 673330 285504 675114 285560
rect 675170 285504 675175 285560
rect 673269 285502 675175 285504
rect 673269 285499 673335 285502
rect 675109 285499 675175 285502
rect 651557 285290 651623 285293
rect 650164 285288 651623 285290
rect 650164 285232 651562 285288
rect 651618 285232 651623 285288
rect 650164 285230 651623 285232
rect 651557 285227 651623 285230
rect 62113 285154 62179 285157
rect 62113 285152 64492 285154
rect 62113 285096 62118 285152
rect 62174 285096 64492 285152
rect 62113 285094 64492 285096
rect 62113 285091 62179 285094
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 675661 282842 675727 282845
rect 675886 282842 675892 282844
rect 675661 282840 675892 282842
rect 675661 282784 675666 282840
rect 675722 282784 675892 282840
rect 675661 282782 675892 282784
rect 675661 282779 675727 282782
rect 675886 282780 675892 282782
rect 675956 282780 675962 282844
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 41965 281484 42031 281485
rect 41965 281480 42012 281484
rect 42076 281482 42082 281484
rect 41965 281424 41970 281480
rect 41965 281420 42012 281424
rect 42076 281422 42122 281482
rect 42076 281420 42082 281422
rect 41965 281419 42031 281420
rect 40902 278700 40908 278764
rect 40972 278762 40978 278764
rect 42517 278762 42583 278765
rect 40972 278760 42583 278762
rect 40972 278704 42522 278760
rect 42578 278704 42583 278760
rect 40972 278702 42583 278704
rect 40972 278700 40978 278702
rect 42517 278699 42583 278702
rect 673085 278764 673151 278765
rect 673085 278760 673132 278764
rect 673196 278762 673202 278764
rect 673085 278704 673090 278760
rect 673085 278700 673132 278704
rect 673196 278702 673242 278762
rect 673196 278700 673202 278702
rect 673085 278699 673151 278700
rect 673862 278564 673868 278628
rect 673932 278564 673938 278628
rect 54477 278082 54543 278085
rect 641989 278082 642055 278085
rect 54477 278080 642055 278082
rect 54477 278024 54482 278080
rect 54538 278024 641994 278080
rect 642050 278024 642055 278080
rect 54477 278022 642055 278024
rect 54477 278019 54543 278022
rect 641989 278019 642055 278022
rect 673870 277676 673930 278564
rect 673862 277612 673868 277676
rect 673932 277612 673938 277676
rect 40718 277340 40724 277404
rect 40788 277402 40794 277404
rect 41781 277402 41847 277405
rect 40788 277400 41847 277402
rect 40788 277344 41786 277400
rect 41842 277344 41847 277400
rect 40788 277342 41847 277344
rect 40788 277340 40794 277342
rect 41781 277339 41847 277342
rect 499573 277402 499639 277405
rect 502333 277402 502399 277405
rect 499573 277400 502399 277402
rect 499573 277344 499578 277400
rect 499634 277344 502338 277400
rect 502394 277344 502399 277400
rect 499573 277342 502399 277344
rect 499573 277339 499639 277342
rect 502333 277339 502399 277342
rect 53465 276994 53531 276997
rect 656893 276994 656959 276997
rect 53465 276992 656959 276994
rect 53465 276936 53470 276992
rect 53526 276936 656898 276992
rect 656954 276936 656959 276992
rect 53465 276934 656959 276936
rect 53465 276931 53531 276934
rect 656893 276931 656959 276934
rect 45001 276722 45067 276725
rect 648705 276722 648771 276725
rect 45001 276720 648771 276722
rect 45001 276664 45006 276720
rect 45062 276664 648710 276720
rect 648766 276664 648771 276720
rect 45001 276662 648771 276664
rect 45001 276659 45067 276662
rect 648705 276659 648771 276662
rect 497457 276450 497523 276453
rect 508865 276450 508931 276453
rect 497457 276448 508931 276450
rect 497457 276392 497462 276448
rect 497518 276392 508870 276448
rect 508926 276392 508931 276448
rect 497457 276390 508931 276392
rect 497457 276387 497523 276390
rect 508865 276387 508931 276390
rect 491845 276178 491911 276181
rect 499205 276178 499271 276181
rect 491845 276176 499271 276178
rect 491845 276120 491850 276176
rect 491906 276120 499210 276176
rect 499266 276120 499271 276176
rect 491845 276118 499271 276120
rect 491845 276115 491911 276118
rect 499205 276115 499271 276118
rect 483013 276042 483079 276045
rect 489913 276042 489979 276045
rect 483013 276040 489979 276042
rect 483013 275984 483018 276040
rect 483074 275984 489918 276040
rect 489974 275984 489979 276040
rect 483013 275982 489979 275984
rect 483013 275979 483079 275982
rect 489913 275979 489979 275982
rect 490097 276042 490163 276045
rect 491477 276042 491543 276045
rect 490097 276040 491543 276042
rect 490097 275984 490102 276040
rect 490158 275984 491482 276040
rect 491538 275984 491543 276040
rect 490097 275982 491543 275984
rect 490097 275979 490163 275982
rect 491477 275979 491543 275982
rect 499389 276042 499455 276045
rect 499757 276042 499823 276045
rect 499389 276040 499823 276042
rect 499389 275984 499394 276040
rect 499450 275984 499762 276040
rect 499818 275984 499823 276040
rect 499389 275982 499823 275984
rect 499389 275979 499455 275982
rect 499757 275979 499823 275982
rect 399661 275770 399727 275773
rect 400765 275770 400831 275773
rect 399661 275768 400831 275770
rect 399661 275712 399666 275768
rect 399722 275712 400770 275768
rect 400826 275712 400831 275768
rect 399661 275710 400831 275712
rect 399661 275707 399727 275710
rect 400765 275707 400831 275710
rect 480161 275770 480227 275773
rect 480345 275770 480411 275773
rect 480161 275768 480411 275770
rect 480161 275712 480166 275768
rect 480222 275712 480350 275768
rect 480406 275712 480411 275768
rect 480161 275710 480411 275712
rect 480161 275707 480227 275710
rect 480345 275707 480411 275710
rect 489729 275770 489795 275773
rect 490005 275770 490071 275773
rect 489729 275768 490071 275770
rect 489729 275712 489734 275768
rect 489790 275712 490010 275768
rect 490066 275712 490071 275768
rect 489729 275710 490071 275712
rect 489729 275707 489795 275710
rect 490005 275707 490071 275710
rect 501137 275770 501203 275773
rect 504725 275770 504791 275773
rect 501137 275768 504791 275770
rect 501137 275712 501142 275768
rect 501198 275712 504730 275768
rect 504786 275712 504791 275768
rect 501137 275710 504791 275712
rect 501137 275707 501203 275710
rect 504725 275707 504791 275710
rect 509233 275770 509299 275773
rect 512177 275770 512243 275773
rect 509233 275768 512243 275770
rect 509233 275712 509238 275768
rect 509294 275712 512182 275768
rect 512238 275712 512243 275768
rect 509233 275710 512243 275712
rect 509233 275707 509299 275710
rect 512177 275707 512243 275710
rect 446213 275498 446279 275501
rect 541065 275498 541131 275501
rect 446213 275496 541131 275498
rect 446213 275440 446218 275496
rect 446274 275440 541070 275496
rect 541126 275440 541131 275496
rect 446213 275438 541131 275440
rect 446213 275435 446279 275438
rect 541065 275435 541131 275438
rect 481449 275226 481515 275229
rect 619081 275226 619147 275229
rect 481449 275224 619147 275226
rect 481449 275168 481454 275224
rect 481510 275168 619086 275224
rect 619142 275168 619147 275224
rect 481449 275166 619147 275168
rect 481449 275163 481515 275166
rect 619081 275163 619147 275166
rect 489913 274954 489979 274957
rect 494973 274954 495039 274957
rect 489913 274952 495039 274954
rect 489913 274896 489918 274952
rect 489974 274896 494978 274952
rect 495034 274896 495039 274952
rect 489913 274894 495039 274896
rect 489913 274891 489979 274894
rect 494973 274891 495039 274894
rect 470225 274682 470291 274685
rect 472157 274682 472223 274685
rect 470225 274680 472223 274682
rect 470225 274624 470230 274680
rect 470286 274624 472162 274680
rect 472218 274624 472223 274680
rect 470225 274622 472223 274624
rect 470225 274619 470291 274622
rect 472157 274619 472223 274622
rect 503621 274682 503687 274685
rect 509325 274682 509391 274685
rect 503621 274680 509391 274682
rect 503621 274624 503626 274680
rect 503682 274624 509330 274680
rect 509386 274624 509391 274680
rect 503621 274622 509391 274624
rect 503621 274619 503687 274622
rect 509325 274619 509391 274622
rect 490465 274546 490531 274549
rect 497181 274546 497247 274549
rect 490465 274544 497247 274546
rect 490465 274488 490470 274544
rect 490526 274488 497186 274544
rect 497242 274488 497247 274544
rect 490465 274486 497247 274488
rect 490465 274483 490531 274486
rect 497181 274483 497247 274486
rect 460933 274410 460999 274413
rect 470409 274410 470475 274413
rect 460933 274408 470475 274410
rect 460933 274352 460938 274408
rect 460994 274352 470414 274408
rect 470470 274352 470475 274408
rect 460933 274350 470475 274352
rect 460933 274347 460999 274350
rect 470409 274347 470475 274350
rect 475837 274410 475903 274413
rect 479793 274410 479859 274413
rect 475837 274408 479859 274410
rect 475837 274352 475842 274408
rect 475898 274352 479798 274408
rect 479854 274352 479859 274408
rect 475837 274350 479859 274352
rect 475837 274347 475903 274350
rect 479793 274347 479859 274350
rect 482553 274410 482619 274413
rect 489729 274410 489795 274413
rect 482553 274408 489795 274410
rect 482553 274352 482558 274408
rect 482614 274352 489734 274408
rect 489790 274352 489795 274408
rect 482553 274350 489795 274352
rect 482553 274347 482619 274350
rect 489729 274347 489795 274350
rect 434345 274138 434411 274141
rect 543457 274138 543523 274141
rect 434345 274136 543523 274138
rect 434345 274080 434350 274136
rect 434406 274080 543462 274136
rect 543518 274080 543523 274136
rect 434345 274078 543523 274080
rect 434345 274075 434411 274078
rect 543457 274075 543523 274078
rect 454861 273866 454927 273869
rect 461025 273866 461091 273869
rect 454861 273864 461091 273866
rect 454861 273808 454866 273864
rect 454922 273808 461030 273864
rect 461086 273808 461091 273864
rect 454861 273806 461091 273808
rect 454861 273803 454927 273806
rect 461025 273803 461091 273806
rect 489453 273866 489519 273869
rect 632145 273866 632211 273869
rect 489453 273864 632211 273866
rect 489453 273808 489458 273864
rect 489514 273808 632150 273864
rect 632206 273808 632211 273864
rect 489453 273806 632211 273808
rect 489453 273803 489519 273806
rect 632145 273803 632211 273806
rect 665173 273730 665239 273733
rect 665725 273732 665791 273733
rect 665398 273730 665404 273732
rect 665173 273728 665404 273730
rect 665173 273672 665178 273728
rect 665234 273672 665404 273728
rect 665173 273670 665404 273672
rect 665173 273667 665239 273670
rect 665398 273668 665404 273670
rect 665468 273668 665474 273732
rect 665725 273730 665772 273732
rect 665680 273728 665772 273730
rect 665680 273672 665730 273728
rect 665680 273670 665772 273672
rect 665725 273668 665772 273670
rect 665836 273668 665842 273732
rect 665725 273667 665791 273668
rect 426249 273594 426315 273597
rect 432045 273594 432111 273597
rect 426249 273592 432111 273594
rect 426249 273536 426254 273592
rect 426310 273536 432050 273592
rect 432106 273536 432111 273592
rect 426249 273534 432111 273536
rect 426249 273531 426315 273534
rect 432045 273531 432111 273534
rect 489729 273594 489795 273597
rect 490097 273594 490163 273597
rect 489729 273592 490163 273594
rect 489729 273536 489734 273592
rect 489790 273536 490102 273592
rect 490158 273536 490163 273592
rect 489729 273534 490163 273536
rect 489729 273531 489795 273534
rect 490097 273531 490163 273534
rect 497641 273594 497707 273597
rect 505277 273594 505343 273597
rect 497641 273592 505343 273594
rect 497641 273536 497646 273592
rect 497702 273536 505282 273592
rect 505338 273536 505343 273592
rect 497641 273534 505343 273536
rect 497641 273531 497707 273534
rect 505277 273531 505343 273534
rect 665541 273460 665607 273461
rect 665541 273458 665588 273460
rect 665496 273456 665588 273458
rect 665496 273400 665546 273456
rect 665496 273398 665588 273400
rect 665541 273396 665588 273398
rect 665652 273396 665658 273460
rect 665541 273395 665607 273396
rect 449709 273186 449775 273189
rect 450997 273186 451063 273189
rect 449709 273184 451063 273186
rect 449709 273128 449714 273184
rect 449770 273128 451002 273184
rect 451058 273128 451063 273184
rect 449709 273126 451063 273128
rect 449709 273123 449775 273126
rect 450997 273123 451063 273126
rect 40534 272988 40540 273052
rect 40604 273050 40610 273052
rect 41781 273050 41847 273053
rect 40604 273048 41847 273050
rect 40604 272992 41786 273048
rect 41842 272992 41847 273048
rect 40604 272990 41847 272992
rect 40604 272988 40610 272990
rect 41781 272987 41847 272990
rect 487797 273050 487863 273053
rect 490649 273050 490715 273053
rect 487797 273048 490715 273050
rect 487797 272992 487802 273048
rect 487858 272992 490654 273048
rect 490710 272992 490715 273048
rect 487797 272990 490715 272992
rect 487797 272987 487863 272990
rect 490649 272987 490715 272990
rect 491201 273050 491267 273053
rect 491201 273048 499590 273050
rect 491201 272992 491206 273048
rect 491262 272992 499590 273048
rect 491201 272990 499590 272992
rect 491201 272987 491267 272990
rect 436921 272914 436987 272917
rect 437933 272914 437999 272917
rect 436921 272912 437999 272914
rect 436921 272856 436926 272912
rect 436982 272856 437938 272912
rect 437994 272856 437999 272912
rect 436921 272854 437999 272856
rect 436921 272851 436987 272854
rect 437933 272851 437999 272854
rect 450537 272914 450603 272917
rect 452101 272914 452167 272917
rect 450537 272912 452167 272914
rect 450537 272856 450542 272912
rect 450598 272856 452106 272912
rect 452162 272856 452167 272912
rect 450537 272854 452167 272856
rect 450537 272851 450603 272854
rect 452101 272851 452167 272854
rect 453757 272914 453823 272917
rect 454677 272914 454743 272917
rect 453757 272912 454743 272914
rect 453757 272856 453762 272912
rect 453818 272856 454682 272912
rect 454738 272856 454743 272912
rect 453757 272854 454743 272856
rect 453757 272851 453823 272854
rect 454677 272851 454743 272854
rect 466269 272778 466335 272781
rect 476021 272778 476087 272781
rect 466269 272776 476087 272778
rect 466269 272720 466274 272776
rect 466330 272720 476026 272776
rect 476082 272720 476087 272776
rect 466269 272718 476087 272720
rect 466269 272715 466335 272718
rect 476021 272715 476087 272718
rect 480069 272778 480135 272781
rect 480989 272778 481055 272781
rect 480069 272776 481055 272778
rect 480069 272720 480074 272776
rect 480130 272720 480994 272776
rect 481050 272720 481055 272776
rect 480069 272718 481055 272720
rect 480069 272715 480135 272718
rect 480989 272715 481055 272718
rect 487613 272778 487679 272781
rect 499205 272778 499271 272781
rect 487613 272776 499271 272778
rect 487613 272720 487618 272776
rect 487674 272720 499210 272776
rect 499266 272720 499271 272776
rect 487613 272718 499271 272720
rect 499530 272778 499590 272990
rect 514109 272778 514175 272781
rect 499530 272776 514175 272778
rect 499530 272720 514114 272776
rect 514170 272720 514175 272776
rect 499530 272718 514175 272720
rect 487613 272715 487679 272718
rect 499205 272715 499271 272718
rect 514109 272715 514175 272718
rect 431861 272506 431927 272509
rect 437565 272506 437631 272509
rect 431861 272504 437631 272506
rect 431861 272448 431866 272504
rect 431922 272448 437570 272504
rect 437626 272448 437631 272504
rect 431861 272446 437631 272448
rect 431861 272443 431927 272446
rect 437565 272443 437631 272446
rect 452101 272506 452167 272509
rect 454401 272506 454467 272509
rect 452101 272504 454467 272506
rect 452101 272448 452106 272504
rect 452162 272448 454406 272504
rect 454462 272448 454467 272504
rect 452101 272446 454467 272448
rect 452101 272443 452167 272446
rect 454401 272443 454467 272446
rect 460841 272506 460907 272509
rect 461761 272506 461827 272509
rect 460841 272504 461827 272506
rect 460841 272448 460846 272504
rect 460902 272448 461766 272504
rect 461822 272448 461827 272504
rect 460841 272446 461827 272448
rect 460841 272443 460907 272446
rect 461761 272443 461827 272446
rect 464889 272506 464955 272509
rect 593137 272506 593203 272509
rect 464889 272504 593203 272506
rect 464889 272448 464894 272504
rect 464950 272448 593142 272504
rect 593198 272448 593203 272504
rect 464889 272446 593203 272448
rect 464889 272443 464955 272446
rect 593137 272443 593203 272446
rect 41781 272372 41847 272373
rect 41781 272368 41828 272372
rect 41892 272370 41898 272372
rect 424501 272370 424567 272373
rect 427261 272370 427327 272373
rect 41781 272312 41786 272368
rect 41781 272308 41828 272312
rect 41892 272310 41938 272370
rect 424501 272368 427327 272370
rect 424501 272312 424506 272368
rect 424562 272312 427266 272368
rect 427322 272312 427327 272368
rect 424501 272310 427327 272312
rect 41892 272308 41898 272310
rect 41781 272307 41847 272308
rect 424501 272307 424567 272310
rect 427261 272307 427327 272310
rect 429285 272234 429351 272237
rect 437105 272234 437171 272237
rect 429285 272232 437171 272234
rect 429285 272176 429290 272232
rect 429346 272176 437110 272232
rect 437166 272176 437171 272232
rect 429285 272174 437171 272176
rect 429285 272171 429351 272174
rect 437105 272171 437171 272174
rect 437381 272234 437447 272237
rect 442441 272234 442507 272237
rect 437381 272232 442507 272234
rect 437381 272176 437386 272232
rect 437442 272176 442446 272232
rect 442502 272176 442507 272232
rect 437381 272174 442507 272176
rect 437381 272171 437447 272174
rect 442441 272171 442507 272174
rect 445385 272234 445451 272237
rect 447869 272234 447935 272237
rect 445385 272232 447935 272234
rect 445385 272176 445390 272232
rect 445446 272176 447874 272232
rect 447930 272176 447935 272232
rect 445385 272174 447935 272176
rect 445385 272171 445451 272174
rect 447869 272171 447935 272174
rect 458633 272234 458699 272237
rect 466269 272234 466335 272237
rect 458633 272232 466335 272234
rect 458633 272176 458638 272232
rect 458694 272176 466274 272232
rect 466330 272176 466335 272232
rect 458633 272174 466335 272176
rect 458633 272171 458699 272174
rect 466269 272171 466335 272174
rect 475653 272234 475719 272237
rect 480069 272234 480135 272237
rect 475653 272232 480135 272234
rect 475653 272176 475658 272232
rect 475714 272176 480074 272232
rect 480130 272176 480135 272232
rect 475653 272174 480135 272176
rect 475653 272171 475719 272174
rect 480069 272171 480135 272174
rect 480989 272234 481055 272237
rect 490005 272234 490071 272237
rect 480989 272232 490071 272234
rect 480989 272176 480994 272232
rect 481050 272176 490010 272232
rect 490066 272176 490071 272232
rect 480989 272174 490071 272176
rect 480989 272171 481055 272174
rect 490005 272171 490071 272174
rect 498837 272234 498903 272237
rect 499849 272234 499915 272237
rect 507853 272234 507919 272237
rect 498837 272232 499682 272234
rect 498837 272176 498842 272232
rect 498898 272176 499682 272232
rect 498837 272174 499682 272176
rect 498837 272171 498903 272174
rect 441521 271962 441587 271965
rect 444189 271962 444255 271965
rect 441521 271960 444255 271962
rect 441521 271904 441526 271960
rect 441582 271904 444194 271960
rect 444250 271904 444255 271960
rect 441521 271902 444255 271904
rect 441521 271899 441587 271902
rect 444189 271899 444255 271902
rect 448329 271962 448395 271965
rect 451089 271962 451155 271965
rect 448329 271960 451155 271962
rect 448329 271904 448334 271960
rect 448390 271904 451094 271960
rect 451150 271904 451155 271960
rect 448329 271902 451155 271904
rect 448329 271899 448395 271902
rect 451089 271899 451155 271902
rect 487613 271962 487679 271965
rect 489637 271962 489703 271965
rect 487613 271960 489703 271962
rect 487613 271904 487618 271960
rect 487674 271904 489642 271960
rect 489698 271904 489703 271960
rect 487613 271902 489703 271904
rect 499622 271962 499682 272174
rect 499849 272232 507919 272234
rect 499849 272176 499854 272232
rect 499910 272176 507858 272232
rect 507914 272176 507919 272232
rect 499849 272174 507919 272176
rect 499849 272171 499915 272174
rect 507853 272171 507919 272174
rect 500217 271962 500283 271965
rect 499622 271960 500283 271962
rect 499622 271904 500222 271960
rect 500278 271904 500283 271960
rect 499622 271902 500283 271904
rect 487613 271899 487679 271902
rect 489637 271899 489703 271902
rect 500217 271899 500283 271902
rect 490005 271826 490071 271829
rect 499389 271826 499455 271829
rect 490005 271824 499455 271826
rect 490005 271768 490010 271824
rect 490066 271768 499394 271824
rect 499450 271768 499455 271824
rect 490005 271766 499455 271768
rect 490005 271763 490071 271766
rect 499389 271763 499455 271766
rect 409689 271690 409755 271693
rect 489862 271690 489868 271692
rect 409689 271688 489868 271690
rect 409689 271632 409694 271688
rect 409750 271632 489868 271688
rect 409689 271630 489868 271632
rect 409689 271627 409755 271630
rect 489862 271628 489868 271630
rect 489932 271628 489938 271692
rect 499757 271690 499823 271693
rect 509417 271690 509483 271693
rect 499757 271688 509483 271690
rect 499757 271632 499762 271688
rect 499818 271632 509422 271688
rect 509478 271632 509483 271688
rect 499757 271630 509483 271632
rect 499757 271627 499823 271630
rect 509417 271627 509483 271630
rect 391749 271554 391815 271557
rect 402605 271554 402671 271557
rect 391749 271552 402671 271554
rect 391749 271496 391754 271552
rect 391810 271496 402610 271552
rect 402666 271496 402671 271552
rect 391749 271494 402671 271496
rect 391749 271491 391815 271494
rect 402605 271491 402671 271494
rect 432965 271418 433031 271421
rect 446029 271418 446095 271421
rect 432965 271416 446095 271418
rect 432965 271360 432970 271416
rect 433026 271360 446034 271416
rect 446090 271360 446095 271416
rect 432965 271358 446095 271360
rect 432965 271355 433031 271358
rect 446029 271355 446095 271358
rect 446305 271418 446371 271421
rect 451365 271418 451431 271421
rect 446305 271416 451431 271418
rect 446305 271360 446310 271416
rect 446366 271360 451370 271416
rect 451426 271360 451431 271416
rect 446305 271358 451431 271360
rect 446305 271355 446371 271358
rect 451365 271355 451431 271358
rect 451549 271418 451615 271421
rect 456885 271418 456951 271421
rect 451549 271416 456951 271418
rect 451549 271360 451554 271416
rect 451610 271360 456890 271416
rect 456946 271360 456951 271416
rect 451549 271358 456951 271360
rect 451549 271355 451615 271358
rect 456885 271355 456951 271358
rect 466453 271418 466519 271421
rect 480529 271418 480595 271421
rect 466453 271416 480595 271418
rect 466453 271360 466458 271416
rect 466514 271360 480534 271416
rect 480590 271360 480595 271416
rect 466453 271358 480595 271360
rect 466453 271355 466519 271358
rect 480529 271355 480595 271358
rect 489269 271418 489335 271421
rect 490097 271418 490163 271421
rect 626165 271418 626231 271421
rect 489269 271416 490163 271418
rect 489269 271360 489274 271416
rect 489330 271360 490102 271416
rect 490158 271360 490163 271416
rect 489269 271358 490163 271360
rect 489269 271355 489335 271358
rect 490097 271355 490163 271358
rect 494654 271416 626231 271418
rect 494654 271360 626170 271416
rect 626226 271360 626231 271416
rect 494654 271358 626231 271360
rect 462497 271282 462563 271285
rect 465349 271282 465415 271285
rect 462497 271280 465415 271282
rect 462497 271224 462502 271280
rect 462558 271224 465354 271280
rect 465410 271224 465415 271280
rect 462497 271222 465415 271224
rect 462497 271219 462563 271222
rect 465349 271219 465415 271222
rect 412909 271146 412975 271149
rect 413921 271146 413987 271149
rect 412909 271144 413987 271146
rect 412909 271088 412914 271144
rect 412970 271088 413926 271144
rect 413982 271088 413987 271144
rect 412909 271086 413987 271088
rect 412909 271083 412975 271086
rect 413921 271083 413987 271086
rect 431493 271146 431559 271149
rect 433609 271146 433675 271149
rect 431493 271144 433675 271146
rect 431493 271088 431498 271144
rect 431554 271088 433614 271144
rect 433670 271088 433675 271144
rect 431493 271086 433675 271088
rect 431493 271083 431559 271086
rect 433609 271083 433675 271086
rect 456747 271146 456813 271149
rect 461761 271146 461827 271149
rect 456747 271144 461827 271146
rect 456747 271088 456752 271144
rect 456808 271088 461766 271144
rect 461822 271088 461827 271144
rect 456747 271086 461827 271088
rect 456747 271083 456813 271086
rect 461761 271083 461827 271086
rect 465993 271146 466059 271149
rect 466545 271146 466611 271149
rect 465993 271144 466611 271146
rect 465993 271088 465998 271144
rect 466054 271088 466550 271144
rect 466606 271088 466611 271144
rect 465993 271086 466611 271088
rect 465993 271083 466059 271086
rect 466545 271083 466611 271086
rect 480437 271146 480503 271149
rect 489637 271146 489703 271149
rect 480437 271144 489703 271146
rect 480437 271088 480442 271144
rect 480498 271088 489642 271144
rect 489698 271088 489703 271144
rect 480437 271086 489703 271088
rect 480437 271083 480503 271086
rect 489637 271083 489703 271086
rect 490281 271146 490347 271149
rect 493041 271146 493107 271149
rect 490281 271144 493107 271146
rect 490281 271088 490286 271144
rect 490342 271088 493046 271144
rect 493102 271088 493107 271144
rect 490281 271086 493107 271088
rect 490281 271083 490347 271086
rect 493041 271083 493107 271086
rect 402973 271010 403039 271013
rect 411253 271010 411319 271013
rect 402973 271008 411319 271010
rect 402973 270952 402978 271008
rect 403034 270952 411258 271008
rect 411314 270952 411319 271008
rect 402973 270950 411319 270952
rect 402973 270947 403039 270950
rect 411253 270947 411319 270950
rect 417693 270874 417759 270877
rect 418153 270874 418219 270877
rect 417693 270872 418219 270874
rect 417693 270816 417698 270872
rect 417754 270816 418158 270872
rect 418214 270816 418219 270872
rect 417693 270814 418219 270816
rect 417693 270811 417759 270814
rect 418153 270811 418219 270814
rect 485589 270874 485655 270877
rect 494654 270874 494714 271358
rect 626165 271355 626231 271358
rect 496721 271146 496787 271149
rect 642725 271146 642791 271149
rect 496721 271144 642791 271146
rect 496721 271088 496726 271144
rect 496782 271088 642730 271144
rect 642786 271088 642791 271144
rect 496721 271086 642791 271088
rect 496721 271083 496787 271086
rect 642725 271083 642791 271086
rect 504541 270874 504607 270877
rect 485589 270872 494714 270874
rect 485589 270816 485594 270872
rect 485650 270816 494714 270872
rect 485589 270814 494714 270816
rect 494838 270872 504607 270874
rect 494838 270816 504546 270872
rect 504602 270816 504607 270872
rect 494838 270814 504607 270816
rect 485589 270811 485655 270814
rect 429101 270738 429167 270741
rect 436277 270738 436343 270741
rect 429101 270736 436343 270738
rect 429101 270680 429106 270736
rect 429162 270680 436282 270736
rect 436338 270680 436343 270736
rect 429101 270678 436343 270680
rect 429101 270675 429167 270678
rect 436277 270675 436343 270678
rect 402789 270602 402855 270605
rect 403065 270602 403131 270605
rect 402789 270600 403131 270602
rect 402789 270544 402794 270600
rect 402850 270544 403070 270600
rect 403126 270544 403131 270600
rect 402789 270542 403131 270544
rect 402789 270539 402855 270542
rect 403065 270539 403131 270542
rect 404169 270602 404235 270605
rect 405917 270602 405983 270605
rect 404169 270600 405983 270602
rect 404169 270544 404174 270600
rect 404230 270544 405922 270600
rect 405978 270544 405983 270600
rect 404169 270542 405983 270544
rect 404169 270539 404235 270542
rect 405917 270539 405983 270542
rect 472249 270602 472315 270605
rect 485773 270602 485839 270605
rect 472249 270600 485839 270602
rect 472249 270544 472254 270600
rect 472310 270544 485778 270600
rect 485834 270544 485839 270600
rect 472249 270542 485839 270544
rect 472249 270539 472315 270542
rect 485773 270539 485839 270542
rect 490046 270540 490052 270604
rect 490116 270602 490122 270604
rect 494838 270602 494898 270814
rect 504541 270811 504607 270814
rect 509233 270738 509299 270741
rect 518341 270738 518407 270741
rect 509233 270736 518407 270738
rect 509233 270680 509238 270736
rect 509294 270680 518346 270736
rect 518402 270680 518407 270736
rect 509233 270678 518407 270680
rect 509233 270675 509299 270678
rect 518341 270675 518407 270678
rect 490116 270542 494898 270602
rect 495065 270602 495131 270605
rect 499665 270602 499731 270605
rect 495065 270600 499731 270602
rect 495065 270544 495070 270600
rect 495126 270544 499670 270600
rect 499726 270544 499731 270600
rect 495065 270542 499731 270544
rect 490116 270540 490122 270542
rect 495065 270539 495131 270542
rect 499665 270539 499731 270542
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 379145 270330 379211 270333
rect 379513 270330 379579 270333
rect 379145 270328 379579 270330
rect 379145 270272 379150 270328
rect 379206 270272 379518 270328
rect 379574 270272 379579 270328
rect 379145 270270 379579 270272
rect 379145 270267 379211 270270
rect 379513 270267 379579 270270
rect 380525 270330 380591 270333
rect 383561 270330 383627 270333
rect 380525 270328 383627 270330
rect 380525 270272 380530 270328
rect 380586 270272 383566 270328
rect 383622 270272 383627 270328
rect 380525 270270 383627 270272
rect 380525 270267 380591 270270
rect 383561 270267 383627 270270
rect 443545 270330 443611 270333
rect 557901 270330 557967 270333
rect 443545 270328 557967 270330
rect 443545 270272 443550 270328
rect 443606 270272 557906 270328
rect 557962 270272 557967 270328
rect 443545 270270 557967 270272
rect 443545 270267 443611 270270
rect 557901 270267 557967 270270
rect 369117 270194 369183 270197
rect 376937 270194 377003 270197
rect 369117 270192 377003 270194
rect 369117 270136 369122 270192
rect 369178 270136 376942 270192
rect 376998 270136 377003 270192
rect 369117 270134 377003 270136
rect 369117 270131 369183 270134
rect 376937 270131 377003 270134
rect 406745 270194 406811 270197
rect 408769 270194 408835 270197
rect 406745 270192 408835 270194
rect 406745 270136 406750 270192
rect 406806 270136 408774 270192
rect 408830 270136 408835 270192
rect 406745 270134 408835 270136
rect 406745 270131 406811 270134
rect 408769 270131 408835 270134
rect 377121 270058 377187 270061
rect 379329 270058 379395 270061
rect 377121 270056 379395 270058
rect 377121 270000 377126 270056
rect 377182 270000 379334 270056
rect 379390 270000 379395 270056
rect 377121 269998 379395 270000
rect 377121 269995 377187 269998
rect 379329 269995 379395 269998
rect 383653 270058 383719 270061
rect 386965 270058 387031 270061
rect 383653 270056 387031 270058
rect 383653 270000 383658 270056
rect 383714 270000 386970 270056
rect 387026 270000 387031 270056
rect 383653 269998 387031 270000
rect 383653 269995 383719 269998
rect 386965 269995 387031 269998
rect 438669 270058 438735 270061
rect 445109 270058 445175 270061
rect 438669 270056 445175 270058
rect 438669 270000 438674 270056
rect 438730 270000 445114 270056
rect 445170 270000 445175 270056
rect 438669 269998 445175 270000
rect 438669 269995 438735 269998
rect 445109 269995 445175 269998
rect 459369 270058 459435 270061
rect 461761 270058 461827 270061
rect 459369 270056 461827 270058
rect 459369 270000 459374 270056
rect 459430 270000 461766 270056
rect 461822 270000 461827 270056
rect 459369 269998 461827 270000
rect 459369 269995 459435 269998
rect 461761 269995 461827 269998
rect 470501 270058 470567 270061
rect 474917 270058 474983 270061
rect 470501 270056 474983 270058
rect 470501 270000 470506 270056
rect 470562 270000 474922 270056
rect 474978 270000 474983 270056
rect 470501 269998 474983 270000
rect 470501 269995 470567 269998
rect 474917 269995 474983 269998
rect 480069 270058 480135 270061
rect 483013 270058 483079 270061
rect 480069 270056 483079 270058
rect 480069 270000 480074 270056
rect 480130 270000 483018 270056
rect 483074 270000 483079 270056
rect 480069 269998 483079 270000
rect 480069 269995 480135 269998
rect 483013 269995 483079 269998
rect 493685 270058 493751 270061
rect 499389 270058 499455 270061
rect 500033 270058 500099 270061
rect 637573 270058 637639 270061
rect 493685 270056 499130 270058
rect 493685 270000 493690 270056
rect 493746 270000 499130 270056
rect 493685 269998 499130 270000
rect 493685 269995 493751 269998
rect 488165 269922 488231 269925
rect 489729 269922 489795 269925
rect 488165 269920 489795 269922
rect 488165 269864 488170 269920
rect 488226 269864 489734 269920
rect 489790 269864 489795 269920
rect 488165 269862 489795 269864
rect 499070 269922 499130 269998
rect 499389 270056 500099 270058
rect 499389 270000 499394 270056
rect 499450 270000 500038 270056
rect 500094 270000 500099 270056
rect 499389 269998 500099 270000
rect 499389 269995 499455 269998
rect 500033 269995 500099 269998
rect 504406 270056 637639 270058
rect 504406 270000 637578 270056
rect 637634 270000 637639 270056
rect 504406 269998 637639 270000
rect 499070 269862 499314 269922
rect 488165 269859 488231 269862
rect 489729 269859 489795 269862
rect 400121 269786 400187 269789
rect 487981 269786 488047 269789
rect 400121 269784 488047 269786
rect 400121 269728 400126 269784
rect 400182 269728 487986 269784
rect 488042 269728 488047 269784
rect 400121 269726 488047 269728
rect 499254 269786 499314 269862
rect 504406 269786 504466 269998
rect 637573 269995 637639 269998
rect 640701 269786 640767 269789
rect 499254 269726 504466 269786
rect 509190 269784 640767 269786
rect 509190 269728 640706 269784
rect 640762 269728 640767 269784
rect 509190 269726 640767 269728
rect 400121 269723 400187 269726
rect 487981 269723 488047 269726
rect 383377 269650 383443 269653
rect 383745 269650 383811 269653
rect 383377 269648 383811 269650
rect 383377 269592 383382 269648
rect 383438 269592 383750 269648
rect 383806 269592 383811 269648
rect 383377 269590 383811 269592
rect 383377 269587 383443 269590
rect 383745 269587 383811 269590
rect 397913 269650 397979 269653
rect 398925 269650 398991 269653
rect 397913 269648 398991 269650
rect 397913 269592 397918 269648
rect 397974 269592 398930 269648
rect 398986 269592 398991 269648
rect 397913 269590 398991 269592
rect 397913 269587 397979 269590
rect 398925 269587 398991 269590
rect 373717 269514 373783 269517
rect 375189 269514 375255 269517
rect 373717 269512 375255 269514
rect 373717 269456 373722 269512
rect 373778 269456 375194 269512
rect 375250 269456 375255 269512
rect 373717 269454 375255 269456
rect 373717 269451 373783 269454
rect 375189 269451 375255 269454
rect 384113 269514 384179 269517
rect 388989 269514 389055 269517
rect 384113 269512 389055 269514
rect 384113 269456 384118 269512
rect 384174 269456 388994 269512
rect 389050 269456 389055 269512
rect 384113 269454 389055 269456
rect 384113 269451 384179 269454
rect 388989 269451 389055 269454
rect 415853 269514 415919 269517
rect 503621 269514 503687 269517
rect 509190 269514 509250 269726
rect 640701 269723 640767 269726
rect 415853 269512 503687 269514
rect 415853 269456 415858 269512
rect 415914 269456 503626 269512
rect 503682 269456 503687 269512
rect 415853 269454 503687 269456
rect 415853 269451 415919 269454
rect 503621 269451 503687 269454
rect 504406 269454 509250 269514
rect 393681 269378 393747 269381
rect 401593 269378 401659 269381
rect 393681 269376 401659 269378
rect 393681 269320 393686 269376
rect 393742 269320 401598 269376
rect 401654 269320 401659 269376
rect 393681 269318 401659 269320
rect 393681 269315 393747 269318
rect 401593 269315 401659 269318
rect 429929 269242 429995 269245
rect 432781 269242 432847 269245
rect 429929 269240 432847 269242
rect 429929 269184 429934 269240
rect 429990 269184 432786 269240
rect 432842 269184 432847 269240
rect 429929 269182 432847 269184
rect 429929 269179 429995 269182
rect 432781 269179 432847 269182
rect 455137 269242 455203 269245
rect 456793 269242 456859 269245
rect 455137 269240 456859 269242
rect 455137 269184 455142 269240
rect 455198 269184 456798 269240
rect 456854 269184 456859 269240
rect 455137 269182 456859 269184
rect 455137 269179 455203 269182
rect 456793 269179 456859 269182
rect 476021 269242 476087 269245
rect 477493 269242 477559 269245
rect 476021 269240 477559 269242
rect 476021 269184 476026 269240
rect 476082 269184 477498 269240
rect 477554 269184 477559 269240
rect 476021 269182 477559 269184
rect 476021 269179 476087 269182
rect 477493 269179 477559 269182
rect 489729 269242 489795 269245
rect 499205 269242 499271 269245
rect 489729 269240 499271 269242
rect 489729 269184 489734 269240
rect 489790 269184 499210 269240
rect 499266 269184 499271 269240
rect 489729 269182 499271 269184
rect 489729 269179 489795 269182
rect 499205 269179 499271 269182
rect 499757 269242 499823 269245
rect 504406 269242 504466 269454
rect 499757 269240 504466 269242
rect 499757 269184 499762 269240
rect 499818 269184 504466 269240
rect 499757 269182 504466 269184
rect 509049 269242 509115 269245
rect 510613 269242 510679 269245
rect 509049 269240 510679 269242
rect 509049 269184 509054 269240
rect 509110 269184 510618 269240
rect 510674 269184 510679 269240
rect 509049 269182 510679 269184
rect 499757 269179 499823 269182
rect 509049 269179 509115 269182
rect 510613 269179 510679 269182
rect 408493 269106 408559 269109
rect 416773 269106 416839 269109
rect 408493 269104 416839 269106
rect 408493 269048 408498 269104
rect 408554 269048 416778 269104
rect 416834 269048 416839 269104
rect 408493 269046 416839 269048
rect 408493 269043 408559 269046
rect 416773 269043 416839 269046
rect 437013 269106 437079 269109
rect 438853 269106 438919 269109
rect 437013 269104 438919 269106
rect 437013 269048 437018 269104
rect 437074 269048 438858 269104
rect 438914 269048 438919 269104
rect 437013 269046 438919 269048
rect 437013 269043 437079 269046
rect 438853 269043 438919 269046
rect 441337 268970 441403 268973
rect 443177 268970 443243 268973
rect 441337 268968 443243 268970
rect 441337 268912 441342 268968
rect 441398 268912 443182 268968
rect 443238 268912 443243 268968
rect 441337 268910 443243 268912
rect 441337 268907 441403 268910
rect 443177 268907 443243 268910
rect 466453 268970 466519 268973
rect 468017 268970 468083 268973
rect 466453 268968 468083 268970
rect 466453 268912 466458 268968
rect 466514 268912 468022 268968
rect 468078 268912 468083 268968
rect 466453 268910 468083 268912
rect 466453 268907 466519 268910
rect 468017 268907 468083 268910
rect 480253 268970 480319 268973
rect 499205 268970 499271 268973
rect 480253 268968 499271 268970
rect 480253 268912 480258 268968
rect 480314 268912 499210 268968
rect 499266 268912 499271 268968
rect 480253 268910 499271 268912
rect 480253 268907 480319 268910
rect 499205 268907 499271 268910
rect 499389 268970 499455 268973
rect 501137 268970 501203 268973
rect 499389 268968 501203 268970
rect 499389 268912 499394 268968
rect 499450 268912 501142 268968
rect 501198 268912 501203 268968
rect 499389 268910 501203 268912
rect 499389 268907 499455 268910
rect 501137 268907 501203 268910
rect 461577 268698 461643 268701
rect 587893 268698 587959 268701
rect 461577 268696 587959 268698
rect 461577 268640 461582 268696
rect 461638 268640 587898 268696
rect 587954 268640 587959 268696
rect 461577 268638 587959 268640
rect 461577 268635 461643 268638
rect 587893 268635 587959 268638
rect 675293 268698 675359 268701
rect 675293 268696 676292 268698
rect 675293 268640 675298 268696
rect 675354 268640 676292 268696
rect 675293 268638 676292 268640
rect 675293 268635 675359 268638
rect 447041 268562 447107 268565
rect 448513 268562 448579 268565
rect 447041 268560 448579 268562
rect 447041 268504 447046 268560
rect 447102 268504 448518 268560
rect 448574 268504 448579 268560
rect 447041 268502 448579 268504
rect 447041 268499 447107 268502
rect 448513 268499 448579 268502
rect 460105 268426 460171 268429
rect 462313 268426 462379 268429
rect 460105 268424 462379 268426
rect 460105 268368 460110 268424
rect 460166 268368 462318 268424
rect 462374 268368 462379 268424
rect 460105 268366 462379 268368
rect 460105 268363 460171 268366
rect 462313 268363 462379 268366
rect 466361 268426 466427 268429
rect 466729 268426 466795 268429
rect 466361 268424 466795 268426
rect 466361 268368 466366 268424
rect 466422 268368 466734 268424
rect 466790 268368 466795 268424
rect 466361 268366 466795 268368
rect 466361 268363 466427 268366
rect 466729 268363 466795 268366
rect 475561 268426 475627 268429
rect 480345 268426 480411 268429
rect 607213 268426 607279 268429
rect 475561 268424 480411 268426
rect 475561 268368 475566 268424
rect 475622 268368 480350 268424
rect 480406 268368 480411 268424
rect 475561 268366 480411 268368
rect 475561 268363 475627 268366
rect 480345 268363 480411 268366
rect 489870 268424 607279 268426
rect 489870 268368 607218 268424
rect 607274 268368 607279 268424
rect 489870 268366 607279 268368
rect 425237 268290 425303 268293
rect 429285 268290 429351 268293
rect 425237 268288 429351 268290
rect 425237 268232 425242 268288
rect 425298 268232 429290 268288
rect 429346 268232 429351 268288
rect 425237 268230 429351 268232
rect 425237 268227 425303 268230
rect 429285 268227 429351 268230
rect 416681 268154 416747 268157
rect 418061 268154 418127 268157
rect 416681 268152 418127 268154
rect 416681 268096 416686 268152
rect 416742 268096 418066 268152
rect 418122 268096 418127 268152
rect 416681 268094 418127 268096
rect 416681 268091 416747 268094
rect 418061 268091 418127 268094
rect 457897 268154 457963 268157
rect 461945 268154 462011 268157
rect 457897 268152 462011 268154
rect 457897 268096 457902 268152
rect 457958 268096 461950 268152
rect 462006 268096 462011 268152
rect 457897 268094 462011 268096
rect 457897 268091 457963 268094
rect 461945 268091 462011 268094
rect 464705 268154 464771 268157
rect 469213 268154 469279 268157
rect 464705 268152 469279 268154
rect 464705 268096 464710 268152
rect 464766 268096 469218 268152
rect 469274 268096 469279 268152
rect 464705 268094 469279 268096
rect 464705 268091 464771 268094
rect 469213 268091 469279 268094
rect 473721 268154 473787 268157
rect 489870 268154 489930 268366
rect 607213 268363 607279 268366
rect 675477 268290 675543 268293
rect 675477 268288 676292 268290
rect 675477 268232 675482 268288
rect 675538 268232 676292 268288
rect 675477 268230 676292 268232
rect 675477 268227 675543 268230
rect 473721 268152 489930 268154
rect 473721 268096 473726 268152
rect 473782 268096 489930 268152
rect 473721 268094 489930 268096
rect 473721 268091 473787 268094
rect 424869 268018 424935 268021
rect 428457 268018 428523 268021
rect 424869 268016 428523 268018
rect 424869 267960 424874 268016
rect 424930 267960 428462 268016
rect 428518 267960 428523 268016
rect 424869 267958 428523 267960
rect 424869 267955 424935 267958
rect 428457 267955 428523 267958
rect 417693 267882 417759 267885
rect 422661 267882 422727 267885
rect 417693 267880 422727 267882
rect 417693 267824 417698 267880
rect 417754 267824 422666 267880
rect 422722 267824 422727 267880
rect 417693 267822 422727 267824
rect 417693 267819 417759 267822
rect 422661 267819 422727 267822
rect 494145 267882 494211 267885
rect 508865 267882 508931 267885
rect 494145 267880 508931 267882
rect 494145 267824 494150 267880
rect 494206 267824 508870 267880
rect 508926 267824 508931 267880
rect 494145 267822 508931 267824
rect 494145 267819 494211 267822
rect 508865 267819 508931 267822
rect 675477 267882 675543 267885
rect 675477 267880 676292 267882
rect 675477 267824 675482 267880
rect 675538 267824 676292 267880
rect 675477 267822 676292 267824
rect 675477 267819 675543 267822
rect 436001 267746 436067 267749
rect 437381 267746 437447 267749
rect 436001 267744 437447 267746
rect 436001 267688 436006 267744
rect 436062 267688 437386 267744
rect 437442 267688 437447 267744
rect 436001 267686 437447 267688
rect 436001 267683 436067 267686
rect 437381 267683 437447 267686
rect 468201 267746 468267 267749
rect 471421 267746 471487 267749
rect 468201 267744 471487 267746
rect 468201 267688 468206 267744
rect 468262 267688 471426 267744
rect 471482 267688 471487 267744
rect 468201 267686 471487 267688
rect 468201 267683 468267 267686
rect 471421 267683 471487 267686
rect 379329 267610 379395 267613
rect 381353 267610 381419 267613
rect 379329 267608 381419 267610
rect 379329 267552 379334 267608
rect 379390 267552 381358 267608
rect 381414 267552 381419 267608
rect 379329 267550 381419 267552
rect 379329 267547 379395 267550
rect 381353 267547 381419 267550
rect 392577 267610 392643 267613
rect 393405 267610 393471 267613
rect 392577 267608 393471 267610
rect 392577 267552 392582 267608
rect 392638 267552 393410 267608
rect 393466 267552 393471 267608
rect 392577 267550 393471 267552
rect 392577 267547 392643 267550
rect 393405 267547 393471 267550
rect 427353 267610 427419 267613
rect 427997 267610 428063 267613
rect 427353 267608 428063 267610
rect 427353 267552 427358 267608
rect 427414 267552 428002 267608
rect 428058 267552 428063 267608
rect 427353 267550 428063 267552
rect 427353 267547 427419 267550
rect 427997 267547 428063 267550
rect 466177 267610 466243 267613
rect 467005 267610 467071 267613
rect 466177 267608 467071 267610
rect 466177 267552 466182 267608
rect 466238 267552 467010 267608
rect 467066 267552 467071 267608
rect 466177 267550 467071 267552
rect 466177 267547 466243 267550
rect 467005 267547 467071 267550
rect 483105 267610 483171 267613
rect 489729 267610 489795 267613
rect 483105 267608 489795 267610
rect 483105 267552 483110 267608
rect 483166 267552 489734 267608
rect 489790 267552 489795 267608
rect 483105 267550 489795 267552
rect 483105 267547 483171 267550
rect 489729 267547 489795 267550
rect 490465 267610 490531 267613
rect 491385 267610 491451 267613
rect 490465 267608 491451 267610
rect 490465 267552 490470 267608
rect 490526 267552 491390 267608
rect 491446 267552 491451 267608
rect 490465 267550 491451 267552
rect 490465 267547 490531 267550
rect 491385 267547 491451 267550
rect 492121 267610 492187 267613
rect 578877 267610 578943 267613
rect 492121 267608 578943 267610
rect 492121 267552 492126 267608
rect 492182 267552 578882 267608
rect 578938 267552 578943 267608
rect 492121 267550 578943 267552
rect 492121 267547 492187 267550
rect 578877 267547 578943 267550
rect 675109 267474 675175 267477
rect 675109 267472 676292 267474
rect 675109 267416 675114 267472
rect 675170 267416 676292 267472
rect 675109 267414 676292 267416
rect 675109 267411 675175 267414
rect 366633 267338 366699 267341
rect 370497 267338 370563 267341
rect 366633 267336 370563 267338
rect 366633 267280 366638 267336
rect 366694 267280 370502 267336
rect 370558 267280 370563 267336
rect 366633 267278 370563 267280
rect 366633 267275 366699 267278
rect 370497 267275 370563 267278
rect 388161 267338 388227 267341
rect 390461 267338 390527 267341
rect 388161 267336 390527 267338
rect 388161 267280 388166 267336
rect 388222 267280 390466 267336
rect 390522 267280 390527 267336
rect 388161 267278 390527 267280
rect 388161 267275 388227 267278
rect 390461 267275 390527 267278
rect 428089 267338 428155 267341
rect 532969 267338 533035 267341
rect 428089 267336 533035 267338
rect 428089 267280 428094 267336
rect 428150 267280 532974 267336
rect 533030 267280 533035 267336
rect 428089 267278 533035 267280
rect 428089 267275 428155 267278
rect 532969 267275 533035 267278
rect 426893 267066 426959 267069
rect 432597 267066 432663 267069
rect 426893 267064 432663 267066
rect 426893 267008 426898 267064
rect 426954 267008 432602 267064
rect 432658 267008 432663 267064
rect 426893 267006 432663 267008
rect 426893 267003 426959 267006
rect 432597 267003 432663 267006
rect 450169 267066 450235 267069
rect 454861 267066 454927 267069
rect 466821 267066 466887 267069
rect 450169 267064 454927 267066
rect 450169 267008 450174 267064
rect 450230 267008 454866 267064
rect 454922 267008 454927 267064
rect 450169 267006 454927 267008
rect 450169 267003 450235 267006
rect 454861 267003 454927 267006
rect 466410 267064 466887 267066
rect 466410 267008 466826 267064
rect 466882 267008 466887 267064
rect 466410 267006 466887 267008
rect 412817 266930 412883 266933
rect 414657 266930 414723 266933
rect 412817 266928 414723 266930
rect 412817 266872 412822 266928
rect 412878 266872 414662 266928
rect 414718 266872 414723 266928
rect 412817 266870 414723 266872
rect 412817 266867 412883 266870
rect 414657 266867 414723 266870
rect 369301 266794 369367 266797
rect 371785 266794 371851 266797
rect 369301 266792 371851 266794
rect 369301 266736 369306 266792
rect 369362 266736 371790 266792
rect 371846 266736 371851 266792
rect 369301 266734 371851 266736
rect 369301 266731 369367 266734
rect 371785 266731 371851 266734
rect 437381 266794 437447 266797
rect 442441 266794 442507 266797
rect 437381 266792 442507 266794
rect 437381 266736 437386 266792
rect 437442 266736 442446 266792
rect 442502 266736 442507 266792
rect 437381 266734 442507 266736
rect 437381 266731 437447 266734
rect 442441 266731 442507 266734
rect 463601 266794 463667 266797
rect 466410 266794 466470 267006
rect 466821 267003 466887 267006
rect 470041 267066 470107 267069
rect 497457 267066 497523 267069
rect 470041 267064 497523 267066
rect 470041 267008 470046 267064
rect 470102 267008 497462 267064
rect 497518 267008 497523 267064
rect 470041 267006 497523 267008
rect 470041 267003 470107 267006
rect 497457 267003 497523 267006
rect 499021 267066 499087 267069
rect 636193 267066 636259 267069
rect 499021 267064 636259 267066
rect 499021 267008 499026 267064
rect 499082 267008 636198 267064
rect 636254 267008 636259 267064
rect 499021 267006 636259 267008
rect 499021 267003 499087 267006
rect 636193 267003 636259 267006
rect 675293 267066 675359 267069
rect 675293 267064 676292 267066
rect 675293 267008 675298 267064
rect 675354 267008 676292 267064
rect 675293 267006 676292 267008
rect 675293 267003 675359 267006
rect 473997 266794 474063 266797
rect 463601 266792 466470 266794
rect 463601 266736 463606 266792
rect 463662 266736 466470 266792
rect 463601 266734 466470 266736
rect 473310 266792 474063 266794
rect 473310 266736 474002 266792
rect 474058 266736 474063 266792
rect 473310 266734 474063 266736
rect 463601 266731 463667 266734
rect 420729 266658 420795 266661
rect 423857 266658 423923 266661
rect 420729 266656 423923 266658
rect 420729 266600 420734 266656
rect 420790 266600 423862 266656
rect 423918 266600 423923 266656
rect 420729 266598 423923 266600
rect 420729 266595 420795 266598
rect 423857 266595 423923 266598
rect 396257 266522 396323 266525
rect 398465 266522 398531 266525
rect 396257 266520 398531 266522
rect 396257 266464 396262 266520
rect 396318 266464 398470 266520
rect 398526 266464 398531 266520
rect 396257 266462 398531 266464
rect 396257 266459 396323 266462
rect 398465 266459 398531 266462
rect 466177 266522 466243 266525
rect 473310 266522 473370 266734
rect 473997 266731 474063 266734
rect 474641 266794 474707 266797
rect 479885 266794 479951 266797
rect 474641 266792 479951 266794
rect 474641 266736 474646 266792
rect 474702 266736 479890 266792
rect 479946 266736 479951 266792
rect 474641 266734 479951 266736
rect 474641 266731 474707 266734
rect 479885 266731 479951 266734
rect 488073 266794 488139 266797
rect 490189 266794 490255 266797
rect 488073 266792 490255 266794
rect 488073 266736 488078 266792
rect 488134 266736 490194 266792
rect 490250 266736 490255 266792
rect 488073 266734 490255 266736
rect 488073 266731 488139 266734
rect 490189 266731 490255 266734
rect 490465 266794 490531 266797
rect 494881 266794 494947 266797
rect 490465 266792 494947 266794
rect 490465 266736 490470 266792
rect 490526 266736 494886 266792
rect 494942 266736 494947 266792
rect 490465 266734 494947 266736
rect 490465 266731 490531 266734
rect 494881 266731 494947 266734
rect 496537 266794 496603 266797
rect 499205 266794 499271 266797
rect 496537 266792 499271 266794
rect 496537 266736 496542 266792
rect 496598 266736 499210 266792
rect 499266 266736 499271 266792
rect 496537 266734 499271 266736
rect 496537 266731 496603 266734
rect 499205 266731 499271 266734
rect 675477 266658 675543 266661
rect 675477 266656 676292 266658
rect 675477 266600 675482 266656
rect 675538 266600 676292 266656
rect 675477 266598 676292 266600
rect 675477 266595 675543 266598
rect 466177 266520 473370 266522
rect 466177 266464 466182 266520
rect 466238 266464 473370 266520
rect 466177 266462 473370 266464
rect 489729 266522 489795 266525
rect 494513 266522 494579 266525
rect 489729 266520 494579 266522
rect 489729 266464 489734 266520
rect 489790 266464 494518 266520
rect 494574 266464 494579 266520
rect 489729 266462 494579 266464
rect 466177 266459 466243 266462
rect 489729 266459 489795 266462
rect 494513 266459 494579 266462
rect 498009 266522 498075 266525
rect 499389 266522 499455 266525
rect 498009 266520 499455 266522
rect 498009 266464 498014 266520
rect 498070 266464 499394 266520
rect 499450 266464 499455 266520
rect 498009 266462 499455 266464
rect 498009 266459 498075 266462
rect 499389 266459 499455 266462
rect 410793 266386 410859 266389
rect 417417 266386 417483 266389
rect 410793 266384 417483 266386
rect 410793 266328 410798 266384
rect 410854 266328 417422 266384
rect 417478 266328 417483 266384
rect 410793 266326 417483 266328
rect 410793 266323 410859 266326
rect 417417 266323 417483 266326
rect 454953 266386 455019 266389
rect 456885 266386 456951 266389
rect 454953 266384 456951 266386
rect 454953 266328 454958 266384
rect 455014 266328 456890 266384
rect 456946 266328 456951 266384
rect 454953 266326 456951 266328
rect 454953 266323 455019 266326
rect 456885 266323 456951 266326
rect 457161 266386 457227 266389
rect 462497 266386 462563 266389
rect 457161 266384 462563 266386
rect 457161 266328 457166 266384
rect 457222 266328 462502 266384
rect 462558 266328 462563 266384
rect 457161 266326 462563 266328
rect 457161 266323 457227 266326
rect 462497 266323 462563 266326
rect 446857 266250 446923 266253
rect 449065 266250 449131 266253
rect 446857 266248 449131 266250
rect 446857 266192 446862 266248
rect 446918 266192 449070 266248
rect 449126 266192 449131 266248
rect 446857 266190 449131 266192
rect 446857 266187 446923 266190
rect 449065 266187 449131 266190
rect 675477 266250 675543 266253
rect 675477 266248 676292 266250
rect 675477 266192 675482 266248
rect 675538 266192 676292 266248
rect 675477 266190 676292 266192
rect 675477 266187 675543 266190
rect 461025 266114 461091 266117
rect 461761 266114 461827 266117
rect 589273 266114 589339 266117
rect 461025 266112 461827 266114
rect 461025 266056 461030 266112
rect 461086 266056 461766 266112
rect 461822 266056 461827 266112
rect 461025 266054 461827 266056
rect 461025 266051 461091 266054
rect 461761 266051 461827 266054
rect 466410 266112 589339 266114
rect 466410 266056 589278 266112
rect 589334 266056 589339 266112
rect 466410 266054 589339 266056
rect 462681 265842 462747 265845
rect 466410 265842 466470 266054
rect 589273 266051 589339 266054
rect 462681 265840 466470 265842
rect 462681 265784 462686 265840
rect 462742 265784 466470 265840
rect 462681 265782 466470 265784
rect 479609 265842 479675 265845
rect 614757 265842 614823 265845
rect 479609 265840 614823 265842
rect 479609 265784 479614 265840
rect 479670 265784 614762 265840
rect 614818 265784 614823 265840
rect 479609 265782 614823 265784
rect 462681 265779 462747 265782
rect 479609 265779 479675 265782
rect 614757 265779 614823 265782
rect 675293 265842 675359 265845
rect 675293 265840 676292 265842
rect 675293 265784 675298 265840
rect 675354 265784 676292 265840
rect 675293 265782 676292 265784
rect 675293 265779 675359 265782
rect 50705 265570 50771 265573
rect 658457 265570 658523 265573
rect 50705 265568 658523 265570
rect 50705 265512 50710 265568
rect 50766 265512 658462 265568
rect 658518 265512 658523 265568
rect 50705 265510 658523 265512
rect 50705 265507 50771 265510
rect 658457 265507 658523 265510
rect 675477 265434 675543 265437
rect 675477 265432 676292 265434
rect 675477 265376 675482 265432
rect 675538 265376 676292 265432
rect 675477 265374 676292 265376
rect 675477 265371 675543 265374
rect 465809 265298 465875 265301
rect 466913 265298 466979 265301
rect 465809 265296 466979 265298
rect 465809 265240 465814 265296
rect 465870 265240 466918 265296
rect 466974 265240 466979 265296
rect 465809 265238 466979 265240
rect 465809 265235 465875 265238
rect 466913 265235 466979 265238
rect 675477 265026 675543 265029
rect 675477 265024 676292 265026
rect 675477 264968 675482 265024
rect 675538 264968 676292 265024
rect 675477 264966 676292 264968
rect 675477 264963 675543 264966
rect 675477 264618 675543 264621
rect 675477 264616 676292 264618
rect 675477 264560 675482 264616
rect 675538 264560 676292 264616
rect 675477 264558 676292 264560
rect 675477 264555 675543 264558
rect 495433 264346 495499 264349
rect 499757 264346 499823 264349
rect 495433 264344 499823 264346
rect 495433 264288 495438 264344
rect 495494 264288 499762 264344
rect 499818 264288 499823 264344
rect 495433 264286 499823 264288
rect 495433 264283 495499 264286
rect 499757 264283 499823 264286
rect 675017 264210 675083 264213
rect 675017 264208 676292 264210
rect 675017 264152 675022 264208
rect 675078 264152 676292 264208
rect 675017 264150 676292 264152
rect 675017 264147 675083 264150
rect 676070 263604 676076 263668
rect 676140 263666 676146 263668
rect 676262 263666 676322 263772
rect 676140 263606 676322 263666
rect 676140 263604 676146 263606
rect 676262 263261 676322 263364
rect 676213 263256 676322 263261
rect 676213 263200 676218 263256
rect 676274 263200 676322 263256
rect 676213 263198 676322 263200
rect 676213 263195 676279 263198
rect 675477 262986 675543 262989
rect 675477 262984 676292 262986
rect 675477 262928 675482 262984
rect 675538 262928 676292 262984
rect 675477 262926 676292 262928
rect 675477 262923 675543 262926
rect 511533 262714 511599 262717
rect 508484 262712 511599 262714
rect 508484 262656 511538 262712
rect 511594 262656 511599 262712
rect 508484 262654 511599 262656
rect 511533 262651 511599 262654
rect 681046 262445 681106 262548
rect 680997 262440 681106 262445
rect 680997 262384 681002 262440
rect 681058 262384 681106 262440
rect 680997 262382 681106 262384
rect 680997 262379 681063 262382
rect 674465 262170 674531 262173
rect 674465 262168 676292 262170
rect 674465 262112 674470 262168
rect 674526 262112 676292 262168
rect 674465 262110 676292 262112
rect 674465 262107 674531 262110
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 675477 261354 675543 261357
rect 675477 261352 676292 261354
rect 675477 261296 675482 261352
rect 675538 261296 676292 261352
rect 675477 261294 676292 261296
rect 675477 261291 675543 261294
rect 676814 260812 676874 260916
rect 676806 260748 676812 260812
rect 676876 260748 676882 260812
rect 675661 260538 675727 260541
rect 675661 260536 676292 260538
rect 675661 260480 675666 260536
rect 675722 260480 676292 260536
rect 675661 260478 676292 260480
rect 675661 260475 675727 260478
rect 511349 260266 511415 260269
rect 508484 260264 511415 260266
rect 508484 260208 511354 260264
rect 511410 260208 511415 260264
rect 508484 260206 511415 260208
rect 511349 260203 511415 260206
rect 675477 260130 675543 260133
rect 675477 260128 676292 260130
rect 675477 260072 675482 260128
rect 675538 260072 676292 260128
rect 675477 260070 676292 260072
rect 675477 260067 675543 260070
rect 675293 259722 675359 259725
rect 675293 259720 676292 259722
rect 675293 259664 675298 259720
rect 675354 259664 676292 259720
rect 675293 259662 676292 259664
rect 675293 259659 675359 259662
rect 39941 259586 40007 259589
rect 46565 259586 46631 259589
rect 39941 259584 46631 259586
rect 39941 259528 39946 259584
rect 40002 259528 46570 259584
rect 46626 259528 46631 259584
rect 39941 259526 46631 259528
rect 39941 259523 40007 259526
rect 46565 259523 46631 259526
rect 675477 259314 675543 259317
rect 675477 259312 676292 259314
rect 675477 259256 675482 259312
rect 675538 259256 676292 259312
rect 675477 259254 676292 259256
rect 675477 259251 675543 259254
rect 674649 258906 674715 258909
rect 674649 258904 676292 258906
rect 674649 258848 674654 258904
rect 674710 258848 676292 258904
rect 674649 258846 676292 258848
rect 674649 258843 674715 258846
rect 675477 258498 675543 258501
rect 675477 258496 676292 258498
rect 675477 258440 675482 258496
rect 675538 258440 676292 258496
rect 675477 258438 676292 258440
rect 675477 258435 675543 258438
rect 35801 258090 35867 258093
rect 35788 258088 35867 258090
rect 35788 258032 35806 258088
rect 35862 258032 35867 258088
rect 35788 258030 35867 258032
rect 35801 258027 35867 258030
rect 511441 257818 511507 257821
rect 508484 257816 511507 257818
rect 508484 257760 511446 257816
rect 511502 257760 511507 257816
rect 508484 257758 511507 257760
rect 511441 257755 511507 257758
rect 35574 257549 35634 257652
rect 683070 257549 683130 258060
rect 35574 257544 35683 257549
rect 35574 257488 35622 257544
rect 35678 257488 35683 257544
rect 35574 257486 35683 257488
rect 35617 257483 35683 257486
rect 39573 257546 39639 257549
rect 43161 257546 43227 257549
rect 39573 257544 43227 257546
rect 39573 257488 39578 257544
rect 39634 257488 43166 257544
rect 43222 257488 43227 257544
rect 39573 257486 43227 257488
rect 683070 257544 683179 257549
rect 683070 257488 683118 257544
rect 683174 257488 683179 257544
rect 683070 257486 683179 257488
rect 39573 257483 39639 257486
rect 43161 257483 43227 257486
rect 683113 257483 683179 257486
rect 675477 257274 675543 257277
rect 675477 257272 676292 257274
rect 35390 257141 35450 257244
rect 675477 257216 675482 257272
rect 675538 257216 676292 257272
rect 675477 257214 676292 257216
rect 675477 257211 675543 257214
rect 35390 257136 35499 257141
rect 35801 257138 35867 257141
rect 35390 257080 35438 257136
rect 35494 257080 35499 257136
rect 35390 257078 35499 257080
rect 35433 257075 35499 257078
rect 35758 257136 35867 257138
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257075 35867 257080
rect 35758 256836 35818 257075
rect 35390 256325 35450 256428
rect 35390 256320 35499 256325
rect 35390 256264 35438 256320
rect 35494 256264 35499 256320
rect 35390 256262 35499 256264
rect 35433 256259 35499 256262
rect 35574 255917 35634 256020
rect 35574 255912 35683 255917
rect 35574 255856 35622 255912
rect 35678 255856 35683 255912
rect 35574 255854 35683 255856
rect 35617 255851 35683 255854
rect 35758 255509 35818 255612
rect 35758 255504 35867 255509
rect 35758 255448 35806 255504
rect 35862 255448 35867 255504
rect 35758 255446 35867 255448
rect 35801 255443 35867 255446
rect 511165 255370 511231 255373
rect 508484 255368 511231 255370
rect 508484 255312 511170 255368
rect 511226 255312 511231 255368
rect 508484 255310 511231 255312
rect 511165 255307 511231 255310
rect 35390 255101 35450 255204
rect 35390 255096 35499 255101
rect 35801 255098 35867 255101
rect 35390 255040 35438 255096
rect 35494 255040 35499 255096
rect 35390 255038 35499 255040
rect 35433 255035 35499 255038
rect 35758 255096 35867 255098
rect 35758 255040 35806 255096
rect 35862 255040 35867 255096
rect 35758 255035 35867 255040
rect 35758 254796 35818 255035
rect 35617 254690 35683 254693
rect 35574 254688 35683 254690
rect 35574 254632 35622 254688
rect 35678 254632 35683 254688
rect 35574 254627 35683 254632
rect 35574 254388 35634 254627
rect 35801 254282 35867 254285
rect 35758 254280 35867 254282
rect 35758 254224 35806 254280
rect 35862 254224 35867 254280
rect 35758 254219 35867 254224
rect 41229 254282 41295 254285
rect 44265 254282 44331 254285
rect 41229 254280 44331 254282
rect 41229 254224 41234 254280
rect 41290 254224 44270 254280
rect 44326 254224 44331 254280
rect 41229 254222 44331 254224
rect 41229 254219 41295 254222
rect 44265 254219 44331 254222
rect 35758 253980 35818 254219
rect 674833 254010 674899 254013
rect 675937 254010 676003 254013
rect 674833 254008 676003 254010
rect 674833 253952 674838 254008
rect 674894 253952 675942 254008
rect 675998 253952 676003 254008
rect 674833 253950 676003 253952
rect 674833 253947 674899 253950
rect 675937 253947 676003 253950
rect 40033 253874 40099 253877
rect 42885 253874 42951 253877
rect 40033 253872 42951 253874
rect 40033 253816 40038 253872
rect 40094 253816 42890 253872
rect 42946 253816 42951 253872
rect 40033 253814 42951 253816
rect 40033 253811 40099 253814
rect 42885 253811 42951 253814
rect 42425 253602 42491 253605
rect 41492 253600 42491 253602
rect 41492 253544 42430 253600
rect 42486 253544 42491 253600
rect 41492 253542 42491 253544
rect 42425 253539 42491 253542
rect 35574 253061 35634 253164
rect 35525 253056 35634 253061
rect 35801 253058 35867 253061
rect 35525 253000 35530 253056
rect 35586 253000 35634 253056
rect 35525 252998 35634 253000
rect 35758 253056 35867 253058
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35525 252995 35591 252998
rect 35758 252995 35867 253000
rect 40401 253058 40467 253061
rect 45369 253058 45435 253061
rect 40401 253056 45435 253058
rect 40401 253000 40406 253056
rect 40462 253000 45374 253056
rect 45430 253000 45435 253056
rect 40401 252998 45435 253000
rect 40401 252995 40467 252998
rect 45369 252995 45435 252998
rect 35758 252756 35818 252995
rect 511901 252922 511967 252925
rect 508484 252920 511967 252922
rect 508484 252864 511906 252920
rect 511962 252864 511967 252920
rect 508484 252862 511967 252864
rect 511901 252859 511967 252862
rect 39757 252650 39823 252653
rect 43437 252650 43503 252653
rect 39757 252648 43503 252650
rect 39757 252592 39762 252648
rect 39818 252592 43442 252648
rect 43498 252592 43503 252648
rect 39757 252590 43503 252592
rect 39757 252587 39823 252590
rect 43437 252587 43503 252590
rect 674966 252588 674972 252652
rect 675036 252650 675042 252652
rect 680997 252650 681063 252653
rect 675036 252648 681063 252650
rect 675036 252592 681002 252648
rect 681058 252592 681063 252648
rect 675036 252590 681063 252592
rect 675036 252588 675042 252590
rect 680997 252587 681063 252590
rect 30974 252245 31034 252348
rect 30974 252240 31083 252245
rect 30974 252184 31022 252240
rect 31078 252184 31083 252240
rect 30974 252182 31083 252184
rect 31017 252179 31083 252182
rect 41689 252242 41755 252245
rect 45553 252242 45619 252245
rect 41689 252240 45619 252242
rect 41689 252184 41694 252240
rect 41750 252184 45558 252240
rect 45614 252184 45619 252240
rect 41689 252182 45619 252184
rect 41689 252179 41755 252182
rect 45553 252179 45619 252182
rect 35574 251837 35634 251940
rect 35525 251832 35634 251837
rect 35801 251834 35867 251837
rect 35525 251776 35530 251832
rect 35586 251776 35634 251832
rect 35525 251774 35634 251776
rect 35758 251832 35867 251834
rect 35758 251776 35806 251832
rect 35862 251776 35867 251832
rect 35525 251771 35591 251774
rect 35758 251771 35867 251776
rect 41505 251834 41571 251837
rect 44541 251834 44607 251837
rect 41505 251832 44607 251834
rect 41505 251776 41510 251832
rect 41566 251776 44546 251832
rect 44602 251776 44607 251832
rect 41505 251774 44607 251776
rect 41505 251771 41571 251774
rect 44541 251771 44607 251774
rect 35758 251532 35818 251771
rect 41689 251426 41755 251429
rect 47025 251426 47091 251429
rect 41689 251424 47091 251426
rect 41689 251368 41694 251424
rect 41750 251368 47030 251424
rect 47086 251368 47091 251424
rect 41689 251366 47091 251368
rect 41689 251363 41755 251366
rect 47025 251363 47091 251366
rect 35390 251021 35450 251124
rect 35390 251016 35499 251021
rect 35390 250960 35438 251016
rect 35494 250960 35499 251016
rect 35390 250958 35499 250960
rect 35433 250955 35499 250958
rect 35574 250613 35634 250716
rect 35574 250608 35683 250613
rect 35574 250552 35622 250608
rect 35678 250552 35683 250608
rect 35574 250550 35683 250552
rect 35617 250547 35683 250550
rect 510613 250474 510679 250477
rect 508484 250472 510679 250474
rect 508484 250416 510618 250472
rect 510674 250416 510679 250472
rect 508484 250414 510679 250416
rect 510613 250411 510679 250414
rect 35758 250205 35818 250308
rect 35758 250200 35867 250205
rect 35758 250144 35806 250200
rect 35862 250144 35867 250200
rect 35758 250142 35867 250144
rect 35801 250139 35867 250142
rect 39389 250202 39455 250205
rect 43253 250202 43319 250205
rect 39389 250200 43319 250202
rect 39389 250144 39394 250200
rect 39450 250144 43258 250200
rect 43314 250144 43319 250200
rect 39389 250142 43319 250144
rect 39389 250139 39455 250142
rect 43253 250139 43319 250142
rect 675753 250202 675819 250205
rect 676990 250202 676996 250204
rect 675753 250200 676996 250202
rect 675753 250144 675758 250200
rect 675814 250144 676996 250200
rect 675753 250142 676996 250144
rect 675753 250139 675819 250142
rect 676990 250140 676996 250142
rect 677060 250140 677066 250204
rect 40542 249796 40602 249900
rect 40534 249732 40540 249796
rect 40604 249732 40610 249796
rect 673913 249660 673979 249661
rect 673862 249658 673868 249660
rect 673822 249598 673868 249658
rect 673932 249656 673979 249660
rect 673974 249600 673979 249656
rect 673862 249596 673868 249598
rect 673932 249596 673979 249600
rect 674782 249596 674788 249660
rect 674852 249658 674858 249660
rect 675109 249658 675175 249661
rect 674852 249656 675175 249658
rect 674852 249600 675114 249656
rect 675170 249600 675175 249656
rect 674852 249598 675175 249600
rect 674852 249596 674858 249598
rect 673913 249595 673979 249596
rect 675109 249595 675175 249598
rect 675293 249658 675359 249661
rect 676070 249658 676076 249660
rect 675293 249656 676076 249658
rect 675293 249600 675298 249656
rect 675354 249600 676076 249656
rect 675293 249598 676076 249600
rect 675293 249595 675359 249598
rect 676070 249596 676076 249598
rect 676140 249596 676146 249660
rect 35390 249389 35450 249492
rect 35390 249384 35499 249389
rect 35390 249328 35438 249384
rect 35494 249328 35499 249384
rect 35390 249326 35499 249328
rect 35433 249323 35499 249326
rect 35574 248981 35634 249084
rect 35574 248976 35683 248981
rect 35574 248920 35622 248976
rect 35678 248920 35683 248976
rect 35574 248918 35683 248920
rect 35617 248915 35683 248918
rect 35758 248573 35818 248676
rect 35758 248568 35867 248573
rect 35758 248512 35806 248568
rect 35862 248512 35867 248568
rect 35758 248510 35867 248512
rect 35801 248507 35867 248510
rect 39113 248570 39179 248573
rect 43805 248570 43871 248573
rect 39113 248568 43871 248570
rect 39113 248512 39118 248568
rect 39174 248512 43810 248568
rect 43866 248512 43871 248568
rect 39113 248510 43871 248512
rect 39113 248507 39179 248510
rect 43805 248507 43871 248510
rect 35758 248165 35818 248268
rect 35758 248160 35867 248165
rect 35758 248104 35806 248160
rect 35862 248104 35867 248160
rect 35758 248102 35867 248104
rect 35801 248099 35867 248102
rect 511073 248026 511139 248029
rect 508484 248024 511139 248026
rect 508484 247968 511078 248024
rect 511134 247968 511139 248024
rect 508484 247966 511139 247968
rect 511073 247963 511139 247966
rect 35574 247757 35634 247860
rect 35574 247752 35683 247757
rect 35574 247696 35622 247752
rect 35678 247696 35683 247752
rect 35574 247694 35683 247696
rect 35617 247691 35683 247694
rect 673269 247754 673335 247757
rect 675477 247754 675543 247757
rect 673269 247752 675543 247754
rect 673269 247696 673274 247752
rect 673330 247696 675482 247752
rect 675538 247696 675543 247752
rect 673269 247694 675543 247696
rect 673269 247691 673335 247694
rect 675477 247691 675543 247694
rect 35758 247349 35818 247452
rect 35758 247344 35867 247349
rect 35758 247288 35806 247344
rect 35862 247288 35867 247344
rect 35758 247286 35867 247288
rect 35801 247283 35867 247286
rect 40401 247346 40467 247349
rect 44173 247346 44239 247349
rect 40401 247344 44239 247346
rect 40401 247288 40406 247344
rect 40462 247288 44178 247344
rect 44234 247288 44239 247344
rect 40401 247286 44239 247288
rect 40401 247283 40467 247286
rect 44173 247283 44239 247286
rect 671797 247074 671863 247077
rect 675477 247074 675543 247077
rect 671797 247072 675543 247074
rect 40726 246940 40786 247044
rect 671797 247016 671802 247072
rect 671858 247016 675482 247072
rect 675538 247016 675543 247072
rect 671797 247014 675543 247016
rect 671797 247011 671863 247014
rect 675477 247011 675543 247014
rect 40718 246876 40724 246940
rect 40788 246876 40794 246940
rect 675753 246666 675819 246669
rect 676806 246666 676812 246668
rect 675753 246664 676812 246666
rect 41462 246530 41522 246636
rect 675753 246608 675758 246664
rect 675814 246608 676812 246664
rect 675753 246606 676812 246608
rect 675753 246603 675819 246606
rect 676806 246604 676812 246606
rect 676876 246604 676882 246668
rect 41462 246470 51090 246530
rect 39849 245714 39915 245717
rect 45737 245714 45803 245717
rect 39849 245712 45803 245714
rect 39849 245656 39854 245712
rect 39910 245656 45742 245712
rect 45798 245656 45803 245712
rect 39849 245654 45803 245656
rect 51030 245714 51090 246470
rect 675477 245988 675543 245989
rect 675477 245984 675524 245988
rect 675588 245986 675594 245988
rect 675477 245928 675482 245984
rect 675477 245924 675524 245928
rect 675588 245926 675634 245986
rect 675588 245924 675594 245926
rect 675477 245923 675543 245924
rect 668158 245788 668164 245852
rect 668228 245850 668234 245852
rect 668393 245850 668459 245853
rect 668228 245848 668459 245850
rect 668228 245792 668398 245848
rect 668454 245792 668459 245848
rect 668228 245790 668459 245792
rect 668228 245788 668234 245790
rect 668393 245787 668459 245790
rect 130377 245714 130443 245717
rect 666737 245716 666803 245717
rect 668025 245716 668091 245717
rect 666686 245714 666692 245716
rect 51030 245712 130443 245714
rect 51030 245656 130382 245712
rect 130438 245656 130443 245712
rect 51030 245654 130443 245656
rect 666646 245654 666692 245714
rect 666756 245712 666803 245716
rect 667974 245714 667980 245716
rect 666798 245656 666803 245712
rect 39849 245651 39915 245654
rect 45737 245651 45803 245654
rect 130377 245651 130443 245654
rect 666686 245652 666692 245654
rect 666756 245652 666803 245656
rect 667934 245654 667980 245714
rect 668044 245712 668091 245716
rect 668086 245656 668091 245712
rect 667974 245652 667980 245654
rect 668044 245652 668091 245656
rect 666737 245651 666803 245652
rect 668025 245651 668091 245652
rect 511809 245578 511875 245581
rect 508484 245576 511875 245578
rect 508484 245520 511814 245576
rect 511870 245520 511875 245576
rect 508484 245518 511875 245520
rect 511809 245515 511875 245518
rect 666502 245380 666508 245444
rect 666572 245442 666578 245444
rect 666737 245442 666803 245445
rect 666572 245440 666803 245442
rect 666572 245384 666742 245440
rect 666798 245384 666803 245440
rect 666572 245382 666803 245384
rect 666572 245380 666578 245382
rect 666737 245379 666803 245382
rect 40125 245170 40191 245173
rect 43069 245170 43135 245173
rect 40125 245168 43135 245170
rect 40125 245112 40130 245168
rect 40186 245112 43074 245168
rect 43130 245112 43135 245168
rect 40125 245110 43135 245112
rect 40125 245107 40191 245110
rect 43069 245107 43135 245110
rect 511257 243130 511323 243133
rect 508484 243128 511323 243130
rect 508484 243072 511262 243128
rect 511318 243072 511323 243128
rect 508484 243070 511323 243072
rect 511257 243067 511323 243070
rect 510705 240682 510771 240685
rect 508484 240680 510771 240682
rect 508484 240624 510710 240680
rect 510766 240624 510771 240680
rect 508484 240622 510771 240624
rect 510705 240619 510771 240622
rect 42057 240138 42123 240141
rect 44541 240138 44607 240141
rect 42057 240136 44607 240138
rect 42057 240080 42062 240136
rect 42118 240080 44546 240136
rect 44602 240080 44607 240136
rect 42057 240078 44607 240080
rect 42057 240075 42123 240078
rect 44541 240075 44607 240078
rect 675385 238644 675451 238645
rect 675334 238642 675340 238644
rect 675294 238582 675340 238642
rect 675404 238640 675451 238644
rect 675446 238584 675451 238640
rect 675334 238580 675340 238582
rect 675404 238580 675451 238584
rect 675385 238579 675451 238580
rect 40718 238444 40724 238508
rect 40788 238506 40794 238508
rect 41781 238506 41847 238509
rect 40788 238504 41847 238506
rect 40788 238448 41786 238504
rect 41842 238448 41847 238504
rect 40788 238446 41847 238448
rect 40788 238444 40794 238446
rect 41781 238443 41847 238446
rect 42057 238370 42123 238373
rect 42609 238370 42675 238373
rect 42057 238368 42675 238370
rect 42057 238312 42062 238368
rect 42118 238312 42614 238368
rect 42670 238312 42675 238368
rect 42057 238310 42675 238312
rect 42057 238307 42123 238310
rect 42609 238307 42675 238310
rect 507534 237965 507594 238204
rect 507485 237960 507594 237965
rect 507485 237904 507490 237960
rect 507546 237904 507594 237960
rect 507485 237902 507594 237904
rect 507485 237899 507551 237902
rect 42006 237628 42012 237692
rect 42076 237690 42082 237692
rect 42241 237690 42307 237693
rect 42076 237688 42307 237690
rect 42076 237632 42246 237688
rect 42302 237632 42307 237688
rect 42076 237630 42307 237632
rect 42076 237628 42082 237630
rect 42241 237627 42307 237630
rect 42425 237420 42491 237421
rect 42374 237418 42380 237420
rect 42334 237358 42380 237418
rect 42444 237416 42491 237420
rect 42486 237360 42491 237416
rect 42374 237356 42380 237358
rect 42444 237356 42491 237360
rect 42425 237355 42491 237356
rect 40534 236540 40540 236604
rect 40604 236602 40610 236604
rect 41781 236602 41847 236605
rect 40604 236600 41847 236602
rect 40604 236544 41786 236600
rect 41842 236544 41847 236600
rect 40604 236542 41847 236544
rect 40604 236540 40610 236542
rect 41781 236539 41847 236542
rect 510889 235786 510955 235789
rect 508484 235784 510955 235786
rect 508484 235728 510894 235784
rect 510950 235728 510955 235784
rect 508484 235726 510955 235728
rect 510889 235723 510955 235726
rect 510613 233338 510679 233341
rect 508484 233336 510679 233338
rect 508484 233280 510618 233336
rect 510674 233280 510679 233336
rect 508484 233278 510679 233280
rect 510613 233275 510679 233278
rect 129181 230890 129247 230893
rect 132585 230890 132651 230893
rect 129181 230888 132651 230890
rect 129181 230832 129186 230888
rect 129242 230832 132590 230888
rect 132646 230832 132651 230888
rect 129181 230830 132651 230832
rect 129181 230827 129247 230830
rect 132585 230827 132651 230830
rect 144637 230890 144703 230893
rect 153837 230890 153903 230893
rect 144637 230888 153903 230890
rect 144637 230832 144642 230888
rect 144698 230832 153842 230888
rect 153898 230832 153903 230888
rect 144637 230830 153903 230832
rect 144637 230827 144703 230830
rect 153837 230827 153903 230830
rect 166809 230890 166875 230893
rect 169293 230890 169359 230893
rect 166809 230888 169359 230890
rect 166809 230832 166814 230888
rect 166870 230832 169298 230888
rect 169354 230832 169359 230888
rect 166809 230830 169359 230832
rect 166809 230827 166875 230830
rect 169293 230827 169359 230830
rect 132493 230618 132559 230621
rect 164325 230618 164391 230621
rect 132493 230616 151830 230618
rect 132493 230560 132498 230616
rect 132554 230560 151830 230616
rect 132493 230558 151830 230560
rect 132493 230555 132559 230558
rect 151770 230482 151830 230558
rect 152230 230616 164391 230618
rect 152230 230560 164330 230616
rect 164386 230560 164391 230616
rect 152230 230558 164391 230560
rect 152230 230482 152290 230558
rect 164325 230555 164391 230558
rect 484761 230618 484827 230621
rect 491385 230618 491451 230621
rect 484761 230616 491451 230618
rect 484761 230560 484766 230616
rect 484822 230560 491390 230616
rect 491446 230560 491451 230616
rect 484761 230558 491451 230560
rect 484761 230555 484827 230558
rect 491385 230555 491451 230558
rect 151770 230422 152290 230482
rect 190269 230482 190335 230485
rect 190453 230482 190519 230485
rect 190269 230480 190519 230482
rect 190269 230424 190274 230480
rect 190330 230424 190458 230480
rect 190514 230424 190519 230480
rect 190269 230422 190519 230424
rect 190269 230419 190335 230422
rect 190453 230419 190519 230422
rect 61377 230346 61443 230349
rect 145833 230346 145899 230349
rect 61377 230344 145899 230346
rect 61377 230288 61382 230344
rect 61438 230288 145838 230344
rect 145894 230288 145899 230344
rect 61377 230286 145899 230288
rect 61377 230283 61443 230286
rect 145833 230283 145899 230286
rect 146017 230346 146083 230349
rect 150525 230346 150591 230349
rect 146017 230344 150591 230346
rect 146017 230288 146022 230344
rect 146078 230288 150530 230344
rect 150586 230288 150591 230344
rect 146017 230286 150591 230288
rect 146017 230283 146083 230286
rect 150525 230283 150591 230286
rect 153745 230346 153811 230349
rect 160461 230346 160527 230349
rect 153745 230344 160527 230346
rect 153745 230288 153750 230344
rect 153806 230288 160466 230344
rect 160522 230288 160527 230344
rect 153745 230286 160527 230288
rect 153745 230283 153811 230286
rect 160461 230283 160527 230286
rect 161473 230346 161539 230349
rect 166993 230346 167059 230349
rect 161473 230344 167059 230346
rect 161473 230288 161478 230344
rect 161534 230288 166998 230344
rect 167054 230288 167059 230344
rect 161473 230286 167059 230288
rect 161473 230283 161539 230286
rect 166993 230283 167059 230286
rect 168833 230346 168899 230349
rect 172053 230346 172119 230349
rect 168833 230344 172119 230346
rect 168833 230288 168838 230344
rect 168894 230288 172058 230344
rect 172114 230288 172119 230344
rect 168833 230286 172119 230288
rect 168833 230283 168899 230286
rect 172053 230283 172119 230286
rect 483289 230346 483355 230349
rect 488441 230346 488507 230349
rect 483289 230344 488507 230346
rect 483289 230288 483294 230344
rect 483350 230288 488446 230344
rect 488502 230288 488507 230344
rect 483289 230286 488507 230288
rect 483289 230283 483355 230286
rect 488441 230283 488507 230286
rect 56041 230074 56107 230077
rect 654133 230074 654199 230077
rect 56041 230072 654199 230074
rect 56041 230016 56046 230072
rect 56102 230016 654138 230072
rect 654194 230016 654199 230072
rect 56041 230014 654199 230016
rect 56041 230011 56107 230014
rect 654133 230011 654199 230014
rect 54661 229802 54727 229805
rect 654317 229802 654383 229805
rect 54661 229800 654383 229802
rect 54661 229744 54666 229800
rect 54722 229744 654322 229800
rect 654378 229744 654383 229800
rect 54661 229742 654383 229744
rect 54661 229739 54727 229742
rect 654317 229739 654383 229742
rect 111057 229530 111123 229533
rect 165153 229530 165219 229533
rect 111057 229528 165219 229530
rect 111057 229472 111062 229528
rect 111118 229472 165158 229528
rect 165214 229472 165219 229528
rect 111057 229470 165219 229472
rect 111057 229467 111123 229470
rect 165153 229467 165219 229470
rect 170029 229530 170095 229533
rect 174997 229530 175063 229533
rect 170029 229528 175063 229530
rect 170029 229472 170034 229528
rect 170090 229472 175002 229528
rect 175058 229472 175063 229528
rect 170029 229470 175063 229472
rect 170029 229467 170095 229470
rect 174997 229467 175063 229470
rect 190913 229530 190979 229533
rect 196065 229530 196131 229533
rect 190913 229528 196131 229530
rect 190913 229472 190918 229528
rect 190974 229472 196070 229528
rect 196126 229472 196131 229528
rect 190913 229470 196131 229472
rect 190913 229467 190979 229470
rect 196065 229467 196131 229470
rect 214097 229530 214163 229533
rect 214649 229530 214715 229533
rect 214097 229528 214715 229530
rect 214097 229472 214102 229528
rect 214158 229472 214654 229528
rect 214710 229472 214715 229528
rect 214097 229470 214715 229472
rect 214097 229467 214163 229470
rect 214649 229467 214715 229470
rect 483289 229530 483355 229533
rect 489177 229530 489243 229533
rect 483289 229528 489243 229530
rect 483289 229472 483294 229528
rect 483350 229472 489182 229528
rect 489238 229472 489243 229528
rect 483289 229470 489243 229472
rect 483289 229467 483355 229470
rect 489177 229467 489243 229470
rect 202597 229394 202663 229397
rect 204529 229394 204595 229397
rect 202597 229392 204595 229394
rect 202597 229336 202602 229392
rect 202658 229336 204534 229392
rect 204590 229336 204595 229392
rect 202597 229334 204595 229336
rect 202597 229331 202663 229334
rect 204529 229331 204595 229334
rect 145833 229258 145899 229261
rect 151905 229258 151971 229261
rect 145833 229256 151971 229258
rect 145833 229200 145838 229256
rect 145894 229200 151910 229256
rect 151966 229200 151971 229256
rect 145833 229198 151971 229200
rect 145833 229195 145899 229198
rect 151905 229195 151971 229198
rect 190637 229258 190703 229261
rect 191557 229258 191623 229261
rect 190637 229256 191623 229258
rect 190637 229200 190642 229256
rect 190698 229200 191562 229256
rect 191618 229200 191623 229256
rect 190637 229198 191623 229200
rect 190637 229195 190703 229198
rect 191557 229195 191623 229198
rect 158437 229122 158503 229125
rect 163773 229122 163839 229125
rect 158437 229120 163839 229122
rect 158437 229064 158442 229120
rect 158498 229064 163778 229120
rect 163834 229064 163839 229120
rect 158437 229062 163839 229064
rect 158437 229059 158503 229062
rect 163773 229059 163839 229062
rect 41965 228988 42031 228989
rect 41965 228984 42012 228988
rect 42076 228986 42082 228988
rect 41965 228928 41970 228984
rect 41965 228924 42012 228928
rect 42076 228926 42122 228986
rect 42076 228924 42082 228926
rect 41965 228923 42031 228924
rect 46381 228850 46447 228853
rect 647325 228850 647391 228853
rect 46381 228848 647391 228850
rect 46381 228792 46386 228848
rect 46442 228792 647330 228848
rect 647386 228792 647391 228848
rect 46381 228790 647391 228792
rect 46381 228787 46447 228790
rect 647325 228787 647391 228790
rect 49141 228578 49207 228581
rect 653029 228578 653095 228581
rect 49141 228576 653095 228578
rect 49141 228520 49146 228576
rect 49202 228520 653034 228576
rect 653090 228520 653095 228576
rect 49141 228518 653095 228520
rect 49141 228515 49207 228518
rect 653029 228515 653095 228518
rect 47761 228306 47827 228309
rect 651557 228306 651623 228309
rect 47761 228304 651623 228306
rect 47761 228248 47766 228304
rect 47822 228248 651562 228304
rect 651618 228248 651623 228304
rect 47761 228246 651623 228248
rect 47761 228243 47827 228246
rect 651557 228243 651623 228246
rect 142889 228034 142955 228037
rect 150801 228034 150867 228037
rect 142889 228032 150867 228034
rect 142889 227976 142894 228032
rect 142950 227976 150806 228032
rect 150862 227976 150867 228032
rect 142889 227974 150867 227976
rect 142889 227971 142955 227974
rect 150801 227971 150867 227974
rect 156597 228034 156663 228037
rect 160185 228034 160251 228037
rect 156597 228032 160251 228034
rect 156597 227976 156602 228032
rect 156658 227976 160190 228032
rect 160246 227976 160251 228032
rect 156597 227974 160251 227976
rect 156597 227971 156663 227974
rect 160185 227971 160251 227974
rect 172329 228034 172395 228037
rect 182357 228034 182423 228037
rect 172329 228032 182423 228034
rect 172329 227976 172334 228032
rect 172390 227976 182362 228032
rect 182418 227976 182423 228032
rect 172329 227974 182423 227976
rect 172329 227971 172395 227974
rect 182357 227971 182423 227974
rect 142153 227762 142219 227765
rect 153285 227762 153351 227765
rect 142153 227760 153351 227762
rect 142153 227704 142158 227760
rect 142214 227704 153290 227760
rect 153346 227704 153351 227760
rect 142153 227702 153351 227704
rect 142153 227699 142219 227702
rect 153285 227699 153351 227702
rect 157425 227762 157491 227765
rect 166533 227762 166599 227765
rect 157425 227760 166599 227762
rect 157425 227704 157430 227760
rect 157486 227704 166538 227760
rect 166594 227704 166599 227760
rect 157425 227702 166599 227704
rect 157425 227699 157491 227702
rect 166533 227699 166599 227702
rect 486417 227762 486483 227765
rect 491569 227762 491635 227765
rect 486417 227760 491635 227762
rect 486417 227704 486422 227760
rect 486478 227704 491574 227760
rect 491630 227704 491635 227760
rect 486417 227702 491635 227704
rect 486417 227699 486483 227702
rect 491569 227699 491635 227702
rect 53281 227490 53347 227493
rect 651097 227490 651163 227493
rect 53281 227488 651163 227490
rect 53281 227432 53286 227488
rect 53342 227432 651102 227488
rect 651158 227432 651163 227488
rect 53281 227430 651163 227432
rect 53281 227427 53347 227430
rect 651097 227427 651163 227430
rect 42057 227354 42123 227357
rect 42374 227354 42380 227356
rect 42057 227352 42380 227354
rect 42057 227296 42062 227352
rect 42118 227296 42380 227352
rect 42057 227294 42380 227296
rect 42057 227291 42123 227294
rect 42374 227292 42380 227294
rect 42444 227292 42450 227356
rect 50337 227218 50403 227221
rect 648061 227218 648127 227221
rect 50337 227216 648127 227218
rect 50337 227160 50342 227216
rect 50398 227160 648066 227216
rect 648122 227160 648127 227216
rect 50337 227158 648127 227160
rect 50337 227155 50403 227158
rect 648061 227155 648127 227158
rect 59997 226946 60063 226949
rect 659837 226946 659903 226949
rect 59997 226944 659903 226946
rect 59997 226888 60002 226944
rect 60058 226888 659842 226944
rect 659898 226888 659903 226944
rect 59997 226886 659903 226888
rect 59997 226883 60063 226886
rect 659837 226883 659903 226886
rect 59261 226674 59327 226677
rect 151353 226674 151419 226677
rect 59261 226672 151419 226674
rect 59261 226616 59266 226672
rect 59322 226616 151358 226672
rect 151414 226616 151419 226672
rect 59261 226614 151419 226616
rect 59261 226611 59327 226614
rect 151353 226611 151419 226614
rect 154297 226674 154363 226677
rect 157793 226674 157859 226677
rect 154297 226672 157859 226674
rect 154297 226616 154302 226672
rect 154358 226616 157798 226672
rect 157854 226616 157859 226672
rect 154297 226614 157859 226616
rect 154297 226611 154363 226614
rect 157793 226611 157859 226614
rect 185945 226674 186011 226677
rect 187969 226674 188035 226677
rect 185945 226672 188035 226674
rect 185945 226616 185950 226672
rect 186006 226616 187974 226672
rect 188030 226616 188035 226672
rect 185945 226614 188035 226616
rect 185945 226611 186011 226614
rect 187969 226611 188035 226614
rect 489913 226674 489979 226677
rect 490925 226674 490991 226677
rect 489913 226672 490991 226674
rect 489913 226616 489918 226672
rect 489974 226616 490930 226672
rect 490986 226616 490991 226672
rect 489913 226614 490991 226616
rect 489913 226611 489979 226614
rect 490925 226611 490991 226614
rect 142337 226504 142403 226507
rect 142110 226502 142403 226504
rect 142110 226446 142342 226502
rect 142398 226446 142403 226502
rect 142110 226444 142403 226446
rect 141693 226402 141759 226405
rect 142110 226402 142170 226444
rect 142337 226441 142403 226444
rect 141693 226400 142170 226402
rect 141693 226344 141698 226400
rect 141754 226344 142170 226400
rect 141693 226342 142170 226344
rect 489545 226402 489611 226405
rect 490005 226402 490071 226405
rect 489545 226400 490071 226402
rect 489545 226344 489550 226400
rect 489606 226344 490010 226400
rect 490066 226344 490071 226400
rect 489545 226342 490071 226344
rect 141693 226339 141759 226342
rect 489545 226339 489611 226342
rect 490005 226339 490071 226342
rect 166993 226266 167059 226269
rect 173617 226266 173683 226269
rect 166993 226264 173683 226266
rect 166993 226208 166998 226264
rect 167054 226208 173622 226264
rect 173678 226208 173683 226264
rect 166993 226206 173683 226208
rect 166993 226203 167059 226206
rect 173617 226203 173683 226206
rect 190269 226266 190335 226269
rect 191373 226266 191439 226269
rect 190269 226264 191439 226266
rect 190269 226208 190274 226264
rect 190330 226208 191378 226264
rect 191434 226208 191439 226264
rect 190269 226206 191439 226208
rect 190269 226203 190335 226206
rect 191373 226203 191439 226206
rect 56869 226130 56935 226133
rect 149145 226130 149211 226133
rect 56869 226128 149211 226130
rect 56869 226072 56874 226128
rect 56930 226072 149150 226128
rect 149206 226072 149211 226128
rect 56869 226070 149211 226072
rect 56869 226067 56935 226070
rect 149145 226067 149211 226070
rect 176469 226130 176535 226133
rect 176745 226130 176811 226133
rect 176469 226128 176811 226130
rect 176469 226072 176474 226128
rect 176530 226072 176750 226128
rect 176806 226072 176811 226128
rect 176469 226070 176811 226072
rect 176469 226067 176535 226070
rect 176745 226067 176811 226070
rect 180793 226130 180859 226133
rect 181345 226130 181411 226133
rect 180793 226128 181411 226130
rect 180793 226072 180798 226128
rect 180854 226072 181350 226128
rect 181406 226072 181411 226128
rect 180793 226070 181411 226072
rect 180793 226067 180859 226070
rect 181345 226067 181411 226070
rect 467557 226130 467623 226133
rect 537477 226130 537543 226133
rect 467557 226128 537543 226130
rect 467557 226072 467562 226128
rect 467618 226072 537482 226128
rect 537538 226072 537543 226128
rect 467557 226070 537543 226072
rect 467557 226067 467623 226070
rect 537477 226067 537543 226070
rect 130377 225858 130443 225861
rect 661493 225858 661559 225861
rect 130377 225856 661559 225858
rect 130377 225800 130382 225856
rect 130438 225800 661498 225856
rect 661554 225800 661559 225856
rect 130377 225798 661559 225800
rect 130377 225795 130443 225798
rect 661493 225795 661559 225798
rect 128997 225586 129063 225589
rect 662413 225586 662479 225589
rect 128997 225584 662479 225586
rect 128997 225528 129002 225584
rect 129058 225528 662418 225584
rect 662474 225528 662479 225584
rect 128997 225526 662479 225528
rect 128997 225523 129063 225526
rect 662413 225523 662479 225526
rect 151445 225314 151511 225317
rect 152733 225314 152799 225317
rect 151445 225312 152799 225314
rect 151445 225256 151450 225312
rect 151506 225256 152738 225312
rect 152794 225256 152799 225312
rect 151445 225254 152799 225256
rect 151445 225251 151511 225254
rect 152733 225251 152799 225254
rect 178125 225314 178191 225317
rect 179873 225314 179939 225317
rect 178125 225312 179939 225314
rect 178125 225256 178130 225312
rect 178186 225256 179878 225312
rect 179934 225256 179939 225312
rect 178125 225254 179939 225256
rect 178125 225251 178191 225254
rect 179873 225251 179939 225254
rect 212349 225314 212415 225317
rect 214741 225314 214807 225317
rect 212349 225312 214807 225314
rect 212349 225256 212354 225312
rect 212410 225256 214746 225312
rect 214802 225256 214807 225312
rect 212349 225254 214807 225256
rect 212349 225251 212415 225254
rect 214741 225251 214807 225254
rect 459369 225314 459435 225317
rect 525057 225314 525123 225317
rect 459369 225312 525123 225314
rect 459369 225256 459374 225312
rect 459430 225256 525062 225312
rect 525118 225256 525123 225312
rect 459369 225254 525123 225256
rect 459369 225251 459435 225254
rect 525057 225251 525123 225254
rect 151629 225042 151695 225045
rect 152181 225042 152247 225045
rect 151629 225040 152247 225042
rect 151629 224984 151634 225040
rect 151690 224984 152186 225040
rect 152242 224984 152247 225040
rect 151629 224982 152247 224984
rect 151629 224979 151695 224982
rect 152181 224979 152247 224982
rect 187049 225042 187115 225045
rect 189993 225042 190059 225045
rect 187049 225040 190059 225042
rect 187049 224984 187054 225040
rect 187110 224984 189998 225040
rect 190054 224984 190059 225040
rect 187049 224982 190059 224984
rect 187049 224979 187115 224982
rect 189993 224979 190059 224982
rect 486785 225042 486851 225045
rect 489729 225042 489795 225045
rect 486785 225040 489795 225042
rect 486785 224984 486790 225040
rect 486846 224984 489734 225040
rect 489790 224984 489795 225040
rect 486785 224982 489795 224984
rect 486785 224979 486851 224982
rect 489729 224979 489795 224982
rect 489913 225042 489979 225045
rect 492765 225042 492831 225045
rect 489913 225040 492831 225042
rect 489913 224984 489918 225040
rect 489974 224984 492770 225040
rect 492826 224984 492831 225040
rect 489913 224982 492831 224984
rect 489913 224979 489979 224982
rect 492765 224979 492831 224982
rect 214373 224906 214439 224909
rect 215569 224906 215635 224909
rect 214373 224904 215635 224906
rect 214373 224848 214378 224904
rect 214434 224848 215574 224904
rect 215630 224848 215635 224904
rect 214373 224846 215635 224848
rect 214373 224843 214439 224846
rect 215569 224843 215635 224846
rect 157333 224770 157399 224773
rect 161473 224770 161539 224773
rect 157333 224768 161539 224770
rect 157333 224712 157338 224768
rect 157394 224712 161478 224768
rect 161534 224712 161539 224768
rect 157333 224710 161539 224712
rect 157333 224707 157399 224710
rect 161473 224707 161539 224710
rect 190361 224770 190427 224773
rect 190637 224770 190703 224773
rect 190361 224768 190703 224770
rect 190361 224712 190366 224768
rect 190422 224712 190642 224768
rect 190698 224712 190703 224768
rect 190361 224710 190703 224712
rect 190361 224707 190427 224710
rect 190637 224707 190703 224710
rect 481081 224634 481147 224637
rect 481449 224634 481515 224637
rect 481081 224632 481515 224634
rect 481081 224576 481086 224632
rect 481142 224576 481454 224632
rect 481510 224576 481515 224632
rect 481081 224574 481515 224576
rect 481081 224571 481147 224574
rect 481449 224571 481515 224574
rect 499573 224634 499639 224637
rect 505185 224634 505251 224637
rect 499573 224632 505251 224634
rect 499573 224576 499578 224632
rect 499634 224576 505190 224632
rect 505246 224576 505251 224632
rect 499573 224574 505251 224576
rect 499573 224571 499639 224574
rect 505185 224571 505251 224574
rect 524229 224634 524295 224637
rect 526345 224634 526411 224637
rect 524229 224632 526411 224634
rect 524229 224576 524234 224632
rect 524290 224576 526350 224632
rect 526406 224576 526411 224632
rect 524229 224574 526411 224576
rect 524229 224571 524295 224574
rect 526345 224571 526411 224574
rect 147029 224498 147095 224501
rect 151905 224498 151971 224501
rect 147029 224496 151971 224498
rect 147029 224440 147034 224496
rect 147090 224440 151910 224496
rect 151966 224440 151971 224496
rect 147029 224438 151971 224440
rect 147029 224435 147095 224438
rect 151905 224435 151971 224438
rect 155033 224498 155099 224501
rect 157425 224498 157491 224501
rect 155033 224496 157491 224498
rect 155033 224440 155038 224496
rect 155094 224440 157430 224496
rect 157486 224440 157491 224496
rect 155033 224438 157491 224440
rect 155033 224435 155099 224438
rect 157425 224435 157491 224438
rect 157793 224498 157859 224501
rect 159909 224498 159975 224501
rect 157793 224496 159975 224498
rect 157793 224440 157798 224496
rect 157854 224440 159914 224496
rect 159970 224440 159975 224496
rect 157793 224438 159975 224440
rect 157793 224435 157859 224438
rect 159909 224435 159975 224438
rect 485221 224498 485287 224501
rect 489085 224498 489151 224501
rect 485221 224496 489151 224498
rect 485221 224440 485226 224496
rect 485282 224440 489090 224496
rect 489146 224440 489151 224496
rect 485221 224438 489151 224440
rect 485221 224435 485287 224438
rect 489085 224435 489151 224438
rect 206829 224362 206895 224365
rect 208761 224362 208827 224365
rect 206829 224360 208827 224362
rect 206829 224304 206834 224360
rect 206890 224304 208766 224360
rect 208822 224304 208827 224360
rect 206829 224302 208827 224304
rect 206829 224299 206895 224302
rect 208761 224299 208827 224302
rect 479977 224362 480043 224365
rect 481081 224362 481147 224365
rect 479977 224360 481147 224362
rect 479977 224304 479982 224360
rect 480038 224304 481086 224360
rect 481142 224304 481147 224360
rect 479977 224302 481147 224304
rect 479977 224299 480043 224302
rect 481081 224299 481147 224302
rect 499297 224362 499363 224365
rect 499665 224362 499731 224365
rect 499297 224360 499731 224362
rect 499297 224304 499302 224360
rect 499358 224304 499670 224360
rect 499726 224304 499731 224360
rect 499297 224302 499731 224304
rect 499297 224299 499363 224302
rect 499665 224299 499731 224302
rect 71681 224226 71747 224229
rect 157977 224226 158043 224229
rect 71681 224224 158043 224226
rect 71681 224168 71686 224224
rect 71742 224168 157982 224224
rect 158038 224168 158043 224224
rect 71681 224166 158043 224168
rect 71681 224163 71747 224166
rect 157977 224163 158043 224166
rect 193489 224226 193555 224229
rect 199193 224226 199259 224229
rect 193489 224224 199259 224226
rect 193489 224168 193494 224224
rect 193550 224168 199198 224224
rect 199254 224168 199259 224224
rect 193489 224166 199259 224168
rect 193489 224163 193555 224166
rect 199193 224163 199259 224166
rect 28533 223954 28599 223957
rect 666737 223954 666803 223957
rect 28533 223952 666803 223954
rect 28533 223896 28538 223952
rect 28594 223896 666742 223952
rect 666798 223896 666803 223952
rect 28533 223894 666803 223896
rect 28533 223891 28599 223894
rect 666737 223891 666803 223894
rect 41689 223682 41755 223685
rect 668945 223682 669011 223685
rect 41689 223680 669011 223682
rect 41689 223624 41694 223680
rect 41750 223624 668950 223680
rect 669006 223624 669011 223680
rect 41689 223622 669011 223624
rect 41689 223619 41755 223622
rect 668945 223619 669011 223622
rect 675109 223546 675175 223549
rect 675109 223544 676292 223546
rect 675109 223488 675114 223544
rect 675170 223488 676292 223544
rect 675109 223486 676292 223488
rect 675109 223483 675175 223486
rect 150157 223410 150223 223413
rect 155585 223410 155651 223413
rect 150157 223408 155651 223410
rect 150157 223352 150162 223408
rect 150218 223352 155590 223408
rect 155646 223352 155651 223408
rect 150157 223350 155651 223352
rect 150157 223347 150223 223350
rect 155585 223347 155651 223350
rect 185025 223410 185091 223413
rect 185577 223410 185643 223413
rect 185025 223408 185643 223410
rect 185025 223352 185030 223408
rect 185086 223352 185582 223408
rect 185638 223352 185643 223408
rect 185025 223350 185643 223352
rect 185025 223347 185091 223350
rect 185577 223347 185643 223350
rect 490833 223410 490899 223413
rect 499527 223410 499593 223413
rect 490833 223408 499593 223410
rect 490833 223352 490838 223408
rect 490894 223352 499532 223408
rect 499588 223352 499593 223408
rect 490833 223350 499593 223352
rect 490833 223347 490899 223350
rect 499527 223347 499593 223350
rect 504725 223410 504791 223413
rect 510061 223410 510127 223413
rect 504725 223408 510127 223410
rect 504725 223352 504730 223408
rect 504786 223352 510066 223408
rect 510122 223352 510127 223408
rect 504725 223350 510127 223352
rect 504725 223347 504791 223350
rect 510061 223347 510127 223350
rect 514569 223410 514635 223413
rect 517421 223410 517487 223413
rect 524229 223410 524295 223413
rect 514569 223408 524295 223410
rect 514569 223352 514574 223408
rect 514630 223352 517426 223408
rect 517482 223352 524234 223408
rect 524290 223352 524295 223408
rect 514569 223350 524295 223352
rect 514569 223347 514635 223350
rect 517421 223347 517487 223350
rect 524229 223347 524295 223350
rect 142153 223138 142219 223141
rect 148317 223138 148383 223141
rect 142153 223136 148383 223138
rect 142153 223080 142158 223136
rect 142214 223080 148322 223136
rect 148378 223080 148383 223136
rect 142153 223078 148383 223080
rect 142153 223075 142219 223078
rect 148317 223075 148383 223078
rect 157149 223138 157215 223141
rect 157425 223138 157491 223141
rect 157149 223136 157491 223138
rect 157149 223080 157154 223136
rect 157210 223080 157430 223136
rect 157486 223080 157491 223136
rect 157149 223078 157491 223080
rect 157149 223075 157215 223078
rect 157425 223075 157491 223078
rect 157977 223138 158043 223141
rect 165705 223138 165771 223141
rect 157977 223136 165771 223138
rect 157977 223080 157982 223136
rect 158038 223080 165710 223136
rect 165766 223080 165771 223136
rect 157977 223078 165771 223080
rect 157977 223075 158043 223078
rect 165705 223075 165771 223078
rect 483381 223138 483447 223141
rect 485865 223138 485931 223141
rect 483381 223136 485931 223138
rect 483381 223080 483386 223136
rect 483442 223080 485870 223136
rect 485926 223080 485931 223136
rect 483381 223078 485931 223080
rect 483381 223075 483447 223078
rect 485865 223075 485931 223078
rect 489269 223138 489335 223141
rect 495249 223138 495315 223141
rect 489269 223136 495315 223138
rect 489269 223080 489274 223136
rect 489330 223080 495254 223136
rect 495310 223080 495315 223136
rect 489269 223078 495315 223080
rect 489269 223075 489335 223078
rect 495249 223075 495315 223078
rect 499297 223138 499363 223141
rect 499665 223138 499731 223141
rect 499297 223136 499731 223138
rect 499297 223080 499302 223136
rect 499358 223080 499670 223136
rect 499726 223080 499731 223136
rect 499297 223078 499731 223080
rect 499297 223075 499363 223078
rect 499665 223075 499731 223078
rect 675477 223138 675543 223141
rect 675477 223136 676292 223138
rect 675477 223080 675482 223136
rect 675538 223080 676292 223136
rect 675477 223078 676292 223080
rect 675477 223075 675543 223078
rect 173065 223002 173131 223005
rect 174077 223002 174143 223005
rect 173065 223000 174143 223002
rect 173065 222944 173070 223000
rect 173126 222944 174082 223000
rect 174138 222944 174143 223000
rect 173065 222942 174143 222944
rect 173065 222939 173131 222942
rect 174077 222939 174143 222942
rect 181161 223002 181227 223005
rect 189625 223002 189691 223005
rect 181161 223000 189691 223002
rect 181161 222944 181166 223000
rect 181222 222944 189630 223000
rect 189686 222944 189691 223000
rect 181161 222942 189691 222944
rect 181161 222939 181227 222942
rect 189625 222939 189691 222942
rect 136541 222866 136607 222869
rect 142613 222866 142679 222869
rect 136541 222864 142679 222866
rect 136541 222808 136546 222864
rect 136602 222808 142618 222864
rect 142674 222808 142679 222864
rect 136541 222806 142679 222808
rect 136541 222803 136607 222806
rect 142613 222803 142679 222806
rect 148961 222866 149027 222869
rect 157333 222866 157399 222869
rect 148961 222864 157399 222866
rect 148961 222808 148966 222864
rect 149022 222808 157338 222864
rect 157394 222808 157399 222864
rect 148961 222806 157399 222808
rect 148961 222803 149027 222806
rect 157333 222803 157399 222806
rect 157517 222866 157583 222869
rect 158345 222866 158411 222869
rect 157517 222864 158411 222866
rect 157517 222808 157522 222864
rect 157578 222808 158350 222864
rect 158406 222808 158411 222864
rect 157517 222806 158411 222808
rect 157517 222803 157583 222806
rect 158345 222803 158411 222806
rect 213361 222866 213427 222869
rect 214741 222866 214807 222869
rect 213361 222864 214807 222866
rect 213361 222808 213366 222864
rect 213422 222808 214746 222864
rect 214802 222808 214807 222864
rect 213361 222806 214807 222808
rect 213361 222803 213427 222806
rect 214741 222803 214807 222806
rect 462773 222866 462839 222869
rect 530393 222866 530459 222869
rect 462773 222864 530459 222866
rect 462773 222808 462778 222864
rect 462834 222808 530398 222864
rect 530454 222808 530459 222864
rect 462773 222806 530459 222808
rect 462773 222803 462839 222806
rect 530393 222803 530459 222806
rect 675293 222730 675359 222733
rect 180750 222670 200130 222730
rect 47577 222594 47643 222597
rect 180750 222594 180810 222670
rect 47577 222592 180810 222594
rect 47577 222536 47582 222592
rect 47638 222536 180810 222592
rect 47577 222534 180810 222536
rect 200070 222594 200130 222670
rect 675293 222728 676292 222730
rect 675293 222672 675298 222728
rect 675354 222672 676292 222728
rect 675293 222670 676292 222672
rect 675293 222667 675359 222670
rect 662873 222594 662939 222597
rect 200070 222592 662939 222594
rect 200070 222536 662878 222592
rect 662934 222536 662939 222592
rect 200070 222534 662939 222536
rect 47577 222531 47643 222534
rect 662873 222531 662939 222534
rect 40677 222322 40743 222325
rect 668393 222322 668459 222325
rect 40677 222320 668459 222322
rect 40677 222264 40682 222320
rect 40738 222264 668398 222320
rect 668454 222264 668459 222320
rect 40677 222262 668459 222264
rect 40677 222259 40743 222262
rect 668393 222259 668459 222262
rect 675477 222322 675543 222325
rect 675477 222320 676292 222322
rect 675477 222264 675482 222320
rect 675538 222264 676292 222320
rect 675477 222262 676292 222264
rect 675477 222259 675543 222262
rect 50337 222050 50403 222053
rect 59997 222050 60063 222053
rect 50337 222048 60063 222050
rect 50337 221992 50342 222048
rect 50398 221992 60002 222048
rect 60058 221992 60063 222048
rect 50337 221990 60063 221992
rect 50337 221987 50403 221990
rect 59997 221987 60063 221990
rect 66713 222050 66779 222053
rect 154757 222050 154823 222053
rect 66713 222048 154823 222050
rect 66713 221992 66718 222048
rect 66774 221992 154762 222048
rect 154818 221992 154823 222048
rect 66713 221990 154823 221992
rect 66713 221987 66779 221990
rect 154757 221987 154823 221990
rect 171133 222050 171199 222053
rect 174813 222050 174879 222053
rect 171133 222048 174879 222050
rect 171133 221992 171138 222048
rect 171194 221992 174818 222048
rect 174874 221992 174879 222048
rect 171133 221990 174879 221992
rect 171133 221987 171199 221990
rect 174813 221987 174879 221990
rect 181989 222050 182055 222053
rect 187785 222050 187851 222053
rect 181989 222048 187851 222050
rect 181989 221992 181994 222048
rect 182050 221992 187790 222048
rect 187846 221992 187851 222048
rect 181989 221990 187851 221992
rect 181989 221987 182055 221990
rect 187785 221987 187851 221990
rect 200113 222050 200179 222053
rect 205909 222050 205975 222053
rect 200113 222048 205975 222050
rect 200113 221992 200118 222048
rect 200174 221992 205914 222048
rect 205970 221992 205975 222048
rect 200113 221990 205975 221992
rect 200113 221987 200179 221990
rect 205909 221987 205975 221990
rect 458081 222050 458147 222053
rect 521653 222050 521719 222053
rect 458081 222048 521719 222050
rect 458081 221992 458086 222048
rect 458142 221992 521658 222048
rect 521714 221992 521719 222048
rect 458081 221990 521719 221992
rect 458081 221987 458147 221990
rect 521653 221987 521719 221990
rect 675109 221914 675175 221917
rect 675109 221912 676292 221914
rect 675109 221856 675114 221912
rect 675170 221856 676292 221912
rect 675109 221854 676292 221856
rect 675109 221851 675175 221854
rect 51717 221778 51783 221781
rect 669129 221778 669195 221781
rect 51717 221776 669195 221778
rect 51717 221720 51722 221776
rect 51778 221720 669134 221776
rect 669190 221720 669195 221776
rect 51717 221718 669195 221720
rect 51717 221715 51783 221718
rect 669129 221715 669195 221718
rect 59997 221506 60063 221509
rect 663793 221506 663859 221509
rect 59997 221504 663859 221506
rect 59997 221448 60002 221504
rect 60058 221448 663798 221504
rect 663854 221448 663859 221504
rect 59997 221446 663859 221448
rect 59997 221443 60063 221446
rect 663793 221443 663859 221446
rect 675477 221506 675543 221509
rect 675477 221504 676292 221506
rect 675477 221448 675482 221504
rect 675538 221448 676292 221504
rect 675477 221446 676292 221448
rect 675477 221443 675543 221446
rect 72877 221234 72943 221237
rect 151629 221234 151695 221237
rect 156229 221234 156295 221237
rect 72877 221232 142170 221234
rect 72877 221176 72882 221232
rect 72938 221176 142170 221232
rect 72877 221174 142170 221176
rect 72877 221171 72943 221174
rect 142110 220962 142170 221174
rect 151629 221232 156295 221234
rect 151629 221176 151634 221232
rect 151690 221176 156234 221232
rect 156290 221176 156295 221232
rect 151629 221174 156295 221176
rect 151629 221171 151695 221174
rect 156229 221171 156295 221174
rect 159817 221234 159883 221237
rect 160921 221234 160987 221237
rect 159817 221232 160987 221234
rect 159817 221176 159822 221232
rect 159878 221176 160926 221232
rect 160982 221176 160987 221232
rect 159817 221174 160987 221176
rect 159817 221171 159883 221174
rect 160921 221171 160987 221174
rect 161105 221234 161171 221237
rect 166625 221234 166691 221237
rect 161105 221232 166691 221234
rect 161105 221176 161110 221232
rect 161166 221176 166630 221232
rect 166686 221176 166691 221232
rect 161105 221174 166691 221176
rect 161105 221171 161171 221174
rect 166625 221171 166691 221174
rect 192293 221234 192359 221237
rect 196341 221234 196407 221237
rect 192293 221232 196407 221234
rect 192293 221176 192298 221232
rect 192354 221176 196346 221232
rect 196402 221176 196407 221232
rect 192293 221174 196407 221176
rect 192293 221171 192359 221174
rect 196341 221171 196407 221174
rect 437289 221234 437355 221237
rect 481449 221234 481515 221237
rect 485865 221234 485931 221237
rect 437289 221232 470610 221234
rect 437289 221176 437294 221232
rect 437350 221176 470610 221232
rect 437289 221174 470610 221176
rect 437289 221171 437355 221174
rect 166809 221098 166875 221101
rect 171225 221098 171291 221101
rect 166809 221096 171291 221098
rect 166809 221040 166814 221096
rect 166870 221040 171230 221096
rect 171286 221040 171291 221096
rect 166809 221038 171291 221040
rect 166809 221035 166875 221038
rect 171225 221035 171291 221038
rect 199469 221098 199535 221101
rect 200297 221098 200363 221101
rect 199469 221096 200363 221098
rect 199469 221040 199474 221096
rect 199530 221040 200302 221096
rect 200358 221040 200363 221096
rect 199469 221038 200363 221040
rect 199469 221035 199535 221038
rect 200297 221035 200363 221038
rect 158897 220962 158963 220965
rect 142110 220960 158963 220962
rect 142110 220904 158902 220960
rect 158958 220904 158963 220960
rect 142110 220902 158963 220904
rect 470550 220962 470610 221174
rect 481449 221232 485931 221234
rect 481449 221176 481454 221232
rect 481510 221176 485870 221232
rect 485926 221176 485931 221232
rect 481449 221174 485931 221176
rect 481449 221171 481515 221174
rect 485865 221171 485931 221174
rect 495249 221234 495315 221237
rect 499757 221234 499823 221237
rect 495249 221232 499823 221234
rect 495249 221176 495254 221232
rect 495310 221176 499762 221232
rect 499818 221176 499823 221232
rect 495249 221174 499823 221176
rect 495249 221171 495315 221174
rect 499757 221171 499823 221174
rect 499941 221234 500007 221237
rect 504725 221234 504791 221237
rect 499941 221232 504791 221234
rect 499941 221176 499946 221232
rect 500002 221176 504730 221232
rect 504786 221176 504791 221232
rect 499941 221174 504791 221176
rect 499941 221171 500007 221174
rect 504725 221171 504791 221174
rect 562317 221098 562383 221101
rect 564065 221098 564131 221101
rect 562317 221096 564131 221098
rect 562317 221040 562322 221096
rect 562378 221040 564070 221096
rect 564126 221040 564131 221096
rect 562317 221038 564131 221040
rect 562317 221035 562383 221038
rect 564065 221035 564131 221038
rect 675293 221098 675359 221101
rect 675293 221096 676292 221098
rect 675293 221040 675298 221096
rect 675354 221040 676292 221096
rect 675293 221038 676292 221040
rect 675293 221035 675359 221038
rect 491661 220962 491727 220965
rect 470550 220960 491727 220962
rect 470550 220904 491666 220960
rect 491722 220904 491727 220960
rect 470550 220902 491727 220904
rect 158897 220899 158963 220902
rect 491661 220899 491727 220902
rect 176561 220826 176627 220829
rect 181437 220826 181503 220829
rect 176561 220824 181503 220826
rect 176561 220768 176566 220824
rect 176622 220768 181442 220824
rect 181498 220768 181503 220824
rect 176561 220766 181503 220768
rect 176561 220763 176627 220766
rect 181437 220763 181503 220766
rect 199653 220826 199719 220829
rect 201953 220826 202019 220829
rect 199653 220824 202019 220826
rect 199653 220768 199658 220824
rect 199714 220768 201958 220824
rect 202014 220768 202019 220824
rect 199653 220766 202019 220768
rect 199653 220763 199719 220766
rect 201953 220763 202019 220766
rect 545757 220826 545823 220829
rect 549345 220826 549411 220829
rect 545757 220824 549411 220826
rect 545757 220768 545762 220824
rect 545818 220768 549350 220824
rect 549406 220768 549411 220824
rect 545757 220766 549411 220768
rect 545757 220763 545823 220766
rect 549345 220763 549411 220766
rect 560569 220826 560635 220829
rect 562133 220826 562199 220829
rect 572437 220826 572503 220829
rect 560569 220824 572503 220826
rect 560569 220768 560574 220824
rect 560630 220768 562138 220824
rect 562194 220768 572442 220824
rect 572498 220768 572503 220824
rect 560569 220766 572503 220768
rect 560569 220763 560635 220766
rect 562133 220763 562199 220766
rect 572437 220763 572503 220766
rect 572621 220826 572687 220829
rect 575105 220826 575171 220829
rect 572621 220824 575171 220826
rect 572621 220768 572626 220824
rect 572682 220768 575110 220824
rect 575166 220768 575171 220824
rect 572621 220766 575171 220768
rect 572621 220763 572687 220766
rect 575105 220763 575171 220766
rect 147673 220690 147739 220693
rect 152089 220690 152155 220693
rect 147673 220688 152155 220690
rect 147673 220632 147678 220688
rect 147734 220632 152094 220688
rect 152150 220632 152155 220688
rect 147673 220630 152155 220632
rect 147673 220627 147739 220630
rect 152089 220627 152155 220630
rect 156873 220690 156939 220693
rect 157793 220690 157859 220693
rect 192477 220690 192543 220693
rect 194041 220690 194107 220693
rect 156873 220688 157859 220690
rect 156873 220632 156878 220688
rect 156934 220632 157798 220688
rect 157854 220632 157859 220688
rect 156873 220630 157859 220632
rect 156873 220627 156939 220630
rect 157793 220627 157859 220630
rect 162166 220630 176026 220690
rect 130193 220418 130259 220421
rect 162166 220418 162226 220630
rect 175966 220554 176026 220630
rect 192477 220688 194107 220690
rect 192477 220632 192482 220688
rect 192538 220632 194046 220688
rect 194102 220632 194107 220688
rect 192477 220630 194107 220632
rect 192477 220627 192543 220630
rect 194041 220627 194107 220630
rect 485865 220690 485931 220693
rect 488533 220690 488599 220693
rect 485865 220688 488599 220690
rect 485865 220632 485870 220688
rect 485926 220632 488538 220688
rect 488594 220632 488599 220688
rect 675293 220690 675359 220693
rect 675293 220688 676292 220690
rect 562961 220656 563027 220659
rect 485865 220630 488599 220632
rect 485865 220627 485931 220630
rect 488533 220627 488599 220630
rect 562918 220654 563027 220656
rect 562918 220598 562966 220654
rect 563022 220598 563027 220654
rect 675293 220632 675298 220688
rect 675354 220632 676292 220688
rect 675293 220630 676292 220632
rect 675293 220627 675359 220630
rect 562918 220593 563027 220598
rect 177849 220554 177915 220557
rect 175966 220552 177915 220554
rect 175966 220496 177854 220552
rect 177910 220496 177915 220552
rect 175966 220494 177915 220496
rect 177849 220491 177915 220494
rect 495249 220554 495315 220557
rect 496813 220554 496879 220557
rect 495249 220552 496879 220554
rect 495249 220496 495254 220552
rect 495310 220496 496818 220552
rect 496874 220496 496879 220552
rect 495249 220494 496879 220496
rect 495249 220491 495315 220494
rect 496813 220491 496879 220494
rect 548149 220554 548215 220557
rect 548885 220554 548951 220557
rect 548149 220552 548951 220554
rect 548149 220496 548154 220552
rect 548210 220496 548890 220552
rect 548946 220496 548951 220552
rect 548149 220494 548951 220496
rect 548149 220491 548215 220494
rect 548885 220491 548951 220494
rect 554957 220554 555023 220557
rect 562918 220554 562978 220593
rect 554957 220552 562978 220554
rect 554957 220496 554962 220552
rect 555018 220496 562978 220552
rect 554957 220494 562978 220496
rect 572529 220554 572595 220557
rect 575841 220554 575907 220557
rect 572529 220552 575907 220554
rect 572529 220496 572534 220552
rect 572590 220496 575846 220552
rect 575902 220496 575907 220552
rect 572529 220494 575907 220496
rect 554957 220491 555023 220494
rect 572529 220491 572595 220494
rect 575841 220491 575907 220494
rect 130193 220416 162226 220418
rect 130193 220360 130198 220416
rect 130254 220360 162226 220416
rect 130193 220358 162226 220360
rect 165981 220418 166047 220421
rect 169017 220418 169083 220421
rect 165981 220416 169083 220418
rect 165981 220360 165986 220416
rect 166042 220360 169022 220416
rect 169078 220360 169083 220416
rect 165981 220358 169083 220360
rect 130193 220355 130259 220358
rect 165981 220355 166047 220358
rect 169017 220355 169083 220358
rect 173433 220418 173499 220421
rect 175825 220418 175891 220421
rect 173433 220416 175891 220418
rect 173433 220360 173438 220416
rect 173494 220360 175830 220416
rect 175886 220360 175891 220416
rect 173433 220358 175891 220360
rect 173433 220355 173499 220358
rect 175825 220355 175891 220358
rect 181161 220418 181227 220421
rect 189901 220418 189967 220421
rect 181161 220416 189967 220418
rect 181161 220360 181166 220416
rect 181222 220360 189906 220416
rect 189962 220360 189967 220416
rect 181161 220358 189967 220360
rect 181161 220355 181227 220358
rect 189901 220355 189967 220358
rect 449893 220418 449959 220421
rect 490281 220418 490347 220421
rect 572253 220418 572319 220421
rect 449893 220416 490347 220418
rect 449893 220360 449898 220416
rect 449954 220360 490286 220416
rect 490342 220360 490347 220416
rect 449893 220358 490347 220360
rect 449893 220355 449959 220358
rect 490281 220355 490347 220358
rect 563102 220416 572319 220418
rect 563102 220360 572258 220416
rect 572314 220360 572319 220416
rect 563102 220358 572319 220360
rect 511993 220282 512059 220285
rect 512637 220282 512703 220285
rect 563102 220282 563162 220358
rect 572253 220355 572319 220358
rect 511993 220280 563162 220282
rect 511993 220224 511998 220280
rect 512054 220224 512642 220280
rect 512698 220224 563162 220280
rect 511993 220222 563162 220224
rect 572437 220282 572503 220285
rect 576025 220282 576091 220285
rect 572437 220280 576091 220282
rect 572437 220224 572442 220280
rect 572498 220224 576030 220280
rect 576086 220224 576091 220280
rect 572437 220222 576091 220224
rect 511993 220219 512059 220222
rect 512637 220219 512703 220222
rect 572437 220219 572503 220222
rect 576025 220219 576091 220222
rect 674649 220282 674715 220285
rect 674649 220280 676292 220282
rect 674649 220224 674654 220280
rect 674710 220224 676292 220280
rect 674649 220222 676292 220224
rect 674649 220219 674715 220222
rect 150341 220146 150407 220149
rect 204345 220146 204411 220149
rect 150341 220144 204411 220146
rect 150341 220088 150346 220144
rect 150402 220088 204350 220144
rect 204406 220088 204411 220144
rect 150341 220086 204411 220088
rect 150341 220083 150407 220086
rect 204345 220083 204411 220086
rect 219341 220146 219407 220149
rect 220077 220146 220143 220149
rect 219341 220144 220143 220146
rect 219341 220088 219346 220144
rect 219402 220088 220082 220144
rect 220138 220088 220143 220144
rect 219341 220086 220143 220088
rect 219341 220083 219407 220086
rect 220077 220083 220143 220086
rect 442901 220146 442967 220149
rect 493317 220146 493383 220149
rect 442901 220144 493383 220146
rect 442901 220088 442906 220144
rect 442962 220088 493322 220144
rect 493378 220088 493383 220144
rect 442901 220086 493383 220088
rect 442901 220083 442967 220086
rect 493317 220083 493383 220086
rect 563240 220086 569970 220146
rect 56501 220010 56567 220013
rect 148041 220010 148107 220013
rect 56501 220008 148107 220010
rect 56501 219952 56506 220008
rect 56562 219952 148046 220008
rect 148102 219952 148107 220008
rect 56501 219950 148107 219952
rect 56501 219947 56567 219950
rect 148041 219947 148107 219950
rect 502333 220010 502399 220013
rect 503478 220010 503484 220012
rect 502333 220008 503484 220010
rect 502333 219952 502338 220008
rect 502394 219952 503484 220008
rect 502333 219950 503484 219952
rect 502333 219947 502399 219950
rect 503478 219948 503484 219950
rect 503548 219948 503554 220012
rect 525057 220010 525123 220013
rect 533521 220010 533587 220013
rect 563240 220010 563300 220086
rect 525057 220008 533354 220010
rect 525057 219952 525062 220008
rect 525118 219952 533354 220008
rect 525057 219950 533354 219952
rect 525057 219947 525123 219950
rect 171041 219874 171107 219877
rect 173249 219874 173315 219877
rect 171041 219872 173315 219874
rect 171041 219816 171046 219872
rect 171102 219816 173254 219872
rect 173310 219816 173315 219872
rect 171041 219814 173315 219816
rect 171041 219811 171107 219814
rect 173249 219811 173315 219814
rect 209681 219874 209747 219877
rect 209865 219874 209931 219877
rect 209681 219872 209931 219874
rect 209681 219816 209686 219872
rect 209742 219816 209870 219872
rect 209926 219816 209931 219872
rect 209681 219814 209931 219816
rect 209681 219811 209747 219814
rect 209865 219811 209931 219814
rect 505093 219874 505159 219877
rect 505093 219872 514770 219874
rect 505093 219816 505098 219872
rect 505154 219816 514770 219872
rect 505093 219814 514770 219816
rect 505093 219811 505159 219814
rect 143073 219738 143139 219741
rect 147765 219738 147831 219741
rect 143073 219736 147831 219738
rect 143073 219680 143078 219736
rect 143134 219680 147770 219736
rect 147826 219680 147831 219736
rect 143073 219678 147831 219680
rect 143073 219675 143139 219678
rect 147765 219675 147831 219678
rect 152825 219738 152891 219741
rect 154665 219738 154731 219741
rect 152825 219736 154731 219738
rect 152825 219680 152830 219736
rect 152886 219680 154670 219736
rect 154726 219680 154731 219736
rect 152825 219678 154731 219680
rect 152825 219675 152891 219678
rect 154665 219675 154731 219678
rect 202321 219738 202387 219741
rect 205909 219738 205975 219741
rect 202321 219736 205975 219738
rect 202321 219680 202326 219736
rect 202382 219680 205914 219736
rect 205970 219680 205975 219736
rect 202321 219678 205975 219680
rect 514710 219738 514770 219814
rect 533061 219738 533127 219741
rect 514710 219736 533127 219738
rect 514710 219680 533066 219736
rect 533122 219680 533127 219736
rect 514710 219678 533127 219680
rect 533294 219738 533354 219950
rect 533521 220008 563300 220010
rect 533521 219952 533526 220008
rect 533582 219952 563300 220008
rect 533521 219950 563300 219952
rect 569910 220010 569970 220086
rect 569910 219950 572730 220010
rect 533521 219947 533587 219950
rect 572437 219738 572503 219741
rect 533294 219736 572503 219738
rect 533294 219680 572442 219736
rect 572498 219680 572503 219736
rect 533294 219678 572503 219680
rect 572670 219738 572730 219950
rect 574134 219948 574140 220012
rect 574204 220010 574210 220012
rect 614021 220010 614087 220013
rect 574204 220008 614087 220010
rect 574204 219952 614026 220008
rect 614082 219952 614087 220008
rect 574204 219950 614087 219952
rect 574204 219948 574210 219950
rect 614021 219947 614087 219950
rect 675477 219874 675543 219877
rect 675477 219872 676292 219874
rect 675477 219816 675482 219872
rect 675538 219816 676292 219872
rect 675477 219814 676292 219816
rect 675477 219811 675543 219814
rect 614941 219738 615007 219741
rect 572670 219736 615007 219738
rect 572670 219680 614946 219736
rect 615002 219680 615007 219736
rect 572670 219678 615007 219680
rect 202321 219675 202387 219678
rect 205909 219675 205975 219678
rect 533061 219675 533127 219678
rect 572437 219675 572503 219678
rect 614941 219675 615007 219678
rect 142061 219602 142127 219605
rect 142245 219602 142311 219605
rect 142061 219600 142311 219602
rect 142061 219544 142066 219600
rect 142122 219544 142250 219600
rect 142306 219544 142311 219600
rect 142061 219542 142311 219544
rect 142061 219539 142127 219542
rect 142245 219539 142311 219542
rect 160921 219602 160987 219605
rect 165613 219602 165679 219605
rect 160921 219600 165679 219602
rect 160921 219544 160926 219600
rect 160982 219544 165618 219600
rect 165674 219544 165679 219600
rect 160921 219542 165679 219544
rect 160921 219539 160987 219542
rect 165613 219539 165679 219542
rect 180517 219602 180583 219605
rect 182173 219602 182239 219605
rect 180517 219600 182239 219602
rect 180517 219544 180522 219600
rect 180578 219544 182178 219600
rect 182234 219544 182239 219600
rect 180517 219542 182239 219544
rect 180517 219539 180583 219542
rect 182173 219539 182239 219542
rect 183277 219602 183343 219605
rect 187969 219602 188035 219605
rect 183277 219600 188035 219602
rect 183277 219544 183282 219600
rect 183338 219544 187974 219600
rect 188030 219544 188035 219600
rect 183277 219542 188035 219544
rect 183277 219539 183343 219542
rect 187969 219539 188035 219542
rect 474457 219602 474523 219605
rect 476573 219602 476639 219605
rect 474457 219600 476639 219602
rect 474457 219544 474462 219600
rect 474518 219544 476578 219600
rect 476634 219544 476639 219600
rect 474457 219542 476639 219544
rect 474457 219539 474523 219542
rect 476573 219539 476639 219542
rect 480345 219602 480411 219605
rect 485865 219602 485931 219605
rect 480345 219600 485931 219602
rect 480345 219544 480350 219600
rect 480406 219544 485870 219600
rect 485926 219544 485931 219600
rect 480345 219542 485931 219544
rect 480345 219539 480411 219542
rect 485865 219539 485931 219542
rect 204989 219466 205055 219469
rect 205633 219466 205699 219469
rect 204989 219464 205699 219466
rect 204989 219408 204994 219464
rect 205050 219408 205638 219464
rect 205694 219408 205699 219464
rect 204989 219406 205699 219408
rect 204989 219403 205055 219406
rect 205633 219403 205699 219406
rect 507761 219466 507827 219469
rect 615493 219466 615559 219469
rect 507761 219464 563070 219466
rect 507761 219408 507766 219464
rect 507822 219408 563070 219464
rect 507761 219406 563070 219408
rect 507761 219403 507827 219406
rect 563010 219364 563070 219406
rect 563240 219464 615559 219466
rect 563240 219408 615498 219464
rect 615554 219408 615559 219464
rect 563240 219406 615559 219408
rect 563240 219364 563300 219406
rect 615493 219403 615559 219406
rect 674465 219466 674531 219469
rect 674465 219464 676292 219466
rect 674465 219408 674470 219464
rect 674526 219408 676292 219464
rect 674465 219406 676292 219408
rect 674465 219403 674531 219406
rect 563010 219304 563300 219364
rect 542537 219194 542603 219197
rect 543457 219194 543523 219197
rect 542537 219192 543523 219194
rect 542537 219136 542542 219192
rect 542598 219136 543462 219192
rect 543518 219136 543523 219192
rect 542537 219134 543523 219136
rect 542537 219131 542603 219134
rect 543457 219131 543523 219134
rect 544377 219194 544443 219197
rect 552657 219194 552723 219197
rect 544377 219192 552723 219194
rect 544377 219136 544382 219192
rect 544438 219136 552662 219192
rect 552718 219136 552723 219192
rect 544377 219134 552723 219136
rect 544377 219131 544443 219134
rect 552657 219131 552723 219134
rect 553485 219194 553551 219197
rect 556981 219194 557047 219197
rect 553485 219192 557047 219194
rect 553485 219136 553490 219192
rect 553546 219136 556986 219192
rect 557042 219136 557047 219192
rect 553485 219134 557047 219136
rect 553485 219131 553551 219134
rect 556981 219131 557047 219134
rect 559782 219132 559788 219196
rect 559852 219194 559858 219196
rect 562501 219194 562567 219197
rect 559852 219192 562567 219194
rect 559852 219136 562506 219192
rect 562562 219136 562567 219192
rect 559852 219134 562567 219136
rect 559852 219132 559858 219134
rect 562501 219131 562567 219134
rect 563421 219194 563487 219197
rect 571926 219194 571932 219196
rect 563421 219192 571932 219194
rect 563421 219136 563426 219192
rect 563482 219136 571932 219192
rect 563421 219134 571932 219136
rect 563421 219131 563487 219134
rect 571926 219132 571932 219134
rect 571996 219132 572002 219196
rect 572161 219194 572227 219197
rect 573725 219194 573791 219197
rect 572161 219192 573791 219194
rect 572161 219136 572166 219192
rect 572222 219136 573730 219192
rect 573786 219136 573791 219192
rect 572161 219134 573791 219136
rect 572161 219131 572227 219134
rect 573725 219131 573791 219134
rect 675150 218996 675156 219060
rect 675220 219058 675226 219060
rect 675220 218998 676292 219058
rect 675220 218996 675226 218998
rect 535361 218922 535427 218925
rect 613377 218922 613443 218925
rect 535361 218920 613443 218922
rect 535361 218864 535366 218920
rect 535422 218864 613382 218920
rect 613438 218864 613443 218920
rect 535361 218862 613443 218864
rect 535361 218859 535427 218862
rect 613377 218859 613443 218862
rect 497457 218650 497523 218653
rect 631041 218650 631107 218653
rect 497457 218648 631107 218650
rect 497457 218592 497462 218648
rect 497518 218592 631046 218648
rect 631102 218592 631107 218648
rect 497457 218590 631107 218592
rect 497457 218587 497523 218590
rect 631041 218587 631107 218590
rect 675518 218588 675524 218652
rect 675588 218650 675594 218652
rect 675588 218590 676292 218650
rect 675588 218588 675594 218590
rect 494789 218378 494855 218381
rect 495065 218378 495131 218381
rect 574645 218378 574711 218381
rect 494789 218376 574711 218378
rect 494789 218320 494794 218376
rect 494850 218320 495070 218376
rect 495126 218320 574650 218376
rect 574706 218320 574711 218376
rect 494789 218318 574711 218320
rect 494789 218315 494855 218318
rect 495065 218315 495131 218318
rect 574645 218315 574711 218318
rect 674833 218242 674899 218245
rect 674833 218240 676292 218242
rect 674833 218184 674838 218240
rect 674894 218184 676292 218240
rect 674833 218182 676292 218184
rect 674833 218179 674899 218182
rect 490281 218106 490347 218109
rect 612273 218106 612339 218109
rect 490281 218104 612339 218106
rect 490281 218048 490286 218104
rect 490342 218048 612278 218104
rect 612334 218048 612339 218104
rect 490281 218046 612339 218048
rect 490281 218043 490347 218046
rect 612273 218043 612339 218046
rect 493317 217834 493383 217837
rect 504173 217834 504239 217837
rect 550633 217834 550699 217837
rect 556797 217834 556863 217837
rect 560109 217836 560175 217837
rect 560109 217834 560156 217836
rect 493317 217832 499590 217834
rect 493317 217776 493322 217832
rect 493378 217776 499590 217832
rect 493317 217774 499590 217776
rect 493317 217771 493383 217774
rect 499530 217562 499590 217774
rect 504173 217832 505110 217834
rect 504173 217776 504178 217832
rect 504234 217776 505110 217832
rect 504173 217774 505110 217776
rect 504173 217771 504239 217774
rect 505050 217562 505110 217774
rect 540930 217774 548626 217834
rect 540930 217562 540990 217774
rect 542077 217666 542143 217667
rect 542077 217664 542124 217666
rect 542032 217662 542124 217664
rect 542032 217606 542082 217662
rect 542032 217604 542124 217606
rect 542077 217602 542124 217604
rect 542188 217602 542194 217666
rect 542077 217601 542143 217602
rect 499530 217502 504466 217562
rect 505050 217502 540990 217562
rect 541157 217564 541223 217565
rect 542491 217564 542557 217565
rect 541157 217560 541204 217564
rect 541268 217562 541274 217564
rect 542486 217562 542492 217564
rect 541157 217504 541162 217560
rect 41505 217290 41571 217293
rect 42057 217290 42123 217293
rect 41505 217288 42123 217290
rect 41505 217232 41510 217288
rect 41566 217232 42062 217288
rect 42118 217232 42123 217288
rect 41505 217230 42123 217232
rect 41505 217227 41571 217230
rect 42057 217227 42123 217230
rect 488165 217290 488231 217293
rect 504173 217290 504239 217293
rect 488165 217288 504239 217290
rect 488165 217232 488170 217288
rect 488226 217232 504178 217288
rect 504234 217232 504239 217288
rect 488165 217230 504239 217232
rect 504406 217290 504466 217502
rect 541157 217500 541204 217504
rect 541268 217502 541314 217562
rect 542400 217502 542492 217562
rect 541268 217500 541274 217502
rect 542486 217500 542492 217502
rect 542556 217500 542562 217564
rect 542670 217500 542676 217564
rect 542740 217562 542746 217564
rect 543641 217562 543707 217565
rect 542740 217560 543707 217562
rect 542740 217504 543646 217560
rect 543702 217504 543707 217560
rect 542740 217502 543707 217504
rect 542740 217500 542746 217502
rect 541157 217499 541223 217500
rect 542491 217499 542557 217500
rect 543641 217499 543707 217502
rect 546125 217562 546191 217565
rect 547965 217562 548031 217565
rect 546125 217560 548031 217562
rect 546125 217504 546130 217560
rect 546186 217504 547970 217560
rect 548026 217504 548031 217560
rect 546125 217502 548031 217504
rect 548566 217562 548626 217774
rect 550633 217832 556863 217834
rect 550633 217776 550638 217832
rect 550694 217776 556802 217832
rect 556858 217776 556863 217832
rect 550633 217774 556863 217776
rect 560064 217832 560156 217834
rect 560064 217776 560114 217832
rect 560064 217774 560156 217776
rect 550633 217771 550699 217774
rect 556797 217771 556863 217774
rect 560109 217772 560156 217774
rect 560220 217772 560226 217836
rect 561029 217834 561095 217837
rect 563145 217834 563211 217837
rect 563421 217836 563487 217837
rect 563421 217834 563468 217836
rect 561029 217832 563211 217834
rect 561029 217776 561034 217832
rect 561090 217776 563150 217832
rect 563206 217776 563211 217832
rect 561029 217774 563211 217776
rect 563376 217832 563468 217834
rect 563376 217776 563426 217832
rect 563376 217774 563468 217776
rect 560109 217771 560175 217772
rect 561029 217771 561095 217774
rect 563145 217771 563211 217774
rect 563421 217772 563468 217774
rect 563532 217772 563538 217836
rect 563697 217834 563763 217837
rect 572621 217834 572687 217837
rect 563697 217832 572687 217834
rect 563697 217776 563702 217832
rect 563758 217776 572626 217832
rect 572682 217776 572687 217832
rect 563697 217774 572687 217776
rect 563421 217771 563487 217772
rect 563697 217771 563763 217774
rect 572621 217771 572687 217774
rect 572846 217772 572852 217836
rect 572916 217834 572922 217836
rect 574461 217834 574527 217837
rect 572916 217832 574527 217834
rect 572916 217776 574466 217832
rect 574522 217776 574527 217832
rect 572916 217774 574527 217776
rect 572916 217772 572922 217774
rect 574461 217771 574527 217774
rect 675334 217772 675340 217836
rect 675404 217834 675410 217836
rect 675404 217774 676292 217834
rect 675404 217772 675410 217774
rect 574461 217562 574527 217565
rect 548566 217560 574527 217562
rect 548566 217504 574466 217560
rect 574522 217504 574527 217560
rect 548566 217502 574527 217504
rect 546125 217499 546191 217502
rect 547965 217499 548031 217502
rect 574461 217499 574527 217502
rect 672625 217426 672691 217429
rect 673310 217426 673316 217428
rect 672625 217424 673316 217426
rect 672625 217368 672630 217424
rect 672686 217368 673316 217424
rect 672625 217366 673316 217368
rect 672625 217363 672691 217366
rect 673310 217364 673316 217366
rect 673380 217364 673386 217428
rect 675293 217426 675359 217429
rect 675293 217424 676292 217426
rect 675293 217368 675298 217424
rect 675354 217368 676292 217424
rect 675293 217366 676292 217368
rect 675293 217363 675359 217366
rect 612825 217290 612891 217293
rect 504406 217288 612891 217290
rect 504406 217232 612830 217288
rect 612886 217232 612891 217288
rect 504406 217230 612891 217232
rect 488165 217227 488231 217230
rect 504173 217227 504239 217230
rect 612825 217227 612891 217230
rect 485773 217018 485839 217021
rect 486877 217018 486943 217021
rect 611721 217018 611787 217021
rect 485773 217016 611787 217018
rect 485773 216960 485778 217016
rect 485834 216960 486882 217016
rect 486938 216960 611726 217016
rect 611782 216960 611787 217016
rect 485773 216958 611787 216960
rect 485773 216955 485839 216958
rect 486877 216955 486943 216958
rect 611721 216955 611787 216958
rect 675477 217018 675543 217021
rect 675477 217016 676292 217018
rect 675477 216960 675482 217016
rect 675538 216960 676292 217016
rect 675477 216958 676292 216960
rect 675477 216955 675543 216958
rect 40309 216746 40375 216749
rect 45277 216746 45343 216749
rect 40309 216744 45343 216746
rect 40309 216688 40314 216744
rect 40370 216688 45282 216744
rect 45338 216688 45343 216744
rect 40309 216686 45343 216688
rect 40309 216683 40375 216686
rect 45277 216683 45343 216686
rect 484853 216746 484919 216749
rect 631593 216746 631659 216749
rect 484853 216744 631659 216746
rect 484853 216688 484858 216744
rect 484914 216688 631598 216744
rect 631654 216688 631659 216744
rect 484853 216686 631659 216688
rect 484853 216683 484919 216686
rect 631593 216683 631659 216686
rect 675702 216548 675708 216612
rect 675772 216610 675778 216612
rect 675772 216550 676292 216610
rect 675772 216548 675778 216550
rect 513833 216474 513899 216477
rect 520641 216474 520707 216477
rect 513833 216472 520707 216474
rect 513833 216416 513838 216472
rect 513894 216416 520646 216472
rect 520702 216416 520707 216472
rect 513833 216414 520707 216416
rect 513833 216411 513899 216414
rect 520641 216411 520707 216414
rect 526069 216474 526135 216477
rect 531221 216474 531287 216477
rect 526069 216472 531287 216474
rect 526069 216416 526074 216472
rect 526130 216416 531226 216472
rect 531282 216416 531287 216472
rect 526069 216414 531287 216416
rect 526069 216411 526135 216414
rect 531221 216411 531287 216414
rect 537385 216474 537451 216477
rect 545665 216474 545731 216477
rect 546769 216476 546835 216477
rect 537385 216472 545731 216474
rect 537385 216416 537390 216472
rect 537446 216416 545670 216472
rect 545726 216416 545731 216472
rect 537385 216414 545731 216416
rect 537385 216411 537451 216414
rect 545665 216411 545731 216414
rect 546718 216412 546724 216476
rect 546788 216474 546835 216476
rect 549437 216474 549503 216477
rect 553945 216474 554011 216477
rect 546788 216472 546880 216474
rect 546830 216416 546880 216472
rect 546788 216414 546880 216416
rect 549437 216472 554011 216474
rect 549437 216416 549442 216472
rect 549498 216416 553950 216472
rect 554006 216416 554011 216472
rect 549437 216414 554011 216416
rect 546788 216412 546835 216414
rect 546769 216411 546835 216412
rect 549437 216411 549503 216414
rect 553945 216411 554011 216414
rect 556981 216474 557047 216477
rect 576761 216474 576827 216477
rect 556981 216472 576827 216474
rect 556981 216416 556986 216472
rect 557042 216416 576766 216472
rect 576822 216416 576827 216472
rect 556981 216414 576827 216416
rect 556981 216411 557047 216414
rect 576761 216411 576827 216414
rect 542486 216140 542492 216204
rect 542556 216202 542562 216204
rect 559782 216202 559788 216204
rect 542556 216142 559788 216202
rect 542556 216140 542562 216142
rect 559782 216140 559788 216142
rect 559852 216140 559858 216204
rect 560150 216140 560156 216204
rect 560220 216202 560226 216204
rect 574001 216202 574067 216205
rect 560220 216200 574067 216202
rect 560220 216144 574006 216200
rect 574062 216144 574067 216200
rect 560220 216142 574067 216144
rect 560220 216140 560226 216142
rect 574001 216139 574067 216142
rect 574461 216202 574527 216205
rect 575473 216202 575539 216205
rect 574461 216200 575539 216202
rect 574461 216144 574466 216200
rect 574522 216144 575478 216200
rect 575534 216144 575539 216200
rect 574461 216142 575539 216144
rect 574461 216139 574527 216142
rect 575473 216139 575539 216142
rect 675109 216202 675175 216205
rect 675109 216200 676292 216202
rect 675109 216144 675114 216200
rect 675170 216144 676292 216200
rect 675109 216142 676292 216144
rect 675109 216139 675175 216142
rect 578693 216066 578759 216069
rect 576350 216064 578759 216066
rect 576350 216008 578698 216064
rect 578754 216008 578759 216064
rect 576350 216006 578759 216008
rect 541198 215868 541204 215932
rect 541268 215930 541274 215932
rect 546718 215930 546724 215932
rect 541268 215870 546724 215930
rect 541268 215868 541274 215870
rect 546718 215868 546724 215870
rect 546788 215868 546794 215932
rect 563462 215868 563468 215932
rect 563532 215930 563538 215932
rect 574553 215930 574619 215933
rect 563532 215928 574619 215930
rect 563532 215872 574558 215928
rect 574614 215872 574619 215928
rect 563532 215870 574619 215872
rect 563532 215868 563538 215870
rect 574553 215867 574619 215870
rect 576350 215764 576410 216006
rect 578693 216003 578759 216006
rect 596265 215930 596331 215933
rect 600497 215930 600563 215933
rect 596265 215928 600563 215930
rect 596265 215872 596270 215928
rect 596326 215872 600502 215928
rect 600558 215872 600563 215928
rect 596265 215870 600563 215872
rect 596265 215867 596331 215870
rect 600497 215867 600563 215870
rect 576577 215794 576643 215797
rect 595805 215794 595871 215797
rect 576577 215792 595871 215794
rect 576577 215736 576582 215792
rect 576638 215736 595810 215792
rect 595866 215736 595871 215792
rect 576577 215734 595871 215736
rect 576577 215731 576643 215734
rect 595805 215731 595871 215734
rect 675477 215794 675543 215797
rect 675477 215792 676292 215794
rect 675477 215736 675482 215792
rect 675538 215736 676292 215792
rect 675477 215734 676292 215736
rect 675477 215731 675543 215734
rect 595989 215658 596055 215661
rect 596633 215658 596699 215661
rect 595989 215656 596699 215658
rect 595989 215600 595994 215656
rect 596050 215600 596638 215656
rect 596694 215600 596699 215656
rect 595989 215598 596699 215600
rect 595989 215595 596055 215598
rect 596633 215595 596699 215598
rect 673494 215596 673500 215660
rect 673564 215658 673570 215660
rect 673913 215658 673979 215661
rect 673564 215656 673979 215658
rect 673564 215600 673918 215656
rect 673974 215600 673979 215656
rect 673564 215598 673979 215600
rect 673564 215596 673570 215598
rect 673913 215595 673979 215598
rect 586697 215522 586763 215525
rect 586470 215520 586763 215522
rect 586470 215464 586702 215520
rect 586758 215464 586763 215520
rect 586470 215462 586763 215464
rect 576025 215386 576091 215389
rect 586470 215386 586530 215462
rect 586697 215459 586763 215462
rect 673729 215388 673795 215389
rect 673678 215386 673684 215388
rect 576025 215384 586530 215386
rect 576025 215328 576030 215384
rect 576086 215328 586530 215384
rect 576025 215326 586530 215328
rect 673638 215326 673684 215386
rect 673748 215384 673795 215388
rect 673790 215328 673795 215384
rect 576025 215323 576091 215326
rect 673678 215324 673684 215326
rect 673748 215324 673795 215328
rect 673729 215323 673795 215324
rect 675293 215386 675359 215389
rect 675293 215384 676292 215386
rect 675293 215328 675298 215384
rect 675354 215328 676292 215384
rect 675293 215326 676292 215328
rect 675293 215323 675359 215326
rect 586605 215250 586671 215253
rect 594057 215250 594123 215253
rect 586605 215248 594123 215250
rect 586605 215192 586610 215248
rect 586666 215192 594062 215248
rect 594118 215192 594123 215248
rect 586605 215190 594123 215192
rect 586605 215187 586671 215190
rect 594057 215187 594123 215190
rect 35801 215114 35867 215117
rect 35758 215112 35867 215114
rect 35758 215056 35806 215112
rect 35862 215056 35867 215112
rect 35758 215051 35867 215056
rect 41505 215114 41571 215117
rect 43161 215114 43227 215117
rect 41505 215112 43227 215114
rect 41505 215056 41510 215112
rect 41566 215056 43166 215112
rect 43222 215056 43227 215112
rect 41505 215054 43227 215056
rect 41505 215051 41571 215054
rect 43161 215051 43227 215054
rect 35758 214948 35818 215051
rect 675886 214916 675892 214980
rect 675956 214978 675962 214980
rect 675956 214918 676292 214978
rect 675956 214916 675962 214918
rect 673085 214572 673151 214573
rect 673085 214568 673132 214572
rect 673196 214570 673202 214572
rect 35758 214301 35818 214540
rect 673085 214512 673090 214568
rect 673085 214508 673132 214512
rect 673196 214510 673242 214570
rect 673196 214508 673202 214510
rect 675886 214508 675892 214572
rect 675956 214570 675962 214572
rect 675956 214510 676292 214570
rect 675956 214508 675962 214510
rect 673085 214507 673151 214508
rect 33041 214298 33107 214301
rect 32998 214296 33107 214298
rect 32998 214240 33046 214296
rect 33102 214240 33107 214296
rect 32998 214235 33107 214240
rect 35758 214296 35867 214301
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214238 35867 214240
rect 35801 214235 35867 214238
rect 39941 214298 40007 214301
rect 43621 214298 43687 214301
rect 579245 214298 579311 214301
rect 39941 214296 43687 214298
rect 39941 214240 39946 214296
rect 40002 214240 43626 214296
rect 43682 214240 43687 214296
rect 39941 214238 43687 214240
rect 576380 214296 579311 214298
rect 576380 214240 579250 214296
rect 579306 214240 579311 214296
rect 576380 214238 579311 214240
rect 39941 214235 40007 214238
rect 43621 214235 43687 214238
rect 579245 214235 579311 214238
rect 32998 214132 33058 214235
rect 675477 214162 675543 214165
rect 675477 214160 676292 214162
rect 675477 214104 675482 214160
rect 675538 214104 676292 214160
rect 675477 214102 676292 214104
rect 675477 214099 675543 214102
rect 39941 213890 40007 213893
rect 45001 213890 45067 213893
rect 39941 213888 45067 213890
rect 39941 213832 39946 213888
rect 40002 213832 45006 213888
rect 45062 213832 45067 213888
rect 39941 213830 45067 213832
rect 39941 213827 40007 213830
rect 45001 213827 45067 213830
rect 675477 213754 675543 213757
rect 675477 213752 676292 213754
rect 35390 213485 35450 213724
rect 675477 213696 675482 213752
rect 675538 213696 676292 213752
rect 675477 213694 676292 213696
rect 675477 213691 675543 213694
rect 35390 213480 35499 213485
rect 35390 213424 35438 213480
rect 35494 213424 35499 213480
rect 35390 213422 35499 213424
rect 35433 213419 35499 213422
rect 675477 213346 675543 213349
rect 675477 213344 676292 213346
rect 35574 213077 35634 213316
rect 675477 213288 675482 213344
rect 675538 213288 676292 213344
rect 675477 213286 676292 213288
rect 675477 213283 675543 213286
rect 35574 213072 35683 213077
rect 35574 213016 35622 213072
rect 35678 213016 35683 213072
rect 35574 213014 35683 213016
rect 35617 213011 35683 213014
rect 35758 212669 35818 212908
rect 578509 212802 578575 212805
rect 576380 212800 578575 212802
rect 576380 212744 578514 212800
rect 578570 212744 578575 212800
rect 576380 212742 578575 212744
rect 578509 212739 578575 212742
rect 28533 212666 28599 212669
rect 28533 212664 28642 212666
rect 28533 212608 28538 212664
rect 28594 212608 28642 212664
rect 28533 212603 28642 212608
rect 35758 212664 35867 212669
rect 35758 212608 35806 212664
rect 35862 212608 35867 212664
rect 35758 212606 35867 212608
rect 35801 212603 35867 212606
rect 670734 212604 670740 212668
rect 670804 212666 670810 212668
rect 671061 212666 671127 212669
rect 670804 212664 671127 212666
rect 670804 212608 671066 212664
rect 671122 212608 671127 212664
rect 670804 212606 671127 212608
rect 670804 212604 670810 212606
rect 671061 212603 671127 212606
rect 28582 212500 28642 212603
rect 683070 212533 683130 212908
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 683113 212467 683179 212470
rect 40953 212258 41019 212261
rect 43345 212258 43411 212261
rect 40953 212256 43411 212258
rect 40953 212200 40958 212256
rect 41014 212200 43350 212256
rect 43406 212200 43411 212256
rect 40953 212198 43411 212200
rect 40953 212195 41019 212198
rect 43345 212195 43411 212198
rect 675477 212122 675543 212125
rect 675477 212120 676292 212122
rect 35758 211853 35818 212092
rect 675477 212064 675482 212120
rect 675538 212064 676292 212120
rect 675477 212062 676292 212064
rect 675477 212059 675543 212062
rect 35758 211848 35867 211853
rect 35758 211792 35806 211848
rect 35862 211792 35867 211848
rect 35758 211790 35867 211792
rect 35801 211787 35867 211790
rect 35574 211445 35634 211684
rect 35574 211440 35683 211445
rect 35574 211384 35622 211440
rect 35678 211384 35683 211440
rect 35574 211382 35683 211384
rect 35617 211379 35683 211382
rect 39665 211442 39731 211445
rect 42885 211442 42951 211445
rect 39665 211440 42951 211442
rect 39665 211384 39670 211440
rect 39726 211384 42890 211440
rect 42946 211384 42951 211440
rect 39665 211382 42951 211384
rect 39665 211379 39731 211382
rect 42885 211379 42951 211382
rect 35758 211037 35818 211276
rect 576380 211246 576870 211306
rect 576810 211170 576870 211246
rect 578877 211170 578943 211173
rect 576810 211168 578943 211170
rect 576810 211112 578882 211168
rect 578938 211112 578943 211168
rect 576810 211110 578943 211112
rect 578877 211107 578943 211110
rect 35758 211032 35867 211037
rect 35758 210976 35806 211032
rect 35862 210976 35867 211032
rect 35758 210974 35867 210976
rect 35801 210971 35867 210974
rect 41505 211034 41571 211037
rect 42333 211034 42399 211037
rect 41505 211032 42399 211034
rect 41505 210976 41510 211032
rect 41566 210976 42338 211032
rect 42394 210976 42399 211032
rect 41505 210974 42399 210976
rect 41505 210971 41571 210974
rect 42333 210971 42399 210974
rect 35574 210629 35634 210868
rect 35574 210624 35683 210629
rect 35574 210568 35622 210624
rect 35678 210568 35683 210624
rect 35574 210566 35683 210568
rect 35617 210563 35683 210566
rect 670877 210492 670943 210493
rect 670877 210490 670924 210492
rect 670832 210488 670924 210490
rect 35758 210221 35818 210460
rect 670832 210432 670882 210488
rect 670832 210430 670924 210432
rect 670877 210428 670924 210430
rect 670988 210428 670994 210492
rect 670877 210427 670943 210428
rect 35758 210216 35867 210221
rect 35758 210160 35806 210216
rect 35862 210160 35867 210216
rect 35758 210158 35867 210160
rect 35801 210155 35867 210158
rect 675150 210156 675156 210220
rect 675220 210218 675226 210220
rect 675886 210218 675892 210220
rect 675220 210158 675892 210218
rect 675220 210156 675226 210158
rect 675886 210156 675892 210158
rect 675956 210156 675962 210220
rect 41822 210082 41828 210084
rect 41492 210022 41828 210082
rect 41822 210020 41828 210022
rect 41892 210020 41898 210084
rect 669313 209946 669379 209949
rect 675845 209946 675911 209949
rect 669313 209944 675911 209946
rect 669313 209888 669318 209944
rect 669374 209888 675850 209944
rect 675906 209888 675911 209944
rect 669313 209886 675911 209888
rect 669313 209883 669379 209886
rect 675845 209883 675911 209886
rect 579245 209810 579311 209813
rect 576380 209808 579311 209810
rect 576380 209752 579250 209808
rect 579306 209752 579311 209808
rect 576380 209750 579311 209752
rect 579245 209747 579311 209750
rect 35758 209405 35818 209644
rect 669814 209612 669820 209676
rect 669884 209674 669890 209676
rect 670785 209674 670851 209677
rect 669884 209672 670851 209674
rect 669884 209616 670790 209672
rect 670846 209616 670851 209672
rect 669884 209614 670851 209616
rect 669884 209612 669890 209614
rect 670785 209611 670851 209614
rect 35758 209400 35867 209405
rect 35758 209344 35806 209400
rect 35862 209344 35867 209400
rect 35758 209342 35867 209344
rect 35801 209339 35867 209342
rect 30238 208997 30298 209236
rect 30238 208992 30347 208997
rect 30238 208936 30286 208992
rect 30342 208936 30347 208992
rect 30238 208934 30347 208936
rect 30281 208931 30347 208934
rect 40033 208994 40099 208997
rect 41454 208994 41460 208996
rect 40033 208992 41460 208994
rect 40033 208936 40038 208992
rect 40094 208936 41460 208992
rect 40033 208934 41460 208936
rect 40033 208931 40099 208934
rect 41454 208932 41460 208934
rect 41524 208932 41530 208996
rect 35758 208589 35818 208828
rect 665582 208796 665588 208860
rect 665652 208858 665658 208860
rect 665652 208798 666570 208858
rect 665652 208796 665658 208798
rect 35758 208584 35867 208589
rect 35758 208528 35806 208584
rect 35862 208528 35867 208584
rect 35758 208526 35867 208528
rect 35801 208523 35867 208526
rect 40910 208180 40970 208420
rect 578417 208314 578483 208317
rect 576380 208312 578483 208314
rect 576380 208256 578422 208312
rect 578478 208256 578483 208312
rect 576380 208254 578483 208256
rect 578417 208251 578483 208254
rect 40902 208116 40908 208180
rect 40972 208116 40978 208180
rect 589457 208178 589523 208181
rect 589457 208176 592050 208178
rect 589457 208120 589462 208176
rect 589518 208120 592050 208176
rect 589457 208118 592050 208120
rect 589457 208115 589523 208118
rect 591990 208110 592050 208118
rect 591990 208050 592572 208110
rect 40542 207772 40602 208012
rect 40534 207708 40540 207772
rect 40604 207708 40610 207772
rect 35574 207365 35634 207604
rect 666510 207498 666570 208798
rect 669589 208316 669655 208317
rect 669589 208312 669636 208316
rect 669700 208314 669706 208316
rect 669589 208256 669594 208312
rect 669589 208252 669636 208256
rect 669700 208254 669746 208314
rect 669700 208252 669706 208254
rect 669589 208251 669655 208252
rect 666510 207438 666754 207498
rect 35525 207360 35634 207365
rect 35801 207362 35867 207365
rect 35525 207304 35530 207360
rect 35586 207304 35634 207360
rect 35525 207302 35634 207304
rect 35758 207360 35867 207362
rect 35758 207304 35806 207360
rect 35862 207304 35867 207360
rect 35525 207299 35591 207302
rect 35758 207299 35867 207304
rect 35758 207196 35818 207299
rect 666694 207226 666754 207438
rect 666356 207166 666754 207226
rect 40125 206954 40191 206957
rect 42885 206954 42951 206957
rect 40125 206952 42951 206954
rect 40125 206896 40130 206952
rect 40186 206896 42890 206952
rect 42946 206896 42951 206952
rect 40125 206894 42951 206896
rect 40125 206891 40191 206894
rect 42885 206891 42951 206894
rect 578693 206818 578759 206821
rect 576380 206816 578759 206818
rect 35758 206549 35818 206788
rect 576380 206760 578698 206816
rect 578754 206760 578759 206816
rect 576380 206758 578759 206760
rect 578693 206755 578759 206758
rect 35758 206544 35867 206549
rect 35758 206488 35806 206544
rect 35862 206488 35867 206544
rect 35758 206486 35867 206488
rect 35801 206483 35867 206486
rect 589457 206546 589523 206549
rect 589457 206544 592050 206546
rect 589457 206488 589462 206544
rect 589518 206488 592050 206544
rect 589457 206486 592050 206488
rect 589457 206483 589523 206486
rect 591990 206478 592050 206486
rect 591990 206418 592572 206478
rect 40726 206140 40786 206380
rect 40718 206076 40724 206140
rect 40788 206076 40794 206140
rect 35758 205733 35818 205972
rect 35758 205728 35867 205733
rect 35758 205672 35806 205728
rect 35862 205672 35867 205728
rect 35758 205670 35867 205672
rect 35801 205667 35867 205670
rect 39941 205730 40007 205733
rect 44173 205730 44239 205733
rect 39941 205728 44239 205730
rect 39941 205672 39946 205728
rect 40002 205672 44178 205728
rect 44234 205672 44239 205728
rect 39941 205670 44239 205672
rect 39941 205667 40007 205670
rect 44173 205667 44239 205670
rect 35574 205325 35634 205564
rect 669262 205396 669268 205460
rect 669332 205458 669338 205460
rect 669630 205458 669636 205460
rect 669332 205398 669636 205458
rect 669332 205396 669338 205398
rect 669630 205396 669636 205398
rect 669700 205396 669706 205460
rect 35574 205320 35683 205325
rect 35574 205264 35622 205320
rect 35678 205264 35683 205320
rect 35574 205262 35683 205264
rect 35617 205259 35683 205262
rect 40953 205322 41019 205325
rect 43253 205322 43319 205325
rect 579061 205322 579127 205325
rect 40953 205320 43319 205322
rect 40953 205264 40958 205320
rect 41014 205264 43258 205320
rect 43314 205264 43319 205320
rect 40953 205262 43319 205264
rect 576380 205320 579127 205322
rect 576380 205264 579066 205320
rect 579122 205264 579127 205320
rect 576380 205262 579127 205264
rect 40953 205259 41019 205262
rect 43253 205259 43319 205262
rect 579061 205259 579127 205262
rect 35758 204917 35818 205156
rect 675753 205050 675819 205053
rect 676254 205050 676260 205052
rect 675753 205048 676260 205050
rect 675753 204992 675758 205048
rect 675814 204992 676260 205048
rect 675753 204990 676260 204992
rect 675753 204987 675819 204990
rect 676254 204988 676260 204990
rect 676324 204988 676330 205052
rect 35758 204912 35867 204917
rect 35758 204856 35806 204912
rect 35862 204856 35867 204912
rect 35758 204854 35867 204856
rect 35801 204851 35867 204854
rect 589457 204914 589523 204917
rect 589457 204912 592050 204914
rect 589457 204856 589462 204912
rect 589518 204856 592050 204912
rect 589457 204854 592050 204856
rect 589457 204851 589523 204854
rect 591990 204846 592050 204854
rect 591990 204786 592572 204846
rect 35574 204509 35634 204748
rect 35525 204504 35634 204509
rect 35801 204506 35867 204509
rect 35525 204448 35530 204504
rect 35586 204448 35634 204504
rect 35525 204446 35634 204448
rect 35758 204504 35867 204506
rect 35758 204448 35806 204504
rect 35862 204448 35867 204504
rect 35525 204443 35591 204446
rect 35758 204443 35867 204448
rect 40769 204506 40835 204509
rect 44541 204506 44607 204509
rect 40769 204504 44607 204506
rect 40769 204448 40774 204504
rect 40830 204448 44546 204504
rect 44602 204448 44607 204504
rect 40769 204446 44607 204448
rect 40769 204443 40835 204446
rect 44541 204443 44607 204446
rect 35758 204340 35818 204443
rect 666502 204172 666508 204236
rect 666572 204234 666578 204236
rect 675661 204234 675727 204237
rect 675886 204234 675892 204236
rect 666572 204174 666754 204234
rect 666572 204172 666578 204174
rect 39757 204098 39823 204101
rect 43805 204098 43871 204101
rect 39757 204096 43871 204098
rect 39757 204040 39762 204096
rect 39818 204040 43810 204096
rect 43866 204040 43871 204096
rect 39757 204038 43871 204040
rect 39757 204035 39823 204038
rect 43805 204035 43871 204038
rect 666694 203962 666754 204174
rect 675661 204232 675892 204234
rect 675661 204176 675666 204232
rect 675722 204176 675892 204232
rect 675661 204174 675892 204176
rect 675661 204171 675727 204174
rect 675886 204172 675892 204174
rect 675956 204172 675962 204236
rect 35574 203693 35634 203932
rect 666356 203902 666754 203962
rect 578693 203826 578759 203829
rect 576380 203824 578759 203826
rect 576380 203768 578698 203824
rect 578754 203768 578759 203824
rect 576380 203766 578759 203768
rect 578693 203763 578759 203766
rect 35574 203688 35683 203693
rect 35574 203632 35622 203688
rect 35678 203632 35683 203688
rect 35574 203630 35683 203632
rect 35617 203627 35683 203630
rect 35758 203285 35818 203524
rect 35758 203280 35867 203285
rect 35758 203224 35806 203280
rect 35862 203224 35867 203280
rect 35758 203222 35867 203224
rect 35801 203219 35867 203222
rect 40033 203282 40099 203285
rect 47577 203282 47643 203285
rect 40033 203280 47643 203282
rect 40033 203224 40038 203280
rect 40094 203224 47582 203280
rect 47638 203224 47643 203280
rect 40033 203222 47643 203224
rect 40033 203219 40099 203222
rect 47577 203219 47643 203222
rect 589457 203282 589523 203285
rect 589457 203280 592050 203282
rect 589457 203224 589462 203280
rect 589518 203224 592050 203280
rect 589457 203222 592050 203224
rect 589457 203219 589523 203222
rect 591990 203214 592050 203222
rect 591990 203154 592572 203214
rect 41781 203010 41847 203013
rect 43621 203010 43687 203013
rect 41781 203008 43687 203010
rect 41781 202952 41786 203008
rect 41842 202952 43626 203008
rect 43682 202952 43687 203008
rect 41781 202950 43687 202952
rect 41781 202947 41847 202950
rect 43621 202947 43687 202950
rect 675385 202740 675451 202741
rect 675334 202738 675340 202740
rect 675294 202678 675340 202738
rect 675404 202736 675451 202740
rect 675446 202680 675451 202736
rect 675334 202676 675340 202678
rect 675404 202676 675451 202680
rect 675385 202675 675451 202676
rect 578233 202330 578299 202333
rect 668158 202330 668164 202332
rect 576380 202328 578299 202330
rect 576380 202272 578238 202328
rect 578294 202272 578299 202328
rect 576380 202270 578299 202272
rect 666356 202270 668164 202330
rect 578233 202267 578299 202270
rect 668158 202268 668164 202270
rect 668228 202268 668234 202332
rect 30281 202194 30347 202197
rect 41638 202194 41644 202196
rect 30281 202192 41644 202194
rect 30281 202136 30286 202192
rect 30342 202136 41644 202192
rect 30281 202134 41644 202136
rect 30281 202131 30347 202134
rect 41638 202132 41644 202134
rect 41708 202132 41714 202196
rect 589365 201650 589431 201653
rect 589365 201648 592050 201650
rect 589365 201592 589370 201648
rect 589426 201592 592050 201648
rect 589365 201590 592050 201592
rect 589365 201587 589431 201590
rect 591990 201582 592050 201590
rect 591990 201522 592572 201582
rect 578509 200834 578575 200837
rect 576380 200832 578575 200834
rect 576380 200776 578514 200832
rect 578570 200776 578575 200832
rect 576380 200774 578575 200776
rect 578509 200771 578575 200774
rect 673269 200834 673335 200837
rect 674782 200834 674788 200836
rect 673269 200832 674788 200834
rect 673269 200776 673274 200832
rect 673330 200776 674788 200832
rect 673269 200774 674788 200776
rect 673269 200771 673335 200774
rect 674782 200772 674788 200774
rect 674852 200772 674858 200836
rect 589457 200018 589523 200021
rect 675753 200018 675819 200021
rect 676438 200018 676444 200020
rect 589457 200016 592050 200018
rect 589457 199960 589462 200016
rect 589518 199960 592050 200016
rect 589457 199958 592050 199960
rect 589457 199955 589523 199958
rect 591990 199950 592050 199958
rect 675753 200016 676444 200018
rect 675753 199960 675758 200016
rect 675814 199960 676444 200016
rect 675753 199958 676444 199960
rect 675753 199955 675819 199958
rect 676438 199956 676444 199958
rect 676508 199956 676514 200020
rect 591990 199890 592572 199950
rect 578877 199338 578943 199341
rect 576380 199336 578943 199338
rect 576380 199280 578882 199336
rect 578938 199280 578943 199336
rect 576380 199278 578943 199280
rect 578877 199275 578943 199278
rect 666502 199276 666508 199340
rect 666572 199338 666578 199340
rect 666572 199278 666754 199338
rect 666572 199276 666578 199278
rect 666694 199134 666754 199278
rect 666356 199074 666754 199134
rect 674465 198658 674531 198661
rect 676806 198658 676812 198660
rect 674465 198656 676812 198658
rect 674465 198600 674470 198656
rect 674526 198600 676812 198656
rect 674465 198598 676812 198600
rect 674465 198595 674531 198598
rect 676806 198596 676812 198598
rect 676876 198596 676882 198660
rect 590377 198386 590443 198389
rect 590377 198384 592050 198386
rect 590377 198328 590382 198384
rect 590438 198328 592050 198384
rect 590377 198326 592050 198328
rect 590377 198323 590443 198326
rect 591990 198318 592050 198326
rect 591990 198258 592572 198318
rect 578325 197842 578391 197845
rect 576380 197840 578391 197842
rect 576380 197784 578330 197840
rect 578386 197784 578391 197840
rect 576380 197782 578391 197784
rect 578325 197779 578391 197782
rect 668209 197434 668275 197437
rect 666356 197432 668275 197434
rect 666356 197376 668214 197432
rect 668270 197376 668275 197432
rect 666356 197374 668275 197376
rect 668209 197371 668275 197374
rect 40902 197100 40908 197164
rect 40972 197162 40978 197164
rect 41781 197162 41847 197165
rect 40972 197160 41847 197162
rect 40972 197104 41786 197160
rect 41842 197104 41847 197160
rect 40972 197102 41847 197104
rect 40972 197100 40978 197102
rect 41781 197099 41847 197102
rect 675753 197162 675819 197165
rect 676622 197162 676628 197164
rect 675753 197160 676628 197162
rect 675753 197104 675758 197160
rect 675814 197104 676628 197160
rect 675753 197102 676628 197104
rect 675753 197099 675819 197102
rect 676622 197100 676628 197102
rect 676692 197100 676698 197164
rect 589457 196754 589523 196757
rect 589457 196752 592050 196754
rect 589457 196696 589462 196752
rect 589518 196696 592050 196752
rect 589457 196694 592050 196696
rect 589457 196691 589523 196694
rect 591990 196686 592050 196694
rect 591990 196626 592572 196686
rect 579245 196346 579311 196349
rect 576380 196344 579311 196346
rect 576380 196288 579250 196344
rect 579306 196288 579311 196344
rect 576380 196286 579311 196288
rect 579245 196283 579311 196286
rect 669262 196148 669268 196212
rect 669332 196210 669338 196212
rect 669630 196210 669636 196212
rect 669332 196150 669636 196210
rect 669332 196148 669338 196150
rect 669630 196148 669636 196150
rect 669700 196148 669706 196212
rect 669262 195876 669268 195940
rect 669332 195938 669338 195940
rect 669630 195938 669636 195940
rect 669332 195878 669636 195938
rect 669332 195876 669338 195878
rect 669630 195876 669636 195878
rect 669700 195876 669706 195940
rect 41781 195260 41847 195261
rect 41781 195256 41828 195260
rect 41892 195258 41898 195260
rect 41781 195200 41786 195256
rect 41781 195196 41828 195200
rect 41892 195198 41938 195258
rect 41892 195196 41898 195198
rect 41781 195195 41847 195196
rect 589457 195122 589523 195125
rect 589457 195120 592050 195122
rect 589457 195064 589462 195120
rect 589518 195064 592050 195120
rect 589457 195062 592050 195064
rect 589457 195059 589523 195062
rect 591990 195054 592050 195062
rect 591990 194994 592572 195054
rect 578877 194850 578943 194853
rect 576380 194848 578943 194850
rect 576380 194792 578882 194848
rect 578938 194792 578943 194848
rect 576380 194790 578943 194792
rect 578877 194787 578943 194790
rect 667974 194170 667980 194172
rect 666356 194110 667980 194170
rect 667974 194108 667980 194110
rect 668044 194108 668050 194172
rect 670601 193626 670667 193629
rect 675518 193626 675524 193628
rect 670601 193624 675524 193626
rect 670601 193568 670606 193624
rect 670662 193568 675524 193624
rect 670601 193566 675524 193568
rect 670601 193563 670667 193566
rect 675518 193564 675524 193566
rect 675588 193564 675594 193628
rect 578509 193490 578575 193493
rect 576350 193488 578575 193490
rect 576350 193432 578514 193488
rect 578570 193432 578575 193488
rect 576350 193430 578575 193432
rect 576350 193324 576410 193430
rect 578509 193427 578575 193430
rect 589457 193490 589523 193493
rect 589457 193488 592050 193490
rect 589457 193432 589462 193488
rect 589518 193432 592050 193488
rect 589457 193430 592050 193432
rect 589457 193427 589523 193430
rect 591990 193422 592050 193430
rect 591990 193362 592572 193422
rect 675753 193218 675819 193221
rect 676070 193218 676076 193220
rect 675753 193216 676076 193218
rect 675753 193160 675758 193216
rect 675814 193160 676076 193216
rect 675753 193158 676076 193160
rect 675753 193155 675819 193158
rect 676070 193156 676076 193158
rect 676140 193156 676146 193220
rect 666870 192606 666876 192608
rect 666356 192546 666876 192606
rect 666870 192544 666876 192546
rect 666940 192544 666946 192608
rect 579521 191858 579587 191861
rect 576380 191856 579587 191858
rect 576380 191800 579526 191856
rect 579582 191800 579587 191856
rect 576380 191798 579587 191800
rect 579521 191795 579587 191798
rect 591990 191730 592572 191790
rect 589641 191722 589707 191725
rect 591990 191722 592050 191730
rect 589641 191720 592050 191722
rect 589641 191664 589646 191720
rect 589702 191664 592050 191720
rect 589641 191662 592050 191664
rect 589641 191659 589707 191662
rect 40718 191524 40724 191588
rect 40788 191586 40794 191588
rect 41781 191586 41847 191589
rect 40788 191584 41847 191586
rect 40788 191528 41786 191584
rect 41842 191528 41847 191584
rect 40788 191526 41847 191528
rect 40788 191524 40794 191526
rect 41781 191523 41847 191526
rect 675477 191588 675543 191589
rect 675477 191584 675524 191588
rect 675588 191586 675594 191588
rect 675477 191528 675482 191584
rect 675477 191524 675524 191528
rect 675588 191526 675634 191586
rect 675588 191524 675594 191526
rect 675477 191523 675543 191524
rect 578233 190362 578299 190365
rect 576380 190360 578299 190362
rect 576380 190304 578238 190360
rect 578294 190304 578299 190360
rect 576380 190302 578299 190304
rect 578233 190299 578299 190302
rect 589457 190226 589523 190229
rect 589457 190224 592050 190226
rect 589457 190168 589462 190224
rect 589518 190168 592050 190224
rect 589457 190166 592050 190168
rect 589457 190163 589523 190166
rect 591990 190158 592050 190166
rect 591990 190098 592572 190158
rect 666686 189342 666692 189344
rect 666356 189282 666692 189342
rect 666686 189280 666692 189282
rect 666756 189280 666762 189344
rect 579245 188866 579311 188869
rect 576380 188864 579311 188866
rect 576380 188808 579250 188864
rect 579306 188808 579311 188864
rect 576380 188806 579311 188808
rect 579245 188803 579311 188806
rect 589457 188594 589523 188597
rect 589457 188592 592050 188594
rect 589457 188536 589462 188592
rect 589518 188536 592050 188592
rect 589457 188534 592050 188536
rect 589457 188531 589523 188534
rect 591990 188526 592050 188534
rect 591990 188466 592572 188526
rect 667013 187642 667079 187645
rect 666356 187640 667079 187642
rect 666356 187584 667018 187640
rect 667074 187584 667079 187640
rect 666356 187582 667079 187584
rect 667013 187579 667079 187582
rect 578509 187370 578575 187373
rect 576380 187368 578575 187370
rect 576380 187312 578514 187368
rect 578570 187312 578575 187368
rect 576380 187310 578575 187312
rect 578509 187307 578575 187310
rect 589365 186962 589431 186965
rect 589365 186960 592050 186962
rect 589365 186904 589370 186960
rect 589426 186904 592050 186960
rect 589365 186902 592050 186904
rect 589365 186899 589431 186902
rect 591990 186894 592050 186902
rect 591990 186834 592572 186894
rect 669262 186356 669268 186420
rect 669332 186418 669338 186420
rect 669630 186418 669636 186420
rect 669332 186358 669636 186418
rect 669332 186356 669338 186358
rect 669630 186356 669636 186358
rect 669700 186356 669706 186420
rect 41781 185876 41847 185877
rect 41781 185872 41828 185876
rect 41892 185874 41898 185876
rect 578325 185874 578391 185877
rect 41781 185816 41786 185872
rect 41781 185812 41828 185816
rect 41892 185814 41938 185874
rect 576380 185872 578391 185874
rect 576380 185816 578330 185872
rect 578386 185816 578391 185872
rect 576380 185814 578391 185816
rect 41892 185812 41898 185814
rect 41781 185811 41847 185812
rect 578325 185811 578391 185814
rect 674782 185812 674788 185876
rect 674852 185874 674858 185876
rect 676029 185874 676095 185877
rect 674852 185872 676095 185874
rect 674852 185816 676034 185872
rect 676090 185816 676095 185872
rect 674852 185814 676095 185816
rect 674852 185812 674858 185814
rect 676029 185811 676095 185814
rect 589457 185330 589523 185333
rect 589457 185328 592050 185330
rect 589457 185272 589462 185328
rect 589518 185272 592050 185328
rect 589457 185270 592050 185272
rect 589457 185267 589523 185270
rect 591990 185262 592050 185270
rect 591990 185202 592572 185262
rect 579521 184378 579587 184381
rect 576380 184376 579587 184378
rect 576380 184320 579526 184376
rect 579582 184320 579587 184376
rect 576380 184318 579587 184320
rect 666356 184318 666570 184378
rect 579521 184315 579587 184318
rect 666510 184245 666570 184318
rect 666510 184240 666619 184245
rect 666510 184184 666558 184240
rect 666614 184184 666619 184240
rect 666510 184182 666619 184184
rect 666553 184179 666619 184182
rect 41454 184044 41460 184108
rect 41524 184106 41530 184108
rect 41781 184106 41847 184109
rect 41524 184104 41847 184106
rect 41524 184048 41786 184104
rect 41842 184048 41847 184104
rect 41524 184046 41847 184048
rect 41524 184044 41530 184046
rect 41781 184043 41847 184046
rect 592174 183570 592572 183630
rect 590377 183562 590443 183565
rect 592174 183562 592234 183570
rect 590377 183560 592234 183562
rect 590377 183504 590382 183560
rect 590438 183504 592234 183560
rect 590377 183502 592234 183504
rect 672533 183562 672599 183565
rect 672942 183562 672948 183564
rect 672533 183560 672948 183562
rect 672533 183504 672538 183560
rect 672594 183504 672948 183560
rect 672533 183502 672948 183504
rect 590377 183499 590443 183502
rect 672533 183499 672599 183502
rect 672942 183500 672948 183502
rect 673012 183500 673018 183564
rect 40534 183364 40540 183428
rect 40604 183426 40610 183428
rect 41781 183426 41847 183429
rect 40604 183424 41847 183426
rect 40604 183368 41786 183424
rect 41842 183368 41847 183424
rect 40604 183366 41847 183368
rect 40604 183364 40610 183366
rect 41781 183363 41847 183366
rect 578877 182882 578943 182885
rect 576380 182880 578943 182882
rect 576380 182824 578882 182880
rect 578938 182824 578943 182880
rect 576380 182822 578943 182824
rect 578877 182819 578943 182822
rect 668577 182746 668643 182749
rect 666356 182744 668643 182746
rect 666356 182688 668582 182744
rect 668638 182688 668643 182744
rect 666356 182686 668643 182688
rect 668577 182683 668643 182686
rect 588537 182066 588603 182069
rect 588537 182064 592050 182066
rect 588537 182008 588542 182064
rect 588598 182008 592050 182064
rect 588537 182006 592050 182008
rect 588537 182003 588603 182006
rect 591990 181998 592050 182006
rect 591990 181938 592572 181998
rect 578509 181386 578575 181389
rect 576380 181384 578575 181386
rect 576380 181328 578514 181384
rect 578570 181328 578575 181384
rect 576380 181326 578575 181328
rect 578509 181323 578575 181326
rect 589457 180434 589523 180437
rect 589457 180432 592050 180434
rect 589457 180376 589462 180432
rect 589518 180376 592050 180432
rect 589457 180374 592050 180376
rect 589457 180371 589523 180374
rect 591990 180366 592050 180374
rect 591990 180306 592572 180366
rect 578969 179890 579035 179893
rect 576380 179888 579035 179890
rect 576380 179832 578974 179888
rect 579030 179832 579035 179888
rect 576380 179830 579035 179832
rect 578969 179827 579035 179830
rect 669446 179482 669452 179484
rect 666356 179422 669452 179482
rect 669446 179420 669452 179422
rect 669516 179420 669522 179484
rect 589549 178802 589615 178805
rect 589549 178800 592050 178802
rect 589549 178744 589554 178800
rect 589610 178744 592050 178800
rect 589549 178742 592050 178744
rect 589549 178739 589615 178742
rect 591990 178734 592050 178742
rect 591990 178674 592572 178734
rect 675477 178530 675543 178533
rect 675477 178528 676292 178530
rect 675477 178472 675482 178528
rect 675538 178472 676292 178528
rect 675477 178470 676292 178472
rect 675477 178467 675543 178470
rect 578601 178394 578667 178397
rect 576380 178392 578667 178394
rect 576380 178336 578606 178392
rect 578662 178336 578667 178392
rect 576380 178334 578667 178336
rect 578601 178331 578667 178334
rect 675477 178122 675543 178125
rect 675477 178120 676292 178122
rect 675477 178064 675482 178120
rect 675538 178064 676292 178120
rect 675477 178062 676292 178064
rect 675477 178059 675543 178062
rect 668577 177850 668643 177853
rect 666356 177848 668643 177850
rect 666356 177792 668582 177848
rect 668638 177792 668643 177848
rect 666356 177790 668643 177792
rect 668577 177787 668643 177790
rect 675477 177714 675543 177717
rect 675477 177712 676292 177714
rect 675477 177656 675482 177712
rect 675538 177656 676292 177712
rect 675477 177654 676292 177656
rect 675477 177651 675543 177654
rect 676029 177306 676095 177309
rect 676029 177304 676292 177306
rect 676029 177248 676034 177304
rect 676090 177248 676292 177304
rect 676029 177246 676292 177248
rect 676029 177243 676095 177246
rect 589457 177170 589523 177173
rect 589457 177168 592050 177170
rect 589457 177112 589462 177168
rect 589518 177112 592050 177168
rect 589457 177110 592050 177112
rect 589457 177107 589523 177110
rect 591990 177102 592050 177110
rect 591990 177042 592572 177102
rect 579521 176898 579587 176901
rect 576380 176896 579587 176898
rect 576380 176840 579526 176896
rect 579582 176840 579587 176896
rect 576380 176838 579587 176840
rect 579521 176835 579587 176838
rect 675477 176898 675543 176901
rect 675477 176896 676292 176898
rect 675477 176840 675482 176896
rect 675538 176840 676292 176896
rect 675477 176838 676292 176840
rect 675477 176835 675543 176838
rect 675477 176490 675543 176493
rect 675477 176488 676292 176490
rect 675477 176432 675482 176488
rect 675538 176432 676292 176488
rect 675477 176430 676292 176432
rect 675477 176427 675543 176430
rect 674465 176082 674531 176085
rect 674465 176080 676292 176082
rect 674465 176024 674470 176080
rect 674526 176024 676292 176080
rect 674465 176022 676292 176024
rect 674465 176019 674531 176022
rect 674649 175674 674715 175677
rect 674649 175672 676292 175674
rect 674649 175616 674654 175672
rect 674710 175616 676292 175672
rect 674649 175614 676292 175616
rect 674649 175611 674715 175614
rect 579429 175538 579495 175541
rect 576350 175536 579495 175538
rect 576350 175480 579434 175536
rect 579490 175480 579495 175536
rect 576350 175478 579495 175480
rect 576350 175372 576410 175478
rect 579429 175475 579495 175478
rect 589457 175538 589523 175541
rect 589457 175536 592050 175538
rect 589457 175480 589462 175536
rect 589518 175480 592050 175536
rect 589457 175478 592050 175480
rect 589457 175475 589523 175478
rect 591990 175470 592050 175478
rect 591990 175410 592572 175470
rect 675477 175266 675543 175269
rect 675477 175264 676292 175266
rect 675477 175208 675482 175264
rect 675538 175208 676292 175264
rect 675477 175206 676292 175208
rect 675477 175203 675543 175206
rect 676170 174798 676292 174858
rect 675886 174660 675892 174724
rect 675956 174722 675962 174724
rect 676170 174722 676230 174798
rect 675956 174662 676230 174722
rect 675956 174660 675962 174662
rect 669446 174586 669452 174588
rect 666356 174526 669452 174586
rect 669446 174524 669452 174526
rect 669516 174524 669522 174588
rect 675477 174450 675543 174453
rect 675477 174448 676292 174450
rect 675477 174392 675482 174448
rect 675538 174392 676292 174448
rect 675477 174390 676292 174392
rect 675477 174387 675543 174390
rect 675017 174042 675083 174045
rect 675017 174040 676292 174042
rect 675017 173984 675022 174040
rect 675078 173984 676292 174040
rect 675017 173982 676292 173984
rect 675017 173979 675083 173982
rect 578325 173906 578391 173909
rect 576380 173904 578391 173906
rect 576380 173848 578330 173904
rect 578386 173848 578391 173904
rect 576380 173846 578391 173848
rect 578325 173843 578391 173846
rect 589273 173906 589339 173909
rect 589273 173904 592050 173906
rect 589273 173848 589278 173904
rect 589334 173848 592050 173904
rect 589273 173846 592050 173848
rect 589273 173843 589339 173846
rect 591990 173838 592050 173846
rect 591990 173778 592572 173838
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 675845 173226 675911 173229
rect 675845 173224 676292 173226
rect 675845 173168 675850 173224
rect 675906 173168 676292 173224
rect 675845 173166 676292 173168
rect 675845 173163 675911 173166
rect 673126 172954 673132 172956
rect 666356 172894 673132 172954
rect 673126 172892 673132 172894
rect 673196 172892 673202 172956
rect 676029 172818 676095 172821
rect 676029 172816 676292 172818
rect 676029 172760 676034 172816
rect 676090 172760 676292 172816
rect 676029 172758 676292 172760
rect 676029 172755 676095 172758
rect 579061 172410 579127 172413
rect 576380 172408 579127 172410
rect 576380 172352 579066 172408
rect 579122 172352 579127 172408
rect 576380 172350 579127 172352
rect 579061 172347 579127 172350
rect 678237 172410 678303 172413
rect 678237 172408 678316 172410
rect 678237 172352 678242 172408
rect 678298 172352 678316 172408
rect 678237 172350 678316 172352
rect 678237 172347 678303 172350
rect 589365 172274 589431 172277
rect 589365 172272 592050 172274
rect 589365 172216 589370 172272
rect 589426 172216 592050 172272
rect 589365 172214 592050 172216
rect 589365 172211 589431 172214
rect 591990 172206 592050 172214
rect 591990 172146 592572 172206
rect 674465 172002 674531 172005
rect 674465 172000 676292 172002
rect 674465 171944 674470 172000
rect 674526 171944 676292 172000
rect 674465 171942 676292 171944
rect 674465 171939 674531 171942
rect 675201 171594 675267 171597
rect 675201 171592 676292 171594
rect 675201 171536 675206 171592
rect 675262 171536 676292 171592
rect 675201 171534 676292 171536
rect 675201 171531 675267 171534
rect 675477 171186 675543 171189
rect 675477 171184 676292 171186
rect 675477 171128 675482 171184
rect 675538 171128 676292 171184
rect 675477 171126 676292 171128
rect 675477 171123 675543 171126
rect 579521 170914 579587 170917
rect 576380 170912 579587 170914
rect 576380 170856 579526 170912
rect 579582 170856 579587 170912
rect 576380 170854 579587 170856
rect 579521 170851 579587 170854
rect 676673 170778 676739 170781
rect 676660 170776 676739 170778
rect 676660 170720 676678 170776
rect 676734 170720 676739 170776
rect 676660 170718 676739 170720
rect 676673 170715 676739 170718
rect 589457 170642 589523 170645
rect 589457 170640 592050 170642
rect 589457 170584 589462 170640
rect 589518 170584 592050 170640
rect 589457 170582 592050 170584
rect 589457 170579 589523 170582
rect 591990 170574 592050 170582
rect 591990 170514 592572 170574
rect 675886 170308 675892 170372
rect 675956 170370 675962 170372
rect 675956 170310 676292 170370
rect 675956 170308 675962 170310
rect 676397 169962 676463 169965
rect 676397 169960 676476 169962
rect 676397 169904 676402 169960
rect 676458 169904 676476 169960
rect 676397 169902 676476 169904
rect 676397 169899 676463 169902
rect 669957 169690 670023 169693
rect 666356 169688 670023 169690
rect 666356 169632 669962 169688
rect 670018 169632 670023 169688
rect 666356 169630 670023 169632
rect 669957 169627 670023 169630
rect 675477 169554 675543 169557
rect 675477 169552 676292 169554
rect 675477 169496 675482 169552
rect 675538 169496 676292 169552
rect 675477 169494 676292 169496
rect 675477 169491 675543 169494
rect 578233 169418 578299 169421
rect 576380 169416 578299 169418
rect 576380 169360 578238 169416
rect 578294 169360 578299 169416
rect 576380 169358 578299 169360
rect 578233 169355 578299 169358
rect 675477 169146 675543 169149
rect 675477 169144 676292 169146
rect 675477 169088 675482 169144
rect 675538 169088 676292 169144
rect 675477 169086 676292 169088
rect 675477 169083 675543 169086
rect 589457 169010 589523 169013
rect 589457 169008 592050 169010
rect 589457 168952 589462 169008
rect 589518 168952 592050 169008
rect 589457 168950 592050 168952
rect 589457 168947 589523 168950
rect 591990 168942 592050 168950
rect 591990 168882 592572 168942
rect 675477 168738 675543 168741
rect 675477 168736 676292 168738
rect 675477 168680 675482 168736
rect 675538 168680 676292 168736
rect 675477 168678 676292 168680
rect 675477 168675 675543 168678
rect 672073 168332 672139 168333
rect 672022 168330 672028 168332
rect 671982 168270 672028 168330
rect 672092 168328 672139 168332
rect 672134 168272 672139 168328
rect 672022 168268 672028 168270
rect 672092 168268 672139 168272
rect 672073 168267 672139 168268
rect 676170 168270 676292 168330
rect 676170 168194 676230 168270
rect 672214 168134 676230 168194
rect 670918 168058 670924 168060
rect 666356 167998 670924 168058
rect 670918 167996 670924 167998
rect 670988 167996 670994 168060
rect 671981 168058 672047 168061
rect 672214 168058 672274 168134
rect 671981 168056 672274 168058
rect 671981 168000 671986 168056
rect 672042 168000 672274 168056
rect 671981 167998 672274 168000
rect 671981 167995 672047 167998
rect 579429 167922 579495 167925
rect 576380 167920 579495 167922
rect 576380 167864 579434 167920
rect 579490 167864 579495 167920
rect 576380 167862 579495 167864
rect 579429 167859 579495 167862
rect 675661 167922 675727 167925
rect 675661 167920 676292 167922
rect 675661 167864 675666 167920
rect 675722 167864 676292 167920
rect 675661 167862 676292 167864
rect 675661 167859 675727 167862
rect 675886 167452 675892 167516
rect 675956 167514 675962 167516
rect 675956 167454 676292 167514
rect 675956 167452 675962 167454
rect 589457 167378 589523 167381
rect 589457 167376 592050 167378
rect 589457 167320 589462 167376
rect 589518 167320 592050 167376
rect 589457 167318 592050 167320
rect 589457 167315 589523 167318
rect 591990 167310 592050 167318
rect 591990 167250 592572 167310
rect 675477 167106 675543 167109
rect 675477 167104 676292 167106
rect 675477 167048 675482 167104
rect 675538 167048 676292 167104
rect 675477 167046 676292 167048
rect 675477 167043 675543 167046
rect 579061 166426 579127 166429
rect 576380 166424 579127 166426
rect 576380 166368 579066 166424
rect 579122 166368 579127 166424
rect 576380 166366 579127 166368
rect 579061 166363 579127 166366
rect 676397 166428 676463 166429
rect 676397 166424 676444 166428
rect 676508 166426 676514 166428
rect 676397 166368 676402 166424
rect 676397 166364 676444 166368
rect 676508 166366 676554 166426
rect 676508 166364 676514 166366
rect 676397 166363 676463 166364
rect 676673 166292 676739 166293
rect 676622 166228 676628 166292
rect 676692 166290 676739 166292
rect 676692 166288 676784 166290
rect 676734 166232 676784 166288
rect 676692 166230 676784 166232
rect 676692 166228 676739 166230
rect 676673 166227 676739 166228
rect 592174 165618 592572 165678
rect 589457 165610 589523 165613
rect 592174 165610 592234 165618
rect 589457 165608 592234 165610
rect 589457 165552 589462 165608
rect 589518 165552 592234 165608
rect 589457 165550 592234 165552
rect 589457 165547 589523 165550
rect 576350 164386 576410 164900
rect 670734 164794 670740 164796
rect 666356 164734 670740 164794
rect 670734 164732 670740 164734
rect 670804 164732 670810 164796
rect 579521 164386 579587 164389
rect 576350 164384 579587 164386
rect 576350 164328 579526 164384
rect 579582 164328 579587 164384
rect 576350 164326 579587 164328
rect 579521 164323 579587 164326
rect 589917 164114 589983 164117
rect 589917 164112 592050 164114
rect 589917 164056 589922 164112
rect 589978 164056 592050 164112
rect 589917 164054 592050 164056
rect 589917 164051 589983 164054
rect 591990 164046 592050 164054
rect 591990 163986 592572 164046
rect 578693 163434 578759 163437
rect 576380 163432 578759 163434
rect 576380 163376 578698 163432
rect 578754 163376 578759 163432
rect 576380 163374 578759 163376
rect 578693 163371 578759 163374
rect 668025 163162 668091 163165
rect 666356 163160 668091 163162
rect 666356 163104 668030 163160
rect 668086 163104 668091 163160
rect 666356 163102 668091 163104
rect 668025 163099 668091 163102
rect 589457 162482 589523 162485
rect 589457 162480 592050 162482
rect 589457 162424 589462 162480
rect 589518 162424 592050 162480
rect 589457 162422 592050 162424
rect 589457 162419 589523 162422
rect 591990 162414 592050 162422
rect 591990 162354 592572 162414
rect 674833 162210 674899 162213
rect 676029 162210 676095 162213
rect 674833 162208 676095 162210
rect 674833 162152 674838 162208
rect 674894 162152 676034 162208
rect 676090 162152 676095 162208
rect 674833 162150 676095 162152
rect 674833 162147 674899 162150
rect 676029 162147 676095 162150
rect 578877 161938 578943 161941
rect 576380 161936 578943 161938
rect 576380 161880 578882 161936
rect 578938 161880 578943 161936
rect 576380 161878 578943 161880
rect 578877 161875 578943 161878
rect 675702 161876 675708 161940
rect 675772 161938 675778 161940
rect 678237 161938 678303 161941
rect 675772 161936 678303 161938
rect 675772 161880 678242 161936
rect 678298 161880 678303 161936
rect 675772 161878 678303 161880
rect 675772 161876 675778 161878
rect 678237 161875 678303 161878
rect 589457 160850 589523 160853
rect 589457 160848 592050 160850
rect 589457 160792 589462 160848
rect 589518 160792 592050 160848
rect 589457 160790 592050 160792
rect 589457 160787 589523 160790
rect 591990 160782 592050 160790
rect 591990 160722 592572 160782
rect 578509 160442 578575 160445
rect 576380 160440 578575 160442
rect 576380 160384 578514 160440
rect 578570 160384 578575 160440
rect 576380 160382 578575 160384
rect 578509 160379 578575 160382
rect 672022 159898 672028 159900
rect 666356 159838 672028 159898
rect 672022 159836 672028 159838
rect 672092 159836 672098 159900
rect 588721 159218 588787 159221
rect 588721 159216 592050 159218
rect 588721 159160 588726 159216
rect 588782 159160 592050 159216
rect 588721 159158 592050 159160
rect 588721 159155 588787 159158
rect 591990 159150 592050 159158
rect 591990 159090 592572 159150
rect 579521 158946 579587 158949
rect 576380 158944 579587 158946
rect 576380 158888 579526 158944
rect 579582 158888 579587 158944
rect 576380 158886 579587 158888
rect 579521 158883 579587 158886
rect 668761 158266 668827 158269
rect 666356 158264 668827 158266
rect 666356 158208 668766 158264
rect 668822 158208 668827 158264
rect 666356 158206 668827 158208
rect 668761 158203 668827 158206
rect 589457 157586 589523 157589
rect 589457 157584 592050 157586
rect 589457 157528 589462 157584
rect 589518 157528 592050 157584
rect 589457 157526 592050 157528
rect 589457 157523 589523 157526
rect 591990 157518 592050 157526
rect 591990 157458 592572 157518
rect 579429 157450 579495 157453
rect 576380 157448 579495 157450
rect 576380 157392 579434 157448
rect 579490 157392 579495 157448
rect 576380 157390 579495 157392
rect 579429 157387 579495 157390
rect 675753 156362 675819 156365
rect 676622 156362 676628 156364
rect 675753 156360 676628 156362
rect 675753 156304 675758 156360
rect 675814 156304 676628 156360
rect 675753 156302 676628 156304
rect 675753 156299 675819 156302
rect 676622 156300 676628 156302
rect 676692 156300 676698 156364
rect 579245 155954 579311 155957
rect 576380 155952 579311 155954
rect 576380 155896 579250 155952
rect 579306 155896 579311 155952
rect 576380 155894 579311 155896
rect 579245 155891 579311 155894
rect 590377 155954 590443 155957
rect 590377 155952 592050 155954
rect 590377 155896 590382 155952
rect 590438 155896 592050 155952
rect 590377 155894 592050 155896
rect 590377 155891 590443 155894
rect 591990 155886 592050 155894
rect 591990 155826 592572 155886
rect 671245 155138 671311 155141
rect 666694 155136 671311 155138
rect 666694 155080 671250 155136
rect 671306 155080 671311 155136
rect 666694 155078 671311 155080
rect 666356 154968 666570 155002
rect 666694 154968 666754 155078
rect 671245 155075 671311 155078
rect 666356 154942 666754 154968
rect 666510 154908 666754 154942
rect 579245 154458 579311 154461
rect 576380 154456 579311 154458
rect 576380 154400 579250 154456
rect 579306 154400 579311 154456
rect 576380 154398 579311 154400
rect 579245 154395 579311 154398
rect 589365 154322 589431 154325
rect 589365 154320 592050 154322
rect 589365 154264 589370 154320
rect 589426 154264 592050 154320
rect 589365 154262 592050 154264
rect 589365 154259 589431 154262
rect 591990 154254 592050 154262
rect 591990 154194 592572 154254
rect 666356 153310 673470 153370
rect 673410 153234 673470 153310
rect 673678 153234 673684 153236
rect 673410 153174 673684 153234
rect 673678 153172 673684 153174
rect 673748 153172 673754 153236
rect 675661 153100 675727 153101
rect 675661 153096 675708 153100
rect 675772 153098 675778 153100
rect 675661 153040 675666 153096
rect 675661 153036 675708 153040
rect 675772 153038 675818 153098
rect 675772 153036 675778 153038
rect 675661 153035 675727 153036
rect 578693 152962 578759 152965
rect 576380 152960 578759 152962
rect 576380 152904 578698 152960
rect 578754 152904 578759 152960
rect 576380 152902 578759 152904
rect 578693 152899 578759 152902
rect 589457 152690 589523 152693
rect 589457 152688 592050 152690
rect 589457 152632 589462 152688
rect 589518 152632 592050 152688
rect 589457 152630 592050 152632
rect 589457 152627 589523 152630
rect 591990 152622 592050 152630
rect 591990 152562 592572 152622
rect 579153 151466 579219 151469
rect 576380 151464 579219 151466
rect 576380 151408 579158 151464
rect 579214 151408 579219 151464
rect 576380 151406 579219 151408
rect 579153 151403 579219 151406
rect 675753 151466 675819 151469
rect 676438 151466 676444 151468
rect 675753 151464 676444 151466
rect 675753 151408 675758 151464
rect 675814 151408 676444 151464
rect 675753 151406 676444 151408
rect 675753 151403 675819 151406
rect 676438 151404 676444 151406
rect 676508 151404 676514 151468
rect 589457 151058 589523 151061
rect 589457 151056 592050 151058
rect 589457 151000 589462 151056
rect 589518 151000 592050 151056
rect 589457 150998 592050 151000
rect 589457 150995 589523 150998
rect 591990 150990 592050 150998
rect 591990 150930 592572 150990
rect 675753 150378 675819 150381
rect 676254 150378 676260 150380
rect 675753 150376 676260 150378
rect 675753 150320 675758 150376
rect 675814 150320 676260 150376
rect 675753 150318 676260 150320
rect 675753 150315 675819 150318
rect 676254 150316 676260 150318
rect 676324 150316 676330 150380
rect 666356 150046 669882 150106
rect 578877 149970 578943 149973
rect 576380 149968 578943 149970
rect 576380 149912 578882 149968
rect 578938 149912 578943 149968
rect 576380 149910 578943 149912
rect 578877 149907 578943 149910
rect 669822 149698 669882 150046
rect 673494 149698 673500 149700
rect 669822 149638 673500 149698
rect 673494 149636 673500 149638
rect 673564 149636 673570 149700
rect 589457 149426 589523 149429
rect 589457 149424 592050 149426
rect 589457 149368 589462 149424
rect 589518 149368 592050 149424
rect 589457 149366 592050 149368
rect 589457 149363 589523 149366
rect 591990 149358 592050 149366
rect 591990 149298 592572 149358
rect 579521 148474 579587 148477
rect 668761 148474 668827 148477
rect 576380 148472 579587 148474
rect 576380 148416 579526 148472
rect 579582 148416 579587 148472
rect 576380 148414 579587 148416
rect 666356 148472 668827 148474
rect 666356 148416 668766 148472
rect 668822 148416 668827 148472
rect 666356 148414 668827 148416
rect 579521 148411 579587 148414
rect 668761 148411 668827 148414
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 592174 147666 592572 147726
rect 589457 147658 589523 147661
rect 592174 147658 592234 147666
rect 589457 147656 592234 147658
rect 589457 147600 589462 147656
rect 589518 147600 592234 147656
rect 589457 147598 592234 147600
rect 675661 147658 675727 147661
rect 675886 147658 675892 147660
rect 675661 147656 675892 147658
rect 675661 147600 675666 147656
rect 675722 147600 675892 147656
rect 675661 147598 675892 147600
rect 589457 147595 589523 147598
rect 675661 147595 675727 147598
rect 675886 147596 675892 147598
rect 675956 147596 675962 147660
rect 579245 146978 579311 146981
rect 576380 146976 579311 146978
rect 576380 146920 579250 146976
rect 579306 146920 579311 146976
rect 576380 146918 579311 146920
rect 579245 146915 579311 146918
rect 588537 146162 588603 146165
rect 588537 146160 592050 146162
rect 588537 146104 588542 146160
rect 588598 146104 592050 146160
rect 588537 146102 592050 146104
rect 588537 146099 588603 146102
rect 591990 146094 592050 146102
rect 591990 146034 592572 146094
rect 579429 145482 579495 145485
rect 576380 145480 579495 145482
rect 576380 145424 579434 145480
rect 579490 145424 579495 145480
rect 576380 145422 579495 145424
rect 579429 145419 579495 145422
rect 668761 145210 668827 145213
rect 666356 145208 668827 145210
rect 666356 145152 668766 145208
rect 668822 145152 668827 145208
rect 666356 145150 668827 145152
rect 668761 145147 668827 145150
rect 589917 144530 589983 144533
rect 589917 144528 592050 144530
rect 589917 144472 589922 144528
rect 589978 144472 592050 144528
rect 589917 144470 592050 144472
rect 589917 144467 589983 144470
rect 591990 144462 592050 144470
rect 591990 144402 592572 144462
rect 578509 143986 578575 143989
rect 576380 143984 578575 143986
rect 576380 143928 578514 143984
rect 578570 143928 578575 143984
rect 576380 143926 578575 143928
rect 578509 143923 578575 143926
rect 668761 143578 668827 143581
rect 666356 143576 668827 143578
rect 666356 143520 668766 143576
rect 668822 143520 668827 143576
rect 666356 143518 668827 143520
rect 668761 143515 668827 143518
rect 590009 142898 590075 142901
rect 590009 142896 592050 142898
rect 590009 142840 590014 142896
rect 590070 142840 592050 142896
rect 590009 142838 592050 142840
rect 590009 142835 590075 142838
rect 591990 142830 592050 142838
rect 591990 142770 592572 142830
rect 579521 142490 579587 142493
rect 576380 142488 579587 142490
rect 576380 142432 579526 142488
rect 579582 142432 579587 142488
rect 576380 142430 579587 142432
rect 579521 142427 579587 142430
rect 589457 141266 589523 141269
rect 589457 141264 592050 141266
rect 589457 141208 589462 141264
rect 589518 141208 592050 141264
rect 589457 141206 592050 141208
rect 589457 141203 589523 141206
rect 591990 141198 592050 141206
rect 591990 141138 592572 141198
rect 578877 140994 578943 140997
rect 576380 140992 578943 140994
rect 576380 140936 578882 140992
rect 578938 140936 578943 140992
rect 576380 140934 578943 140936
rect 578877 140931 578943 140934
rect 668761 140314 668827 140317
rect 666356 140312 668827 140314
rect 666356 140256 668766 140312
rect 668822 140256 668827 140312
rect 666356 140254 668827 140256
rect 668761 140251 668827 140254
rect 589457 139634 589523 139637
rect 589457 139632 592050 139634
rect 589457 139576 589462 139632
rect 589518 139576 592050 139632
rect 589457 139574 592050 139576
rect 589457 139571 589523 139574
rect 591990 139566 592050 139574
rect 591990 139506 592572 139566
rect 579521 139498 579587 139501
rect 576380 139496 579587 139498
rect 576380 139440 579526 139496
rect 579582 139440 579587 139496
rect 576380 139438 579587 139440
rect 579521 139435 579587 139438
rect 668761 138682 668827 138685
rect 666356 138680 668827 138682
rect 666356 138624 668766 138680
rect 668822 138624 668827 138680
rect 666356 138622 668827 138624
rect 668761 138619 668827 138622
rect 579245 138002 579311 138005
rect 576380 138000 579311 138002
rect 576380 137944 579250 138000
rect 579306 137944 579311 138000
rect 576380 137942 579311 137944
rect 579245 137939 579311 137942
rect 589457 138002 589523 138005
rect 589457 138000 592050 138002
rect 589457 137944 589462 138000
rect 589518 137944 592050 138000
rect 589457 137942 592050 137944
rect 589457 137939 589523 137942
rect 591990 137934 592050 137942
rect 591990 137874 592572 137934
rect 579061 136506 579127 136509
rect 576380 136504 579127 136506
rect 576380 136448 579066 136504
rect 579122 136448 579127 136504
rect 576380 136446 579127 136448
rect 579061 136443 579127 136446
rect 589365 136370 589431 136373
rect 589365 136368 592050 136370
rect 589365 136312 589370 136368
rect 589426 136312 592050 136368
rect 589365 136310 592050 136312
rect 589365 136307 589431 136310
rect 591990 136302 592050 136310
rect 591990 136242 592572 136302
rect 668209 135418 668275 135421
rect 666356 135416 668275 135418
rect 666356 135360 668214 135416
rect 668270 135360 668275 135416
rect 666356 135358 668275 135360
rect 668209 135355 668275 135358
rect 578233 135010 578299 135013
rect 576380 135008 578299 135010
rect 576380 134952 578238 135008
rect 578294 134952 578299 135008
rect 576380 134950 578299 134952
rect 578233 134947 578299 134950
rect 588721 134738 588787 134741
rect 588721 134736 592050 134738
rect 588721 134680 588726 134736
rect 588782 134680 592050 134736
rect 588721 134678 592050 134680
rect 588721 134675 588787 134678
rect 591990 134670 592050 134678
rect 591990 134610 592572 134670
rect 669221 133786 669287 133789
rect 666356 133784 669287 133786
rect 666356 133728 669226 133784
rect 669282 133728 669287 133784
rect 666356 133726 669287 133728
rect 669221 133723 669287 133726
rect 578509 133514 578575 133517
rect 576380 133512 578575 133514
rect 576380 133456 578514 133512
rect 578570 133456 578575 133512
rect 576380 133454 578575 133456
rect 578509 133451 578575 133454
rect 675477 133378 675543 133381
rect 675477 133376 676292 133378
rect 675477 133320 675482 133376
rect 675538 133320 676292 133376
rect 675477 133318 676292 133320
rect 675477 133315 675543 133318
rect 590377 133106 590443 133109
rect 590377 133104 592050 133106
rect 590377 133048 590382 133104
rect 590438 133048 592050 133104
rect 590377 133046 592050 133048
rect 590377 133043 590443 133046
rect 591990 133038 592050 133046
rect 591990 132978 592572 133038
rect 675477 132970 675543 132973
rect 675477 132968 676292 132970
rect 675477 132912 675482 132968
rect 675538 132912 676292 132968
rect 675477 132910 676292 132912
rect 675477 132907 675543 132910
rect 675477 132562 675543 132565
rect 675477 132560 676292 132562
rect 675477 132504 675482 132560
rect 675538 132504 676292 132560
rect 675477 132502 676292 132504
rect 675477 132499 675543 132502
rect 675477 132154 675543 132157
rect 675477 132152 676292 132154
rect 675477 132096 675482 132152
rect 675538 132096 676292 132152
rect 675477 132094 676292 132096
rect 675477 132091 675543 132094
rect 578417 132018 578483 132021
rect 576380 132016 578483 132018
rect 576380 131960 578422 132016
rect 578478 131960 578483 132016
rect 576380 131958 578483 131960
rect 578417 131955 578483 131958
rect 675477 131746 675543 131749
rect 675477 131744 676292 131746
rect 675477 131688 675482 131744
rect 675538 131688 676292 131744
rect 675477 131686 676292 131688
rect 675477 131683 675543 131686
rect 589457 131474 589523 131477
rect 589457 131472 592050 131474
rect 589457 131416 589462 131472
rect 589518 131416 592050 131472
rect 589457 131414 592050 131416
rect 589457 131411 589523 131414
rect 591990 131406 592050 131414
rect 591990 131346 592572 131406
rect 674649 131338 674715 131341
rect 674649 131336 676292 131338
rect 674649 131280 674654 131336
rect 674710 131280 676292 131336
rect 674649 131278 676292 131280
rect 674649 131275 674715 131278
rect 675477 130930 675543 130933
rect 675477 130928 676292 130930
rect 675477 130872 675482 130928
rect 675538 130872 676292 130928
rect 675477 130870 676292 130872
rect 675477 130867 675543 130870
rect 578601 130522 578667 130525
rect 668301 130522 668367 130525
rect 576380 130520 578667 130522
rect 576380 130464 578606 130520
rect 578662 130464 578667 130520
rect 576380 130462 578667 130464
rect 666356 130520 668367 130522
rect 666356 130464 668306 130520
rect 668362 130464 668367 130520
rect 666356 130462 668367 130464
rect 578601 130459 578667 130462
rect 668301 130459 668367 130462
rect 675477 130522 675543 130525
rect 675477 130520 676292 130522
rect 675477 130464 675482 130520
rect 675538 130464 676292 130520
rect 675477 130462 676292 130464
rect 675477 130459 675543 130462
rect 675477 130114 675543 130117
rect 675477 130112 676292 130114
rect 675477 130056 675482 130112
rect 675538 130056 676292 130112
rect 675477 130054 676292 130056
rect 675477 130051 675543 130054
rect 592174 129714 592572 129774
rect 589457 129706 589523 129709
rect 592174 129706 592234 129714
rect 589457 129704 592234 129706
rect 589457 129648 589462 129704
rect 589518 129648 592234 129704
rect 589457 129646 592234 129648
rect 675477 129706 675543 129709
rect 675477 129704 676292 129706
rect 675477 129648 675482 129704
rect 675538 129648 676292 129704
rect 675477 129646 676292 129648
rect 589457 129643 589523 129646
rect 675477 129643 675543 129646
rect 675477 129298 675543 129301
rect 675477 129296 676292 129298
rect 675477 129240 675482 129296
rect 675538 129240 676292 129296
rect 675477 129238 676292 129240
rect 675477 129235 675543 129238
rect 579429 129026 579495 129029
rect 576380 129024 579495 129026
rect 576380 128968 579434 129024
rect 579490 128968 579495 129024
rect 576380 128966 579495 128968
rect 579429 128963 579495 128966
rect 669221 128890 669287 128893
rect 666356 128888 669287 128890
rect 666356 128832 669226 128888
rect 669282 128832 669287 128888
rect 666356 128830 669287 128832
rect 669221 128827 669287 128830
rect 676262 128620 676322 128860
rect 676254 128556 676260 128620
rect 676324 128556 676330 128620
rect 676262 128213 676322 128452
rect 589457 128210 589523 128213
rect 589457 128208 592050 128210
rect 589457 128152 589462 128208
rect 589518 128152 592050 128208
rect 589457 128150 592050 128152
rect 589457 128147 589523 128150
rect 591990 128142 592050 128150
rect 676213 128208 676322 128213
rect 676213 128152 676218 128208
rect 676274 128152 676322 128208
rect 676213 128150 676322 128152
rect 676213 128147 676279 128150
rect 591990 128082 592572 128142
rect 676446 127805 676506 128044
rect 676397 127800 676506 127805
rect 676397 127744 676402 127800
rect 676458 127744 676506 127800
rect 676397 127742 676506 127744
rect 676397 127739 676463 127742
rect 674833 127666 674899 127669
rect 674833 127664 676292 127666
rect 674833 127608 674838 127664
rect 674894 127608 676292 127664
rect 674833 127606 676292 127608
rect 674833 127603 674899 127606
rect 578325 127530 578391 127533
rect 576380 127528 578391 127530
rect 576380 127472 578330 127528
rect 578386 127472 578391 127528
rect 576380 127470 578391 127472
rect 578325 127467 578391 127470
rect 675886 127196 675892 127260
rect 675956 127258 675962 127260
rect 675956 127198 676292 127258
rect 675956 127196 675962 127198
rect 589733 126578 589799 126581
rect 682886 126578 682946 126820
rect 683113 126578 683179 126581
rect 589733 126576 592050 126578
rect 589733 126520 589738 126576
rect 589794 126520 592050 126576
rect 589733 126518 592050 126520
rect 682886 126576 683179 126578
rect 682886 126520 683118 126576
rect 683174 126520 683179 126576
rect 682886 126518 683179 126520
rect 589733 126515 589799 126518
rect 591990 126510 592050 126518
rect 683113 126515 683179 126518
rect 591990 126450 592572 126510
rect 679574 126173 679634 126412
rect 679574 126168 679683 126173
rect 679574 126112 679622 126168
rect 679678 126112 679683 126168
rect 679574 126110 679683 126112
rect 679617 126107 679683 126110
rect 578509 126034 578575 126037
rect 576380 126032 578575 126034
rect 576380 125976 578514 126032
rect 578570 125976 578575 126032
rect 576380 125974 578575 125976
rect 578509 125971 578575 125974
rect 675477 126034 675543 126037
rect 675477 126032 676292 126034
rect 675477 125976 675482 126032
rect 675538 125976 676292 126032
rect 675477 125974 676292 125976
rect 675477 125971 675543 125974
rect 668209 125626 668275 125629
rect 666356 125624 668275 125626
rect 666356 125568 668214 125624
rect 668270 125568 668275 125624
rect 666356 125566 668275 125568
rect 668209 125563 668275 125566
rect 675477 125626 675543 125629
rect 675477 125624 676292 125626
rect 675477 125568 675482 125624
rect 675538 125568 676292 125624
rect 675477 125566 676292 125568
rect 675477 125563 675543 125566
rect 674373 125218 674439 125221
rect 674373 125216 676292 125218
rect 674373 125160 674378 125216
rect 674434 125160 676292 125216
rect 674373 125158 676292 125160
rect 674373 125155 674439 125158
rect 589917 124946 589983 124949
rect 589917 124944 592050 124946
rect 589917 124888 589922 124944
rect 589978 124888 592050 124944
rect 589917 124886 592050 124888
rect 589917 124883 589983 124886
rect 591990 124878 592050 124886
rect 591990 124818 592572 124878
rect 674189 124810 674255 124813
rect 674189 124808 676292 124810
rect 674189 124752 674194 124808
rect 674250 124752 676292 124808
rect 674189 124750 676292 124752
rect 674189 124747 674255 124750
rect 578877 124538 578943 124541
rect 576380 124536 578943 124538
rect 576380 124480 578882 124536
rect 578938 124480 578943 124536
rect 576380 124478 578943 124480
rect 578877 124475 578943 124478
rect 676806 124476 676812 124540
rect 676876 124538 676882 124540
rect 683113 124538 683179 124541
rect 676876 124536 683179 124538
rect 676876 124480 683118 124536
rect 683174 124480 683179 124536
rect 676876 124478 683179 124480
rect 676876 124476 676882 124478
rect 683113 124475 683179 124478
rect 676998 124132 677058 124372
rect 676990 124068 676996 124132
rect 677060 124068 677066 124132
rect 668025 123994 668091 123997
rect 666356 123992 668091 123994
rect 666356 123936 668030 123992
rect 668086 123936 668091 123992
rect 666356 123934 668091 123936
rect 668025 123931 668091 123934
rect 675477 123994 675543 123997
rect 675477 123992 676292 123994
rect 675477 123936 675482 123992
rect 675538 123936 676292 123992
rect 675477 123934 676292 123936
rect 675477 123931 675543 123934
rect 674649 123586 674715 123589
rect 674649 123584 676292 123586
rect 674649 123528 674654 123584
rect 674710 123528 676292 123584
rect 674649 123526 676292 123528
rect 674649 123523 674715 123526
rect 589457 123314 589523 123317
rect 589457 123312 592050 123314
rect 589457 123256 589462 123312
rect 589518 123256 592050 123312
rect 589457 123254 592050 123256
rect 589457 123251 589523 123254
rect 591990 123246 592050 123254
rect 591990 123186 592572 123246
rect 675477 123178 675543 123181
rect 675477 123176 676292 123178
rect 675477 123120 675482 123176
rect 675538 123120 676292 123176
rect 675477 123118 676292 123120
rect 675477 123115 675543 123118
rect 578877 123042 578943 123045
rect 576380 123040 578943 123042
rect 576380 122984 578882 123040
rect 578938 122984 578943 123040
rect 576380 122982 578943 122984
rect 578877 122979 578943 122982
rect 675702 122844 675708 122908
rect 675772 122906 675778 122908
rect 676213 122906 676279 122909
rect 675772 122904 676279 122906
rect 675772 122848 676218 122904
rect 676274 122848 676279 122904
rect 675772 122846 676279 122848
rect 675772 122844 675778 122846
rect 676213 122843 676279 122846
rect 675477 122498 675543 122501
rect 676446 122498 676506 122740
rect 675477 122496 676506 122498
rect 675477 122440 675482 122496
rect 675538 122440 676506 122496
rect 675477 122438 676506 122440
rect 675477 122435 675543 122438
rect 677550 122093 677610 122332
rect 677550 122088 677659 122093
rect 677550 122032 677598 122088
rect 677654 122032 677659 122088
rect 677550 122030 677659 122032
rect 677593 122027 677659 122030
rect 675477 121954 675543 121957
rect 675477 121952 676292 121954
rect 675477 121896 675482 121952
rect 675538 121896 676292 121952
rect 675477 121894 676292 121896
rect 675477 121891 675543 121894
rect 590377 121682 590443 121685
rect 590377 121680 592050 121682
rect 590377 121624 590382 121680
rect 590438 121624 592050 121680
rect 590377 121622 592050 121624
rect 590377 121619 590443 121622
rect 591990 121614 592050 121622
rect 591990 121554 592572 121614
rect 579521 121546 579587 121549
rect 576380 121544 579587 121546
rect 576380 121488 579526 121544
rect 579582 121488 579587 121544
rect 576380 121486 579587 121488
rect 579521 121483 579587 121486
rect 669681 120730 669747 120733
rect 666356 120728 669747 120730
rect 666356 120672 669686 120728
rect 669742 120672 669747 120728
rect 666356 120670 669747 120672
rect 669681 120667 669747 120670
rect 675702 120260 675708 120324
rect 675772 120322 675778 120324
rect 676070 120322 676076 120324
rect 675772 120262 676076 120322
rect 675772 120260 675778 120262
rect 676070 120260 676076 120262
rect 676140 120260 676146 120324
rect 579245 120050 579311 120053
rect 576380 120048 579311 120050
rect 576380 119992 579250 120048
rect 579306 119992 579311 120048
rect 576380 119990 579311 119992
rect 579245 119987 579311 119990
rect 589457 120050 589523 120053
rect 589457 120048 592050 120050
rect 589457 119992 589462 120048
rect 589518 119992 592050 120048
rect 589457 119990 592050 119992
rect 589457 119987 589523 119990
rect 591990 119982 592050 119990
rect 591990 119922 592572 119982
rect 669221 119098 669287 119101
rect 666356 119096 669287 119098
rect 666356 119040 669226 119096
rect 669282 119040 669287 119096
rect 666356 119038 669287 119040
rect 669221 119035 669287 119038
rect 579061 118554 579127 118557
rect 576380 118552 579127 118554
rect 576380 118496 579066 118552
rect 579122 118496 579127 118552
rect 576380 118494 579127 118496
rect 579061 118491 579127 118494
rect 588537 118418 588603 118421
rect 588537 118416 592050 118418
rect 588537 118360 588542 118416
rect 588598 118360 592050 118416
rect 588537 118358 592050 118360
rect 588537 118355 588603 118358
rect 591990 118350 592050 118358
rect 591990 118290 592572 118350
rect 669957 117466 670023 117469
rect 666356 117464 670023 117466
rect 666356 117408 669962 117464
rect 670018 117408 670023 117464
rect 666356 117406 670023 117408
rect 669957 117403 670023 117406
rect 578325 117058 578391 117061
rect 576380 117056 578391 117058
rect 576380 117000 578330 117056
rect 578386 117000 578391 117056
rect 576380 116998 578391 117000
rect 578325 116995 578391 116998
rect 589457 116786 589523 116789
rect 589457 116784 592050 116786
rect 589457 116728 589462 116784
rect 589518 116728 592050 116784
rect 589457 116726 592050 116728
rect 589457 116723 589523 116726
rect 591990 116718 592050 116726
rect 591990 116658 592572 116718
rect 675702 116044 675708 116108
rect 675772 116106 675778 116108
rect 677593 116106 677659 116109
rect 675772 116104 677659 116106
rect 675772 116048 677598 116104
rect 677654 116048 677659 116104
rect 675772 116046 677659 116048
rect 675772 116044 675778 116046
rect 677593 116043 677659 116046
rect 669221 115834 669287 115837
rect 666356 115832 669287 115834
rect 666356 115776 669226 115832
rect 669282 115776 669287 115832
rect 666356 115774 669287 115776
rect 669221 115771 669287 115774
rect 589273 115154 589339 115157
rect 589273 115152 592050 115154
rect 589273 115096 589278 115152
rect 589334 115096 592050 115152
rect 589273 115094 592050 115096
rect 589273 115091 589339 115094
rect 591990 115086 592050 115094
rect 591990 115026 592572 115086
rect 669221 114202 669287 114205
rect 666356 114200 669287 114202
rect 666356 114144 669226 114200
rect 669282 114144 669287 114200
rect 666356 114142 669287 114144
rect 669221 114139 669287 114142
rect 675753 114202 675819 114205
rect 676254 114202 676260 114204
rect 675753 114200 676260 114202
rect 675753 114144 675758 114200
rect 675814 114144 676260 114200
rect 675753 114142 676260 114144
rect 675753 114139 675819 114142
rect 676254 114140 676260 114142
rect 676324 114140 676330 114204
rect 589457 113522 589523 113525
rect 589457 113520 592050 113522
rect 589457 113464 589462 113520
rect 589518 113464 592050 113520
rect 589457 113462 592050 113464
rect 589457 113459 589523 113462
rect 591990 113454 592050 113462
rect 591990 113394 592572 113454
rect 668301 112570 668367 112573
rect 666356 112568 668367 112570
rect 666356 112512 668306 112568
rect 668362 112512 668367 112568
rect 666356 112510 668367 112512
rect 668301 112507 668367 112510
rect 592174 111762 592572 111822
rect 589457 111754 589523 111757
rect 592174 111754 592234 111762
rect 589457 111752 592234 111754
rect 589457 111696 589462 111752
rect 589518 111696 592234 111752
rect 589457 111694 592234 111696
rect 589457 111691 589523 111694
rect 669037 110938 669103 110941
rect 666356 110936 669103 110938
rect 666356 110880 669042 110936
rect 669098 110880 669103 110936
rect 666356 110878 669103 110880
rect 669037 110875 669103 110878
rect 675753 110394 675819 110397
rect 676990 110394 676996 110396
rect 675753 110392 676996 110394
rect 675753 110336 675758 110392
rect 675814 110336 676996 110392
rect 675753 110334 676996 110336
rect 675753 110331 675819 110334
rect 676990 110332 676996 110334
rect 677060 110332 677066 110396
rect 589917 110258 589983 110261
rect 589917 110256 592050 110258
rect 589917 110200 589922 110256
rect 589978 110200 592050 110256
rect 589917 110198 592050 110200
rect 589917 110195 589983 110198
rect 591990 110190 592050 110198
rect 591990 110130 592572 110190
rect 666737 109374 666803 109377
rect 666356 109372 666803 109374
rect 666356 109316 666742 109372
rect 666798 109316 666803 109372
rect 666356 109314 666803 109316
rect 666737 109311 666803 109314
rect 589457 108626 589523 108629
rect 589457 108624 592050 108626
rect 589457 108568 589462 108624
rect 589518 108568 592050 108624
rect 589457 108566 592050 108568
rect 589457 108563 589523 108566
rect 591990 108558 592050 108566
rect 591990 108498 592572 108558
rect 675661 108082 675727 108085
rect 675886 108082 675892 108084
rect 675661 108080 675892 108082
rect 675661 108024 675666 108080
rect 675722 108024 675892 108080
rect 675661 108022 675892 108024
rect 675661 108019 675727 108022
rect 675886 108020 675892 108022
rect 675956 108020 675962 108084
rect 669129 107674 669195 107677
rect 666356 107672 669195 107674
rect 666356 107616 669134 107672
rect 669190 107616 669195 107672
rect 666356 107614 669195 107616
rect 669129 107611 669195 107614
rect 589365 106994 589431 106997
rect 589365 106992 592050 106994
rect 589365 106936 589370 106992
rect 589426 106936 592050 106992
rect 589365 106934 592050 106936
rect 589365 106931 589431 106934
rect 591990 106926 592050 106934
rect 591990 106866 592572 106926
rect 668761 106042 668827 106045
rect 666356 106040 668827 106042
rect 666356 105984 668766 106040
rect 668822 105984 668827 106040
rect 666356 105982 668827 105984
rect 668761 105979 668827 105982
rect 589273 105362 589339 105365
rect 589273 105360 592050 105362
rect 589273 105304 589278 105360
rect 589334 105304 592050 105360
rect 589273 105302 592050 105304
rect 589273 105299 589339 105302
rect 591990 105294 592050 105302
rect 591990 105234 592572 105294
rect 668945 104410 669011 104413
rect 666356 104408 669011 104410
rect 666356 104352 668950 104408
rect 669006 104352 669011 104408
rect 666356 104350 669011 104352
rect 668945 104347 669011 104350
rect 589365 103730 589431 103733
rect 589365 103728 592050 103730
rect 589365 103672 589370 103728
rect 589426 103672 592050 103728
rect 589365 103670 592050 103672
rect 589365 103667 589431 103670
rect 591990 103662 592050 103670
rect 591990 103602 592572 103662
rect 675753 103186 675819 103189
rect 676070 103186 676076 103188
rect 675753 103184 676076 103186
rect 675753 103128 675758 103184
rect 675814 103128 676076 103184
rect 675753 103126 676076 103128
rect 675753 103123 675819 103126
rect 676070 103124 676076 103126
rect 676140 103124 676146 103188
rect 668577 102778 668643 102781
rect 666356 102776 668643 102778
rect 666356 102720 668582 102776
rect 668638 102720 668643 102776
rect 666356 102718 668643 102720
rect 668577 102715 668643 102718
rect 675661 102644 675727 102645
rect 675661 102640 675708 102644
rect 675772 102642 675778 102644
rect 675661 102584 675666 102640
rect 675661 102580 675708 102584
rect 675772 102582 675818 102642
rect 675772 102580 675778 102582
rect 675661 102579 675727 102580
rect 589457 102098 589523 102101
rect 589457 102096 592050 102098
rect 589457 102040 589462 102096
rect 589518 102040 592050 102096
rect 589457 102038 592050 102040
rect 589457 102035 589523 102038
rect 591990 102030 592050 102038
rect 591990 101970 592572 102030
rect 675753 101418 675819 101421
rect 676806 101418 676812 101420
rect 675753 101416 676812 101418
rect 675753 101360 675758 101416
rect 675814 101360 676812 101416
rect 675753 101358 676812 101360
rect 675753 101355 675819 101358
rect 676806 101356 676812 101358
rect 676876 101356 676882 101420
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 634670 95644 634676 95708
rect 634740 95706 634746 95708
rect 635917 95706 635983 95709
rect 634740 95704 635983 95706
rect 634740 95648 635922 95704
rect 635978 95648 635983 95704
rect 634740 95646 635983 95648
rect 634740 95644 634746 95646
rect 635917 95643 635983 95646
rect 626441 95434 626507 95437
rect 626441 95432 628268 95434
rect 626441 95376 626446 95432
rect 626502 95376 628268 95432
rect 626441 95374 628268 95376
rect 626441 95371 626507 95374
rect 642633 95162 642699 95165
rect 642590 95160 642699 95162
rect 642590 95104 642638 95160
rect 642694 95104 642699 95160
rect 642590 95099 642699 95104
rect 642590 94588 642650 95099
rect 626073 94482 626139 94485
rect 626073 94480 628268 94482
rect 626073 94424 626078 94480
rect 626134 94424 628268 94480
rect 626073 94422 628268 94424
rect 626073 94419 626139 94422
rect 653949 94210 654015 94213
rect 653949 94208 656788 94210
rect 653949 94152 653954 94208
rect 654010 94152 656788 94208
rect 653949 94150 656788 94152
rect 653949 94147 654015 94150
rect 626441 93530 626507 93533
rect 626441 93528 628268 93530
rect 626441 93472 626446 93528
rect 626502 93472 628268 93528
rect 626441 93470 628268 93472
rect 626441 93467 626507 93470
rect 654317 93394 654383 93397
rect 665173 93394 665239 93397
rect 654317 93392 656788 93394
rect 654317 93336 654322 93392
rect 654378 93336 656788 93392
rect 654317 93334 656788 93336
rect 663596 93392 665239 93394
rect 663596 93336 665178 93392
rect 665234 93336 665239 93392
rect 663596 93334 665239 93336
rect 654317 93331 654383 93334
rect 665173 93331 665239 93334
rect 663241 93122 663307 93125
rect 663198 93120 663307 93122
rect 663198 93064 663246 93120
rect 663302 93064 663307 93120
rect 663198 93059 663307 93064
rect 626257 92578 626323 92581
rect 654133 92578 654199 92581
rect 626257 92576 628268 92578
rect 626257 92520 626262 92576
rect 626318 92520 628268 92576
rect 626257 92518 628268 92520
rect 654133 92576 656788 92578
rect 654133 92520 654138 92576
rect 654194 92520 656788 92576
rect 663198 92548 663258 93059
rect 654133 92518 656788 92520
rect 626257 92515 626323 92518
rect 654133 92515 654199 92518
rect 644473 92170 644539 92173
rect 642988 92168 644539 92170
rect 642988 92112 644478 92168
rect 644534 92112 644539 92168
rect 642988 92110 644539 92112
rect 644473 92107 644539 92110
rect 665357 91762 665423 91765
rect 663596 91760 665423 91762
rect 663596 91704 665362 91760
rect 665418 91704 665423 91760
rect 663596 91702 665423 91704
rect 665357 91699 665423 91702
rect 625429 91626 625495 91629
rect 625429 91624 628268 91626
rect 625429 91568 625434 91624
rect 625490 91568 628268 91624
rect 625429 91566 628268 91568
rect 625429 91563 625495 91566
rect 654317 91490 654383 91493
rect 654317 91488 656788 91490
rect 654317 91432 654322 91488
rect 654378 91432 656788 91488
rect 654317 91430 656788 91432
rect 654317 91427 654383 91430
rect 626441 90674 626507 90677
rect 654133 90674 654199 90677
rect 665541 90674 665607 90677
rect 626441 90672 628268 90674
rect 626441 90616 626446 90672
rect 626502 90616 628268 90672
rect 626441 90614 628268 90616
rect 654133 90672 656788 90674
rect 654133 90616 654138 90672
rect 654194 90616 656788 90672
rect 654133 90614 656788 90616
rect 663596 90672 665607 90674
rect 663596 90616 665546 90672
rect 665602 90616 665607 90672
rect 663596 90614 665607 90616
rect 626441 90611 626507 90614
rect 654133 90611 654199 90614
rect 665541 90611 665607 90614
rect 663793 90402 663859 90405
rect 663566 90400 663859 90402
rect 663566 90344 663798 90400
rect 663854 90344 663859 90400
rect 663566 90342 663859 90344
rect 655789 89858 655855 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 663566 89828 663626 90342
rect 663793 90339 663859 90342
rect 655789 89798 656788 89800
rect 655789 89795 655855 89798
rect 626441 89722 626507 89725
rect 644749 89722 644815 89725
rect 626441 89720 628268 89722
rect 626441 89664 626446 89720
rect 626502 89664 628268 89720
rect 626441 89662 628268 89664
rect 642988 89720 644815 89722
rect 642988 89664 644754 89720
rect 644810 89664 644815 89720
rect 642988 89662 644815 89664
rect 626441 89659 626507 89662
rect 644749 89659 644815 89662
rect 663977 89042 664043 89045
rect 663596 89040 664043 89042
rect 663596 88984 663982 89040
rect 664038 88984 664043 89040
rect 663596 88982 664043 88984
rect 663977 88979 664043 88982
rect 624969 88362 625035 88365
rect 628238 88362 628298 88876
rect 624969 88360 628298 88362
rect 624969 88304 624974 88360
rect 625030 88304 628298 88360
rect 624969 88302 628298 88304
rect 624969 88299 625035 88302
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 643553 87138 643619 87141
rect 642988 87136 643619 87138
rect 642988 87080 643558 87136
rect 643614 87080 643619 87136
rect 642988 87078 643619 87080
rect 643553 87075 643619 87078
rect 625613 87002 625679 87005
rect 625613 87000 628268 87002
rect 625613 86944 625618 87000
rect 625674 86944 628268 87000
rect 625613 86942 628268 86944
rect 625613 86939 625679 86942
rect 626441 86050 626507 86053
rect 626441 86048 628268 86050
rect 626441 85992 626446 86048
rect 626502 85992 628268 86048
rect 626441 85990 628268 85992
rect 626441 85987 626507 85990
rect 626441 85098 626507 85101
rect 626441 85096 628268 85098
rect 626441 85040 626446 85096
rect 626502 85040 628268 85096
rect 626441 85038 628268 85040
rect 626441 85035 626507 85038
rect 643369 84690 643435 84693
rect 642988 84688 643435 84690
rect 642988 84632 643374 84688
rect 643430 84632 643435 84688
rect 642988 84630 643435 84632
rect 643369 84627 643435 84630
rect 626441 84146 626507 84149
rect 626441 84144 628268 84146
rect 626441 84088 626446 84144
rect 626502 84088 628268 84144
rect 626441 84086 628268 84088
rect 626441 84083 626507 84086
rect 626257 83194 626323 83197
rect 626257 83192 628268 83194
rect 626257 83136 626262 83192
rect 626318 83136 628268 83192
rect 626257 83134 628268 83136
rect 626257 83131 626323 83134
rect 643093 82786 643159 82789
rect 642774 82784 643159 82786
rect 642774 82728 643098 82784
rect 643154 82728 643159 82784
rect 642774 82726 643159 82728
rect 642774 82212 642834 82726
rect 643093 82723 643159 82726
rect 628606 81701 628666 82212
rect 628557 81696 628666 81701
rect 628557 81640 628562 81696
rect 628618 81640 628666 81696
rect 628557 81638 628666 81640
rect 628557 81635 628623 81638
rect 628790 80882 628850 81396
rect 629201 80882 629267 80885
rect 628790 80880 629267 80882
rect 628790 80824 629206 80880
rect 629262 80824 629267 80880
rect 628790 80822 629267 80824
rect 629201 80819 629267 80822
rect 637113 78572 637179 78573
rect 637062 78570 637068 78572
rect 637022 78510 637068 78570
rect 637132 78568 637179 78572
rect 637174 78512 637179 78568
rect 637062 78508 637068 78510
rect 637132 78508 637179 78512
rect 637113 78507 637179 78508
rect 633893 77754 633959 77757
rect 634670 77754 634676 77756
rect 633893 77752 634676 77754
rect 633893 77696 633898 77752
rect 633954 77696 634676 77752
rect 633893 77694 634676 77696
rect 633893 77691 633959 77694
rect 634670 77692 634676 77694
rect 634740 77692 634746 77756
rect 646865 74490 646931 74493
rect 646668 74488 646931 74490
rect 646668 74432 646870 74488
rect 646926 74432 646931 74488
rect 646668 74430 646931 74432
rect 646865 74427 646931 74430
rect 647417 72994 647483 72997
rect 646668 72992 647483 72994
rect 646668 72936 647422 72992
rect 647478 72936 647483 72992
rect 646668 72934 647483 72936
rect 647417 72931 647483 72934
rect 646129 71770 646195 71773
rect 646086 71768 646195 71770
rect 646086 71712 646134 71768
rect 646190 71712 646195 71768
rect 646086 71707 646195 71712
rect 646086 71468 646146 71707
rect 646313 70410 646379 70413
rect 646270 70408 646379 70410
rect 646270 70352 646318 70408
rect 646374 70352 646379 70408
rect 646270 70347 646379 70352
rect 646270 69972 646330 70347
rect 647601 68506 647667 68509
rect 646668 68504 647667 68506
rect 646668 68448 647606 68504
rect 647662 68448 647667 68504
rect 646668 68446 647667 68448
rect 647601 68443 647667 68446
rect 649165 67010 649231 67013
rect 646668 67008 649231 67010
rect 646668 66952 649170 67008
rect 649226 66952 649231 67008
rect 646668 66950 649231 66952
rect 649165 66947 649231 66950
rect 646129 66058 646195 66061
rect 646086 66056 646195 66058
rect 646086 66000 646134 66056
rect 646190 66000 646195 66056
rect 646086 65995 646195 66000
rect 646086 65484 646146 65995
rect 648797 64018 648863 64021
rect 646668 64016 648863 64018
rect 646668 63960 648802 64016
rect 648858 63960 648863 64016
rect 646668 63958 648863 63960
rect 648797 63955 648863 63958
rect 464838 51716 464844 51780
rect 464908 51778 464914 51780
rect 603073 51778 603139 51781
rect 464908 51776 603139 51778
rect 464908 51720 603078 51776
rect 603134 51720 603139 51776
rect 464908 51718 603139 51720
rect 464908 51716 464914 51718
rect 603073 51715 603139 51718
rect 497549 50554 497615 50557
rect 525742 50554 525748 50556
rect 497549 50552 525748 50554
rect 497549 50496 497554 50552
rect 497610 50496 525748 50552
rect 497549 50494 525748 50496
rect 497549 50491 497615 50494
rect 525742 50492 525748 50494
rect 525812 50492 525818 50556
rect 131021 50282 131087 50285
rect 150382 50282 150388 50284
rect 131021 50280 150388 50282
rect 131021 50224 131026 50280
rect 131082 50224 150388 50280
rect 131021 50222 150388 50224
rect 131021 50219 131087 50222
rect 150382 50220 150388 50222
rect 150452 50220 150458 50284
rect 445201 50282 445267 50285
rect 517462 50282 517468 50284
rect 445201 50280 517468 50282
rect 445201 50224 445206 50280
rect 445262 50224 517468 50280
rect 445201 50222 517468 50224
rect 445201 50219 445267 50222
rect 517462 50220 517468 50222
rect 517532 50220 517538 50284
rect 529790 50220 529796 50284
rect 529860 50282 529866 50284
rect 549253 50282 549319 50285
rect 529860 50280 549319 50282
rect 529860 50224 549258 50280
rect 549314 50224 549319 50280
rect 529860 50222 549319 50224
rect 529860 50220 529866 50222
rect 549253 50219 549319 50222
rect 78581 49740 78647 49741
rect 78581 49736 78628 49740
rect 78692 49738 78698 49740
rect 78581 49680 78586 49736
rect 78581 49676 78628 49680
rect 78692 49678 78738 49738
rect 78692 49676 78698 49678
rect 78581 49675 78647 49676
rect 411110 49132 411116 49196
rect 411180 49194 411186 49196
rect 600313 49194 600379 49197
rect 411180 49192 600379 49194
rect 411180 49136 600318 49192
rect 600374 49136 600379 49192
rect 411180 49134 600379 49136
rect 411180 49132 411186 49134
rect 600313 49131 600379 49134
rect 365478 48860 365484 48924
rect 365548 48922 365554 48924
rect 596173 48922 596239 48925
rect 365548 48920 596239 48922
rect 365548 48864 596178 48920
rect 596234 48864 596239 48920
rect 365548 48862 596239 48864
rect 365548 48860 365554 48862
rect 596173 48859 596239 48862
rect 661266 48245 661326 48482
rect 661217 48240 661326 48245
rect 661217 48184 661222 48240
rect 661278 48184 661326 48240
rect 661217 48182 661326 48184
rect 661217 48179 661283 48182
rect 415209 48106 415275 48109
rect 595437 48106 595503 48109
rect 415209 48104 595503 48106
rect 415209 48048 415214 48104
rect 415270 48048 595442 48104
rect 595498 48048 595503 48104
rect 415209 48046 595503 48048
rect 415209 48043 415275 48046
rect 595437 48043 595503 48046
rect 310462 47772 310468 47836
rect 310532 47834 310538 47836
rect 597553 47834 597619 47837
rect 310532 47832 597619 47834
rect 310532 47776 597558 47832
rect 597614 47776 597619 47832
rect 661585 47791 661651 47794
rect 310532 47774 597619 47776
rect 310532 47772 310538 47774
rect 597553 47771 597619 47774
rect 661388 47789 661651 47791
rect 661388 47733 661590 47789
rect 661646 47733 661651 47789
rect 661388 47731 661651 47733
rect 661585 47728 661651 47731
rect 150382 47500 150388 47564
rect 150452 47562 150458 47564
rect 150452 47502 171150 47562
rect 150452 47500 150458 47502
rect 78622 47228 78628 47292
rect 78692 47290 78698 47292
rect 151905 47290 151971 47293
rect 78692 47230 122850 47290
rect 78692 47228 78698 47230
rect 122790 47018 122850 47230
rect 145238 47288 151971 47290
rect 145238 47232 151910 47288
rect 151966 47232 151971 47288
rect 145238 47230 151971 47232
rect 171090 47290 171150 47502
rect 187550 47500 187556 47564
rect 187620 47562 187626 47564
rect 591297 47562 591363 47565
rect 187620 47560 591363 47562
rect 187620 47504 591302 47560
rect 591358 47504 591363 47560
rect 187620 47502 591363 47504
rect 187620 47500 187626 47502
rect 591297 47499 591363 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 451273 47290 451339 47293
rect 171090 47288 451339 47290
rect 171090 47232 451278 47288
rect 451334 47232 451339 47288
rect 171090 47230 451339 47232
rect 145238 47018 145298 47230
rect 151905 47227 151971 47230
rect 451273 47227 451339 47230
rect 451457 47290 451523 47293
rect 461025 47290 461091 47293
rect 451457 47288 461091 47290
rect 451457 47232 451462 47288
rect 451518 47232 461030 47288
rect 461086 47232 461091 47288
rect 451457 47230 461091 47232
rect 451457 47227 451523 47230
rect 461025 47227 461091 47230
rect 461209 47290 461275 47293
rect 470593 47290 470659 47293
rect 461209 47288 470659 47290
rect 461209 47232 461214 47288
rect 461270 47232 470598 47288
rect 470654 47232 470659 47288
rect 461209 47230 470659 47232
rect 461209 47227 461275 47230
rect 470593 47227 470659 47230
rect 470777 47290 470843 47293
rect 480437 47290 480503 47293
rect 470777 47288 480503 47290
rect 470777 47232 470782 47288
rect 470838 47232 480442 47288
rect 480498 47232 480503 47288
rect 470777 47230 480503 47232
rect 470777 47227 470843 47230
rect 480437 47227 480503 47230
rect 480621 47290 480687 47293
rect 490005 47290 490071 47293
rect 480621 47288 490071 47290
rect 480621 47232 480626 47288
rect 480682 47232 490010 47288
rect 490066 47232 490071 47288
rect 480621 47230 490071 47232
rect 480621 47227 480687 47230
rect 490005 47227 490071 47230
rect 490189 47290 490255 47293
rect 499757 47290 499823 47293
rect 490189 47288 499823 47290
rect 490189 47232 490194 47288
rect 490250 47232 499762 47288
rect 499818 47232 499823 47288
rect 490189 47230 499823 47232
rect 490189 47227 490255 47230
rect 499757 47227 499823 47230
rect 499941 47290 500007 47293
rect 513741 47290 513807 47293
rect 598933 47290 598999 47293
rect 499941 47288 513807 47290
rect 499941 47232 499946 47288
rect 500002 47232 513746 47288
rect 513802 47232 513807 47288
rect 499941 47230 513807 47232
rect 499941 47227 500007 47230
rect 513741 47227 513807 47230
rect 513974 47288 598999 47290
rect 513974 47232 598938 47288
rect 598994 47232 598999 47288
rect 513974 47230 598999 47232
rect 122790 46958 145298 47018
rect 238710 46958 267750 47018
rect 151905 45930 151971 45933
rect 238710 45930 238770 46958
rect 151905 45928 238770 45930
rect 151905 45872 151910 45928
rect 151966 45872 238770 45928
rect 151905 45870 238770 45872
rect 267690 45930 267750 46958
rect 416630 46956 416636 47020
rect 416700 47018 416706 47020
rect 513974 47018 514034 47230
rect 598933 47227 598999 47230
rect 416700 46958 514034 47018
rect 514201 47018 514267 47021
rect 521694 47018 521700 47020
rect 514201 47016 521700 47018
rect 514201 46960 514206 47016
rect 514262 46960 521700 47016
rect 514201 46958 521700 46960
rect 416700 46956 416706 46958
rect 514201 46955 514267 46958
rect 521694 46956 521700 46958
rect 521764 46956 521770 47020
rect 451273 46746 451339 46749
rect 461209 46746 461275 46749
rect 451273 46744 461275 46746
rect 451273 46688 451278 46744
rect 451334 46688 461214 46744
rect 461270 46688 461275 46744
rect 451273 46686 461275 46688
rect 451273 46683 451339 46686
rect 461209 46683 461275 46686
rect 465717 46746 465783 46749
rect 600957 46746 601023 46749
rect 465717 46744 601023 46746
rect 465717 46688 465722 46744
rect 465778 46688 600962 46744
rect 601018 46688 601023 46744
rect 465717 46686 601023 46688
rect 465717 46683 465783 46686
rect 600957 46683 601023 46686
rect 361982 46412 361988 46476
rect 362052 46474 362058 46476
rect 594057 46474 594123 46477
rect 362052 46472 594123 46474
rect 362052 46416 594062 46472
rect 594118 46416 594123 46472
rect 362052 46414 594123 46416
rect 362052 46412 362058 46414
rect 594057 46411 594123 46414
rect 306966 46140 306972 46204
rect 307036 46202 307042 46204
rect 592677 46202 592743 46205
rect 307036 46200 592743 46202
rect 307036 46144 592682 46200
rect 592738 46144 592743 46200
rect 307036 46142 592743 46144
rect 307036 46140 307042 46142
rect 592677 46139 592743 46142
rect 451457 45930 451523 45933
rect 267690 45928 451523 45930
rect 267690 45872 451462 45928
rect 451518 45872 451523 45928
rect 267690 45870 451523 45872
rect 151905 45867 151971 45870
rect 451457 45867 451523 45870
rect 465901 45930 465967 45933
rect 470777 45930 470843 45933
rect 465901 45928 470843 45930
rect 465901 45872 465906 45928
rect 465962 45872 470782 45928
rect 470838 45872 470843 45928
rect 465901 45870 470843 45872
rect 465901 45867 465967 45870
rect 470777 45867 470843 45870
rect 470961 45930 471027 45933
rect 480253 45930 480319 45933
rect 470961 45928 480319 45930
rect 470961 45872 470966 45928
rect 471022 45872 480258 45928
rect 480314 45872 480319 45928
rect 470961 45870 480319 45872
rect 470961 45867 471027 45870
rect 480253 45867 480319 45870
rect 480437 45930 480503 45933
rect 490189 45930 490255 45933
rect 480437 45928 490255 45930
rect 480437 45872 480442 45928
rect 480498 45872 490194 45928
rect 490250 45872 490255 45928
rect 480437 45870 490255 45872
rect 480437 45867 480503 45870
rect 490189 45867 490255 45870
rect 490373 45930 490439 45933
rect 499573 45930 499639 45933
rect 490373 45928 499639 45930
rect 490373 45872 490378 45928
rect 490434 45872 499578 45928
rect 499634 45872 499639 45928
rect 490373 45870 499639 45872
rect 490373 45867 490439 45870
rect 499573 45867 499639 45870
rect 499757 45930 499823 45933
rect 514702 45930 514708 45932
rect 499757 45928 514708 45930
rect 499757 45872 499762 45928
rect 499818 45872 514708 45928
rect 499757 45870 514708 45872
rect 499757 45867 499823 45870
rect 514702 45868 514708 45870
rect 514772 45868 514778 45932
rect 460606 45732 460612 45796
rect 460676 45794 460682 45796
rect 465717 45794 465783 45797
rect 460676 45792 465783 45794
rect 460676 45736 465722 45792
rect 465778 45736 465783 45792
rect 460676 45734 465783 45736
rect 460676 45732 460682 45734
rect 465717 45731 465783 45734
rect 406377 45114 406443 45117
rect 520406 45114 520412 45116
rect 406377 45112 520412 45114
rect 406377 45056 406382 45112
rect 406438 45056 520412 45112
rect 406377 45054 520412 45056
rect 406377 45051 406443 45054
rect 520406 45052 520412 45054
rect 520476 45052 520482 45116
rect 471646 44780 471652 44844
rect 471716 44842 471722 44844
rect 601693 44842 601759 44845
rect 471716 44840 601759 44842
rect 471716 44784 601698 44840
rect 601754 44784 601759 44840
rect 471716 44782 601759 44784
rect 471716 44780 471722 44782
rect 601693 44779 601759 44782
rect 474457 43482 474523 43485
rect 604453 43482 604519 43485
rect 474457 43480 604519 43482
rect 474457 43424 474462 43480
rect 474518 43424 604458 43480
rect 604514 43424 604519 43480
rect 474457 43422 604519 43424
rect 474457 43419 474523 43422
rect 604453 43419 604519 43422
rect 411069 42804 411135 42805
rect 416589 42804 416655 42805
rect 464889 42804 464955 42805
rect 411069 42800 411116 42804
rect 411180 42802 411186 42804
rect 416589 42802 416636 42804
rect 411069 42744 411074 42800
rect 411069 42740 411116 42744
rect 411180 42742 411226 42802
rect 416544 42800 416636 42802
rect 416544 42744 416594 42800
rect 416544 42742 416636 42744
rect 411180 42740 411186 42742
rect 416589 42740 416636 42742
rect 416700 42740 416706 42804
rect 464838 42802 464844 42804
rect 464798 42742 464844 42802
rect 464908 42800 464955 42804
rect 464950 42744 464955 42800
rect 464838 42740 464844 42742
rect 464908 42740 464955 42744
rect 411069 42739 411135 42740
rect 416589 42739 416655 42740
rect 464889 42739 464955 42740
rect 306971 42396 307037 42397
rect 306966 42394 306972 42396
rect 306880 42334 306972 42394
rect 306966 42332 306972 42334
rect 307036 42332 307042 42396
rect 517462 42332 517468 42396
rect 517532 42394 517538 42396
rect 518525 42394 518591 42397
rect 517532 42392 518591 42394
rect 517532 42336 518530 42392
rect 518586 42336 518591 42392
rect 517532 42334 518591 42336
rect 517532 42332 517538 42334
rect 306971 42331 307037 42332
rect 518525 42331 518591 42334
rect 187509 42124 187575 42125
rect 310421 42124 310487 42125
rect 361941 42124 362007 42125
rect 187509 42122 187556 42124
rect 187464 42120 187556 42122
rect 187464 42064 187514 42120
rect 187464 42062 187556 42064
rect 187509 42060 187556 42062
rect 187620 42060 187626 42124
rect 310421 42122 310468 42124
rect 310376 42120 310468 42122
rect 310376 42064 310426 42120
rect 310376 42062 310468 42064
rect 310421 42060 310468 42062
rect 310532 42060 310538 42124
rect 361941 42122 361988 42124
rect 361896 42120 361988 42122
rect 361896 42064 361946 42120
rect 361896 42062 361988 42064
rect 361941 42060 361988 42062
rect 362052 42060 362058 42124
rect 365161 42122 365227 42125
rect 460565 42124 460631 42125
rect 471605 42124 471671 42125
rect 365478 42122 365484 42124
rect 365161 42120 365484 42122
rect 365161 42064 365166 42120
rect 365222 42064 365484 42120
rect 365161 42062 365484 42064
rect 187509 42059 187575 42060
rect 310421 42059 310487 42060
rect 361941 42059 362007 42060
rect 365161 42059 365227 42062
rect 365478 42060 365484 42062
rect 365548 42060 365554 42124
rect 460565 42122 460612 42124
rect 460520 42120 460612 42122
rect 460520 42064 460570 42120
rect 460520 42062 460612 42064
rect 460565 42060 460612 42062
rect 460676 42060 460682 42124
rect 471605 42122 471652 42124
rect 471560 42120 471652 42122
rect 471560 42064 471610 42120
rect 471560 42062 471652 42064
rect 471605 42060 471652 42062
rect 471716 42060 471722 42124
rect 514702 42060 514708 42124
rect 514772 42122 514778 42124
rect 514937 42122 515003 42125
rect 520457 42124 520523 42125
rect 525793 42124 525859 42125
rect 514772 42120 515003 42122
rect 514772 42064 514942 42120
rect 514998 42064 515003 42120
rect 514772 42062 515003 42064
rect 514772 42060 514778 42062
rect 460565 42059 460631 42060
rect 471605 42059 471671 42060
rect 514937 42059 515003 42062
rect 520406 42060 520412 42124
rect 520476 42122 520523 42124
rect 520476 42120 520568 42122
rect 520518 42064 520568 42120
rect 520476 42062 520568 42064
rect 520476 42060 520523 42062
rect 525742 42060 525748 42124
rect 525812 42122 525859 42124
rect 529565 42122 529631 42125
rect 529790 42122 529796 42124
rect 525812 42120 525904 42122
rect 525854 42064 525904 42120
rect 525812 42062 525904 42064
rect 529565 42120 529796 42122
rect 529565 42064 529570 42120
rect 529626 42064 529796 42120
rect 529565 42062 529796 42064
rect 525812 42060 525859 42062
rect 520457 42059 520523 42060
rect 525793 42059 525859 42060
rect 529565 42059 529631 42062
rect 529790 42060 529796 42062
rect 529860 42060 529866 42124
rect 521653 41988 521719 41989
rect 521653 41986 521700 41988
rect 521608 41984 521700 41986
rect 521608 41928 521658 41984
rect 521608 41926 521700 41928
rect 521653 41924 521700 41926
rect 521764 41924 521770 41988
rect 521653 41923 521719 41924
<< via3 >>
rect 383332 997656 383396 997660
rect 383332 997600 383346 997656
rect 383346 997600 383396 997656
rect 383332 997596 383396 997600
rect 194364 997188 194428 997252
rect 389036 997188 389100 997252
rect 138060 996916 138124 996980
rect 90220 996372 90284 996436
rect 86908 995964 86972 996028
rect 86908 995420 86972 995484
rect 90220 995480 90284 995484
rect 90220 995424 90234 995480
rect 90234 995424 90284 995480
rect 90220 995420 90284 995424
rect 138060 995692 138124 995756
rect 189396 995752 189460 995756
rect 189396 995696 189410 995752
rect 189410 995696 189460 995752
rect 189396 995692 189460 995696
rect 242572 996780 242636 996844
rect 295012 996372 295076 996436
rect 243860 996100 243924 996164
rect 239628 995752 239692 995756
rect 239628 995696 239642 995752
rect 239642 995696 239692 995752
rect 239628 995692 239692 995696
rect 243308 995752 243372 995756
rect 243308 995696 243322 995752
rect 243322 995696 243372 995752
rect 243308 995692 243372 995696
rect 295012 995752 295076 995756
rect 295012 995696 295062 995752
rect 295062 995696 295076 995752
rect 295012 995692 295076 995696
rect 243860 995616 243924 995620
rect 243860 995560 243874 995616
rect 243874 995560 243924 995616
rect 243860 995556 243924 995560
rect 274588 995556 274652 995620
rect 473308 996644 473372 996708
rect 388116 995692 388180 995756
rect 389036 995692 389100 995756
rect 473308 995752 473372 995756
rect 529612 996644 529676 996708
rect 627132 996644 627196 996708
rect 473308 995696 473358 995752
rect 473358 995696 473372 995752
rect 473308 995692 473372 995696
rect 630812 996372 630876 996436
rect 529612 995692 529676 995756
rect 536604 995752 536668 995756
rect 536604 995696 536618 995752
rect 536618 995696 536668 995752
rect 536604 995692 536668 995696
rect 627132 995752 627196 995756
rect 627132 995696 627182 995752
rect 627182 995696 627196 995752
rect 627132 995692 627196 995696
rect 630812 995480 630876 995484
rect 630812 995424 630862 995480
rect 630862 995424 630876 995480
rect 630812 995420 630876 995424
rect 573220 989436 573284 989500
rect 41460 968764 41524 968828
rect 42012 967192 42076 967196
rect 42012 967136 42026 967192
rect 42026 967136 42076 967192
rect 42012 967132 42076 967136
rect 675340 966512 675404 966516
rect 675340 966456 675390 966512
rect 675390 966456 675404 966512
rect 675340 966452 675404 966456
rect 676076 965092 676140 965156
rect 675156 963384 675220 963388
rect 675156 963328 675206 963384
rect 675206 963328 675220 963384
rect 675156 963324 675220 963328
rect 41828 962160 41892 962164
rect 41828 962104 41842 962160
rect 41842 962104 41892 962160
rect 41828 962100 41892 962104
rect 676628 961964 676692 962028
rect 675156 959380 675220 959444
rect 41276 959108 41340 959172
rect 676996 958292 677060 958356
rect 40724 956524 40788 956588
rect 676812 956388 676876 956452
rect 40540 955436 40604 955500
rect 41644 952444 41708 952508
rect 41460 952172 41524 952236
rect 41276 951628 41340 951692
rect 42012 951628 42076 951692
rect 676628 951492 676692 951556
rect 676076 949996 676140 950060
rect 675340 948908 675404 948972
rect 41828 938980 41892 939044
rect 41828 936532 41892 936596
rect 676812 931908 676876 931972
rect 676996 930684 677060 930748
rect 676076 877100 676140 877164
rect 676812 876420 676876 876484
rect 675340 874032 675404 874036
rect 675340 873976 675390 874032
rect 675390 873976 675404 874032
rect 675340 873972 675404 873976
rect 675892 869620 675956 869684
rect 675340 869484 675404 869548
rect 42012 813180 42076 813244
rect 40540 810698 40604 810762
rect 42012 808284 42076 808348
rect 40724 805292 40788 805356
rect 40908 805020 40972 805084
rect 42012 805020 42076 805084
rect 41644 804748 41708 804812
rect 41828 803796 41892 803860
rect 42380 801136 42444 801140
rect 42380 801080 42394 801136
rect 42394 801080 42444 801136
rect 42380 801076 42444 801080
rect 41092 800940 41156 801004
rect 40356 800668 40420 800732
rect 40356 796180 40420 796244
rect 41092 794412 41156 794476
rect 40908 793460 40972 793524
rect 42380 792916 42444 792980
rect 40724 791964 40788 792028
rect 40540 790060 40604 790124
rect 41644 789108 41708 789172
rect 41828 788428 41892 788492
rect 41460 788156 41524 788220
rect 674236 784212 674300 784276
rect 674604 783940 674668 784004
rect 676076 772652 676140 772716
rect 41460 769796 41524 769860
rect 675892 768708 675956 768772
rect 675708 766532 675772 766596
rect 40908 765716 40972 765780
rect 40540 765308 40604 765372
rect 40724 764900 40788 764964
rect 41644 759596 41708 759660
rect 42196 758432 42260 758436
rect 42196 758376 42246 758432
rect 42246 758376 42260 758432
rect 42196 758372 42260 758376
rect 41828 757692 41892 757756
rect 42012 757012 42076 757076
rect 675892 757012 675956 757076
rect 42012 755440 42076 755444
rect 42012 755384 42026 755440
rect 42026 755384 42076 755440
rect 42012 755380 42076 755384
rect 42196 754896 42260 754900
rect 42196 754840 42210 754896
rect 42210 754840 42260 754896
rect 42196 754836 42260 754840
rect 675892 752388 675956 752452
rect 40724 752116 40788 752180
rect 40908 751028 40972 751092
rect 40540 749396 40604 749460
rect 41460 746540 41524 746604
rect 41644 746268 41708 746332
rect 41828 745044 41892 745108
rect 674420 738108 674484 738172
rect 677180 732940 677244 733004
rect 676260 728044 676324 728108
rect 674236 727772 674300 727836
rect 41828 725792 41892 725796
rect 41828 725736 41842 725792
rect 41842 725736 41892 725792
rect 41828 725732 41892 725736
rect 40724 721708 40788 721772
rect 40908 721708 40972 721772
rect 41644 721708 41708 721772
rect 676076 721516 676140 721580
rect 40540 718524 40604 718588
rect 41828 716756 41892 716820
rect 42564 714716 42628 714780
rect 41092 714172 41156 714236
rect 676812 713488 676876 713492
rect 676812 713432 676826 713488
rect 676826 713432 676876 713488
rect 676812 713428 676876 713432
rect 42564 711588 42628 711652
rect 41092 709820 41156 709884
rect 674604 708732 674668 708796
rect 40908 708460 40972 708524
rect 40724 707372 40788 707436
rect 673316 706284 673380 706348
rect 40540 706148 40604 706212
rect 41460 703700 41524 703764
rect 41644 702340 41708 702404
rect 41828 701796 41892 701860
rect 674604 698532 674668 698596
rect 675340 696824 675404 696828
rect 675340 696768 675390 696824
rect 675390 696768 675404 696824
rect 675340 696764 675404 696768
rect 676812 694044 676876 694108
rect 675340 685204 675404 685268
rect 41828 682408 41892 682412
rect 41828 682352 41842 682408
rect 41842 682352 41892 682408
rect 41828 682348 41892 682352
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 41828 678872 41892 678876
rect 41828 678816 41842 678872
rect 41842 678816 41892 678872
rect 41828 678812 41892 678816
rect 676076 678268 676140 678332
rect 674420 674052 674484 674116
rect 41828 672692 41892 672756
rect 41092 672480 41156 672484
rect 41092 672424 41142 672480
rect 41142 672424 41156 672480
rect 41092 672420 41156 672424
rect 42196 672208 42260 672212
rect 42196 672152 42246 672208
rect 42246 672152 42260 672208
rect 42196 672148 42260 672152
rect 41092 669020 41156 669084
rect 42196 667388 42260 667452
rect 676996 665348 677060 665412
rect 40724 664124 40788 664188
rect 40540 662764 40604 662828
rect 41460 660316 41524 660380
rect 41644 658820 41708 658884
rect 41828 658548 41892 658612
rect 675524 652896 675588 652900
rect 675524 652840 675574 652896
rect 675574 652840 675588 652896
rect 675524 652836 675588 652840
rect 674420 648620 674484 648684
rect 675340 645824 675404 645828
rect 675340 645768 675354 645824
rect 675354 645768 675404 645824
rect 675340 645764 675404 645768
rect 41460 640596 41524 640660
rect 675340 637800 675404 637804
rect 675340 637744 675354 637800
rect 675354 637744 675404 637800
rect 675340 637740 675404 637744
rect 675524 637664 675588 637668
rect 675524 637608 675574 637664
rect 675574 637608 675588 637664
rect 675524 637604 675588 637608
rect 41644 637332 41708 637396
rect 40540 636924 40604 636988
rect 40908 636108 40972 636172
rect 40724 635700 40788 635764
rect 41828 635292 41892 635356
rect 676076 631348 676140 631412
rect 40908 625364 40972 625428
rect 672948 625092 673012 625156
rect 674604 621012 674668 621076
rect 40724 619788 40788 619852
rect 676812 619108 676876 619172
rect 40540 618972 40604 619036
rect 41828 618700 41892 618764
rect 41460 615980 41524 616044
rect 41828 612776 41892 612780
rect 41828 612720 41842 612776
rect 41842 612720 41892 612776
rect 41828 612716 41892 612720
rect 674236 607820 674300 607884
rect 677180 607276 677244 607340
rect 674604 602924 674668 602988
rect 674972 597680 675036 597684
rect 674972 597624 674986 597680
rect 674986 597624 675036 597680
rect 674972 597620 675036 597624
rect 42196 596396 42260 596460
rect 42012 595716 42076 595780
rect 41828 593948 41892 594012
rect 674972 592452 675036 592516
rect 40724 589656 40788 589660
rect 40724 589600 40774 589656
rect 40774 589600 40788 589656
rect 40724 589596 40788 589600
rect 40908 589460 40972 589524
rect 676076 589188 676140 589252
rect 41828 587148 41892 587212
rect 42196 586604 42260 586668
rect 672948 586196 673012 586260
rect 676076 586196 676140 586260
rect 41092 585788 41156 585852
rect 41276 585516 41340 585580
rect 42380 585440 42444 585444
rect 42380 585384 42430 585440
rect 42430 585384 42444 585440
rect 42380 585380 42444 585384
rect 40356 584564 40420 584628
rect 41276 582524 41340 582588
rect 42380 581632 42444 581636
rect 42380 581576 42430 581632
rect 42430 581576 42444 581632
rect 42380 581572 42444 581576
rect 41092 581436 41156 581500
rect 40908 580076 40972 580140
rect 40356 579804 40420 579868
rect 40724 579532 40788 579596
rect 42380 579532 42444 579596
rect 42196 577008 42260 577012
rect 42196 576952 42210 577008
rect 42210 576952 42260 577008
rect 42196 576948 42260 576952
rect 40540 575588 40604 575652
rect 42380 574636 42444 574700
rect 674420 573276 674484 573340
rect 41460 572732 41524 572796
rect 41644 572052 41708 572116
rect 41828 570208 41892 570212
rect 41828 570152 41842 570208
rect 41842 570152 41892 570208
rect 41828 570148 41892 570152
rect 675340 561912 675404 561916
rect 675340 561856 675390 561912
rect 675390 561856 675404 561912
rect 675340 561852 675404 561856
rect 675524 559464 675588 559468
rect 675524 559408 675538 559464
rect 675538 559408 675588 559464
rect 675524 559404 675588 559408
rect 676812 558996 676876 559060
rect 42196 553964 42260 554028
rect 42380 552740 42444 552804
rect 676996 552060 677060 552124
rect 42012 550292 42076 550356
rect 675524 549672 675588 549676
rect 675524 549616 675538 549672
rect 675538 549616 675588 549672
rect 675524 549612 675588 549616
rect 675340 547844 675404 547908
rect 677180 547572 677244 547636
rect 674236 547028 674300 547092
rect 676076 546756 676140 546820
rect 41644 546348 41708 546412
rect 42380 546348 42444 546412
rect 41828 545804 41892 545868
rect 40724 545532 40788 545596
rect 40540 545260 40604 545324
rect 40908 538188 40972 538252
rect 40724 535196 40788 535260
rect 40540 533292 40604 533356
rect 41460 530164 41524 530228
rect 41828 529756 41892 529820
rect 41828 529408 41892 529412
rect 41828 529352 41842 529408
rect 41842 529352 41892 529408
rect 41828 529348 41892 529352
rect 674604 527036 674668 527100
rect 673868 524452 673932 524516
rect 675892 484740 675956 484804
rect 675892 483924 675956 483988
rect 673316 474812 673380 474876
rect 41828 426396 41892 426460
rect 41828 425580 41892 425644
rect 40724 422248 40788 422312
rect 42012 421908 42076 421972
rect 41828 421152 41892 421156
rect 41828 421096 41842 421152
rect 41842 421096 41892 421152
rect 41828 421092 41892 421096
rect 40540 418644 40604 418708
rect 42012 418644 42076 418708
rect 40724 407492 40788 407556
rect 40540 403820 40604 403884
rect 41828 401976 41892 401980
rect 41828 401920 41842 401976
rect 41842 401920 41892 401976
rect 41828 401916 41892 401920
rect 41460 400012 41524 400076
rect 41828 398848 41892 398852
rect 41828 398792 41878 398848
rect 41878 398792 41892 398848
rect 41828 398788 41892 398792
rect 676076 398788 676140 398852
rect 676260 396748 676324 396812
rect 676628 395116 676692 395180
rect 676444 394708 676508 394772
rect 672948 393212 673012 393276
rect 675892 388452 675956 388516
rect 675708 387636 675772 387700
rect 676260 383556 676324 383620
rect 41460 382196 41524 382260
rect 675708 382256 675772 382260
rect 675708 382200 675758 382256
rect 675758 382200 675772 382256
rect 675708 382196 675772 382200
rect 676444 380564 676508 380628
rect 41644 380156 41708 380220
rect 40908 379340 40972 379404
rect 41828 378932 41892 378996
rect 40540 378524 40604 378588
rect 675892 378524 675956 378588
rect 40724 378116 40788 378180
rect 674788 377708 674852 377772
rect 676628 377300 676692 377364
rect 676076 374988 676140 375052
rect 674788 372540 674852 372604
rect 40908 365604 40972 365668
rect 40724 363700 40788 363764
rect 40540 360572 40604 360636
rect 41828 358728 41892 358732
rect 41828 358672 41878 358728
rect 41878 358672 41892 358728
rect 41828 358668 41892 358672
rect 41460 356900 41524 356964
rect 42012 355736 42076 355740
rect 42012 355680 42026 355736
rect 42026 355680 42076 355736
rect 42012 355676 42076 355680
rect 675340 354180 675404 354244
rect 675524 352956 675588 353020
rect 675708 352140 675772 352204
rect 675892 351868 675956 351932
rect 676444 346564 676508 346628
rect 676628 346488 676692 346492
rect 676628 346432 676642 346488
rect 676642 346432 676692 346488
rect 676628 346428 676692 346432
rect 676260 340172 676324 340236
rect 41460 339764 41524 339828
rect 41828 339492 41892 339556
rect 675340 339008 675404 339012
rect 675340 338952 675390 339008
rect 675390 338952 675404 339008
rect 675340 338948 675404 338952
rect 41644 338540 41708 338604
rect 675892 337724 675956 337788
rect 40540 337316 40604 337380
rect 40724 336092 40788 336156
rect 676444 335276 676508 335340
rect 676628 331196 676692 331260
rect 676076 326844 676140 326908
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 40724 322764 40788 322828
rect 41828 315616 41892 315620
rect 41828 315560 41842 315616
rect 41842 315560 41892 315616
rect 41828 315556 41892 315560
rect 41460 313652 41524 313716
rect 40540 312972 40604 313036
rect 675524 308756 675588 308820
rect 675708 305900 675772 305964
rect 676076 302968 676140 302972
rect 676076 302912 676090 302968
rect 676090 302912 676140 302968
rect 676076 302908 676140 302912
rect 676628 301548 676692 301612
rect 675892 299372 675956 299436
rect 675708 297332 675772 297396
rect 41828 296788 41892 296852
rect 42012 296380 42076 296444
rect 40540 292588 40604 292592
rect 40540 292532 40554 292588
rect 40554 292532 40604 292588
rect 40540 292528 40604 292532
rect 40724 292528 40788 292592
rect 40908 292528 40972 292592
rect 41828 292088 41892 292092
rect 41828 292032 41842 292088
rect 41842 292032 41892 292088
rect 41828 292028 41892 292032
rect 676444 291484 676508 291548
rect 676260 290940 676324 291004
rect 676628 286996 676692 287060
rect 676076 283596 676140 283660
rect 675892 282780 675956 282844
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 42012 281480 42076 281484
rect 42012 281424 42026 281480
rect 42026 281424 42076 281480
rect 42012 281420 42076 281424
rect 40908 278700 40972 278764
rect 673132 278760 673196 278764
rect 673132 278704 673146 278760
rect 673146 278704 673196 278760
rect 673132 278700 673196 278704
rect 673868 278564 673932 278628
rect 673868 277612 673932 277676
rect 40724 277340 40788 277404
rect 665404 273668 665468 273732
rect 665772 273728 665836 273732
rect 665772 273672 665786 273728
rect 665786 273672 665836 273728
rect 665772 273668 665836 273672
rect 665588 273456 665652 273460
rect 665588 273400 665602 273456
rect 665602 273400 665652 273456
rect 665588 273396 665652 273400
rect 40540 272988 40604 273052
rect 41828 272368 41892 272372
rect 41828 272312 41842 272368
rect 41842 272312 41892 272368
rect 41828 272308 41892 272312
rect 489868 271628 489932 271692
rect 490052 270540 490116 270604
rect 41460 270404 41524 270468
rect 676076 263604 676140 263668
rect 676996 261564 677060 261628
rect 676812 260748 676876 260812
rect 674972 252588 675036 252652
rect 676996 250140 677060 250204
rect 40540 249732 40604 249796
rect 673868 249656 673932 249660
rect 673868 249600 673918 249656
rect 673918 249600 673932 249656
rect 673868 249596 673932 249600
rect 674788 249596 674852 249660
rect 676076 249596 676140 249660
rect 40724 246876 40788 246940
rect 676812 246604 676876 246668
rect 675524 245984 675588 245988
rect 675524 245928 675538 245984
rect 675538 245928 675588 245984
rect 675524 245924 675588 245928
rect 668164 245788 668228 245852
rect 666692 245712 666756 245716
rect 666692 245656 666742 245712
rect 666742 245656 666756 245712
rect 666692 245652 666756 245656
rect 667980 245712 668044 245716
rect 667980 245656 668030 245712
rect 668030 245656 668044 245712
rect 667980 245652 668044 245656
rect 666508 245380 666572 245444
rect 675340 238640 675404 238644
rect 675340 238584 675390 238640
rect 675390 238584 675404 238640
rect 675340 238580 675404 238584
rect 40724 238444 40788 238508
rect 42012 237628 42076 237692
rect 42380 237416 42444 237420
rect 42380 237360 42430 237416
rect 42430 237360 42444 237416
rect 42380 237356 42444 237360
rect 40540 236540 40604 236604
rect 42012 228984 42076 228988
rect 42012 228928 42026 228984
rect 42026 228928 42076 228984
rect 42012 228924 42076 228928
rect 42380 227292 42444 227356
rect 503484 219948 503548 220012
rect 574140 219948 574204 220012
rect 559788 219132 559852 219196
rect 571932 219132 571996 219196
rect 675156 218996 675220 219060
rect 675524 218588 675588 218652
rect 542124 217662 542188 217666
rect 542124 217606 542138 217662
rect 542138 217606 542188 217662
rect 542124 217602 542188 217606
rect 541204 217560 541268 217564
rect 541204 217504 541218 217560
rect 541218 217504 541268 217560
rect 541204 217500 541268 217504
rect 542492 217560 542556 217564
rect 542492 217504 542496 217560
rect 542496 217504 542552 217560
rect 542552 217504 542556 217560
rect 542492 217500 542556 217504
rect 542676 217500 542740 217564
rect 560156 217832 560220 217836
rect 560156 217776 560170 217832
rect 560170 217776 560220 217832
rect 560156 217772 560220 217776
rect 563468 217832 563532 217836
rect 563468 217776 563482 217832
rect 563482 217776 563532 217832
rect 563468 217772 563532 217776
rect 572852 217772 572916 217836
rect 675340 217772 675404 217836
rect 673316 217364 673380 217428
rect 675708 216548 675772 216612
rect 546724 216472 546788 216476
rect 546724 216416 546774 216472
rect 546774 216416 546788 216472
rect 546724 216412 546788 216416
rect 542492 216140 542556 216204
rect 559788 216140 559852 216204
rect 560156 216140 560220 216204
rect 541204 215868 541268 215932
rect 546724 215868 546788 215932
rect 563468 215868 563532 215932
rect 673500 215596 673564 215660
rect 673684 215384 673748 215388
rect 673684 215328 673734 215384
rect 673734 215328 673748 215384
rect 673684 215324 673748 215328
rect 675892 214916 675956 214980
rect 673132 214568 673196 214572
rect 673132 214512 673146 214568
rect 673146 214512 673196 214568
rect 673132 214508 673196 214512
rect 675892 214508 675956 214572
rect 670740 212604 670804 212668
rect 670924 210488 670988 210492
rect 670924 210432 670938 210488
rect 670938 210432 670988 210488
rect 670924 210428 670988 210432
rect 675156 210156 675220 210220
rect 675892 210156 675956 210220
rect 41828 210020 41892 210084
rect 669820 209612 669884 209676
rect 41460 208932 41524 208996
rect 665588 208796 665652 208860
rect 40908 208116 40972 208180
rect 40540 207708 40604 207772
rect 669636 208312 669700 208316
rect 669636 208256 669650 208312
rect 669650 208256 669700 208312
rect 669636 208252 669700 208256
rect 40724 206076 40788 206140
rect 669268 205396 669332 205460
rect 669636 205396 669700 205460
rect 676260 204988 676324 205052
rect 666508 204172 666572 204236
rect 675892 204172 675956 204236
rect 675340 202736 675404 202740
rect 675340 202680 675390 202736
rect 675390 202680 675404 202736
rect 675340 202676 675404 202680
rect 668164 202268 668228 202332
rect 41644 202132 41708 202196
rect 674788 200772 674852 200836
rect 676444 199956 676508 200020
rect 666508 199276 666572 199340
rect 676812 198596 676876 198660
rect 40908 197100 40972 197164
rect 676628 197100 676692 197164
rect 669268 196148 669332 196212
rect 669636 196148 669700 196212
rect 669268 195876 669332 195940
rect 669636 195876 669700 195940
rect 41828 195256 41892 195260
rect 41828 195200 41842 195256
rect 41842 195200 41892 195256
rect 41828 195196 41892 195200
rect 667980 194108 668044 194172
rect 675524 193564 675588 193628
rect 676076 193156 676140 193220
rect 666876 192544 666940 192608
rect 40724 191524 40788 191588
rect 675524 191584 675588 191588
rect 675524 191528 675538 191584
rect 675538 191528 675588 191584
rect 675524 191524 675588 191528
rect 666692 189280 666756 189344
rect 669268 186356 669332 186420
rect 669636 186356 669700 186420
rect 41828 185872 41892 185876
rect 41828 185816 41842 185872
rect 41842 185816 41892 185872
rect 41828 185812 41892 185816
rect 674788 185812 674852 185876
rect 41460 184044 41524 184108
rect 672948 183500 673012 183564
rect 40540 183364 40604 183428
rect 669452 179420 669516 179484
rect 675892 174660 675956 174724
rect 669452 174524 669516 174588
rect 675708 173572 675772 173636
rect 673132 172892 673196 172956
rect 675892 170308 675956 170372
rect 672028 168328 672092 168332
rect 672028 168272 672078 168328
rect 672078 168272 672092 168328
rect 672028 168268 672092 168272
rect 670924 167996 670988 168060
rect 675892 167452 675956 167516
rect 676444 166424 676508 166428
rect 676444 166368 676458 166424
rect 676458 166368 676508 166424
rect 676444 166364 676508 166368
rect 676628 166288 676692 166292
rect 676628 166232 676678 166288
rect 676678 166232 676692 166288
rect 676628 166228 676692 166232
rect 670740 164732 670804 164796
rect 675708 161876 675772 161940
rect 672028 159836 672092 159900
rect 676628 156300 676692 156364
rect 673684 153172 673748 153236
rect 675708 153096 675772 153100
rect 675708 153040 675722 153096
rect 675722 153040 675772 153096
rect 675708 153036 675772 153040
rect 676444 151404 676508 151468
rect 676260 150316 676324 150380
rect 673500 149636 673564 149700
rect 676076 148412 676140 148476
rect 675892 147596 675956 147660
rect 676260 128556 676324 128620
rect 675892 127196 675956 127260
rect 676812 124476 676876 124540
rect 676996 124068 677060 124132
rect 675708 122844 675772 122908
rect 675708 120260 675772 120324
rect 676076 120260 676140 120324
rect 675708 116044 675772 116108
rect 676260 114140 676324 114204
rect 676996 110332 677060 110396
rect 675892 108020 675956 108084
rect 676076 103124 676140 103188
rect 675708 102640 675772 102644
rect 675708 102584 675722 102640
rect 675722 102584 675772 102640
rect 675708 102580 675772 102584
rect 676812 101356 676876 101420
rect 637252 96868 637316 96932
rect 634676 95644 634740 95708
rect 637068 78568 637132 78572
rect 637068 78512 637118 78568
rect 637118 78512 637132 78568
rect 637068 78508 637132 78512
rect 634676 77692 634740 77756
rect 464844 51716 464908 51780
rect 525748 50492 525812 50556
rect 150388 50220 150452 50284
rect 517468 50220 517532 50284
rect 529796 50220 529860 50284
rect 78628 49736 78692 49740
rect 78628 49680 78642 49736
rect 78642 49680 78692 49736
rect 78628 49676 78692 49680
rect 411116 49132 411180 49196
rect 365484 48860 365548 48924
rect 310468 47772 310532 47836
rect 150388 47500 150452 47564
rect 78628 47228 78692 47292
rect 187556 47500 187620 47564
rect 416636 46956 416700 47020
rect 521700 46956 521764 47020
rect 361988 46412 362052 46476
rect 306972 46140 307036 46204
rect 514708 45868 514772 45932
rect 460612 45732 460676 45796
rect 520412 45052 520476 45116
rect 471652 44780 471716 44844
rect 411116 42800 411180 42804
rect 411116 42744 411130 42800
rect 411130 42744 411180 42800
rect 411116 42740 411180 42744
rect 416636 42800 416700 42804
rect 416636 42744 416650 42800
rect 416650 42744 416700 42800
rect 416636 42740 416700 42744
rect 464844 42800 464908 42804
rect 464844 42744 464894 42800
rect 464894 42744 464908 42800
rect 464844 42740 464908 42744
rect 306972 42392 307036 42396
rect 306972 42336 306976 42392
rect 306976 42336 307032 42392
rect 307032 42336 307036 42392
rect 306972 42332 307036 42336
rect 517468 42332 517532 42396
rect 187556 42120 187620 42124
rect 187556 42064 187570 42120
rect 187570 42064 187620 42120
rect 187556 42060 187620 42064
rect 310468 42120 310532 42124
rect 310468 42064 310482 42120
rect 310482 42064 310532 42120
rect 310468 42060 310532 42064
rect 361988 42120 362052 42124
rect 361988 42064 362002 42120
rect 362002 42064 362052 42120
rect 361988 42060 362052 42064
rect 365484 42060 365548 42124
rect 460612 42120 460676 42124
rect 460612 42064 460626 42120
rect 460626 42064 460676 42120
rect 460612 42060 460676 42064
rect 471652 42120 471716 42124
rect 471652 42064 471666 42120
rect 471666 42064 471716 42120
rect 471652 42060 471716 42064
rect 514708 42060 514772 42124
rect 520412 42120 520476 42124
rect 520412 42064 520462 42120
rect 520462 42064 520476 42120
rect 520412 42060 520476 42064
rect 525748 42120 525812 42124
rect 525748 42064 525798 42120
rect 525798 42064 525812 42120
rect 525748 42060 525812 42064
rect 529796 42060 529860 42124
rect 521700 41984 521764 41988
rect 521700 41928 521714 41984
rect 521714 41928 521764 41984
rect 521700 41924 521764 41928
<< metal4 >>
rect 383331 997660 383397 997661
rect 383331 997596 383332 997660
rect 383396 997596 383397 997660
rect 383331 997595 383397 997596
rect 383334 997338 383394 997595
rect 389035 997252 389101 997253
rect 389035 997188 389036 997252
rect 389100 997188 389101 997252
rect 389035 997187 389101 997188
rect 138059 996980 138125 996981
rect 138059 996916 138060 996980
rect 138124 996916 138125 996980
rect 138059 996915 138125 996916
rect 90219 996436 90285 996437
rect 90219 996372 90220 996436
rect 90284 996372 90285 996436
rect 90219 996371 90285 996372
rect 86907 996028 86973 996029
rect 86907 995964 86908 996028
rect 86972 995964 86973 996028
rect 86907 995963 86973 995964
rect 86910 995485 86970 995963
rect 90222 995485 90282 996371
rect 138062 995757 138122 996915
rect 189398 995757 189458 997102
rect 239630 995757 239690 997102
rect 242574 996845 242634 997102
rect 242571 996844 242637 996845
rect 242571 996780 242572 996844
rect 242636 996780 242637 996844
rect 242571 996779 242637 996780
rect 243310 995757 243370 997102
rect 243859 996164 243925 996165
rect 243859 996100 243860 996164
rect 243924 996100 243925 996164
rect 243859 996099 243925 996100
rect 138059 995756 138125 995757
rect 138059 995692 138060 995756
rect 138124 995692 138125 995756
rect 138059 995691 138125 995692
rect 189395 995756 189461 995757
rect 189395 995692 189396 995756
rect 189460 995692 189461 995756
rect 189395 995691 189461 995692
rect 239627 995756 239693 995757
rect 239627 995692 239628 995756
rect 239692 995692 239693 995756
rect 239627 995691 239693 995692
rect 243307 995756 243373 995757
rect 243307 995692 243308 995756
rect 243372 995692 243373 995756
rect 243307 995691 243373 995692
rect 243862 995621 243922 996099
rect 274590 995621 274650 997102
rect 295011 996436 295077 996437
rect 295011 996372 295012 996436
rect 295076 996372 295077 996436
rect 295011 996371 295077 996372
rect 295014 995757 295074 996371
rect 388118 995757 388178 997102
rect 389038 995757 389098 997187
rect 473307 996708 473373 996709
rect 473307 996644 473308 996708
rect 473372 996644 473373 996708
rect 473307 996643 473373 996644
rect 529611 996708 529677 996709
rect 529611 996644 529612 996708
rect 529676 996644 529677 996708
rect 529611 996643 529677 996644
rect 473310 995757 473370 996643
rect 529614 995757 529674 996643
rect 536606 995757 536666 997102
rect 295011 995756 295077 995757
rect 295011 995692 295012 995756
rect 295076 995692 295077 995756
rect 295011 995691 295077 995692
rect 388115 995756 388181 995757
rect 388115 995692 388116 995756
rect 388180 995692 388181 995756
rect 388115 995691 388181 995692
rect 389035 995756 389101 995757
rect 389035 995692 389036 995756
rect 389100 995692 389101 995756
rect 389035 995691 389101 995692
rect 473307 995756 473373 995757
rect 473307 995692 473308 995756
rect 473372 995692 473373 995756
rect 473307 995691 473373 995692
rect 529611 995756 529677 995757
rect 529611 995692 529612 995756
rect 529676 995692 529677 995756
rect 529611 995691 529677 995692
rect 536603 995756 536669 995757
rect 536603 995692 536604 995756
rect 536668 995692 536669 995756
rect 536603 995691 536669 995692
rect 243859 995620 243925 995621
rect 243859 995556 243860 995620
rect 243924 995556 243925 995620
rect 243859 995555 243925 995556
rect 274587 995620 274653 995621
rect 274587 995556 274588 995620
rect 274652 995556 274653 995620
rect 274587 995555 274653 995556
rect 86907 995484 86973 995485
rect 86907 995420 86908 995484
rect 86972 995420 86973 995484
rect 86907 995419 86973 995420
rect 90219 995484 90285 995485
rect 90219 995420 90220 995484
rect 90284 995420 90285 995484
rect 90219 995419 90285 995420
rect 573222 989501 573282 997102
rect 627131 996708 627197 996709
rect 627131 996644 627132 996708
rect 627196 996644 627197 996708
rect 627131 996643 627197 996644
rect 627134 995757 627194 996643
rect 630811 996436 630877 996437
rect 630811 996372 630812 996436
rect 630876 996372 630877 996436
rect 630811 996371 630877 996372
rect 627131 995756 627197 995757
rect 627131 995692 627132 995756
rect 627196 995692 627197 995756
rect 627131 995691 627197 995692
rect 630814 995485 630874 996371
rect 630811 995484 630877 995485
rect 630811 995420 630812 995484
rect 630876 995420 630877 995484
rect 630811 995419 630877 995420
rect 573219 989500 573285 989501
rect 573219 989436 573220 989500
rect 573284 989436 573285 989500
rect 573219 989435 573285 989436
rect 41459 968828 41525 968829
rect 41459 968764 41460 968828
rect 41524 968764 41525 968828
rect 41459 968763 41525 968764
rect 41275 959172 41341 959173
rect 41275 959108 41276 959172
rect 41340 959108 41341 959172
rect 41275 959107 41341 959108
rect 40723 956588 40789 956589
rect 40723 956524 40724 956588
rect 40788 956524 40789 956588
rect 40723 956523 40789 956524
rect 40539 955500 40605 955501
rect 40539 955436 40540 955500
rect 40604 955436 40605 955500
rect 40539 955435 40605 955436
rect 40542 937050 40602 955435
rect 40726 939450 40786 956523
rect 41278 951693 41338 959107
rect 41462 952237 41522 968763
rect 42011 967196 42077 967197
rect 42011 967132 42012 967196
rect 42076 967132 42077 967196
rect 42011 967131 42077 967132
rect 41827 962164 41893 962165
rect 41827 962100 41828 962164
rect 41892 962100 41893 962164
rect 41827 962099 41893 962100
rect 41830 953610 41890 962099
rect 41646 953550 41890 953610
rect 41646 952509 41706 953550
rect 41643 952508 41709 952509
rect 41643 952444 41644 952508
rect 41708 952444 41709 952508
rect 41643 952443 41709 952444
rect 41459 952236 41525 952237
rect 41459 952172 41460 952236
rect 41524 952172 41525 952236
rect 41459 952171 41525 952172
rect 42014 951693 42074 967131
rect 675339 966516 675405 966517
rect 675339 966452 675340 966516
rect 675404 966452 675405 966516
rect 675339 966451 675405 966452
rect 675155 963388 675221 963389
rect 675155 963324 675156 963388
rect 675220 963324 675221 963388
rect 675155 963323 675221 963324
rect 675158 959445 675218 963323
rect 675155 959444 675221 959445
rect 675155 959380 675156 959444
rect 675220 959380 675221 959444
rect 675155 959379 675221 959380
rect 41275 951692 41341 951693
rect 41275 951628 41276 951692
rect 41340 951628 41341 951692
rect 41275 951627 41341 951628
rect 42011 951692 42077 951693
rect 42011 951628 42012 951692
rect 42076 951628 42077 951692
rect 42011 951627 42077 951628
rect 675342 948973 675402 966451
rect 676075 965156 676141 965157
rect 676075 965092 676076 965156
rect 676140 965092 676141 965156
rect 676075 965091 676141 965092
rect 676078 950061 676138 965091
rect 676627 962028 676693 962029
rect 676627 961964 676628 962028
rect 676692 961964 676693 962028
rect 676627 961963 676693 961964
rect 676630 951557 676690 961963
rect 676995 958356 677061 958357
rect 676995 958292 676996 958356
rect 677060 958292 677061 958356
rect 676995 958291 677061 958292
rect 676811 956452 676877 956453
rect 676811 956388 676812 956452
rect 676876 956388 676877 956452
rect 676811 956387 676877 956388
rect 676627 951556 676693 951557
rect 676627 951492 676628 951556
rect 676692 951492 676693 951556
rect 676627 951491 676693 951492
rect 676075 950060 676141 950061
rect 676075 949996 676076 950060
rect 676140 949996 676141 950060
rect 676075 949995 676141 949996
rect 675339 948972 675405 948973
rect 675339 948908 675340 948972
rect 675404 948908 675405 948972
rect 675339 948907 675405 948908
rect 40726 939390 41890 939450
rect 41830 939045 41890 939390
rect 41827 939044 41893 939045
rect 41827 938980 41828 939044
rect 41892 938980 41893 939044
rect 41827 938979 41893 938980
rect 40542 936990 41890 937050
rect 41830 936597 41890 936990
rect 41827 936596 41893 936597
rect 41827 936532 41828 936596
rect 41892 936532 41893 936596
rect 41827 936531 41893 936532
rect 676814 931973 676874 956387
rect 676811 931972 676877 931973
rect 676811 931908 676812 931972
rect 676876 931908 676877 931972
rect 676811 931907 676877 931908
rect 676998 930749 677058 958291
rect 676995 930748 677061 930749
rect 676995 930684 676996 930748
rect 677060 930684 677061 930748
rect 676995 930683 677061 930684
rect 676075 877164 676141 877165
rect 676075 877100 676076 877164
rect 676140 877100 676141 877164
rect 676075 877099 676141 877100
rect 675339 874036 675405 874037
rect 675339 873972 675340 874036
rect 675404 873972 675405 874036
rect 675339 873971 675405 873972
rect 675342 869549 675402 873971
rect 675891 869684 675957 869685
rect 675891 869620 675892 869684
rect 675956 869620 675957 869684
rect 675891 869619 675957 869620
rect 675339 869548 675405 869549
rect 675339 869484 675340 869548
rect 675404 869484 675405 869548
rect 675339 869483 675405 869484
rect 42011 813244 42077 813245
rect 42011 813180 42012 813244
rect 42076 813180 42077 813244
rect 42011 813179 42077 813180
rect 40539 810762 40605 810763
rect 40539 810698 40540 810762
rect 40604 810698 40605 810762
rect 40539 810697 40605 810698
rect 40355 800732 40421 800733
rect 40355 800668 40356 800732
rect 40420 800668 40421 800732
rect 40355 800667 40421 800668
rect 40358 796245 40418 800667
rect 40355 796244 40421 796245
rect 40355 796180 40356 796244
rect 40420 796180 40421 796244
rect 40355 796179 40421 796180
rect 40542 790125 40602 810697
rect 42014 809570 42074 813179
rect 41462 809510 42074 809570
rect 40723 805356 40789 805357
rect 40723 805292 40724 805356
rect 40788 805292 40789 805356
rect 40723 805291 40789 805292
rect 40726 792029 40786 805291
rect 40907 805084 40973 805085
rect 40907 805020 40908 805084
rect 40972 805020 40973 805084
rect 40907 805019 40973 805020
rect 40910 793525 40970 805019
rect 41091 801004 41157 801005
rect 41091 800940 41092 801004
rect 41156 800940 41157 801004
rect 41091 800939 41157 800940
rect 41094 794477 41154 800939
rect 41091 794476 41157 794477
rect 41091 794412 41092 794476
rect 41156 794412 41157 794476
rect 41091 794411 41157 794412
rect 40907 793524 40973 793525
rect 40907 793460 40908 793524
rect 40972 793460 40973 793524
rect 40907 793459 40973 793460
rect 40723 792028 40789 792029
rect 40723 791964 40724 792028
rect 40788 791964 40789 792028
rect 40723 791963 40789 791964
rect 40539 790124 40605 790125
rect 40539 790060 40540 790124
rect 40604 790060 40605 790124
rect 40539 790059 40605 790060
rect 41462 788221 41522 809510
rect 42011 808348 42077 808349
rect 42011 808284 42012 808348
rect 42076 808284 42077 808348
rect 42011 808283 42077 808284
rect 42014 805085 42074 808283
rect 42011 805084 42077 805085
rect 42011 805020 42012 805084
rect 42076 805020 42077 805084
rect 42011 805019 42077 805020
rect 41643 804812 41709 804813
rect 41643 804748 41644 804812
rect 41708 804748 41709 804812
rect 41643 804747 41709 804748
rect 41646 789173 41706 804747
rect 41827 803860 41893 803861
rect 41827 803796 41828 803860
rect 41892 803796 41893 803860
rect 41827 803795 41893 803796
rect 41643 789172 41709 789173
rect 41643 789108 41644 789172
rect 41708 789108 41709 789172
rect 41643 789107 41709 789108
rect 41830 788493 41890 803795
rect 42379 801140 42445 801141
rect 42379 801076 42380 801140
rect 42444 801076 42445 801140
rect 42379 801075 42445 801076
rect 42382 792981 42442 801075
rect 42379 792980 42445 792981
rect 42379 792916 42380 792980
rect 42444 792916 42445 792980
rect 42379 792915 42445 792916
rect 41827 788492 41893 788493
rect 41827 788428 41828 788492
rect 41892 788428 41893 788492
rect 41827 788427 41893 788428
rect 41459 788220 41525 788221
rect 41459 788156 41460 788220
rect 41524 788156 41525 788220
rect 41459 788155 41525 788156
rect 674235 784276 674301 784277
rect 674235 784212 674236 784276
rect 674300 784212 674301 784276
rect 674235 784211 674301 784212
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40907 765780 40973 765781
rect 40907 765716 40908 765780
rect 40972 765716 40973 765780
rect 40907 765715 40973 765716
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40542 749461 40602 765307
rect 40723 764964 40789 764965
rect 40723 764900 40724 764964
rect 40788 764900 40789 764964
rect 40723 764899 40789 764900
rect 40726 752181 40786 764899
rect 40723 752180 40789 752181
rect 40723 752116 40724 752180
rect 40788 752116 40789 752180
rect 40723 752115 40789 752116
rect 40910 751093 40970 765715
rect 40907 751092 40973 751093
rect 40907 751028 40908 751092
rect 40972 751028 40973 751092
rect 40907 751027 40973 751028
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 41462 746605 41522 769795
rect 41643 759660 41709 759661
rect 41643 759596 41644 759660
rect 41708 759596 41709 759660
rect 41643 759595 41709 759596
rect 41459 746604 41525 746605
rect 41459 746540 41460 746604
rect 41524 746540 41525 746604
rect 41459 746539 41525 746540
rect 41646 746333 41706 759595
rect 42195 758436 42261 758437
rect 42195 758372 42196 758436
rect 42260 758372 42261 758436
rect 42195 758371 42261 758372
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41643 746332 41709 746333
rect 41643 746268 41644 746332
rect 41708 746268 41709 746332
rect 41643 746267 41709 746268
rect 41830 745109 41890 757691
rect 42011 757076 42077 757077
rect 42011 757012 42012 757076
rect 42076 757012 42077 757076
rect 42011 757011 42077 757012
rect 42014 755445 42074 757011
rect 42011 755444 42077 755445
rect 42011 755380 42012 755444
rect 42076 755380 42077 755444
rect 42011 755379 42077 755380
rect 42198 754901 42258 758371
rect 42195 754900 42261 754901
rect 42195 754836 42196 754900
rect 42260 754836 42261 754900
rect 42195 754835 42261 754836
rect 41827 745108 41893 745109
rect 41827 745044 41828 745108
rect 41892 745044 41893 745108
rect 41827 745043 41893 745044
rect 674238 727837 674298 784211
rect 674603 784004 674669 784005
rect 674603 783940 674604 784004
rect 674668 783940 674669 784004
rect 674603 783939 674669 783940
rect 674419 738172 674485 738173
rect 674419 738108 674420 738172
rect 674484 738108 674485 738172
rect 674419 738107 674485 738108
rect 674235 727836 674301 727837
rect 674235 727772 674236 727836
rect 674300 727772 674301 727836
rect 674235 727771 674301 727772
rect 41827 725796 41893 725797
rect 41827 725732 41828 725796
rect 41892 725732 41893 725796
rect 41827 725731 41893 725732
rect 41830 725250 41890 725731
rect 41462 725190 41890 725250
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40907 721772 40973 721773
rect 40907 721708 40908 721772
rect 40972 721708 40973 721772
rect 40907 721707 40973 721708
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40542 706213 40602 718523
rect 40726 707437 40786 721707
rect 40910 708525 40970 721707
rect 41091 714236 41157 714237
rect 41091 714172 41092 714236
rect 41156 714172 41157 714236
rect 41091 714171 41157 714172
rect 41094 709885 41154 714171
rect 41091 709884 41157 709885
rect 41091 709820 41092 709884
rect 41156 709820 41157 709884
rect 41091 709819 41157 709820
rect 40907 708524 40973 708525
rect 40907 708460 40908 708524
rect 40972 708460 40973 708524
rect 40907 708459 40973 708460
rect 40723 707436 40789 707437
rect 40723 707372 40724 707436
rect 40788 707372 40789 707436
rect 40723 707371 40789 707372
rect 40539 706212 40605 706213
rect 40539 706148 40540 706212
rect 40604 706148 40605 706212
rect 40539 706147 40605 706148
rect 41462 703765 41522 725190
rect 41643 721772 41709 721773
rect 41643 721708 41644 721772
rect 41708 721708 41709 721772
rect 41643 721707 41709 721708
rect 41459 703764 41525 703765
rect 41459 703700 41460 703764
rect 41524 703700 41525 703764
rect 41459 703699 41525 703700
rect 41646 702405 41706 721707
rect 41827 716820 41893 716821
rect 41827 716756 41828 716820
rect 41892 716756 41893 716820
rect 41827 716755 41893 716756
rect 41643 702404 41709 702405
rect 41643 702340 41644 702404
rect 41708 702340 41709 702404
rect 41643 702339 41709 702340
rect 41830 701861 41890 716755
rect 42563 714780 42629 714781
rect 42563 714716 42564 714780
rect 42628 714716 42629 714780
rect 42563 714715 42629 714716
rect 42566 711653 42626 714715
rect 42563 711652 42629 711653
rect 42563 711588 42564 711652
rect 42628 711588 42629 711652
rect 42563 711587 42629 711588
rect 673315 706348 673381 706349
rect 673315 706284 673316 706348
rect 673380 706284 673381 706348
rect 673315 706283 673381 706284
rect 41827 701860 41893 701861
rect 41827 701796 41828 701860
rect 41892 701796 41893 701860
rect 41827 701795 41893 701796
rect 41827 682412 41893 682413
rect 41827 682410 41828 682412
rect 41646 682350 41828 682410
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 41646 678990 41706 682350
rect 41827 682348 41828 682350
rect 41892 682348 41893 682412
rect 41827 682347 41893 682348
rect 40723 678927 40789 678928
rect 41462 678930 41706 678990
rect 40542 662829 40602 678927
rect 40726 664189 40786 678927
rect 41091 672484 41157 672485
rect 41091 672420 41092 672484
rect 41156 672420 41157 672484
rect 41091 672419 41157 672420
rect 41094 669085 41154 672419
rect 41091 669084 41157 669085
rect 41091 669020 41092 669084
rect 41156 669020 41157 669084
rect 41091 669019 41157 669020
rect 40723 664188 40789 664189
rect 40723 664124 40724 664188
rect 40788 664124 40789 664188
rect 40723 664123 40789 664124
rect 40539 662828 40605 662829
rect 40539 662764 40540 662828
rect 40604 662764 40605 662828
rect 40539 662763 40605 662764
rect 41462 660381 41522 678930
rect 41827 678876 41893 678877
rect 41827 678812 41828 678876
rect 41892 678812 41893 678876
rect 41827 678811 41893 678812
rect 41830 678330 41890 678811
rect 41646 678270 41890 678330
rect 41459 660380 41525 660381
rect 41459 660316 41460 660380
rect 41524 660316 41525 660380
rect 41459 660315 41525 660316
rect 41646 658885 41706 678270
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41643 658884 41709 658885
rect 41643 658820 41644 658884
rect 41708 658820 41709 658884
rect 41643 658819 41709 658820
rect 41830 658613 41890 672691
rect 42195 672212 42261 672213
rect 42195 672148 42196 672212
rect 42260 672148 42261 672212
rect 42195 672147 42261 672148
rect 42198 667453 42258 672147
rect 42195 667452 42261 667453
rect 42195 667388 42196 667452
rect 42260 667388 42261 667452
rect 42195 667387 42261 667388
rect 41827 658612 41893 658613
rect 41827 658548 41828 658612
rect 41892 658548 41893 658612
rect 41827 658547 41893 658548
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40539 636988 40605 636989
rect 40539 636924 40540 636988
rect 40604 636924 40605 636988
rect 40539 636923 40605 636924
rect 40542 619037 40602 636923
rect 40907 636172 40973 636173
rect 40907 636108 40908 636172
rect 40972 636108 40973 636172
rect 40907 636107 40973 636108
rect 40723 635764 40789 635765
rect 40723 635700 40724 635764
rect 40788 635700 40789 635764
rect 40723 635699 40789 635700
rect 40726 619853 40786 635699
rect 40910 625429 40970 636107
rect 40907 625428 40973 625429
rect 40907 625364 40908 625428
rect 40972 625364 40973 625428
rect 40907 625363 40973 625364
rect 40723 619852 40789 619853
rect 40723 619788 40724 619852
rect 40788 619788 40789 619852
rect 40723 619787 40789 619788
rect 40539 619036 40605 619037
rect 40539 618972 40540 619036
rect 40604 618972 40605 619036
rect 40539 618971 40605 618972
rect 41462 616045 41522 640595
rect 41643 637396 41709 637397
rect 41643 637332 41644 637396
rect 41708 637332 41709 637396
rect 41643 637331 41709 637332
rect 41646 618270 41706 637331
rect 41827 635356 41893 635357
rect 41827 635292 41828 635356
rect 41892 635292 41893 635356
rect 41827 635291 41893 635292
rect 41830 618765 41890 635291
rect 672947 625156 673013 625157
rect 672947 625092 672948 625156
rect 673012 625092 673013 625156
rect 672947 625091 673013 625092
rect 41827 618764 41893 618765
rect 41827 618700 41828 618764
rect 41892 618700 41893 618764
rect 41827 618699 41893 618700
rect 41646 618210 41890 618270
rect 41459 616044 41525 616045
rect 41459 615980 41460 616044
rect 41524 615980 41525 616044
rect 41459 615979 41525 615980
rect 41830 612781 41890 618210
rect 41827 612780 41893 612781
rect 41827 612716 41828 612780
rect 41892 612716 41893 612780
rect 41827 612715 41893 612716
rect 42195 596460 42261 596461
rect 42195 596396 42196 596460
rect 42260 596396 42261 596460
rect 42195 596395 42261 596396
rect 42011 595780 42077 595781
rect 42011 595716 42012 595780
rect 42076 595716 42077 595780
rect 42011 595715 42077 595716
rect 41827 594012 41893 594013
rect 41827 594010 41828 594012
rect 40542 593950 41828 594010
rect 40355 584628 40421 584629
rect 40355 584564 40356 584628
rect 40420 584564 40421 584628
rect 40355 584563 40421 584564
rect 40358 579869 40418 584563
rect 40355 579868 40421 579869
rect 40355 579804 40356 579868
rect 40420 579804 40421 579868
rect 40355 579803 40421 579804
rect 40542 575653 40602 593950
rect 41827 593948 41828 593950
rect 41892 593948 41893 594012
rect 41827 593947 41893 593948
rect 42014 593330 42074 595715
rect 41462 593270 42074 593330
rect 40723 589660 40789 589661
rect 40723 589596 40724 589660
rect 40788 589596 40789 589660
rect 40723 589595 40789 589596
rect 40726 579597 40786 589595
rect 40907 589524 40973 589525
rect 40907 589460 40908 589524
rect 40972 589460 40973 589524
rect 40907 589459 40973 589460
rect 40910 580141 40970 589459
rect 41091 585852 41157 585853
rect 41091 585788 41092 585852
rect 41156 585788 41157 585852
rect 41091 585787 41157 585788
rect 41094 581501 41154 585787
rect 41275 585580 41341 585581
rect 41275 585516 41276 585580
rect 41340 585516 41341 585580
rect 41275 585515 41341 585516
rect 41278 582589 41338 585515
rect 41275 582588 41341 582589
rect 41275 582524 41276 582588
rect 41340 582524 41341 582588
rect 41275 582523 41341 582524
rect 41091 581500 41157 581501
rect 41091 581436 41092 581500
rect 41156 581436 41157 581500
rect 41091 581435 41157 581436
rect 40907 580140 40973 580141
rect 40907 580076 40908 580140
rect 40972 580076 40973 580140
rect 40907 580075 40973 580076
rect 40723 579596 40789 579597
rect 40723 579532 40724 579596
rect 40788 579532 40789 579596
rect 40723 579531 40789 579532
rect 40539 575652 40605 575653
rect 40539 575588 40540 575652
rect 40604 575588 40605 575652
rect 40539 575587 40605 575588
rect 41462 572797 41522 593270
rect 42198 589290 42258 596395
rect 41646 589230 42258 589290
rect 41459 572796 41525 572797
rect 41459 572732 41460 572796
rect 41524 572732 41525 572796
rect 41459 572731 41525 572732
rect 41646 572117 41706 589230
rect 41827 587212 41893 587213
rect 41827 587148 41828 587212
rect 41892 587148 41893 587212
rect 41827 587147 41893 587148
rect 41643 572116 41709 572117
rect 41643 572052 41644 572116
rect 41708 572052 41709 572116
rect 41643 572051 41709 572052
rect 41830 570213 41890 587147
rect 42195 586668 42261 586669
rect 42195 586604 42196 586668
rect 42260 586604 42261 586668
rect 42195 586603 42261 586604
rect 42198 577013 42258 586603
rect 672950 586261 673010 625091
rect 672947 586260 673013 586261
rect 672947 586196 672948 586260
rect 673012 586196 673013 586260
rect 672947 586195 673013 586196
rect 42379 585444 42445 585445
rect 42379 585380 42380 585444
rect 42444 585380 42445 585444
rect 42379 585379 42445 585380
rect 42382 581637 42442 585379
rect 42379 581636 42445 581637
rect 42379 581572 42380 581636
rect 42444 581572 42445 581636
rect 42379 581571 42445 581572
rect 42379 579596 42445 579597
rect 42379 579532 42380 579596
rect 42444 579532 42445 579596
rect 42379 579531 42445 579532
rect 42195 577012 42261 577013
rect 42195 576948 42196 577012
rect 42260 576948 42261 577012
rect 42195 576947 42261 576948
rect 42382 574701 42442 579531
rect 42379 574700 42445 574701
rect 42379 574636 42380 574700
rect 42444 574636 42445 574700
rect 42379 574635 42445 574636
rect 41827 570212 41893 570213
rect 41827 570148 41828 570212
rect 41892 570148 41893 570212
rect 41827 570147 41893 570148
rect 42195 554028 42261 554029
rect 42195 553964 42196 554028
rect 42260 553964 42261 554028
rect 42195 553963 42261 553964
rect 42011 550356 42077 550357
rect 42011 550292 42012 550356
rect 42076 550292 42077 550356
rect 42011 550291 42077 550292
rect 42014 549130 42074 550291
rect 40910 549070 42074 549130
rect 40723 545596 40789 545597
rect 40723 545532 40724 545596
rect 40788 545532 40789 545596
rect 40723 545531 40789 545532
rect 40539 545324 40605 545325
rect 40539 545260 40540 545324
rect 40604 545260 40605 545324
rect 40539 545259 40605 545260
rect 40542 533357 40602 545259
rect 40726 535261 40786 545531
rect 40910 538253 40970 549070
rect 42198 548450 42258 553963
rect 42379 552804 42445 552805
rect 42379 552740 42380 552804
rect 42444 552740 42445 552804
rect 42379 552739 42445 552740
rect 41462 548390 42258 548450
rect 40907 538252 40973 538253
rect 40907 538188 40908 538252
rect 40972 538188 40973 538252
rect 40907 538187 40973 538188
rect 40723 535260 40789 535261
rect 40723 535196 40724 535260
rect 40788 535196 40789 535260
rect 40723 535195 40789 535196
rect 40539 533356 40605 533357
rect 40539 533292 40540 533356
rect 40604 533292 40605 533356
rect 40539 533291 40605 533292
rect 41462 530229 41522 548390
rect 42382 546413 42442 552739
rect 41643 546412 41709 546413
rect 41643 546348 41644 546412
rect 41708 546348 41709 546412
rect 41643 546347 41709 546348
rect 42379 546412 42445 546413
rect 42379 546348 42380 546412
rect 42444 546348 42445 546412
rect 42379 546347 42445 546348
rect 41459 530228 41525 530229
rect 41459 530164 41460 530228
rect 41524 530164 41525 530228
rect 41459 530163 41525 530164
rect 41646 529410 41706 546347
rect 41827 545868 41893 545869
rect 41827 545804 41828 545868
rect 41892 545804 41893 545868
rect 41827 545803 41893 545804
rect 41830 529821 41890 545803
rect 41827 529820 41893 529821
rect 41827 529756 41828 529820
rect 41892 529756 41893 529820
rect 41827 529755 41893 529756
rect 41827 529412 41893 529413
rect 41827 529410 41828 529412
rect 41646 529350 41828 529410
rect 41827 529348 41828 529350
rect 41892 529348 41893 529412
rect 41827 529347 41893 529348
rect 673318 474877 673378 706283
rect 674422 674117 674482 738107
rect 674606 708797 674666 783939
rect 675894 768773 675954 869619
rect 676078 772717 676138 877099
rect 676811 876484 676877 876485
rect 676811 876420 676812 876484
rect 676876 876420 676877 876484
rect 676811 876419 676877 876420
rect 676075 772716 676141 772717
rect 676075 772652 676076 772716
rect 676140 772652 676141 772716
rect 676075 772651 676141 772652
rect 675891 768772 675957 768773
rect 675891 768708 675892 768772
rect 675956 768708 675957 768772
rect 675891 768707 675957 768708
rect 675707 766596 675773 766597
rect 675707 766532 675708 766596
rect 675772 766532 675773 766596
rect 675707 766531 675773 766532
rect 675710 746610 675770 766531
rect 676814 761790 676874 876419
rect 675894 761730 676874 761790
rect 675894 757077 675954 761730
rect 675891 757076 675957 757077
rect 675891 757012 675892 757076
rect 675956 757012 675957 757076
rect 675891 757011 675957 757012
rect 675891 752452 675957 752453
rect 675891 752388 675892 752452
rect 675956 752450 675957 752452
rect 675956 752390 676322 752450
rect 675956 752388 675957 752390
rect 675891 752387 675957 752388
rect 676262 746610 676322 752390
rect 675710 746550 676138 746610
rect 676262 746550 676874 746610
rect 676078 730010 676138 746550
rect 676078 729950 676322 730010
rect 676262 728109 676322 729950
rect 676259 728108 676325 728109
rect 676259 728044 676260 728108
rect 676324 728044 676325 728108
rect 676259 728043 676325 728044
rect 676075 721580 676141 721581
rect 676075 721516 676076 721580
rect 676140 721516 676141 721580
rect 676075 721515 676141 721516
rect 674603 708796 674669 708797
rect 674603 708732 674604 708796
rect 674668 708732 674669 708796
rect 674603 708731 674669 708732
rect 674603 698596 674669 698597
rect 674603 698532 674604 698596
rect 674668 698532 674669 698596
rect 674603 698531 674669 698532
rect 674419 674116 674485 674117
rect 674419 674052 674420 674116
rect 674484 674052 674485 674116
rect 674419 674051 674485 674052
rect 674419 648684 674485 648685
rect 674419 648620 674420 648684
rect 674484 648620 674485 648684
rect 674419 648619 674485 648620
rect 674235 607884 674301 607885
rect 674235 607820 674236 607884
rect 674300 607820 674301 607884
rect 674235 607819 674301 607820
rect 674238 547093 674298 607819
rect 674422 573341 674482 648619
rect 674606 621077 674666 698531
rect 675339 696828 675405 696829
rect 675339 696764 675340 696828
rect 675404 696764 675405 696828
rect 675339 696763 675405 696764
rect 675342 685269 675402 696763
rect 675339 685268 675405 685269
rect 675339 685204 675340 685268
rect 675404 685204 675405 685268
rect 675339 685203 675405 685204
rect 676078 678333 676138 721515
rect 676814 713493 676874 746550
rect 677179 733004 677245 733005
rect 677179 732940 677180 733004
rect 677244 732940 677245 733004
rect 677179 732939 677245 732940
rect 677182 717630 677242 732939
rect 676998 717570 677242 717630
rect 676811 713492 676877 713493
rect 676811 713428 676812 713492
rect 676876 713428 676877 713492
rect 676811 713427 676877 713428
rect 676811 694108 676877 694109
rect 676811 694044 676812 694108
rect 676876 694044 676877 694108
rect 676811 694043 676877 694044
rect 676075 678332 676141 678333
rect 676075 678268 676076 678332
rect 676140 678268 676141 678332
rect 676075 678267 676141 678268
rect 675523 652900 675589 652901
rect 675523 652836 675524 652900
rect 675588 652836 675589 652900
rect 675523 652835 675589 652836
rect 675339 645828 675405 645829
rect 675339 645764 675340 645828
rect 675404 645764 675405 645828
rect 675339 645763 675405 645764
rect 675342 637805 675402 645763
rect 675339 637804 675405 637805
rect 675339 637740 675340 637804
rect 675404 637740 675405 637804
rect 675339 637739 675405 637740
rect 675526 637669 675586 652835
rect 675523 637668 675589 637669
rect 675523 637604 675524 637668
rect 675588 637604 675589 637668
rect 675523 637603 675589 637604
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 674603 621076 674669 621077
rect 674603 621012 674604 621076
rect 674668 621012 674669 621076
rect 674603 621011 674669 621012
rect 674603 602988 674669 602989
rect 674603 602924 674604 602988
rect 674668 602924 674669 602988
rect 674603 602923 674669 602924
rect 674419 573340 674485 573341
rect 674419 573276 674420 573340
rect 674484 573276 674485 573340
rect 674419 573275 674485 573276
rect 674235 547092 674301 547093
rect 674235 547028 674236 547092
rect 674300 547028 674301 547092
rect 674235 547027 674301 547028
rect 674606 527101 674666 602923
rect 674971 597684 675037 597685
rect 674971 597620 674972 597684
rect 675036 597620 675037 597684
rect 674971 597619 675037 597620
rect 674974 592517 675034 597619
rect 674971 592516 675037 592517
rect 674971 592452 674972 592516
rect 675036 592452 675037 592516
rect 674971 592451 675037 592452
rect 676078 589253 676138 631347
rect 676814 619173 676874 694043
rect 676998 665413 677058 717570
rect 676995 665412 677061 665413
rect 676995 665348 676996 665412
rect 677060 665348 677061 665412
rect 676995 665347 677061 665348
rect 676811 619172 676877 619173
rect 676811 619108 676812 619172
rect 676876 619108 676877 619172
rect 676811 619107 676877 619108
rect 677179 607340 677245 607341
rect 677179 607276 677180 607340
rect 677244 607276 677245 607340
rect 677179 607275 677245 607276
rect 676075 589252 676141 589253
rect 676075 589188 676076 589252
rect 676140 589188 676141 589252
rect 676075 589187 676141 589188
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675339 561916 675405 561917
rect 675339 561852 675340 561916
rect 675404 561852 675405 561916
rect 675339 561851 675405 561852
rect 675342 547909 675402 561851
rect 675523 559468 675589 559469
rect 675523 559404 675524 559468
rect 675588 559404 675589 559468
rect 675523 559403 675589 559404
rect 675526 549677 675586 559403
rect 675523 549676 675589 549677
rect 675523 549612 675524 549676
rect 675588 549612 675589 549676
rect 675523 549611 675589 549612
rect 675339 547908 675405 547909
rect 675339 547844 675340 547908
rect 675404 547844 675405 547908
rect 675339 547843 675405 547844
rect 676078 546821 676138 586195
rect 676811 559060 676877 559061
rect 676811 558996 676812 559060
rect 676876 558996 676877 559060
rect 676811 558995 676877 558996
rect 676075 546820 676141 546821
rect 676075 546756 676076 546820
rect 676140 546756 676141 546820
rect 676075 546755 676141 546756
rect 674603 527100 674669 527101
rect 674603 527036 674604 527100
rect 674668 527036 674669 527100
rect 674603 527035 674669 527036
rect 673867 524516 673933 524517
rect 673867 524452 673868 524516
rect 673932 524452 673933 524516
rect 673867 524451 673933 524452
rect 673315 474876 673381 474877
rect 673315 474812 673316 474876
rect 673380 474812 673381 474876
rect 673315 474811 673381 474812
rect 41827 426460 41893 426461
rect 41827 426396 41828 426460
rect 41892 426396 41893 426460
rect 41827 426395 41893 426396
rect 41830 426050 41890 426395
rect 41462 425990 41890 426050
rect 40723 422312 40789 422313
rect 40723 422248 40724 422312
rect 40788 422248 40789 422312
rect 40723 422247 40789 422248
rect 40539 418708 40605 418709
rect 40539 418644 40540 418708
rect 40604 418644 40605 418708
rect 40539 418643 40605 418644
rect 40542 403885 40602 418643
rect 40726 407557 40786 422247
rect 40723 407556 40789 407557
rect 40723 407492 40724 407556
rect 40788 407492 40789 407556
rect 40723 407491 40789 407492
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 400077 41522 425990
rect 41827 425644 41893 425645
rect 41827 425580 41828 425644
rect 41892 425580 41893 425644
rect 41827 425579 41893 425580
rect 41830 425370 41890 425579
rect 41646 425310 41890 425370
rect 41459 400076 41525 400077
rect 41459 400012 41460 400076
rect 41524 400012 41525 400076
rect 41459 400011 41525 400012
rect 41646 398850 41706 425310
rect 42011 421972 42077 421973
rect 42011 421908 42012 421972
rect 42076 421908 42077 421972
rect 42011 421907 42077 421908
rect 41827 421156 41893 421157
rect 41827 421092 41828 421156
rect 41892 421092 41893 421156
rect 41827 421091 41893 421092
rect 41830 401981 41890 421091
rect 42014 418709 42074 421907
rect 42011 418708 42077 418709
rect 42011 418644 42012 418708
rect 42076 418644 42077 418708
rect 42011 418643 42077 418644
rect 41827 401980 41893 401981
rect 41827 401916 41828 401980
rect 41892 401916 41893 401980
rect 41827 401915 41893 401916
rect 41827 398852 41893 398853
rect 41827 398850 41828 398852
rect 41646 398790 41828 398850
rect 41827 398788 41828 398790
rect 41892 398788 41893 398852
rect 41827 398787 41893 398788
rect 672947 393276 673013 393277
rect 672947 393212 672948 393276
rect 673012 393212 673013 393276
rect 672947 393211 673013 393212
rect 41459 382260 41525 382261
rect 41459 382196 41460 382260
rect 41524 382196 41525 382260
rect 41459 382195 41525 382196
rect 40907 379404 40973 379405
rect 40907 379340 40908 379404
rect 40972 379340 40973 379404
rect 40907 379339 40973 379340
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40542 360637 40602 378523
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363765 40786 378115
rect 40910 365669 40970 379339
rect 40907 365668 40973 365669
rect 40907 365604 40908 365668
rect 40972 365604 40973 365668
rect 40907 365603 40973 365604
rect 40723 363764 40789 363765
rect 40723 363700 40724 363764
rect 40788 363700 40789 363764
rect 40723 363699 40789 363700
rect 40539 360636 40605 360637
rect 40539 360572 40540 360636
rect 40604 360572 40605 360636
rect 40539 360571 40605 360572
rect 41462 356965 41522 382195
rect 41643 380220 41709 380221
rect 41643 380156 41644 380220
rect 41708 380156 41709 380220
rect 41643 380155 41709 380156
rect 41646 358730 41706 380155
rect 41827 378996 41893 378997
rect 41827 378932 41828 378996
rect 41892 378932 41893 378996
rect 41827 378931 41893 378932
rect 41830 364350 41890 378931
rect 41830 364290 42074 364350
rect 41827 358732 41893 358733
rect 41827 358730 41828 358732
rect 41646 358670 41828 358730
rect 41827 358668 41828 358670
rect 41892 358668 41893 358732
rect 41827 358667 41893 358668
rect 41459 356964 41525 356965
rect 41459 356900 41460 356964
rect 41524 356900 41525 356964
rect 41459 356899 41525 356900
rect 42014 355741 42074 364290
rect 42011 355740 42077 355741
rect 42011 355676 42012 355740
rect 42076 355676 42077 355740
rect 42011 355675 42077 355676
rect 41459 339828 41525 339829
rect 41459 339764 41460 339828
rect 41524 339764 41525 339828
rect 41459 339763 41525 339764
rect 40539 337380 40605 337381
rect 40539 337316 40540 337380
rect 40604 337316 40605 337380
rect 40539 337315 40605 337316
rect 40542 313037 40602 337315
rect 40723 336156 40789 336157
rect 40723 336092 40724 336156
rect 40788 336092 40789 336156
rect 40723 336091 40789 336092
rect 40726 322829 40786 336091
rect 40723 322828 40789 322829
rect 40723 322764 40724 322828
rect 40788 322764 40789 322828
rect 40723 322763 40789 322764
rect 41462 313717 41522 339763
rect 41827 339556 41893 339557
rect 41827 339492 41828 339556
rect 41892 339492 41893 339556
rect 41827 339491 41893 339492
rect 41643 338604 41709 338605
rect 41643 338540 41644 338604
rect 41708 338540 41709 338604
rect 41643 338539 41709 338540
rect 41646 316050 41706 338539
rect 41830 324869 41890 339491
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41646 315990 41890 316050
rect 41830 315621 41890 315990
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 41459 313716 41525 313717
rect 41459 313652 41460 313716
rect 41524 313652 41525 313716
rect 41459 313651 41525 313652
rect 40539 313036 40605 313037
rect 40539 312972 40540 313036
rect 40604 312972 40605 313036
rect 40539 312971 40605 312972
rect 41827 296852 41893 296853
rect 41827 296788 41828 296852
rect 41892 296788 41893 296852
rect 41827 296787 41893 296788
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40723 292592 40789 292593
rect 40723 292528 40724 292592
rect 40788 292528 40789 292592
rect 40723 292527 40789 292528
rect 40907 292592 40973 292593
rect 40907 292528 40908 292592
rect 40972 292528 40973 292592
rect 41830 292590 41890 296787
rect 42011 296444 42077 296445
rect 42011 296380 42012 296444
rect 42076 296380 42077 296444
rect 42011 296379 42077 296380
rect 40907 292527 40973 292528
rect 41462 292530 41890 292590
rect 40542 273053 40602 292527
rect 40726 277405 40786 292527
rect 40910 278765 40970 292527
rect 40907 278764 40973 278765
rect 40907 278700 40908 278764
rect 40972 278700 40973 278764
rect 40907 278699 40973 278700
rect 40723 277404 40789 277405
rect 40723 277340 40724 277404
rect 40788 277340 40789 277404
rect 40723 277339 40789 277340
rect 40539 273052 40605 273053
rect 40539 272988 40540 273052
rect 40604 272988 40605 273052
rect 40539 272987 40605 272988
rect 41462 270469 41522 292530
rect 41827 292092 41893 292093
rect 41827 292028 41828 292092
rect 41892 292028 41893 292092
rect 41827 292027 41893 292028
rect 41830 272373 41890 292027
rect 42014 281485 42074 296379
rect 672950 287070 673010 393211
rect 672950 287010 673194 287070
rect 42011 281484 42077 281485
rect 42011 281420 42012 281484
rect 42076 281420 42077 281484
rect 42011 281419 42077 281420
rect 673134 278765 673194 287010
rect 673131 278764 673197 278765
rect 673131 278700 673132 278764
rect 673196 278700 673197 278764
rect 673131 278699 673197 278700
rect 673870 278629 673930 524451
rect 676814 485210 676874 558995
rect 676995 552124 677061 552125
rect 676995 552060 676996 552124
rect 677060 552060 677061 552124
rect 676995 552059 677061 552060
rect 675894 485150 676874 485210
rect 675894 484805 675954 485150
rect 675891 484804 675957 484805
rect 675891 484740 675892 484804
rect 675956 484740 675957 484804
rect 675891 484739 675957 484740
rect 676998 484530 677058 552059
rect 677182 547637 677242 607275
rect 677179 547636 677245 547637
rect 677179 547572 677180 547636
rect 677244 547572 677245 547636
rect 677179 547571 677245 547572
rect 675894 484470 677058 484530
rect 675894 483989 675954 484470
rect 675891 483988 675957 483989
rect 675891 483924 675892 483988
rect 675956 483924 675957 483988
rect 675891 483923 675957 483924
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 388516 675957 388517
rect 675891 388452 675892 388516
rect 675956 388452 675957 388516
rect 675891 388451 675957 388452
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675710 382261 675770 387635
rect 675707 382260 675773 382261
rect 675707 382196 675708 382260
rect 675772 382196 675773 382260
rect 675707 382195 675773 382196
rect 675894 378589 675954 388451
rect 675891 378588 675957 378589
rect 675891 378524 675892 378588
rect 675956 378524 675957 378588
rect 675891 378523 675957 378524
rect 674787 377772 674853 377773
rect 674787 377708 674788 377772
rect 674852 377708 674853 377772
rect 674787 377707 674853 377708
rect 674790 372605 674850 377707
rect 676078 375053 676138 398787
rect 676259 396812 676325 396813
rect 676259 396748 676260 396812
rect 676324 396748 676325 396812
rect 676259 396747 676325 396748
rect 676262 383621 676322 396747
rect 676627 395180 676693 395181
rect 676627 395116 676628 395180
rect 676692 395116 676693 395180
rect 676627 395115 676693 395116
rect 676443 394772 676509 394773
rect 676443 394708 676444 394772
rect 676508 394708 676509 394772
rect 676443 394707 676509 394708
rect 676259 383620 676325 383621
rect 676259 383556 676260 383620
rect 676324 383556 676325 383620
rect 676259 383555 676325 383556
rect 676446 380629 676506 394707
rect 676443 380628 676509 380629
rect 676443 380564 676444 380628
rect 676508 380564 676509 380628
rect 676443 380563 676509 380564
rect 676630 377365 676690 395115
rect 676627 377364 676693 377365
rect 676627 377300 676628 377364
rect 676692 377300 676693 377364
rect 676627 377299 676693 377300
rect 676075 375052 676141 375053
rect 676075 374988 676076 375052
rect 676140 374988 676141 375052
rect 676075 374987 676141 374988
rect 674787 372604 674853 372605
rect 674787 372540 674788 372604
rect 674852 372540 674853 372604
rect 674787 372539 674853 372540
rect 675339 354244 675405 354245
rect 675339 354180 675340 354244
rect 675404 354180 675405 354244
rect 675339 354179 675405 354180
rect 675342 339013 675402 354179
rect 675523 353020 675589 353021
rect 675523 352956 675524 353020
rect 675588 352956 675589 353020
rect 675523 352955 675589 352956
rect 675526 340890 675586 352955
rect 675707 352204 675773 352205
rect 675707 352140 675708 352204
rect 675772 352140 675773 352204
rect 675707 352139 675773 352140
rect 675710 350550 675770 352139
rect 675891 351932 675957 351933
rect 675891 351868 675892 351932
rect 675956 351930 675957 351932
rect 675956 351870 676322 351930
rect 675956 351868 675957 351870
rect 675891 351867 675957 351868
rect 675710 350490 676138 350550
rect 675526 340830 675954 340890
rect 675339 339012 675405 339013
rect 675339 338948 675340 339012
rect 675404 338948 675405 339012
rect 675339 338947 675405 338948
rect 675894 337789 675954 340830
rect 675891 337788 675957 337789
rect 675891 337724 675892 337788
rect 675956 337724 675957 337788
rect 675891 337723 675957 337724
rect 676078 326909 676138 350490
rect 676262 340237 676322 351870
rect 676443 346628 676509 346629
rect 676443 346564 676444 346628
rect 676508 346564 676509 346628
rect 676443 346563 676509 346564
rect 676259 340236 676325 340237
rect 676259 340172 676260 340236
rect 676324 340172 676325 340236
rect 676259 340171 676325 340172
rect 676446 335341 676506 346563
rect 676627 346492 676693 346493
rect 676627 346428 676628 346492
rect 676692 346428 676693 346492
rect 676627 346427 676693 346428
rect 676443 335340 676509 335341
rect 676443 335276 676444 335340
rect 676508 335276 676509 335340
rect 676443 335275 676509 335276
rect 676630 331261 676690 346427
rect 676627 331260 676693 331261
rect 676627 331196 676628 331260
rect 676692 331196 676693 331260
rect 676627 331195 676693 331196
rect 676075 326908 676141 326909
rect 676075 326844 676076 326908
rect 676140 326844 676141 326908
rect 676075 326843 676141 326844
rect 675523 308820 675589 308821
rect 675523 308756 675524 308820
rect 675588 308756 675589 308820
rect 675523 308755 675589 308756
rect 675526 302250 675586 308755
rect 675707 305964 675773 305965
rect 675707 305900 675708 305964
rect 675772 305900 675773 305964
rect 675707 305899 675773 305900
rect 675710 304330 675770 305899
rect 675710 304270 676506 304330
rect 676075 302972 676141 302973
rect 676075 302908 676076 302972
rect 676140 302970 676141 302972
rect 676140 302910 676322 302970
rect 676140 302908 676141 302910
rect 676075 302907 676141 302908
rect 675526 302190 676138 302250
rect 675891 299436 675957 299437
rect 675891 299372 675892 299436
rect 675956 299372 675957 299436
rect 675891 299371 675957 299372
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 675710 281621 675770 297331
rect 675894 282845 675954 299371
rect 676078 283661 676138 302190
rect 676262 291005 676322 302910
rect 676446 291549 676506 304270
rect 676627 301612 676693 301613
rect 676627 301548 676628 301612
rect 676692 301548 676693 301612
rect 676627 301547 676693 301548
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676259 291004 676325 291005
rect 676259 290940 676260 291004
rect 676324 290940 676325 291004
rect 676259 290939 676325 290940
rect 676630 287061 676690 301547
rect 676627 287060 676693 287061
rect 676627 286996 676628 287060
rect 676692 286996 676693 287060
rect 676627 286995 676693 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 282844 675957 282845
rect 675891 282780 675892 282844
rect 675956 282780 675957 282844
rect 675891 282779 675957 282780
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 673867 278628 673933 278629
rect 673867 278564 673868 278628
rect 673932 278564 673933 278628
rect 673867 278563 673933 278564
rect 673867 277676 673933 277677
rect 673867 277612 673868 277676
rect 673932 277612 673933 277676
rect 673867 277611 673933 277612
rect 665403 273732 665469 273733
rect 665403 273668 665404 273732
rect 665468 273668 665469 273732
rect 665403 273667 665469 273668
rect 665771 273732 665837 273733
rect 665771 273668 665772 273732
rect 665836 273668 665837 273732
rect 665771 273667 665837 273668
rect 41827 272372 41893 272373
rect 41827 272308 41828 272372
rect 41892 272308 41893 272372
rect 41827 272307 41893 272308
rect 489867 271692 489933 271693
rect 489867 271628 489868 271692
rect 489932 271690 489933 271692
rect 489932 271630 490114 271690
rect 489932 271628 489933 271630
rect 489867 271627 489933 271628
rect 490054 270605 490114 271630
rect 490051 270604 490117 270605
rect 490051 270540 490052 270604
rect 490116 270540 490117 270604
rect 490051 270539 490117 270540
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 40539 249796 40605 249797
rect 40539 249732 40540 249796
rect 40604 249732 40605 249796
rect 40539 249731 40605 249732
rect 40542 236605 40602 249731
rect 40723 246940 40789 246941
rect 40723 246876 40724 246940
rect 40788 246876 40789 246940
rect 40723 246875 40789 246876
rect 40726 238509 40786 246875
rect 40723 238508 40789 238509
rect 40723 238444 40724 238508
rect 40788 238444 40789 238508
rect 40723 238443 40789 238444
rect 42011 237692 42077 237693
rect 42011 237628 42012 237692
rect 42076 237628 42077 237692
rect 42011 237627 42077 237628
rect 40539 236604 40605 236605
rect 40539 236540 40540 236604
rect 40604 236540 40605 236604
rect 40539 236539 40605 236540
rect 42014 228989 42074 237627
rect 42379 237420 42445 237421
rect 42379 237356 42380 237420
rect 42444 237356 42445 237420
rect 42379 237355 42445 237356
rect 42011 228988 42077 228989
rect 42011 228924 42012 228988
rect 42076 228924 42077 228988
rect 42011 228923 42077 228924
rect 42382 227357 42442 237355
rect 42379 227356 42445 227357
rect 42379 227292 42380 227356
rect 42444 227292 42445 227356
rect 42379 227291 42445 227292
rect 559787 219196 559853 219197
rect 559787 219132 559788 219196
rect 559852 219132 559853 219196
rect 559787 219131 559853 219132
rect 571931 219196 571997 219197
rect 571931 219132 571932 219196
rect 571996 219132 571997 219196
rect 571931 219131 571997 219132
rect 542126 217910 542738 217970
rect 542126 217667 542186 217910
rect 542123 217666 542189 217667
rect 542123 217602 542124 217666
rect 542188 217602 542189 217666
rect 542123 217601 542189 217602
rect 542678 217565 542738 217910
rect 541203 217564 541269 217565
rect 541203 217500 541204 217564
rect 541268 217500 541269 217564
rect 541203 217499 541269 217500
rect 542491 217564 542557 217565
rect 542491 217500 542492 217564
rect 542556 217500 542557 217564
rect 542491 217499 542557 217500
rect 542675 217564 542741 217565
rect 542675 217500 542676 217564
rect 542740 217500 542741 217564
rect 542675 217499 542741 217500
rect 541206 215933 541266 217499
rect 542494 216205 542554 217499
rect 546723 216476 546789 216477
rect 546723 216412 546724 216476
rect 546788 216412 546789 216476
rect 546723 216411 546789 216412
rect 542491 216204 542557 216205
rect 542491 216140 542492 216204
rect 542556 216140 542557 216204
rect 542491 216139 542557 216140
rect 546726 215933 546786 216411
rect 559790 216205 559850 219131
rect 571934 218650 571994 219131
rect 571934 218590 572914 218650
rect 572854 217837 572914 218590
rect 560155 217836 560221 217837
rect 560155 217772 560156 217836
rect 560220 217772 560221 217836
rect 560155 217771 560221 217772
rect 563467 217836 563533 217837
rect 563467 217772 563468 217836
rect 563532 217772 563533 217836
rect 563467 217771 563533 217772
rect 572851 217836 572917 217837
rect 572851 217772 572852 217836
rect 572916 217772 572917 217836
rect 572851 217771 572917 217772
rect 560158 216205 560218 217771
rect 559787 216204 559853 216205
rect 559787 216140 559788 216204
rect 559852 216140 559853 216204
rect 559787 216139 559853 216140
rect 560155 216204 560221 216205
rect 560155 216140 560156 216204
rect 560220 216140 560221 216204
rect 560155 216139 560221 216140
rect 563470 215933 563530 217771
rect 541203 215932 541269 215933
rect 541203 215868 541204 215932
rect 541268 215868 541269 215932
rect 541203 215867 541269 215868
rect 546723 215932 546789 215933
rect 546723 215868 546724 215932
rect 546788 215868 546789 215932
rect 546723 215867 546789 215868
rect 563467 215932 563533 215933
rect 563467 215868 563468 215932
rect 563532 215868 563533 215932
rect 563467 215867 563533 215868
rect 41827 210084 41893 210085
rect 41827 210020 41828 210084
rect 41892 210020 41893 210084
rect 41827 210019 41893 210020
rect 41459 208996 41525 208997
rect 41459 208932 41460 208996
rect 41524 208932 41525 208996
rect 41459 208931 41525 208932
rect 40907 208180 40973 208181
rect 40907 208116 40908 208180
rect 40972 208116 40973 208180
rect 40907 208115 40973 208116
rect 40539 207772 40605 207773
rect 40539 207708 40540 207772
rect 40604 207708 40605 207772
rect 40539 207707 40605 207708
rect 40542 183429 40602 207707
rect 40723 206140 40789 206141
rect 40723 206076 40724 206140
rect 40788 206076 40789 206140
rect 40723 206075 40789 206076
rect 40726 191589 40786 206075
rect 40910 197165 40970 208115
rect 40907 197164 40973 197165
rect 40907 197100 40908 197164
rect 40972 197100 40973 197164
rect 40907 197099 40973 197100
rect 40723 191588 40789 191589
rect 40723 191524 40724 191588
rect 40788 191524 40789 191588
rect 40723 191523 40789 191524
rect 41462 184109 41522 208931
rect 41643 202196 41709 202197
rect 41643 202132 41644 202196
rect 41708 202132 41709 202196
rect 41643 202131 41709 202132
rect 41646 186330 41706 202131
rect 41830 195261 41890 210019
rect 665406 205650 665466 273667
rect 665587 273460 665653 273461
rect 665587 273396 665588 273460
rect 665652 273396 665653 273460
rect 665587 273395 665653 273396
rect 665590 208861 665650 273395
rect 665774 229110 665834 273667
rect 673870 249661 673930 277611
rect 676075 263668 676141 263669
rect 676075 263604 676076 263668
rect 676140 263604 676141 263668
rect 676075 263603 676141 263604
rect 674971 252652 675037 252653
rect 674971 252588 674972 252652
rect 675036 252588 675037 252652
rect 674971 252587 675037 252588
rect 674974 251190 675034 252587
rect 674790 251130 675034 251190
rect 674790 249661 674850 251130
rect 676078 249661 676138 263603
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 260812 676877 260813
rect 676811 260748 676812 260812
rect 676876 260748 676877 260812
rect 676811 260747 676877 260748
rect 673867 249660 673933 249661
rect 673867 249596 673868 249660
rect 673932 249596 673933 249660
rect 673867 249595 673933 249596
rect 674787 249660 674853 249661
rect 674787 249596 674788 249660
rect 674852 249596 674853 249660
rect 674787 249595 674853 249596
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 676814 246669 676874 260747
rect 676998 250205 677058 261563
rect 676995 250204 677061 250205
rect 676995 250140 676996 250204
rect 677060 250140 677061 250204
rect 676995 250139 677061 250140
rect 676811 246668 676877 246669
rect 676811 246604 676812 246668
rect 676876 246604 676877 246668
rect 676811 246603 676877 246604
rect 675523 245988 675589 245989
rect 675523 245924 675524 245988
rect 675588 245924 675589 245988
rect 675523 245923 675589 245924
rect 668163 245852 668229 245853
rect 668163 245788 668164 245852
rect 668228 245788 668229 245852
rect 668163 245787 668229 245788
rect 666691 245716 666757 245717
rect 666691 245652 666692 245716
rect 666756 245652 666757 245716
rect 666691 245651 666757 245652
rect 667979 245716 668045 245717
rect 667979 245652 667980 245716
rect 668044 245652 668045 245716
rect 667979 245651 668045 245652
rect 666507 245444 666573 245445
rect 666507 245380 666508 245444
rect 666572 245380 666573 245444
rect 666507 245379 666573 245380
rect 665774 229050 666202 229110
rect 665587 208860 665653 208861
rect 665587 208796 665588 208860
rect 665652 208796 665653 208860
rect 665587 208795 665653 208796
rect 665406 205590 666018 205650
rect 665958 202330 666018 205590
rect 666142 205050 666202 229050
rect 666510 205650 666570 245379
rect 666694 209790 666754 245651
rect 666694 209730 666938 209790
rect 666510 205590 666754 205650
rect 666142 204990 666570 205050
rect 666510 204237 666570 204990
rect 666507 204236 666573 204237
rect 666507 204172 666508 204236
rect 666572 204172 666573 204236
rect 666507 204171 666573 204172
rect 665958 202270 666570 202330
rect 666510 199341 666570 202270
rect 666507 199340 666573 199341
rect 666507 199276 666508 199340
rect 666572 199276 666573 199340
rect 666507 199275 666573 199276
rect 41827 195260 41893 195261
rect 41827 195196 41828 195260
rect 41892 195196 41893 195260
rect 41827 195195 41893 195196
rect 666694 189345 666754 205590
rect 666878 192609 666938 209730
rect 667982 194173 668042 245651
rect 668166 202333 668226 245787
rect 675526 241530 675586 245923
rect 675342 241470 675586 241530
rect 675342 238645 675402 241470
rect 675339 238644 675405 238645
rect 675339 238580 675340 238644
rect 675404 238580 675405 238644
rect 675339 238579 675405 238580
rect 675155 219060 675221 219061
rect 675155 218996 675156 219060
rect 675220 218996 675221 219060
rect 675155 218995 675221 218996
rect 673315 217428 673381 217429
rect 673315 217364 673316 217428
rect 673380 217364 673381 217428
rect 673315 217363 673381 217364
rect 673131 214572 673197 214573
rect 673131 214570 673132 214572
rect 672950 214510 673132 214570
rect 670739 212668 670805 212669
rect 670739 212604 670740 212668
rect 670804 212604 670805 212668
rect 670739 212603 670805 212604
rect 669819 209676 669885 209677
rect 669819 209612 669820 209676
rect 669884 209612 669885 209676
rect 669819 209611 669885 209612
rect 669635 208316 669701 208317
rect 669635 208252 669636 208316
rect 669700 208252 669701 208316
rect 669635 208251 669701 208252
rect 669638 206410 669698 208251
rect 669270 206350 669698 206410
rect 669270 205461 669330 206350
rect 669822 205730 669882 209611
rect 669454 205670 669882 205730
rect 669267 205460 669333 205461
rect 669267 205396 669268 205460
rect 669332 205396 669333 205460
rect 669267 205395 669333 205396
rect 668163 202332 668229 202333
rect 668163 202268 668164 202332
rect 668228 202268 668229 202332
rect 668163 202267 668229 202268
rect 669267 196212 669333 196213
rect 669267 196148 669268 196212
rect 669332 196148 669333 196212
rect 669267 196147 669333 196148
rect 669270 195941 669330 196147
rect 669267 195940 669333 195941
rect 669267 195876 669268 195940
rect 669332 195876 669333 195940
rect 669267 195875 669333 195876
rect 667979 194172 668045 194173
rect 667979 194108 667980 194172
rect 668044 194108 668045 194172
rect 667979 194107 668045 194108
rect 666875 192608 666941 192609
rect 666875 192544 666876 192608
rect 666940 192544 666941 192608
rect 666875 192543 666941 192544
rect 666691 189344 666757 189345
rect 666691 189280 666692 189344
rect 666756 189280 666757 189344
rect 666691 189279 666757 189280
rect 669267 186420 669333 186421
rect 669267 186356 669268 186420
rect 669332 186356 669333 186420
rect 669267 186355 669333 186356
rect 41646 186270 41890 186330
rect 41830 185877 41890 186270
rect 41827 185876 41893 185877
rect 41827 185812 41828 185876
rect 41892 185812 41893 185876
rect 41827 185811 41893 185812
rect 41459 184108 41525 184109
rect 41459 184044 41460 184108
rect 41524 184044 41525 184108
rect 41459 184043 41525 184044
rect 40539 183428 40605 183429
rect 40539 183364 40540 183428
rect 40604 183364 40605 183428
rect 40539 183363 40605 183364
rect 669270 176670 669330 186355
rect 669454 179485 669514 205670
rect 669635 205460 669701 205461
rect 669635 205396 669636 205460
rect 669700 205396 669701 205460
rect 669635 205395 669701 205396
rect 669638 196213 669698 205395
rect 669635 196212 669701 196213
rect 669635 196148 669636 196212
rect 669700 196148 669701 196212
rect 669635 196147 669701 196148
rect 669635 195940 669701 195941
rect 669635 195876 669636 195940
rect 669700 195876 669701 195940
rect 669635 195875 669701 195876
rect 669638 186421 669698 195875
rect 669635 186420 669701 186421
rect 669635 186356 669636 186420
rect 669700 186356 669701 186420
rect 669635 186355 669701 186356
rect 669451 179484 669517 179485
rect 669451 179420 669452 179484
rect 669516 179420 669517 179484
rect 669451 179419 669517 179420
rect 669270 176610 669514 176670
rect 669454 174589 669514 176610
rect 669451 174588 669517 174589
rect 669451 174524 669452 174588
rect 669516 174524 669517 174588
rect 669451 174523 669517 174524
rect 670742 164797 670802 212603
rect 670923 210492 670989 210493
rect 670923 210428 670924 210492
rect 670988 210428 670989 210492
rect 670923 210427 670989 210428
rect 670926 168061 670986 210427
rect 672950 183565 673010 214510
rect 673131 214508 673132 214510
rect 673196 214508 673197 214572
rect 673131 214507 673197 214508
rect 673318 212550 673378 217363
rect 673499 215660 673565 215661
rect 673499 215596 673500 215660
rect 673564 215596 673565 215660
rect 673499 215595 673565 215596
rect 673134 212490 673378 212550
rect 672947 183564 673013 183565
rect 672947 183500 672948 183564
rect 673012 183500 673013 183564
rect 672947 183499 673013 183500
rect 673134 172957 673194 212490
rect 673131 172956 673197 172957
rect 673131 172892 673132 172956
rect 673196 172892 673197 172956
rect 673131 172891 673197 172892
rect 672027 168332 672093 168333
rect 672027 168268 672028 168332
rect 672092 168268 672093 168332
rect 672027 168267 672093 168268
rect 670923 168060 670989 168061
rect 670923 167996 670924 168060
rect 670988 167996 670989 168060
rect 670923 167995 670989 167996
rect 670739 164796 670805 164797
rect 670739 164732 670740 164796
rect 670804 164732 670805 164796
rect 670739 164731 670805 164732
rect 672030 159901 672090 168267
rect 672027 159900 672093 159901
rect 672027 159836 672028 159900
rect 672092 159836 672093 159900
rect 672027 159835 672093 159836
rect 673502 149701 673562 215595
rect 673683 215388 673749 215389
rect 673683 215324 673684 215388
rect 673748 215324 673749 215388
rect 673683 215323 673749 215324
rect 673686 153237 673746 215323
rect 675158 210221 675218 218995
rect 675523 218652 675589 218653
rect 675523 218588 675524 218652
rect 675588 218588 675589 218652
rect 675523 218587 675589 218588
rect 675339 217836 675405 217837
rect 675339 217772 675340 217836
rect 675404 217772 675405 217836
rect 675339 217771 675405 217772
rect 675155 210220 675221 210221
rect 675155 210156 675156 210220
rect 675220 210156 675221 210220
rect 675155 210155 675221 210156
rect 675342 202741 675402 217771
rect 675526 210490 675586 218587
rect 675707 216612 675773 216613
rect 675707 216548 675708 216612
rect 675772 216548 675773 216612
rect 675707 216547 675773 216548
rect 675710 213890 675770 216547
rect 675894 215190 676690 215250
rect 675894 214981 675954 215190
rect 675891 214980 675957 214981
rect 675891 214916 675892 214980
rect 675956 214916 675957 214980
rect 675891 214915 675957 214916
rect 675891 214572 675957 214573
rect 675891 214508 675892 214572
rect 675956 214570 675957 214572
rect 675956 214510 676506 214570
rect 675956 214508 675957 214510
rect 675891 214507 675957 214508
rect 675710 213830 676322 213890
rect 675526 210430 676138 210490
rect 675891 210220 675957 210221
rect 675891 210156 675892 210220
rect 675956 210156 675957 210220
rect 675891 210155 675957 210156
rect 675894 204237 675954 210155
rect 675891 204236 675957 204237
rect 675891 204172 675892 204236
rect 675956 204172 675957 204236
rect 675891 204171 675957 204172
rect 675339 202740 675405 202741
rect 675339 202676 675340 202740
rect 675404 202676 675405 202740
rect 675339 202675 675405 202676
rect 674787 200836 674853 200837
rect 674787 200772 674788 200836
rect 674852 200772 674853 200836
rect 674787 200771 674853 200772
rect 674790 185877 674850 200771
rect 675523 193628 675589 193629
rect 675523 193564 675524 193628
rect 675588 193564 675589 193628
rect 675523 193563 675589 193564
rect 675526 191589 675586 193563
rect 676078 193221 676138 210430
rect 676262 205053 676322 213830
rect 676259 205052 676325 205053
rect 676259 204988 676260 205052
rect 676324 204988 676325 205052
rect 676259 204987 676325 204988
rect 676446 200021 676506 214510
rect 676443 200020 676509 200021
rect 676443 199956 676444 200020
rect 676508 199956 676509 200020
rect 676443 199955 676509 199956
rect 676630 197165 676690 215190
rect 676811 198660 676877 198661
rect 676811 198596 676812 198660
rect 676876 198596 676877 198660
rect 676811 198595 676877 198596
rect 676627 197164 676693 197165
rect 676627 197100 676628 197164
rect 676692 197100 676693 197164
rect 676627 197099 676693 197100
rect 676075 193220 676141 193221
rect 676075 193156 676076 193220
rect 676140 193156 676141 193220
rect 676075 193155 676141 193156
rect 675523 191588 675589 191589
rect 675523 191524 675524 191588
rect 675588 191524 675589 191588
rect 675523 191523 675589 191524
rect 674787 185876 674853 185877
rect 674787 185812 674788 185876
rect 674852 185812 674853 185876
rect 674787 185811 674853 185812
rect 676814 183570 676874 198595
rect 676262 183510 676874 183570
rect 675891 174724 675957 174725
rect 675891 174660 675892 174724
rect 675956 174660 675957 174724
rect 675891 174659 675957 174660
rect 675894 174450 675954 174659
rect 676262 174450 676322 183510
rect 675894 174390 676322 174450
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675710 169690 675770 173571
rect 675891 170372 675957 170373
rect 675891 170308 675892 170372
rect 675956 170370 675957 170372
rect 675956 170310 676322 170370
rect 675956 170308 675957 170310
rect 675891 170307 675957 170308
rect 675710 169630 676138 169690
rect 675891 167516 675957 167517
rect 675891 167452 675892 167516
rect 675956 167452 675957 167516
rect 675891 167451 675957 167452
rect 675707 161940 675773 161941
rect 675707 161876 675708 161940
rect 675772 161876 675773 161940
rect 675707 161875 675773 161876
rect 673683 153236 673749 153237
rect 673683 153172 673684 153236
rect 673748 153172 673749 153236
rect 673683 153171 673749 153172
rect 675710 153101 675770 161875
rect 675707 153100 675773 153101
rect 675707 153036 675708 153100
rect 675772 153036 675773 153100
rect 675707 153035 675773 153036
rect 673499 149700 673565 149701
rect 673499 149636 673500 149700
rect 673564 149636 673565 149700
rect 673499 149635 673565 149636
rect 675894 147661 675954 167451
rect 676078 148477 676138 169630
rect 676262 150381 676322 170310
rect 676443 166428 676509 166429
rect 676443 166364 676444 166428
rect 676508 166364 676509 166428
rect 676443 166363 676509 166364
rect 676446 151469 676506 166363
rect 676627 166292 676693 166293
rect 676627 166228 676628 166292
rect 676692 166228 676693 166292
rect 676627 166227 676693 166228
rect 676630 156365 676690 166227
rect 676627 156364 676693 156365
rect 676627 156300 676628 156364
rect 676692 156300 676693 156364
rect 676627 156299 676693 156300
rect 676443 151468 676509 151469
rect 676443 151404 676444 151468
rect 676508 151404 676509 151468
rect 676443 151403 676509 151404
rect 676259 150380 676325 150381
rect 676259 150316 676260 150380
rect 676324 150316 676325 150380
rect 676259 150315 676325 150316
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675891 147660 675957 147661
rect 675891 147596 675892 147660
rect 675956 147596 675957 147660
rect 675891 147595 675957 147596
rect 676259 128620 676325 128621
rect 676259 128556 676260 128620
rect 676324 128556 676325 128620
rect 676259 128555 676325 128556
rect 675891 127260 675957 127261
rect 675891 127196 675892 127260
rect 675956 127196 675957 127260
rect 675891 127195 675957 127196
rect 675707 122908 675773 122909
rect 675707 122844 675708 122908
rect 675772 122844 675773 122908
rect 675707 122843 675773 122844
rect 675710 120325 675770 122843
rect 675707 120324 675773 120325
rect 675707 120260 675708 120324
rect 675772 120260 675773 120324
rect 675707 120259 675773 120260
rect 675707 116108 675773 116109
rect 675707 116044 675708 116108
rect 675772 116044 675773 116108
rect 675707 116043 675773 116044
rect 675710 102645 675770 116043
rect 675894 108085 675954 127195
rect 676075 120324 676141 120325
rect 676075 120260 676076 120324
rect 676140 120260 676141 120324
rect 676075 120259 676141 120260
rect 675891 108084 675957 108085
rect 675891 108020 675892 108084
rect 675956 108020 675957 108084
rect 675891 108019 675957 108020
rect 676078 103189 676138 120259
rect 676262 114205 676322 128555
rect 676811 124540 676877 124541
rect 676811 124476 676812 124540
rect 676876 124476 676877 124540
rect 676811 124475 676877 124476
rect 676259 114204 676325 114205
rect 676259 114140 676260 114204
rect 676324 114140 676325 114204
rect 676259 114139 676325 114140
rect 676075 103188 676141 103189
rect 676075 103124 676076 103188
rect 676140 103124 676141 103188
rect 676075 103123 676141 103124
rect 675707 102644 675773 102645
rect 675707 102580 675708 102644
rect 675772 102580 675773 102644
rect 675707 102579 675773 102580
rect 676814 101421 676874 124475
rect 676995 124132 677061 124133
rect 676995 124068 676996 124132
rect 677060 124068 677061 124132
rect 676995 124067 677061 124068
rect 676998 110397 677058 124067
rect 676995 110396 677061 110397
rect 676995 110332 676996 110396
rect 677060 110332 677061 110396
rect 676995 110331 677061 110332
rect 676811 101420 676877 101421
rect 676811 101356 676812 101420
rect 676876 101356 676877 101420
rect 676811 101355 676877 101356
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 634675 95708 634741 95709
rect 634675 95644 634676 95708
rect 634740 95644 634741 95708
rect 634675 95643 634741 95644
rect 634678 77757 634738 95643
rect 637254 84210 637314 96867
rect 637070 84150 637314 84210
rect 637070 78573 637130 84150
rect 637067 78572 637133 78573
rect 637067 78508 637068 78572
rect 637132 78508 637133 78572
rect 637067 78507 637133 78508
rect 634675 77756 634741 77757
rect 634675 77692 634676 77756
rect 634740 77692 634741 77756
rect 634675 77691 634741 77692
rect 464843 51780 464909 51781
rect 464843 51716 464844 51780
rect 464908 51716 464909 51780
rect 464843 51715 464909 51716
rect 150387 50284 150453 50285
rect 150387 50220 150388 50284
rect 150452 50220 150453 50284
rect 150387 50219 150453 50220
rect 78627 49740 78693 49741
rect 78627 49676 78628 49740
rect 78692 49676 78693 49740
rect 78627 49675 78693 49676
rect 78630 47293 78690 49675
rect 150390 47565 150450 50219
rect 411115 49196 411181 49197
rect 411115 49132 411116 49196
rect 411180 49132 411181 49196
rect 411115 49131 411181 49132
rect 365483 48924 365549 48925
rect 365483 48860 365484 48924
rect 365548 48860 365549 48924
rect 365483 48859 365549 48860
rect 310467 47836 310533 47837
rect 310467 47772 310468 47836
rect 310532 47772 310533 47836
rect 310467 47771 310533 47772
rect 150387 47564 150453 47565
rect 150387 47500 150388 47564
rect 150452 47500 150453 47564
rect 150387 47499 150453 47500
rect 187555 47564 187621 47565
rect 187555 47500 187556 47564
rect 187620 47500 187621 47564
rect 187555 47499 187621 47500
rect 78627 47292 78693 47293
rect 78627 47228 78628 47292
rect 78692 47228 78693 47292
rect 78627 47227 78693 47228
rect 187558 42125 187618 47499
rect 306971 46204 307037 46205
rect 306971 46140 306972 46204
rect 307036 46140 307037 46204
rect 306971 46139 307037 46140
rect 306974 42397 307034 46139
rect 306971 42396 307037 42397
rect 306971 42332 306972 42396
rect 307036 42332 307037 42396
rect 306971 42331 307037 42332
rect 310470 42125 310530 47771
rect 361987 46476 362053 46477
rect 361987 46412 361988 46476
rect 362052 46412 362053 46476
rect 361987 46411 362053 46412
rect 361990 42125 362050 46411
rect 365486 42125 365546 48859
rect 411118 42805 411178 49131
rect 416635 47020 416701 47021
rect 416635 46956 416636 47020
rect 416700 46956 416701 47020
rect 416635 46955 416701 46956
rect 416638 42805 416698 46955
rect 460611 45796 460677 45797
rect 460611 45732 460612 45796
rect 460676 45732 460677 45796
rect 460611 45731 460677 45732
rect 411115 42804 411181 42805
rect 411115 42740 411116 42804
rect 411180 42740 411181 42804
rect 411115 42739 411181 42740
rect 416635 42804 416701 42805
rect 416635 42740 416636 42804
rect 416700 42740 416701 42804
rect 416635 42739 416701 42740
rect 460614 42125 460674 45731
rect 464846 42805 464906 51715
rect 525747 50556 525813 50557
rect 525747 50492 525748 50556
rect 525812 50492 525813 50556
rect 525747 50491 525813 50492
rect 517467 50284 517533 50285
rect 517467 50220 517468 50284
rect 517532 50220 517533 50284
rect 517467 50219 517533 50220
rect 514707 45932 514773 45933
rect 514707 45868 514708 45932
rect 514772 45868 514773 45932
rect 514707 45867 514773 45868
rect 471651 44844 471717 44845
rect 471651 44780 471652 44844
rect 471716 44780 471717 44844
rect 471651 44779 471717 44780
rect 464843 42804 464909 42805
rect 464843 42740 464844 42804
rect 464908 42740 464909 42804
rect 464843 42739 464909 42740
rect 471654 42125 471714 44779
rect 514710 42125 514770 45867
rect 517470 42397 517530 50219
rect 521699 47020 521765 47021
rect 521699 46956 521700 47020
rect 521764 46956 521765 47020
rect 521699 46955 521765 46956
rect 520411 45116 520477 45117
rect 520411 45052 520412 45116
rect 520476 45052 520477 45116
rect 520411 45051 520477 45052
rect 517467 42396 517533 42397
rect 517467 42332 517468 42396
rect 517532 42332 517533 42396
rect 517467 42331 517533 42332
rect 520414 42125 520474 45051
rect 187555 42124 187621 42125
rect 187555 42060 187556 42124
rect 187620 42060 187621 42124
rect 187555 42059 187621 42060
rect 310467 42124 310533 42125
rect 310467 42060 310468 42124
rect 310532 42060 310533 42124
rect 310467 42059 310533 42060
rect 361987 42124 362053 42125
rect 361987 42060 361988 42124
rect 362052 42060 362053 42124
rect 361987 42059 362053 42060
rect 365483 42124 365549 42125
rect 365483 42060 365484 42124
rect 365548 42060 365549 42124
rect 365483 42059 365549 42060
rect 460611 42124 460677 42125
rect 460611 42060 460612 42124
rect 460676 42060 460677 42124
rect 460611 42059 460677 42060
rect 471651 42124 471717 42125
rect 471651 42060 471652 42124
rect 471716 42060 471717 42124
rect 471651 42059 471717 42060
rect 514707 42124 514773 42125
rect 514707 42060 514708 42124
rect 514772 42060 514773 42124
rect 514707 42059 514773 42060
rect 520411 42124 520477 42125
rect 520411 42060 520412 42124
rect 520476 42060 520477 42124
rect 520411 42059 520477 42060
rect 521702 41989 521762 46955
rect 525750 42125 525810 50491
rect 529795 50284 529861 50285
rect 529795 50220 529796 50284
rect 529860 50220 529861 50284
rect 529795 50219 529861 50220
rect 529798 42125 529858 50219
rect 525747 42124 525813 42125
rect 525747 42060 525748 42124
rect 525812 42060 525813 42124
rect 525747 42059 525813 42060
rect 529795 42124 529861 42125
rect 529795 42060 529796 42124
rect 529860 42060 529861 42124
rect 529795 42059 529861 42060
rect 521699 41988 521765 41989
rect 521699 41924 521700 41988
rect 521764 41924 521765 41988
rect 521699 41923 521765 41924
<< via4 >>
rect 189310 997102 189546 997338
rect 194278 997252 194514 997338
rect 194278 997188 194364 997252
rect 194364 997188 194428 997252
rect 194428 997188 194514 997252
rect 194278 997102 194514 997188
rect 239542 997102 239778 997338
rect 242486 997102 242722 997338
rect 243222 997102 243458 997338
rect 274502 997102 274738 997338
rect 383246 997102 383482 997338
rect 388030 997102 388266 997338
rect 536518 997102 536754 997338
rect 573134 997102 573370 997338
rect 503398 220012 503634 220098
rect 503398 219948 503484 220012
rect 503484 219948 503548 220012
rect 503548 219948 503634 220012
rect 503398 219862 503634 219948
rect 574054 220012 574290 220098
rect 574054 219948 574140 220012
rect 574140 219948 574204 220012
rect 574204 219948 574290 220012
rect 574054 219862 574290 219948
<< metal5 >>
rect 189268 997338 194556 997380
rect 189268 997102 189310 997338
rect 189546 997102 194278 997338
rect 194514 997102 194556 997338
rect 189268 997060 194556 997102
rect 239500 997338 242764 997380
rect 239500 997102 239542 997338
rect 239778 997102 242486 997338
rect 242722 997102 242764 997338
rect 239500 997060 242764 997102
rect 243180 997338 274780 997380
rect 243180 997102 243222 997338
rect 243458 997102 274502 997338
rect 274738 997102 274780 997338
rect 243180 997060 274780 997102
rect 383204 997338 388308 997380
rect 383204 997102 383246 997338
rect 383482 997102 388030 997338
rect 388266 997102 388308 997338
rect 383204 997060 388308 997102
rect 536476 997338 573412 997380
rect 536476 997102 536518 997338
rect 536754 997102 573134 997338
rect 573370 997102 573412 997338
rect 536476 997060 573412 997102
rect 503356 220098 574332 220140
rect 503356 219862 503398 220098
rect 503634 219862 574054 220098
rect 574290 219862 574332 220098
rect 503356 219820 574332 219862
use user_id_programming  user_id_value
timestamp 1665401783
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1665401783
transform 1 0 52034 0 1 53002
box 844 -400 524400 164400
use xres_buf  rstb_level
timestamp 1665401783
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use simple_por  por
timestamp 1665401783
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use digital_pll  pll
timestamp 1665401783
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use housekeeping  housekeeping
timestamp 1665401783
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1665401783
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1665401783
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use caravel_clocking  clock_ctrl
timestamp 1665401783
transform 1 0 626764 0 1 63284
box -38 -48 20000 12000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1665401783
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1665401783
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1665401783
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1665401783
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1665401783
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1665401783
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1665401783
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1665401783
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1665401783
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use mgmt_protect  mgmt_buffers
timestamp 1665401783
transform 1 0 128180 0 1 232036
box 1066 -400 380400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1665401783
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1665401783
transform 1 0 89351 0 1 248673
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1665401783
transform 1 0 575145 0 1 246987
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1665401783
transform 1 0 613558 0 1 245856
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1665401783
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1665401783
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1665401783
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1665401783
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1665401783
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1665401783
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1665401783
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1665401783
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1665401783
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1665401783
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1665401783
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1665401783
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1665401783
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1665401783
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1665401783
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1665401783
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1665401783
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1665401783
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1665401783
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1665401783
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1665401783
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1665401783
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1665401783
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1665401783
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1665401783
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1665401783
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1665401783
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1665401783
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1665401783
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1665401783
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1665401783
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1665401783
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1665401783
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1665401783
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1665401783
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1665401783
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1665401783
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1665401783
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1665401783
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1665401783
transform -1 0 710203 0 1 749200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1665401783
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1665401783
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1665401783
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1665401783
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1665401783
transform 1 0 7631 0 1 931200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1665401783
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1665401783
transform -1 0 710203 0 1 927600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1665401783
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1665401783
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1665401783
transform 0 1 97200 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1665401783
transform 0 1 148600 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1665401783
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1665401783
transform 0 1 200000 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1665401783
transform 0 1 251400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1665401783
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1665401783
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1665401783
transform 0 1 303000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1665401783
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1665401783
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1665401783
transform 0 1 420800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1665401783
transform 0 1 353400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1665401783
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1665401783
transform 0 1 497800 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1665401783
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1665401783
transform 0 1 549200 -1 0 1030077
box 872 416 34000 13000
use caravel_power_routing  caravel_power_routing
timestamp 1665401783
transform 1 0 6022 0 1 33900
box 0 0 705792 997796
use user_project_wrapper  mprj
timestamp 1665401783
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1665401783
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
