VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_motto
  CLASS BLOCK ;
  FOREIGN caravel_motto ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 25.000 ;
END caravel_motto
END LIBRARY

