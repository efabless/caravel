magic
tech sky130A
magscale 1 2
timestamp 1636108275
<< nwell >>
rect -38 1893 5006 2214
rect -38 805 5006 1371
<< obsli1 >>
rect 0 527 4968 2193
<< obsm1 >>
rect 0 496 4968 2224
<< metal2 >>
rect 202 0 258 400
rect 570 0 626 400
rect 938 0 994 400
rect 1306 0 1362 400
rect 1674 0 1730 400
rect 2042 0 2098 400
rect 2410 0 2466 400
rect 2870 0 2926 400
rect 3238 0 3294 400
rect 3606 0 3662 400
rect 3974 0 4030 400
rect 4342 0 4398 400
rect 4710 0 4766 400
<< obsm2 >>
rect 78 2200 322 2224
rect 1478 2200 1722 2224
rect 2878 2200 3122 2224
rect 4278 2200 4522 2224
rect 78 456 4764 2200
rect 78 326 146 456
rect 314 326 514 456
rect 682 326 882 456
rect 1050 326 1250 456
rect 1418 326 1618 456
rect 1786 326 1986 456
rect 2154 326 2354 456
rect 2522 326 2814 456
rect 2982 326 3182 456
rect 3350 326 3550 456
rect 3718 326 3918 456
rect 4086 326 4286 456
rect 4454 326 4654 456
<< obsm3 >>
rect 60 2200 340 2209
rect 1460 2200 1740 2209
rect 2860 2200 3140 2209
rect 4260 2200 4540 2209
rect 60 511 4540 2200
<< metal4 >>
rect 60 496 340 2224
rect 760 496 1040 2224
rect 1460 496 1740 2224
rect 2160 496 2440 2224
rect 2860 496 3140 2224
rect 3560 496 3840 2224
rect 4260 496 4540 2224
<< metal5 >>
rect 0 1436 4968 1756
rect 0 736 4968 1056
<< labels >>
rlabel metal5 s 0 1436 4968 1756 6 VGND
port 1 nsew ground input
rlabel metal4 s 760 496 1040 2224 6 VGND
port 1 nsew ground input
rlabel metal4 s 2160 496 2440 2224 6 VGND
port 1 nsew ground input
rlabel metal4 s 3560 496 3840 2224 6 VGND
port 1 nsew ground input
rlabel metal5 s 0 736 4968 1056 6 VPWR
port 2 nsew power input
rlabel metal4 s 60 496 340 2224 6 VPWR
port 2 nsew power input
rlabel metal4 s 1460 496 1740 2224 6 VPWR
port 2 nsew power input
rlabel metal4 s 2860 496 3140 2224 6 VPWR
port 2 nsew power input
rlabel metal4 s 4260 496 4540 2224 6 VPWR
port 2 nsew power input
rlabel metal2 s 202 0 258 400 6 gpio_defaults[0]
port 3 nsew signal output
rlabel metal2 s 3974 0 4030 400 6 gpio_defaults[10]
port 4 nsew signal output
rlabel metal2 s 4342 0 4398 400 6 gpio_defaults[11]
port 5 nsew signal output
rlabel metal2 s 4710 0 4766 400 6 gpio_defaults[12]
port 6 nsew signal output
rlabel metal2 s 570 0 626 400 6 gpio_defaults[1]
port 7 nsew signal output
rlabel metal2 s 938 0 994 400 6 gpio_defaults[2]
port 8 nsew signal output
rlabel metal2 s 1306 0 1362 400 6 gpio_defaults[3]
port 9 nsew signal output
rlabel metal2 s 1674 0 1730 400 6 gpio_defaults[4]
port 10 nsew signal output
rlabel metal2 s 2042 0 2098 400 6 gpio_defaults[5]
port 11 nsew signal output
rlabel metal2 s 2410 0 2466 400 6 gpio_defaults[6]
port 12 nsew signal output
rlabel metal2 s 2870 0 2926 400 6 gpio_defaults[7]
port 13 nsew signal output
rlabel metal2 s 3238 0 3294 400 6 gpio_defaults[8]
port 14 nsew signal output
rlabel metal2 s 3606 0 3662 400 6 gpio_defaults[9]
port 15 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 5000 2200
string LEFview TRUE
string GDS_FILE ../gds/gpio_defaults_block.gds
string GDS_END 47838
string GDS_START 20982
<< end >>

