VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan_power_routing
  CLASS BLOCK ;
  FOREIGN caravan_power_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  OBS
      LAYER met1 ;
        RECT 3240.520 233.690 3248.350 235.940 ;
        RECT 3240.520 232.990 3250.800 233.690 ;
        RECT 3240.520 232.950 3248.350 232.990 ;
      LAYER via ;
        RECT 3240.830 233.300 3248.040 235.620 ;
      LAYER met2 ;
        RECT 3240.520 232.950 3248.350 235.940 ;
      LAYER via2 ;
        RECT 3240.830 233.300 3248.040 235.620 ;
      LAYER met3 ;
        RECT 2878.500 4975.160 2902.395 4988.390 ;
        RECT 2928.390 4975.160 2952.290 4988.390 ;
        RECT 2878.810 4974.420 2901.920 4975.160 ;
        RECT 2928.790 4974.490 2951.900 4975.160 ;
        RECT 3376.330 4511.910 3559.020 4517.910 ;
        RECT 3358.050 4503.910 3552.950 4509.910 ;
        RECT 3429.570 4495.500 3499.990 4501.500 ;
        RECT 3396.620 4487.500 3494.020 4493.500 ;
        RECT 199.260 4188.390 250.010 4212.290 ;
        RECT 199.260 4138.495 250.010 4162.395 ;
        RECT 3335.860 4142.605 3389.090 4166.505 ;
        RECT 30.110 4114.910 277.300 4120.910 ;
        RECT 36.180 4106.910 269.080 4112.910 ;
        RECT 89.140 4098.500 158.310 4104.500 ;
        RECT 95.110 4090.500 191.260 4096.500 ;
        RECT 3335.860 4092.710 3389.090 4116.610 ;
        RECT 30.110 3898.910 277.300 3904.910 ;
        RECT 36.180 3890.910 269.080 3896.910 ;
        RECT 89.140 3882.500 158.310 3888.500 ;
        RECT 95.110 3874.500 191.260 3880.500 ;
        RECT 30.110 3682.910 277.300 3688.910 ;
        RECT 36.180 3674.910 269.080 3680.910 ;
        RECT 89.140 3666.500 158.310 3672.500 ;
        RECT 95.110 3658.500 191.260 3664.500 ;
        RECT 3376.380 3608.910 3559.070 3614.910 ;
        RECT 3358.100 3600.910 3553.000 3606.910 ;
        RECT 3429.620 3592.500 3500.040 3598.500 ;
        RECT 3396.670 3584.500 3494.070 3590.500 ;
        RECT 30.110 3466.910 277.300 3472.910 ;
        RECT 36.180 3458.910 269.080 3464.910 ;
        RECT 89.140 3450.500 158.310 3456.500 ;
        RECT 95.110 3442.500 191.260 3448.500 ;
        RECT 3376.380 3382.910 3559.070 3388.910 ;
        RECT 3358.100 3374.910 3553.000 3380.910 ;
        RECT 3429.620 3366.500 3500.040 3372.500 ;
        RECT 3396.670 3358.500 3494.070 3364.500 ;
        RECT 30.110 3250.910 277.300 3256.910 ;
        RECT 36.180 3242.910 269.080 3248.910 ;
        RECT 89.140 3234.500 158.310 3240.500 ;
        RECT 95.110 3226.500 191.260 3232.500 ;
        RECT 3376.380 3157.910 3559.070 3163.910 ;
        RECT 3358.100 3149.910 3553.000 3155.910 ;
        RECT 3429.620 3141.500 3500.040 3147.500 ;
        RECT 3396.670 3133.500 3494.070 3139.500 ;
        RECT 30.110 3034.910 277.300 3040.910 ;
        RECT 36.180 3026.910 269.080 3032.910 ;
        RECT 89.140 3018.500 158.310 3024.500 ;
        RECT 95.110 3010.500 191.260 3016.500 ;
        RECT 3376.380 2931.910 3559.070 2937.910 ;
        RECT 3358.100 2923.910 3553.000 2929.910 ;
        RECT 3429.620 2915.500 3500.040 2921.500 ;
        RECT 3396.670 2907.500 3494.070 2913.500 ;
        RECT 30.110 2818.910 277.300 2824.910 ;
        RECT 36.180 2810.910 269.080 2816.910 ;
        RECT 89.140 2802.500 158.310 2808.500 ;
        RECT 95.110 2794.500 191.260 2800.500 ;
        RECT 3376.380 2706.910 3559.070 2712.910 ;
        RECT 3358.100 2698.910 3553.000 2704.910 ;
        RECT 3429.620 2690.500 3500.040 2696.500 ;
        RECT 3396.670 2682.500 3494.070 2688.500 ;
        RECT 3335.310 2569.605 3388.500 2593.505 ;
        RECT 3335.310 2519.710 3388.500 2543.610 ;
        RECT 199.620 2465.390 261.460 2489.290 ;
        RECT 3376.380 2486.910 3559.070 2492.910 ;
        RECT 3358.100 2478.910 3553.000 2484.910 ;
        RECT 3429.620 2470.500 3500.040 2476.500 ;
        RECT 3396.670 2462.500 3494.070 2468.500 ;
        RECT 199.620 2415.495 261.460 2439.395 ;
        RECT 30.110 2180.910 277.300 2186.910 ;
        RECT 36.180 2172.910 269.080 2178.910 ;
        RECT 89.140 2164.500 158.310 2170.500 ;
        RECT 95.110 2156.500 191.260 2162.500 ;
        RECT 3319.570 2128.740 3388.560 2152.505 ;
        RECT 3319.570 2127.810 3335.550 2128.740 ;
        RECT 3319.570 2078.710 3388.560 2102.610 ;
        RECT 3376.380 2045.910 3559.070 2051.910 ;
        RECT 3358.100 2037.910 3553.000 2043.910 ;
        RECT 3429.620 2029.500 3500.040 2035.500 ;
        RECT 3396.670 2021.500 3494.070 2027.500 ;
        RECT 30.110 1964.910 277.300 1970.910 ;
        RECT 36.180 1956.910 269.080 1962.910 ;
        RECT 89.140 1948.500 158.310 1954.500 ;
        RECT 95.110 1940.500 191.260 1946.500 ;
        RECT 3376.380 1819.910 3559.070 1825.910 ;
        RECT 3358.100 1811.910 3553.000 1817.910 ;
        RECT 3429.620 1803.500 3500.040 1809.500 ;
        RECT 3396.670 1795.500 3494.070 1801.500 ;
        RECT 30.110 1748.910 277.300 1754.910 ;
        RECT 36.180 1740.910 269.080 1746.910 ;
        RECT 89.140 1732.500 158.310 1738.500 ;
        RECT 95.110 1724.500 191.260 1730.500 ;
        RECT 3376.380 1594.910 3559.070 1600.910 ;
        RECT 3358.100 1586.910 3553.000 1592.910 ;
        RECT 3429.620 1578.500 3500.040 1584.500 ;
        RECT 3396.670 1570.500 3494.070 1576.500 ;
        RECT 30.110 1532.910 277.300 1538.910 ;
        RECT 36.180 1524.910 269.080 1530.910 ;
        RECT 89.140 1516.500 158.310 1522.500 ;
        RECT 95.110 1508.500 191.260 1514.500 ;
        RECT 3376.380 1369.910 3559.070 1375.910 ;
        RECT 3358.100 1361.910 3553.000 1367.910 ;
        RECT 3429.620 1353.500 3500.040 1359.500 ;
        RECT 3396.670 1345.500 3494.070 1351.500 ;
        RECT 30.110 1316.910 277.300 1322.910 ;
        RECT 36.180 1308.910 269.080 1314.910 ;
        RECT 89.140 1300.500 158.310 1306.500 ;
        RECT 95.110 1292.500 191.260 1298.500 ;
        RECT 3376.380 1143.910 3559.070 1149.910 ;
        RECT 3358.100 1135.910 3553.000 1141.910 ;
        RECT 3429.620 1127.500 3500.040 1133.500 ;
        RECT 3396.670 1119.500 3494.070 1125.500 ;
        RECT 30.110 1100.910 277.300 1106.910 ;
        RECT 36.180 1092.910 269.080 1098.910 ;
        RECT 89.140 1084.500 158.310 1090.500 ;
        RECT 95.110 1076.500 191.260 1082.500 ;
        RECT 3376.380 918.910 3559.070 924.910 ;
        RECT 3358.100 910.910 3553.000 916.910 ;
        RECT 3429.620 902.500 3500.040 908.500 ;
        RECT 3396.670 894.500 3494.070 900.500 ;
        RECT 3376.380 692.910 3559.070 698.910 ;
        RECT 3358.100 684.910 3553.000 690.910 ;
        RECT 3429.620 676.500 3500.040 682.500 ;
        RECT 3396.670 668.500 3494.070 674.500 ;
        RECT 197.280 390.755 229.220 413.720 ;
        RECT 197.280 341.280 229.220 364.500 ;
        RECT 740.340 169.500 744.630 203.910 ;
        RECT 748.000 175.570 752.290 206.035 ;
        RECT 1208.450 197.130 1230.245 233.430 ;
        RECT 1256.500 197.130 1278.510 233.430 ;
        RECT 3240.520 232.950 3248.350 235.940 ;
        RECT 3209.770 169.600 3218.470 220.130 ;
        RECT 3267.310 179.040 3284.550 225.780 ;
      LAYER via3 ;
        RECT 3376.990 4512.240 3382.400 4517.730 ;
        RECT 3554.870 4512.120 3558.370 4517.690 ;
        RECT 3358.460 4504.150 3363.870 4509.640 ;
        RECT 3548.880 4504.140 3552.380 4509.710 ;
        RECT 3430.010 4495.770 3433.780 4501.160 ;
        RECT 3495.950 4495.680 3499.700 4501.340 ;
        RECT 3397.280 4487.900 3401.090 4493.320 ;
        RECT 3489.930 4487.690 3493.680 4493.350 ;
        RECT 239.540 4189.000 248.470 4211.620 ;
        RECT 239.540 4139.340 248.470 4161.960 ;
        RECT 3336.420 4143.150 3348.660 4166.030 ;
        RECT 30.760 4115.120 34.260 4120.690 ;
        RECT 271.230 4115.240 276.640 4120.730 ;
        RECT 36.750 4107.140 40.250 4112.710 ;
        RECT 263.260 4107.150 268.670 4112.640 ;
        RECT 89.430 4098.680 93.180 4104.340 ;
        RECT 154.100 4098.770 157.870 4104.160 ;
        RECT 95.450 4090.690 99.200 4096.350 ;
        RECT 186.790 4090.900 190.600 4096.320 ;
        RECT 3336.350 4093.180 3348.590 4116.060 ;
        RECT 30.760 3899.120 34.260 3904.690 ;
        RECT 271.230 3899.240 276.640 3904.730 ;
        RECT 36.750 3891.140 40.250 3896.710 ;
        RECT 263.260 3891.150 268.670 3896.640 ;
        RECT 89.430 3882.680 93.180 3888.340 ;
        RECT 154.100 3882.770 157.870 3888.160 ;
        RECT 95.450 3874.690 99.200 3880.350 ;
        RECT 186.790 3874.900 190.600 3880.320 ;
        RECT 30.760 3683.120 34.260 3688.690 ;
        RECT 271.230 3683.240 276.640 3688.730 ;
        RECT 36.750 3675.140 40.250 3680.710 ;
        RECT 263.260 3675.150 268.670 3680.640 ;
        RECT 89.430 3666.680 93.180 3672.340 ;
        RECT 154.100 3666.770 157.870 3672.160 ;
        RECT 95.450 3658.690 99.200 3664.350 ;
        RECT 186.790 3658.900 190.600 3664.320 ;
        RECT 3377.040 3609.240 3382.450 3614.730 ;
        RECT 3554.920 3609.120 3558.420 3614.690 ;
        RECT 3358.510 3601.150 3363.920 3606.640 ;
        RECT 3548.930 3601.140 3552.430 3606.710 ;
        RECT 3430.060 3592.770 3433.830 3598.160 ;
        RECT 3496.000 3592.680 3499.750 3598.340 ;
        RECT 3397.330 3584.900 3401.140 3590.320 ;
        RECT 3489.980 3584.690 3493.730 3590.350 ;
        RECT 30.760 3467.120 34.260 3472.690 ;
        RECT 271.230 3467.240 276.640 3472.730 ;
        RECT 36.750 3459.140 40.250 3464.710 ;
        RECT 263.260 3459.150 268.670 3464.640 ;
        RECT 89.430 3450.680 93.180 3456.340 ;
        RECT 154.100 3450.770 157.870 3456.160 ;
        RECT 95.450 3442.690 99.200 3448.350 ;
        RECT 186.790 3442.900 190.600 3448.320 ;
        RECT 3377.040 3383.240 3382.450 3388.730 ;
        RECT 3554.920 3383.120 3558.420 3388.690 ;
        RECT 3358.510 3375.150 3363.920 3380.640 ;
        RECT 3548.930 3375.140 3552.430 3380.710 ;
        RECT 3430.060 3366.770 3433.830 3372.160 ;
        RECT 3496.000 3366.680 3499.750 3372.340 ;
        RECT 3397.330 3358.900 3401.140 3364.320 ;
        RECT 3489.980 3358.690 3493.730 3364.350 ;
        RECT 30.760 3251.120 34.260 3256.690 ;
        RECT 271.230 3251.240 276.640 3256.730 ;
        RECT 36.750 3243.140 40.250 3248.710 ;
        RECT 263.260 3243.150 268.670 3248.640 ;
        RECT 89.430 3234.680 93.180 3240.340 ;
        RECT 154.100 3234.770 157.870 3240.160 ;
        RECT 95.450 3226.690 99.200 3232.350 ;
        RECT 186.790 3226.900 190.600 3232.320 ;
        RECT 3377.040 3158.240 3382.450 3163.730 ;
        RECT 3554.920 3158.120 3558.420 3163.690 ;
        RECT 3358.510 3150.150 3363.920 3155.640 ;
        RECT 3548.930 3150.140 3552.430 3155.710 ;
        RECT 3430.060 3141.770 3433.830 3147.160 ;
        RECT 3496.000 3141.680 3499.750 3147.340 ;
        RECT 3397.330 3133.900 3401.140 3139.320 ;
        RECT 3489.980 3133.690 3493.730 3139.350 ;
        RECT 30.760 3035.120 34.260 3040.690 ;
        RECT 271.230 3035.240 276.640 3040.730 ;
        RECT 36.750 3027.140 40.250 3032.710 ;
        RECT 263.260 3027.150 268.670 3032.640 ;
        RECT 89.430 3018.680 93.180 3024.340 ;
        RECT 154.100 3018.770 157.870 3024.160 ;
        RECT 95.450 3010.690 99.200 3016.350 ;
        RECT 186.790 3010.900 190.600 3016.320 ;
        RECT 3377.040 2932.240 3382.450 2937.730 ;
        RECT 3554.920 2932.120 3558.420 2937.690 ;
        RECT 3358.510 2924.150 3363.920 2929.640 ;
        RECT 3548.930 2924.140 3552.430 2929.710 ;
        RECT 3430.060 2915.770 3433.830 2921.160 ;
        RECT 3496.000 2915.680 3499.750 2921.340 ;
        RECT 3397.330 2907.900 3401.140 2913.320 ;
        RECT 3489.980 2907.690 3493.730 2913.350 ;
        RECT 30.760 2819.120 34.260 2824.690 ;
        RECT 271.230 2819.240 276.640 2824.730 ;
        RECT 36.750 2811.140 40.250 2816.710 ;
        RECT 263.260 2811.150 268.670 2816.640 ;
        RECT 89.430 2802.680 93.180 2808.340 ;
        RECT 154.100 2802.770 157.870 2808.160 ;
        RECT 95.450 2794.690 99.200 2800.350 ;
        RECT 186.790 2794.900 190.600 2800.320 ;
        RECT 3377.040 2707.240 3382.450 2712.730 ;
        RECT 3554.920 2707.120 3558.420 2712.690 ;
        RECT 3358.510 2699.150 3363.920 2704.640 ;
        RECT 3548.930 2699.140 3552.430 2704.710 ;
        RECT 3430.060 2690.770 3433.830 2696.160 ;
        RECT 3496.000 2690.680 3499.750 2696.340 ;
        RECT 3397.330 2682.900 3401.140 2688.320 ;
        RECT 3489.980 2682.690 3493.730 2688.350 ;
        RECT 3336.680 2570.280 3348.530 2592.910 ;
        RECT 3336.750 2520.330 3348.600 2542.960 ;
        RECT 251.820 2466.250 260.460 2488.660 ;
        RECT 3377.040 2487.240 3382.450 2492.730 ;
        RECT 3554.920 2487.120 3558.420 2492.690 ;
        RECT 3358.510 2479.150 3363.920 2484.640 ;
        RECT 3548.930 2479.140 3552.430 2484.710 ;
        RECT 3430.060 2470.770 3433.830 2476.160 ;
        RECT 3496.000 2470.680 3499.750 2476.340 ;
        RECT 3397.330 2462.900 3401.140 2468.320 ;
        RECT 3489.980 2462.690 3493.730 2468.350 ;
        RECT 251.760 2416.300 260.400 2438.710 ;
        RECT 30.760 2181.120 34.260 2186.690 ;
        RECT 271.230 2181.240 276.640 2186.730 ;
        RECT 36.750 2173.140 40.250 2178.710 ;
        RECT 263.260 2173.150 268.670 2178.640 ;
        RECT 89.430 2164.680 93.180 2170.340 ;
        RECT 154.100 2164.770 157.870 2170.160 ;
        RECT 95.450 2156.690 99.200 2162.350 ;
        RECT 186.790 2156.900 190.600 2162.320 ;
        RECT 3320.670 2128.420 3332.700 2151.950 ;
        RECT 3320.560 2079.280 3332.640 2102.310 ;
        RECT 3377.040 2046.240 3382.450 2051.730 ;
        RECT 3554.920 2046.120 3558.420 2051.690 ;
        RECT 3358.510 2038.150 3363.920 2043.640 ;
        RECT 3548.930 2038.140 3552.430 2043.710 ;
        RECT 3430.060 2029.770 3433.830 2035.160 ;
        RECT 3496.000 2029.680 3499.750 2035.340 ;
        RECT 3397.330 2021.900 3401.140 2027.320 ;
        RECT 3489.980 2021.690 3493.730 2027.350 ;
        RECT 30.760 1965.120 34.260 1970.690 ;
        RECT 271.230 1965.240 276.640 1970.730 ;
        RECT 36.750 1957.140 40.250 1962.710 ;
        RECT 263.260 1957.150 268.670 1962.640 ;
        RECT 89.430 1948.680 93.180 1954.340 ;
        RECT 154.100 1948.770 157.870 1954.160 ;
        RECT 95.450 1940.690 99.200 1946.350 ;
        RECT 186.790 1940.900 190.600 1946.320 ;
        RECT 3377.040 1820.240 3382.450 1825.730 ;
        RECT 3554.920 1820.120 3558.420 1825.690 ;
        RECT 3358.510 1812.150 3363.920 1817.640 ;
        RECT 3548.930 1812.140 3552.430 1817.710 ;
        RECT 3430.060 1803.770 3433.830 1809.160 ;
        RECT 3496.000 1803.680 3499.750 1809.340 ;
        RECT 3397.330 1795.900 3401.140 1801.320 ;
        RECT 3489.980 1795.690 3493.730 1801.350 ;
        RECT 30.760 1749.120 34.260 1754.690 ;
        RECT 271.230 1749.240 276.640 1754.730 ;
        RECT 36.750 1741.140 40.250 1746.710 ;
        RECT 263.260 1741.150 268.670 1746.640 ;
        RECT 89.430 1732.680 93.180 1738.340 ;
        RECT 154.100 1732.770 157.870 1738.160 ;
        RECT 95.450 1724.690 99.200 1730.350 ;
        RECT 186.790 1724.900 190.600 1730.320 ;
        RECT 3377.040 1595.240 3382.450 1600.730 ;
        RECT 3554.920 1595.120 3558.420 1600.690 ;
        RECT 3358.510 1587.150 3363.920 1592.640 ;
        RECT 3548.930 1587.140 3552.430 1592.710 ;
        RECT 3430.060 1578.770 3433.830 1584.160 ;
        RECT 3496.000 1578.680 3499.750 1584.340 ;
        RECT 3397.330 1570.900 3401.140 1576.320 ;
        RECT 3489.980 1570.690 3493.730 1576.350 ;
        RECT 30.760 1533.120 34.260 1538.690 ;
        RECT 271.230 1533.240 276.640 1538.730 ;
        RECT 36.750 1525.140 40.250 1530.710 ;
        RECT 263.260 1525.150 268.670 1530.640 ;
        RECT 89.430 1516.680 93.180 1522.340 ;
        RECT 154.100 1516.770 157.870 1522.160 ;
        RECT 95.450 1508.690 99.200 1514.350 ;
        RECT 186.790 1508.900 190.600 1514.320 ;
        RECT 3377.040 1370.240 3382.450 1375.730 ;
        RECT 3554.920 1370.120 3558.420 1375.690 ;
        RECT 3358.510 1362.150 3363.920 1367.640 ;
        RECT 3548.930 1362.140 3552.430 1367.710 ;
        RECT 3430.060 1353.770 3433.830 1359.160 ;
        RECT 3496.000 1353.680 3499.750 1359.340 ;
        RECT 3397.330 1345.900 3401.140 1351.320 ;
        RECT 3489.980 1345.690 3493.730 1351.350 ;
        RECT 30.760 1317.120 34.260 1322.690 ;
        RECT 271.230 1317.240 276.640 1322.730 ;
        RECT 36.750 1309.140 40.250 1314.710 ;
        RECT 263.260 1309.150 268.670 1314.640 ;
        RECT 89.430 1300.680 93.180 1306.340 ;
        RECT 154.100 1300.770 157.870 1306.160 ;
        RECT 95.450 1292.690 99.200 1298.350 ;
        RECT 186.790 1292.900 190.600 1298.320 ;
        RECT 3377.040 1144.240 3382.450 1149.730 ;
        RECT 3554.920 1144.120 3558.420 1149.690 ;
        RECT 3358.510 1136.150 3363.920 1141.640 ;
        RECT 3548.930 1136.140 3552.430 1141.710 ;
        RECT 3430.060 1127.770 3433.830 1133.160 ;
        RECT 3496.000 1127.680 3499.750 1133.340 ;
        RECT 3397.330 1119.900 3401.140 1125.320 ;
        RECT 3489.980 1119.690 3493.730 1125.350 ;
        RECT 30.760 1101.120 34.260 1106.690 ;
        RECT 271.230 1101.240 276.640 1106.730 ;
        RECT 36.750 1093.140 40.250 1098.710 ;
        RECT 263.260 1093.150 268.670 1098.640 ;
        RECT 89.430 1084.680 93.180 1090.340 ;
        RECT 154.100 1084.770 157.870 1090.160 ;
        RECT 95.450 1076.690 99.200 1082.350 ;
        RECT 186.790 1076.900 190.600 1082.320 ;
        RECT 3377.040 919.240 3382.450 924.730 ;
        RECT 3554.920 919.120 3558.420 924.690 ;
        RECT 3358.510 911.150 3363.920 916.640 ;
        RECT 3548.930 911.140 3552.430 916.710 ;
        RECT 3430.060 902.770 3433.830 908.160 ;
        RECT 3496.000 902.680 3499.750 908.340 ;
        RECT 3397.330 894.900 3401.140 900.320 ;
        RECT 3489.980 894.690 3493.730 900.350 ;
        RECT 3377.040 693.240 3382.450 698.730 ;
        RECT 3554.920 693.120 3558.420 698.690 ;
        RECT 3358.510 685.150 3363.920 690.640 ;
        RECT 3548.930 685.140 3552.430 690.710 ;
        RECT 3430.060 676.770 3433.830 682.160 ;
        RECT 3496.000 676.680 3499.750 682.340 ;
        RECT 3397.330 668.900 3401.140 674.320 ;
        RECT 3489.980 668.690 3493.730 674.350 ;
        RECT 209.730 391.210 228.360 413.530 ;
        RECT 209.610 341.690 228.240 364.010 ;
        RECT 1208.700 214.210 1229.930 233.080 ;
        RECT 748.090 204.940 752.200 205.740 ;
        RECT 740.430 202.960 744.540 203.760 ;
        RECT 1256.960 214.280 1278.190 233.150 ;
        RECT 3240.830 233.300 3248.040 235.620 ;
        RECT 3209.970 210.990 3218.300 219.940 ;
        RECT 748.160 175.830 752.180 179.980 ;
        RECT 740.490 169.790 744.510 173.940 ;
        RECT 3267.890 213.170 3283.860 225.130 ;
        RECT 3210.130 169.940 3218.170 173.800 ;
      LAYER met4 ;
        RECT 2878.400 4974.020 2902.390 4987.310 ;
        RECT 2928.350 4974.020 2952.340 4987.310 ;
        RECT 3376.680 4511.870 3382.710 4517.940 ;
        RECT 3358.200 4503.870 3364.230 4509.940 ;
        RECT 3430.010 4495.770 3433.780 4501.160 ;
        RECT 3397.280 4487.900 3401.090 4493.320 ;
        RECT 3489.780 4429.740 3493.780 4494.660 ;
        RECT 3495.780 4438.110 3499.780 4501.550 ;
        RECT 3548.600 4443.380 3552.600 4510.210 ;
        RECT 3554.600 4434.730 3558.600 4518.350 ;
        RECT 238.960 4188.290 249.110 4212.310 ;
        RECT 238.960 4138.510 249.110 4162.530 ;
        RECT 3336.010 4142.600 3349.010 4166.550 ;
        RECT 30.530 4037.730 34.530 4121.350 ;
        RECT 270.920 4114.870 276.950 4120.940 ;
        RECT 36.530 4046.380 40.530 4113.210 ;
        RECT 262.900 4106.870 268.930 4112.940 ;
        RECT 89.350 4041.110 93.350 4104.550 ;
        RECT 154.100 4098.770 157.870 4104.160 ;
        RECT 95.350 4032.740 99.350 4097.660 ;
        RECT 186.790 4090.900 190.600 4096.320 ;
        RECT 3336.070 4092.730 3349.070 4116.680 ;
        RECT 30.530 3821.730 34.530 3905.350 ;
        RECT 270.920 3898.870 276.950 3904.940 ;
        RECT 36.530 3830.380 40.530 3897.210 ;
        RECT 262.900 3890.870 268.930 3896.940 ;
        RECT 89.350 3825.110 93.350 3888.550 ;
        RECT 154.100 3882.770 157.870 3888.160 ;
        RECT 95.350 3816.740 99.350 3881.660 ;
        RECT 186.790 3874.900 190.600 3880.320 ;
        RECT 30.530 3605.730 34.530 3689.350 ;
        RECT 270.920 3682.870 276.950 3688.940 ;
        RECT 36.530 3614.380 40.530 3681.210 ;
        RECT 262.900 3674.870 268.930 3680.940 ;
        RECT 89.350 3609.110 93.350 3672.550 ;
        RECT 154.100 3666.770 157.870 3672.160 ;
        RECT 95.350 3600.740 99.350 3665.660 ;
        RECT 186.790 3658.900 190.600 3664.320 ;
        RECT 3376.730 3608.870 3382.760 3614.940 ;
        RECT 3358.250 3600.870 3364.280 3606.940 ;
        RECT 3430.060 3592.770 3433.830 3598.160 ;
        RECT 3397.330 3584.900 3401.140 3590.320 ;
        RECT 3489.830 3526.740 3493.830 3591.660 ;
        RECT 3495.830 3535.110 3499.830 3598.550 ;
        RECT 3548.650 3540.380 3552.650 3607.210 ;
        RECT 3554.650 3531.730 3558.650 3615.350 ;
        RECT 30.530 3389.730 34.530 3473.350 ;
        RECT 270.920 3466.870 276.950 3472.940 ;
        RECT 36.530 3398.380 40.530 3465.210 ;
        RECT 262.900 3458.870 268.930 3464.940 ;
        RECT 89.350 3393.110 93.350 3456.550 ;
        RECT 154.100 3450.770 157.870 3456.160 ;
        RECT 95.350 3384.740 99.350 3449.660 ;
        RECT 186.790 3442.900 190.600 3448.320 ;
        RECT 3376.730 3382.870 3382.760 3388.940 ;
        RECT 3358.250 3374.870 3364.280 3380.940 ;
        RECT 3430.060 3366.770 3433.830 3372.160 ;
        RECT 3397.330 3358.900 3401.140 3364.320 ;
        RECT 3489.830 3300.740 3493.830 3365.660 ;
        RECT 3495.830 3309.110 3499.830 3372.550 ;
        RECT 3548.650 3314.380 3552.650 3381.210 ;
        RECT 3554.650 3305.730 3558.650 3389.350 ;
        RECT 30.530 3173.730 34.530 3257.350 ;
        RECT 270.920 3250.870 276.950 3256.940 ;
        RECT 36.530 3182.380 40.530 3249.210 ;
        RECT 262.900 3242.870 268.930 3248.940 ;
        RECT 89.350 3177.110 93.350 3240.550 ;
        RECT 154.100 3234.770 157.870 3240.160 ;
        RECT 95.350 3168.740 99.350 3233.660 ;
        RECT 186.790 3226.900 190.600 3232.320 ;
        RECT 3376.730 3157.870 3382.760 3163.940 ;
        RECT 3358.250 3149.870 3364.280 3155.940 ;
        RECT 3430.060 3141.770 3433.830 3147.160 ;
        RECT 3397.330 3133.900 3401.140 3139.320 ;
        RECT 3489.830 3075.740 3493.830 3140.660 ;
        RECT 3495.830 3084.110 3499.830 3147.550 ;
        RECT 3548.650 3089.380 3552.650 3156.210 ;
        RECT 3554.650 3080.730 3558.650 3164.350 ;
        RECT 30.530 2957.730 34.530 3041.350 ;
        RECT 270.920 3034.870 276.950 3040.940 ;
        RECT 36.530 2966.380 40.530 3033.210 ;
        RECT 262.900 3026.870 268.930 3032.940 ;
        RECT 89.350 2961.110 93.350 3024.550 ;
        RECT 154.100 3018.770 157.870 3024.160 ;
        RECT 95.350 2952.740 99.350 3017.660 ;
        RECT 186.790 3010.900 190.600 3016.320 ;
        RECT 3376.730 2931.870 3382.760 2937.940 ;
        RECT 3358.250 2923.870 3364.280 2929.940 ;
        RECT 3430.060 2915.770 3433.830 2921.160 ;
        RECT 3397.330 2907.900 3401.140 2913.320 ;
        RECT 3489.830 2849.740 3493.830 2914.660 ;
        RECT 3495.830 2858.110 3499.830 2921.550 ;
        RECT 3548.650 2863.380 3552.650 2930.210 ;
        RECT 3554.650 2854.730 3558.650 2938.350 ;
        RECT 30.530 2741.730 34.530 2825.350 ;
        RECT 270.920 2818.870 276.950 2824.940 ;
        RECT 36.530 2750.380 40.530 2817.210 ;
        RECT 262.900 2810.870 268.930 2816.940 ;
        RECT 89.350 2745.110 93.350 2808.550 ;
        RECT 154.100 2802.770 157.870 2808.160 ;
        RECT 95.350 2736.740 99.350 2801.660 ;
        RECT 186.790 2794.900 190.600 2800.320 ;
        RECT 3376.730 2706.870 3382.760 2712.940 ;
        RECT 3358.250 2698.870 3364.280 2704.940 ;
        RECT 3430.060 2690.770 3433.830 2696.160 ;
        RECT 3397.330 2682.900 3401.140 2688.320 ;
        RECT 3489.830 2624.740 3493.830 2689.660 ;
        RECT 3495.830 2633.110 3499.830 2696.550 ;
        RECT 3548.650 2638.380 3552.650 2705.210 ;
        RECT 3554.650 2629.730 3558.650 2713.350 ;
        RECT 3336.030 2569.600 3349.070 2593.480 ;
        RECT 3336.090 2519.750 3349.130 2543.630 ;
        RECT 250.860 2465.420 260.980 2489.370 ;
        RECT 3376.730 2486.870 3382.760 2492.940 ;
        RECT 3358.250 2478.870 3364.280 2484.940 ;
        RECT 3430.060 2470.770 3433.830 2476.160 ;
        RECT 3397.330 2462.900 3401.140 2468.320 ;
        RECT 250.990 2415.470 261.110 2439.420 ;
        RECT 3489.830 2404.740 3493.830 2469.660 ;
        RECT 3495.830 2413.110 3499.830 2476.550 ;
        RECT 3548.650 2418.380 3552.650 2485.210 ;
        RECT 3554.650 2409.730 3558.650 2493.350 ;
        RECT 30.530 2103.730 34.530 2187.350 ;
        RECT 270.920 2180.870 276.950 2186.940 ;
        RECT 36.530 2112.380 40.530 2179.210 ;
        RECT 262.900 2172.870 268.930 2178.940 ;
        RECT 89.350 2107.110 93.350 2170.550 ;
        RECT 154.100 2164.770 157.870 2170.160 ;
        RECT 95.350 2098.740 99.350 2163.660 ;
        RECT 186.790 2156.900 190.600 2162.320 ;
        RECT 3320.040 2127.860 3333.060 2152.450 ;
        RECT 3320.090 2078.800 3333.170 2102.620 ;
        RECT 3376.730 2045.870 3382.760 2051.940 ;
        RECT 3358.250 2037.870 3364.280 2043.940 ;
        RECT 3430.060 2029.770 3433.830 2035.160 ;
        RECT 3397.330 2021.900 3401.140 2027.320 ;
        RECT 30.530 1887.730 34.530 1971.350 ;
        RECT 270.920 1964.870 276.950 1970.940 ;
        RECT 3489.830 1963.740 3493.830 2028.660 ;
        RECT 3495.830 1972.110 3499.830 2035.550 ;
        RECT 3548.650 1977.380 3552.650 2044.210 ;
        RECT 3554.650 1968.730 3558.650 2052.350 ;
        RECT 36.530 1896.380 40.530 1963.210 ;
        RECT 262.900 1956.870 268.930 1962.940 ;
        RECT 89.350 1891.110 93.350 1954.550 ;
        RECT 154.100 1948.770 157.870 1954.160 ;
        RECT 95.350 1882.740 99.350 1947.660 ;
        RECT 186.790 1940.900 190.600 1946.320 ;
        RECT 3376.730 1819.870 3382.760 1825.940 ;
        RECT 3358.250 1811.870 3364.280 1817.940 ;
        RECT 3430.060 1803.770 3433.830 1809.160 ;
        RECT 3397.330 1795.900 3401.140 1801.320 ;
        RECT 30.530 1671.730 34.530 1755.350 ;
        RECT 270.920 1748.870 276.950 1754.940 ;
        RECT 36.530 1680.380 40.530 1747.210 ;
        RECT 262.900 1740.870 268.930 1746.940 ;
        RECT 89.350 1675.110 93.350 1738.550 ;
        RECT 154.100 1732.770 157.870 1738.160 ;
        RECT 3489.830 1737.740 3493.830 1802.660 ;
        RECT 3495.830 1746.110 3499.830 1809.550 ;
        RECT 3548.650 1751.380 3552.650 1818.210 ;
        RECT 3554.650 1742.730 3558.650 1826.350 ;
        RECT 95.350 1666.740 99.350 1731.660 ;
        RECT 186.790 1724.900 190.600 1730.320 ;
        RECT 3376.730 1594.870 3382.760 1600.940 ;
        RECT 3358.250 1586.870 3364.280 1592.940 ;
        RECT 3430.060 1578.770 3433.830 1584.160 ;
        RECT 3397.330 1570.900 3401.140 1576.320 ;
        RECT 30.530 1455.730 34.530 1539.350 ;
        RECT 270.920 1532.870 276.950 1538.940 ;
        RECT 36.530 1464.380 40.530 1531.210 ;
        RECT 262.900 1524.870 268.930 1530.940 ;
        RECT 89.350 1459.110 93.350 1522.550 ;
        RECT 154.100 1516.770 157.870 1522.160 ;
        RECT 95.350 1450.740 99.350 1515.660 ;
        RECT 186.790 1508.900 190.600 1514.320 ;
        RECT 3489.830 1512.740 3493.830 1577.660 ;
        RECT 3495.830 1521.110 3499.830 1584.550 ;
        RECT 3548.650 1526.380 3552.650 1593.210 ;
        RECT 3554.650 1517.730 3558.650 1601.350 ;
        RECT 3376.730 1369.870 3382.760 1375.940 ;
        RECT 3358.250 1361.870 3364.280 1367.940 ;
        RECT 3430.060 1353.770 3433.830 1359.160 ;
        RECT 1967.210 1332.370 1971.140 1347.350 ;
        RECT 3397.330 1345.900 3401.140 1351.320 ;
        RECT 30.530 1239.730 34.530 1323.350 ;
        RECT 270.920 1316.870 276.950 1322.940 ;
        RECT 36.530 1248.380 40.530 1315.210 ;
        RECT 262.900 1308.870 268.930 1314.940 ;
        RECT 1970.220 1311.040 1971.120 1332.370 ;
        RECT 2045.470 1327.310 2046.370 1327.380 ;
        RECT 2042.330 1314.270 2046.370 1327.310 ;
        RECT 2045.470 1311.220 2046.370 1314.270 ;
        RECT 89.350 1243.110 93.350 1306.550 ;
        RECT 154.100 1300.770 157.870 1306.160 ;
        RECT 95.350 1234.740 99.350 1299.660 ;
        RECT 186.790 1292.900 190.600 1298.320 ;
        RECT 238.850 1292.330 297.350 1307.330 ;
        RECT 1972.520 1292.340 1977.030 1307.250 ;
        RECT 3489.830 1287.740 3493.830 1352.660 ;
        RECT 3495.830 1296.110 3499.830 1359.550 ;
        RECT 3548.650 1301.380 3552.650 1368.210 ;
        RECT 3554.650 1292.730 3558.650 1376.350 ;
        RECT 250.850 1272.330 302.940 1287.330 ;
        RECT 2048.430 1272.260 2054.040 1287.350 ;
        RECT 262.890 1252.330 316.460 1267.330 ;
        RECT 1058.560 1252.350 1063.050 1267.360 ;
        RECT 1209.060 1252.350 1213.550 1267.360 ;
        RECT 1361.160 1252.350 1363.100 1267.360 ;
        RECT 1510.810 1252.350 1513.570 1267.360 ;
        RECT 1660.560 1252.350 1665.050 1267.360 ;
        RECT 1811.060 1252.350 1815.550 1267.360 ;
        RECT 1962.860 1252.350 1965.550 1267.360 ;
        RECT 983.380 1232.340 988.090 1247.320 ;
        RECT 1133.880 1232.340 1138.590 1247.320 ;
        RECT 1284.380 1232.340 1289.090 1247.320 ;
        RECT 1435.780 1233.950 1438.290 1247.320 ;
        RECT 1586.770 1232.340 1589.010 1246.620 ;
        RECT 1735.880 1232.340 1740.590 1247.320 ;
        RECT 1885.880 1232.340 1890.590 1247.320 ;
        RECT 2035.880 1232.340 2040.590 1247.320 ;
        RECT 3334.450 1232.330 3383.350 1247.380 ;
        RECT 204.920 1212.330 317.170 1227.330 ;
        RECT 204.920 1191.330 218.060 1212.330 ;
        RECT 1062.840 1212.320 1067.700 1227.310 ;
        RECT 1213.340 1212.320 1218.200 1227.310 ;
        RECT 1364.910 1212.320 1366.570 1227.310 ;
        RECT 1515.840 1212.320 1517.300 1227.310 ;
        RECT 1664.840 1212.320 1669.700 1227.310 ;
        RECT 1815.340 1212.320 1820.200 1227.310 ;
        RECT 1966.050 1212.320 1969.000 1227.310 ;
        RECT 220.980 1192.330 317.170 1207.330 ;
        RECT 987.710 1192.400 991.990 1207.350 ;
        RECT 1138.210 1192.400 1142.490 1207.350 ;
        RECT 1288.710 1192.400 1292.990 1207.350 ;
        RECT 1440.340 1192.400 1442.830 1207.350 ;
        RECT 1591.130 1192.400 1592.870 1207.350 ;
        RECT 1740.210 1192.400 1744.490 1207.350 ;
        RECT 1890.210 1192.400 1894.490 1207.350 ;
        RECT 2042.050 1192.400 2043.670 1207.350 ;
        RECT 220.980 1172.330 234.010 1192.330 ;
        RECT 238.930 1172.330 316.250 1187.330 ;
        RECT 1054.330 1172.240 1059.070 1187.370 ;
        RECT 1204.830 1172.240 1209.570 1187.370 ;
        RECT 1356.720 1172.240 1360.070 1187.370 ;
        RECT 1507.570 1172.240 1510.570 1186.450 ;
        RECT 1657.070 1172.240 1661.070 1187.370 ;
        RECT 1806.830 1172.240 1811.570 1187.370 ;
        RECT 1959.170 1172.240 1961.570 1187.370 ;
        RECT 220.930 1152.330 315.800 1167.330 ;
        RECT 448.880 1161.930 450.480 1168.010 ;
        RECT 468.880 1161.930 470.480 1168.010 ;
        RECT 448.880 1156.330 470.480 1161.930 ;
        RECT 848.880 1161.690 850.480 1168.190 ;
        RECT 868.880 1161.690 870.480 1168.060 ;
        RECT 848.880 1156.510 870.480 1161.690 ;
        RECT 979.940 1152.330 983.080 1167.320 ;
        RECT 1130.440 1152.330 1133.580 1167.320 ;
        RECT 1280.940 1152.330 1284.080 1167.320 ;
        RECT 1431.440 1152.330 1434.580 1167.320 ;
        RECT 1581.940 1152.330 1585.080 1167.320 ;
        RECT 1732.440 1152.330 1735.580 1167.320 ;
        RECT 1882.440 1152.330 1885.580 1167.320 ;
        RECT 2033.300 1152.330 2035.580 1167.320 ;
        RECT 2148.880 1162.600 2150.480 1168.060 ;
        RECT 2168.880 1162.600 2170.480 1168.060 ;
        RECT 2148.880 1156.960 2170.480 1162.600 ;
        RECT 30.530 1023.730 34.530 1107.350 ;
        RECT 36.530 1032.380 40.530 1099.210 ;
        RECT 89.350 1027.110 93.350 1090.550 ;
        RECT 154.100 1084.770 157.870 1090.160 ;
        RECT 95.350 1018.740 99.350 1083.660 ;
        RECT 186.790 1076.900 190.600 1082.320 ;
        RECT 220.990 987.490 233.990 1152.330 ;
        RECT 3376.730 1143.870 3382.760 1149.940 ;
        RECT 3358.250 1135.870 3364.280 1141.940 ;
        RECT 3430.060 1127.770 3433.830 1133.160 ;
        RECT 3397.330 1119.900 3401.140 1125.320 ;
        RECT 270.920 1100.870 276.950 1106.940 ;
        RECT 262.900 1092.870 268.930 1098.940 ;
        RECT 2991.840 1047.520 3054.810 1062.520 ;
        RECT 3205.220 1047.640 3210.540 1062.300 ;
        RECT 3489.830 1061.740 3493.830 1126.660 ;
        RECT 3495.830 1070.110 3499.830 1133.550 ;
        RECT 3548.650 1075.380 3552.650 1142.210 ;
        RECT 3554.650 1066.730 3558.650 1150.350 ;
        RECT 2981.310 1039.310 3026.940 1042.510 ;
        RECT 3053.210 1038.460 3054.810 1047.520 ;
        RECT 3206.810 1038.420 3208.410 1047.640 ;
        RECT 2992.480 987.640 3005.870 989.380 ;
        RECT 220.990 984.290 261.720 987.490 ;
        RECT 2992.480 986.040 3034.880 987.640 ;
        RECT 2992.480 984.960 3005.870 986.040 ;
        RECT 220.990 883.710 233.990 984.290 ;
        RECT 2980.360 919.310 3026.940 922.510 ;
        RECT 3376.730 918.870 3382.760 924.940 ;
        RECT 3358.250 910.870 3364.280 916.940 ;
        RECT 3430.060 902.770 3433.830 908.160 ;
        RECT 3397.330 894.900 3401.140 900.320 ;
        RECT 209.320 865.630 233.990 883.710 ;
        RECT 213.230 854.290 261.230 857.490 ;
        RECT 3489.830 836.740 3493.830 901.660 ;
        RECT 3495.830 845.110 3499.830 908.550 ;
        RECT 3548.650 850.380 3552.650 917.210 ;
        RECT 3554.650 841.730 3558.650 925.350 ;
        RECT 2992.480 834.460 3005.870 836.180 ;
        RECT 2992.480 832.860 3034.880 834.460 ;
        RECT 2992.480 831.760 3005.870 832.860 ;
        RECT 2970.360 789.310 3026.940 792.510 ;
        RECT 212.890 724.290 260.890 727.490 ;
        RECT 3376.730 692.870 3382.760 698.940 ;
        RECT 3358.250 684.870 3364.280 690.940 ;
        RECT 2992.480 681.280 3005.870 682.980 ;
        RECT 2992.480 679.680 3034.880 681.280 ;
        RECT 2992.480 678.560 3005.870 679.680 ;
        RECT 3430.060 676.770 3433.830 682.160 ;
        RECT 3397.330 668.900 3401.140 674.320 ;
        RECT 2970.360 659.310 3026.940 662.510 ;
        RECT 3489.830 610.740 3493.830 675.660 ;
        RECT 3495.830 619.110 3499.830 682.550 ;
        RECT 3548.650 624.380 3552.650 691.210 ;
        RECT 3554.650 615.730 3558.650 699.350 ;
        RECT 212.890 594.290 260.890 597.490 ;
        RECT 2970.360 529.310 3026.940 532.510 ;
        RECT 2992.480 528.100 3005.870 528.380 ;
        RECT 2992.480 526.500 3034.880 528.100 ;
        RECT 2992.480 523.960 3005.870 526.500 ;
        RECT 3130.010 493.800 3131.610 511.580 ;
        RECT 3283.610 494.020 3285.210 511.190 ;
        RECT 3127.210 479.780 3134.260 493.800 ;
        RECT 3180.400 482.170 3184.970 493.790 ;
        RECT 3181.770 472.240 3183.370 482.170 ;
        RECT 3281.420 480.250 3288.010 494.020 ;
        RECT 212.890 464.290 260.890 467.490 ;
        RECT 209.320 390.770 228.890 413.970 ;
        RECT 3161.770 404.620 3163.370 410.310 ;
        RECT 3201.770 405.080 3203.370 410.000 ;
        RECT 2970.360 399.310 3026.940 402.510 ;
        RECT 3160.360 390.990 3165.050 404.620 ;
        RECT 3200.490 390.670 3204.610 405.080 ;
        RECT 3123.940 372.140 3125.540 388.490 ;
        RECT 3131.690 372.140 3133.290 388.490 ;
        RECT 3139.440 372.140 3141.040 388.490 ;
        RECT 3147.190 372.140 3148.790 388.490 ;
        RECT 3154.940 372.140 3156.540 388.490 ;
        RECT 3162.690 372.140 3164.290 388.490 ;
        RECT 3170.440 372.140 3172.040 388.490 ;
        RECT 3178.190 372.140 3179.790 388.490 ;
        RECT 3185.940 372.140 3187.540 388.490 ;
        RECT 3193.690 372.140 3195.290 388.490 ;
        RECT 209.290 341.250 228.860 364.450 ;
        RECT 209.310 334.290 261.810 337.490 ;
        RECT 209.370 241.110 292.680 260.610 ;
        RECT 716.620 249.680 723.690 253.440 ;
        RECT 719.300 248.190 720.200 249.680 ;
        RECT 3209.680 238.135 3251.010 240.135 ;
        RECT 712.800 226.980 713.700 236.280 ;
        RECT 708.880 226.970 714.330 226.980 ;
        RECT 706.880 220.650 714.330 226.970 ;
        RECT 717.200 203.810 718.100 236.480 ;
        RECT 723.700 205.790 724.600 236.700 ;
        RECT 1208.400 213.920 1230.280 233.460 ;
        RECT 1256.510 213.940 1278.500 233.420 ;
        RECT 3209.680 210.820 3218.590 238.135 ;
        RECT 3240.520 232.950 3248.350 235.940 ;
        RECT 3267.160 212.440 3284.560 235.270 ;
        RECT 3306.350 234.955 3347.130 236.600 ;
        RECT 723.700 204.890 752.580 205.790 ;
        RECT 717.200 202.910 744.700 203.810 ;
        RECT 748.160 175.830 752.180 179.980 ;
        RECT 740.490 169.790 744.510 173.940 ;
        RECT 3210.130 169.940 3218.170 173.800 ;
      LAYER via4 ;
        RECT 2878.810 4974.420 2901.920 4986.570 ;
        RECT 2928.790 4974.490 2951.900 4986.640 ;
        RECT 3376.990 4512.240 3382.400 4517.730 ;
        RECT 3358.460 4504.150 3363.870 4509.640 ;
        RECT 3495.900 4496.280 3499.680 4497.690 ;
        RECT 3489.900 4492.760 3493.680 4494.170 ;
        RECT 3489.860 4463.780 3493.720 4465.220 ;
        RECT 3489.840 4446.880 3493.700 4448.320 ;
        RECT 3495.840 4472.230 3499.700 4473.670 ;
        RECT 3495.870 4455.320 3499.730 4456.760 ;
        RECT 3548.680 4477.500 3552.510 4478.850 ;
        RECT 3548.690 4460.580 3552.520 4461.930 ;
        RECT 3548.680 4443.640 3552.550 4445.130 ;
        RECT 3554.690 4469.020 3558.520 4470.370 ;
        RECT 3554.660 4452.220 3558.490 4453.570 ;
        RECT 3495.860 4438.410 3499.720 4439.850 ;
        RECT 3554.650 4435.200 3558.520 4436.690 ;
        RECT 3489.840 4429.980 3493.700 4431.420 ;
        RECT 239.540 4189.000 248.470 4211.620 ;
        RECT 239.540 4139.340 248.470 4161.960 ;
        RECT 3336.420 4143.150 3348.660 4166.030 ;
        RECT 271.230 4115.240 276.640 4120.730 ;
        RECT 30.580 4072.030 34.440 4073.420 ;
        RECT 30.600 4055.200 34.480 4056.590 ;
        RECT 263.260 4107.150 268.670 4112.640 ;
        RECT 36.590 4080.440 40.460 4081.930 ;
        RECT 36.600 4063.590 40.460 4064.980 ;
        RECT 36.580 4046.640 40.450 4048.130 ;
        RECT 89.450 4099.280 93.230 4100.690 ;
        RECT 89.430 4075.230 93.290 4076.670 ;
        RECT 89.400 4058.320 93.260 4059.760 ;
        RECT 89.410 4041.410 93.270 4042.850 ;
        RECT 95.450 4095.760 99.230 4097.170 ;
        RECT 3336.350 4093.180 3348.590 4116.060 ;
        RECT 95.410 4066.780 99.270 4068.220 ;
        RECT 95.430 4049.880 99.290 4051.320 ;
        RECT 30.610 4038.200 34.480 4039.690 ;
        RECT 95.430 4032.980 99.290 4034.420 ;
        RECT 271.230 3899.240 276.640 3904.730 ;
        RECT 30.580 3856.030 34.440 3857.420 ;
        RECT 30.600 3839.200 34.480 3840.590 ;
        RECT 263.260 3891.150 268.670 3896.640 ;
        RECT 36.590 3864.440 40.460 3865.930 ;
        RECT 36.600 3847.590 40.460 3848.980 ;
        RECT 36.580 3830.640 40.450 3832.130 ;
        RECT 89.450 3883.280 93.230 3884.690 ;
        RECT 89.430 3859.230 93.290 3860.670 ;
        RECT 89.400 3842.320 93.260 3843.760 ;
        RECT 89.410 3825.410 93.270 3826.850 ;
        RECT 95.450 3879.760 99.230 3881.170 ;
        RECT 95.410 3850.780 99.270 3852.220 ;
        RECT 95.430 3833.880 99.290 3835.320 ;
        RECT 30.610 3822.200 34.480 3823.690 ;
        RECT 95.430 3816.980 99.290 3818.420 ;
        RECT 271.230 3683.240 276.640 3688.730 ;
        RECT 30.580 3640.030 34.440 3641.420 ;
        RECT 30.600 3623.200 34.480 3624.590 ;
        RECT 263.260 3675.150 268.670 3680.640 ;
        RECT 36.590 3648.440 40.460 3649.930 ;
        RECT 36.600 3631.590 40.460 3632.980 ;
        RECT 36.580 3614.640 40.450 3616.130 ;
        RECT 89.450 3667.280 93.230 3668.690 ;
        RECT 89.430 3643.230 93.290 3644.670 ;
        RECT 89.400 3626.320 93.260 3627.760 ;
        RECT 89.410 3609.410 93.270 3610.850 ;
        RECT 95.450 3663.760 99.230 3665.170 ;
        RECT 95.410 3634.780 99.270 3636.220 ;
        RECT 95.430 3617.880 99.290 3619.320 ;
        RECT 30.610 3606.200 34.480 3607.690 ;
        RECT 3377.040 3609.240 3382.450 3614.730 ;
        RECT 95.430 3600.980 99.290 3602.420 ;
        RECT 3358.510 3601.150 3363.920 3606.640 ;
        RECT 3495.950 3593.280 3499.730 3594.690 ;
        RECT 3489.950 3589.760 3493.730 3591.170 ;
        RECT 3489.910 3560.780 3493.770 3562.220 ;
        RECT 3489.890 3543.880 3493.750 3545.320 ;
        RECT 3495.890 3569.230 3499.750 3570.670 ;
        RECT 3495.920 3552.320 3499.780 3553.760 ;
        RECT 3548.730 3574.500 3552.560 3575.850 ;
        RECT 3548.740 3557.580 3552.570 3558.930 ;
        RECT 3548.730 3540.640 3552.600 3542.130 ;
        RECT 3554.740 3566.020 3558.570 3567.370 ;
        RECT 3554.710 3549.220 3558.540 3550.570 ;
        RECT 3495.910 3535.410 3499.770 3536.850 ;
        RECT 3554.700 3532.200 3558.570 3533.690 ;
        RECT 3489.890 3526.980 3493.750 3528.420 ;
        RECT 271.230 3467.240 276.640 3472.730 ;
        RECT 30.580 3424.030 34.440 3425.420 ;
        RECT 30.600 3407.200 34.480 3408.590 ;
        RECT 263.260 3459.150 268.670 3464.640 ;
        RECT 36.590 3432.440 40.460 3433.930 ;
        RECT 36.600 3415.590 40.460 3416.980 ;
        RECT 36.580 3398.640 40.450 3400.130 ;
        RECT 89.450 3451.280 93.230 3452.690 ;
        RECT 89.430 3427.230 93.290 3428.670 ;
        RECT 89.400 3410.320 93.260 3411.760 ;
        RECT 89.410 3393.410 93.270 3394.850 ;
        RECT 95.450 3447.760 99.230 3449.170 ;
        RECT 95.410 3418.780 99.270 3420.220 ;
        RECT 95.430 3401.880 99.290 3403.320 ;
        RECT 30.610 3390.200 34.480 3391.690 ;
        RECT 95.430 3384.980 99.290 3386.420 ;
        RECT 3377.040 3383.240 3382.450 3388.730 ;
        RECT 3358.510 3375.150 3363.920 3380.640 ;
        RECT 3495.950 3367.280 3499.730 3368.690 ;
        RECT 3489.950 3363.760 3493.730 3365.170 ;
        RECT 3489.910 3334.780 3493.770 3336.220 ;
        RECT 3489.890 3317.880 3493.750 3319.320 ;
        RECT 3495.890 3343.230 3499.750 3344.670 ;
        RECT 3495.920 3326.320 3499.780 3327.760 ;
        RECT 3548.730 3348.500 3552.560 3349.850 ;
        RECT 3548.740 3331.580 3552.570 3332.930 ;
        RECT 3548.730 3314.640 3552.600 3316.130 ;
        RECT 3554.740 3340.020 3558.570 3341.370 ;
        RECT 3554.710 3323.220 3558.540 3324.570 ;
        RECT 3495.910 3309.410 3499.770 3310.850 ;
        RECT 3554.700 3306.200 3558.570 3307.690 ;
        RECT 3489.890 3300.980 3493.750 3302.420 ;
        RECT 271.230 3251.240 276.640 3256.730 ;
        RECT 30.580 3208.030 34.440 3209.420 ;
        RECT 30.600 3191.200 34.480 3192.590 ;
        RECT 263.260 3243.150 268.670 3248.640 ;
        RECT 36.590 3216.440 40.460 3217.930 ;
        RECT 36.600 3199.590 40.460 3200.980 ;
        RECT 36.580 3182.640 40.450 3184.130 ;
        RECT 89.450 3235.280 93.230 3236.690 ;
        RECT 89.430 3211.230 93.290 3212.670 ;
        RECT 89.400 3194.320 93.260 3195.760 ;
        RECT 89.410 3177.410 93.270 3178.850 ;
        RECT 95.450 3231.760 99.230 3233.170 ;
        RECT 95.410 3202.780 99.270 3204.220 ;
        RECT 95.430 3185.880 99.290 3187.320 ;
        RECT 30.610 3174.200 34.480 3175.690 ;
        RECT 95.430 3168.980 99.290 3170.420 ;
        RECT 3377.040 3158.240 3382.450 3163.730 ;
        RECT 3358.510 3150.150 3363.920 3155.640 ;
        RECT 3495.950 3142.280 3499.730 3143.690 ;
        RECT 3489.950 3138.760 3493.730 3140.170 ;
        RECT 3489.910 3109.780 3493.770 3111.220 ;
        RECT 3489.890 3092.880 3493.750 3094.320 ;
        RECT 3495.890 3118.230 3499.750 3119.670 ;
        RECT 3495.920 3101.320 3499.780 3102.760 ;
        RECT 3548.730 3123.500 3552.560 3124.850 ;
        RECT 3548.740 3106.580 3552.570 3107.930 ;
        RECT 3548.730 3089.640 3552.600 3091.130 ;
        RECT 3554.740 3115.020 3558.570 3116.370 ;
        RECT 3554.710 3098.220 3558.540 3099.570 ;
        RECT 3495.910 3084.410 3499.770 3085.850 ;
        RECT 3554.700 3081.200 3558.570 3082.690 ;
        RECT 3489.890 3075.980 3493.750 3077.420 ;
        RECT 271.230 3035.240 276.640 3040.730 ;
        RECT 30.580 2992.030 34.440 2993.420 ;
        RECT 30.600 2975.200 34.480 2976.590 ;
        RECT 263.260 3027.150 268.670 3032.640 ;
        RECT 36.590 3000.440 40.460 3001.930 ;
        RECT 36.600 2983.590 40.460 2984.980 ;
        RECT 36.580 2966.640 40.450 2968.130 ;
        RECT 89.450 3019.280 93.230 3020.690 ;
        RECT 89.430 2995.230 93.290 2996.670 ;
        RECT 89.400 2978.320 93.260 2979.760 ;
        RECT 89.410 2961.410 93.270 2962.850 ;
        RECT 95.450 3015.760 99.230 3017.170 ;
        RECT 95.410 2986.780 99.270 2988.220 ;
        RECT 95.430 2969.880 99.290 2971.320 ;
        RECT 30.610 2958.200 34.480 2959.690 ;
        RECT 95.430 2952.980 99.290 2954.420 ;
        RECT 3377.040 2932.240 3382.450 2937.730 ;
        RECT 3358.510 2924.150 3363.920 2929.640 ;
        RECT 3495.950 2916.280 3499.730 2917.690 ;
        RECT 3489.950 2912.760 3493.730 2914.170 ;
        RECT 3489.910 2883.780 3493.770 2885.220 ;
        RECT 3489.890 2866.880 3493.750 2868.320 ;
        RECT 3495.890 2892.230 3499.750 2893.670 ;
        RECT 3495.920 2875.320 3499.780 2876.760 ;
        RECT 3548.730 2897.500 3552.560 2898.850 ;
        RECT 3548.740 2880.580 3552.570 2881.930 ;
        RECT 3548.730 2863.640 3552.600 2865.130 ;
        RECT 3554.740 2889.020 3558.570 2890.370 ;
        RECT 3554.710 2872.220 3558.540 2873.570 ;
        RECT 3495.910 2858.410 3499.770 2859.850 ;
        RECT 3554.700 2855.200 3558.570 2856.690 ;
        RECT 3489.890 2849.980 3493.750 2851.420 ;
        RECT 271.230 2819.240 276.640 2824.730 ;
        RECT 30.580 2776.030 34.440 2777.420 ;
        RECT 30.600 2759.200 34.480 2760.590 ;
        RECT 263.260 2811.150 268.670 2816.640 ;
        RECT 36.590 2784.440 40.460 2785.930 ;
        RECT 36.600 2767.590 40.460 2768.980 ;
        RECT 36.580 2750.640 40.450 2752.130 ;
        RECT 89.450 2803.280 93.230 2804.690 ;
        RECT 89.430 2779.230 93.290 2780.670 ;
        RECT 89.400 2762.320 93.260 2763.760 ;
        RECT 89.410 2745.410 93.270 2746.850 ;
        RECT 95.450 2799.760 99.230 2801.170 ;
        RECT 95.410 2770.780 99.270 2772.220 ;
        RECT 95.430 2753.880 99.290 2755.320 ;
        RECT 30.610 2742.200 34.480 2743.690 ;
        RECT 95.430 2736.980 99.290 2738.420 ;
        RECT 3377.040 2707.240 3382.450 2712.730 ;
        RECT 3358.510 2699.150 3363.920 2704.640 ;
        RECT 3495.950 2691.280 3499.730 2692.690 ;
        RECT 3489.950 2687.760 3493.730 2689.170 ;
        RECT 3489.910 2658.780 3493.770 2660.220 ;
        RECT 3489.890 2641.880 3493.750 2643.320 ;
        RECT 3495.890 2667.230 3499.750 2668.670 ;
        RECT 3495.920 2650.320 3499.780 2651.760 ;
        RECT 3548.730 2672.500 3552.560 2673.850 ;
        RECT 3548.740 2655.580 3552.570 2656.930 ;
        RECT 3548.730 2638.640 3552.600 2640.130 ;
        RECT 3554.740 2664.020 3558.570 2665.370 ;
        RECT 3554.710 2647.220 3558.540 2648.570 ;
        RECT 3495.910 2633.410 3499.770 2634.850 ;
        RECT 3554.700 2630.200 3558.570 2631.690 ;
        RECT 3489.890 2624.980 3493.750 2626.420 ;
        RECT 3336.680 2570.280 3348.530 2592.910 ;
        RECT 3336.750 2520.330 3348.600 2542.960 ;
        RECT 251.820 2466.250 260.460 2488.660 ;
        RECT 3377.040 2487.240 3382.450 2492.730 ;
        RECT 3358.510 2479.150 3363.920 2484.640 ;
        RECT 3495.950 2471.280 3499.730 2472.690 ;
        RECT 3489.950 2467.760 3493.730 2469.170 ;
        RECT 251.760 2416.300 260.400 2438.710 ;
        RECT 3489.910 2438.780 3493.770 2440.220 ;
        RECT 3489.890 2421.880 3493.750 2423.320 ;
        RECT 3495.890 2447.230 3499.750 2448.670 ;
        RECT 3495.920 2430.320 3499.780 2431.760 ;
        RECT 3548.730 2452.500 3552.560 2453.850 ;
        RECT 3548.740 2435.580 3552.570 2436.930 ;
        RECT 3548.730 2418.640 3552.600 2420.130 ;
        RECT 3554.740 2444.020 3558.570 2445.370 ;
        RECT 3554.710 2427.220 3558.540 2428.570 ;
        RECT 3495.910 2413.410 3499.770 2414.850 ;
        RECT 3554.700 2410.200 3558.570 2411.690 ;
        RECT 3489.890 2404.980 3493.750 2406.420 ;
        RECT 271.230 2181.240 276.640 2186.730 ;
        RECT 30.580 2138.030 34.440 2139.420 ;
        RECT 30.600 2121.200 34.480 2122.590 ;
        RECT 263.260 2173.150 268.670 2178.640 ;
        RECT 36.590 2146.440 40.460 2147.930 ;
        RECT 36.600 2129.590 40.460 2130.980 ;
        RECT 36.580 2112.640 40.450 2114.130 ;
        RECT 89.450 2165.280 93.230 2166.690 ;
        RECT 89.430 2141.230 93.290 2142.670 ;
        RECT 89.400 2124.320 93.260 2125.760 ;
        RECT 89.410 2107.410 93.270 2108.850 ;
        RECT 95.450 2161.760 99.230 2163.170 ;
        RECT 95.410 2132.780 99.270 2134.220 ;
        RECT 3320.670 2128.420 3332.700 2151.950 ;
        RECT 95.430 2115.880 99.290 2117.320 ;
        RECT 30.610 2104.200 34.480 2105.690 ;
        RECT 95.430 2098.980 99.290 2100.420 ;
        RECT 3320.560 2079.280 3332.640 2102.310 ;
        RECT 3377.040 2046.240 3382.450 2051.730 ;
        RECT 3358.510 2038.150 3363.920 2043.640 ;
        RECT 3495.950 2030.280 3499.730 2031.690 ;
        RECT 3489.950 2026.760 3493.730 2028.170 ;
        RECT 3489.910 1997.780 3493.770 1999.220 ;
        RECT 3489.890 1980.880 3493.750 1982.320 ;
        RECT 271.230 1965.240 276.640 1970.730 ;
        RECT 3495.890 2006.230 3499.750 2007.670 ;
        RECT 3495.920 1989.320 3499.780 1990.760 ;
        RECT 3548.730 2011.500 3552.560 2012.850 ;
        RECT 3548.740 1994.580 3552.570 1995.930 ;
        RECT 3548.730 1977.640 3552.600 1979.130 ;
        RECT 3554.740 2003.020 3558.570 2004.370 ;
        RECT 3554.710 1986.220 3558.540 1987.570 ;
        RECT 3495.910 1972.410 3499.770 1973.850 ;
        RECT 3554.700 1969.200 3558.570 1970.690 ;
        RECT 3489.890 1963.980 3493.750 1965.420 ;
        RECT 30.580 1922.030 34.440 1923.420 ;
        RECT 30.600 1905.200 34.480 1906.590 ;
        RECT 263.260 1957.150 268.670 1962.640 ;
        RECT 36.590 1930.440 40.460 1931.930 ;
        RECT 36.600 1913.590 40.460 1914.980 ;
        RECT 36.580 1896.640 40.450 1898.130 ;
        RECT 89.450 1949.280 93.230 1950.690 ;
        RECT 89.430 1925.230 93.290 1926.670 ;
        RECT 89.400 1908.320 93.260 1909.760 ;
        RECT 89.410 1891.410 93.270 1892.850 ;
        RECT 95.450 1945.760 99.230 1947.170 ;
        RECT 95.410 1916.780 99.270 1918.220 ;
        RECT 95.430 1899.880 99.290 1901.320 ;
        RECT 30.610 1888.200 34.480 1889.690 ;
        RECT 95.430 1882.980 99.290 1884.420 ;
        RECT 3377.040 1820.240 3382.450 1825.730 ;
        RECT 3358.510 1812.150 3363.920 1817.640 ;
        RECT 3495.950 1804.280 3499.730 1805.690 ;
        RECT 3489.950 1800.760 3493.730 1802.170 ;
        RECT 3489.910 1771.780 3493.770 1773.220 ;
        RECT 271.230 1749.240 276.640 1754.730 ;
        RECT 3489.890 1754.880 3493.750 1756.320 ;
        RECT 30.580 1706.030 34.440 1707.420 ;
        RECT 30.600 1689.200 34.480 1690.590 ;
        RECT 263.260 1741.150 268.670 1746.640 ;
        RECT 3495.890 1780.230 3499.750 1781.670 ;
        RECT 3495.920 1763.320 3499.780 1764.760 ;
        RECT 3548.730 1785.500 3552.560 1786.850 ;
        RECT 3548.740 1768.580 3552.570 1769.930 ;
        RECT 3548.730 1751.640 3552.600 1753.130 ;
        RECT 3554.740 1777.020 3558.570 1778.370 ;
        RECT 3554.710 1760.220 3558.540 1761.570 ;
        RECT 3495.910 1746.410 3499.770 1747.850 ;
        RECT 3554.700 1743.200 3558.570 1744.690 ;
        RECT 36.590 1714.440 40.460 1715.930 ;
        RECT 36.600 1697.590 40.460 1698.980 ;
        RECT 36.580 1680.640 40.450 1682.130 ;
        RECT 89.450 1733.280 93.230 1734.690 ;
        RECT 3489.890 1737.980 3493.750 1739.420 ;
        RECT 89.430 1709.230 93.290 1710.670 ;
        RECT 89.400 1692.320 93.260 1693.760 ;
        RECT 89.410 1675.410 93.270 1676.850 ;
        RECT 95.450 1729.760 99.230 1731.170 ;
        RECT 95.410 1700.780 99.270 1702.220 ;
        RECT 95.430 1683.880 99.290 1685.320 ;
        RECT 30.610 1672.200 34.480 1673.690 ;
        RECT 95.430 1666.980 99.290 1668.420 ;
        RECT 3377.040 1595.240 3382.450 1600.730 ;
        RECT 3358.510 1587.150 3363.920 1592.640 ;
        RECT 3495.950 1579.280 3499.730 1580.690 ;
        RECT 3489.950 1575.760 3493.730 1577.170 ;
        RECT 3489.910 1546.780 3493.770 1548.220 ;
        RECT 271.230 1533.240 276.640 1538.730 ;
        RECT 30.580 1490.030 34.440 1491.420 ;
        RECT 30.600 1473.200 34.480 1474.590 ;
        RECT 263.260 1525.150 268.670 1530.640 ;
        RECT 3489.890 1529.880 3493.750 1531.320 ;
        RECT 36.590 1498.440 40.460 1499.930 ;
        RECT 36.600 1481.590 40.460 1482.980 ;
        RECT 36.580 1464.640 40.450 1466.130 ;
        RECT 89.450 1517.280 93.230 1518.690 ;
        RECT 89.430 1493.230 93.290 1494.670 ;
        RECT 89.400 1476.320 93.260 1477.760 ;
        RECT 89.410 1459.410 93.270 1460.850 ;
        RECT 95.450 1513.760 99.230 1515.170 ;
        RECT 3495.890 1555.230 3499.750 1556.670 ;
        RECT 3495.920 1538.320 3499.780 1539.760 ;
        RECT 3548.730 1560.500 3552.560 1561.850 ;
        RECT 3548.740 1543.580 3552.570 1544.930 ;
        RECT 3548.730 1526.640 3552.600 1528.130 ;
        RECT 3554.740 1552.020 3558.570 1553.370 ;
        RECT 3554.710 1535.220 3558.540 1536.570 ;
        RECT 3495.910 1521.410 3499.770 1522.850 ;
        RECT 3554.700 1518.200 3558.570 1519.690 ;
        RECT 3489.890 1512.980 3493.750 1514.420 ;
        RECT 95.410 1484.780 99.270 1486.220 ;
        RECT 95.430 1467.880 99.290 1469.320 ;
        RECT 30.610 1456.200 34.480 1457.690 ;
        RECT 95.430 1450.980 99.290 1452.420 ;
        RECT 3377.040 1370.240 3382.450 1375.730 ;
        RECT 3358.510 1362.150 3363.920 1367.640 ;
        RECT 3495.950 1354.280 3499.730 1355.690 ;
        RECT 1967.680 1332.780 1970.710 1346.850 ;
        RECT 3489.950 1350.760 3493.730 1352.170 ;
        RECT 271.230 1317.240 276.640 1322.730 ;
        RECT 30.580 1274.030 34.440 1275.420 ;
        RECT 30.600 1257.200 34.480 1258.590 ;
        RECT 263.260 1309.150 268.670 1314.640 ;
        RECT 2042.690 1314.630 2045.960 1326.670 ;
        RECT 3489.910 1321.780 3493.770 1323.220 ;
        RECT 36.590 1282.440 40.460 1283.930 ;
        RECT 36.600 1265.590 40.460 1266.980 ;
        RECT 36.580 1248.640 40.450 1250.130 ;
        RECT 89.450 1301.280 93.230 1302.690 ;
        RECT 89.430 1277.230 93.290 1278.670 ;
        RECT 89.400 1260.320 93.260 1261.760 ;
        RECT 89.410 1243.410 93.270 1244.850 ;
        RECT 95.450 1297.760 99.230 1299.170 ;
        RECT 240.250 1293.380 248.040 1306.690 ;
        RECT 282.770 1293.300 296.760 1306.160 ;
        RECT 1972.950 1292.830 1976.600 1306.680 ;
        RECT 3489.890 1304.880 3493.750 1306.320 ;
        RECT 3495.890 1330.230 3499.750 1331.670 ;
        RECT 3495.920 1313.320 3499.780 1314.760 ;
        RECT 3548.730 1335.500 3552.560 1336.850 ;
        RECT 3548.740 1318.580 3552.570 1319.930 ;
        RECT 3548.730 1301.640 3552.600 1303.130 ;
        RECT 3554.740 1327.020 3558.570 1328.370 ;
        RECT 3554.710 1310.220 3558.540 1311.570 ;
        RECT 3495.910 1296.410 3499.770 1297.850 ;
        RECT 3554.700 1293.200 3558.570 1294.690 ;
        RECT 3489.890 1287.980 3493.750 1289.420 ;
        RECT 252.250 1273.380 260.040 1286.690 ;
        RECT 282.770 1273.300 301.650 1286.160 ;
        RECT 2048.930 1272.790 2053.600 1286.890 ;
        RECT 95.410 1268.780 99.270 1270.220 ;
        RECT 95.430 1251.880 99.290 1253.320 ;
        RECT 263.270 1252.690 268.730 1267.010 ;
        RECT 281.020 1252.740 316.080 1266.980 ;
        RECT 1059.000 1252.860 1062.590 1266.920 ;
        RECT 1209.500 1252.860 1213.090 1266.920 ;
        RECT 1361.160 1252.860 1363.100 1266.920 ;
        RECT 1510.810 1252.860 1513.570 1266.920 ;
        RECT 1661.000 1252.860 1664.590 1266.920 ;
        RECT 1811.500 1252.860 1815.090 1266.920 ;
        RECT 1962.860 1252.860 1965.090 1266.920 ;
        RECT 30.610 1240.200 34.480 1241.690 ;
        RECT 95.430 1234.980 99.290 1236.420 ;
        RECT 983.830 1232.770 987.600 1246.920 ;
        RECT 1134.330 1232.770 1138.100 1246.920 ;
        RECT 1284.830 1232.770 1288.600 1246.920 ;
        RECT 1586.770 1232.770 1589.010 1246.620 ;
        RECT 1736.330 1232.770 1740.100 1246.920 ;
        RECT 1886.330 1232.770 1890.100 1246.920 ;
        RECT 2036.330 1232.770 2040.100 1246.920 ;
        RECT 3335.290 1233.310 3348.210 1246.440 ;
        RECT 3370.780 1233.080 3382.260 1246.480 ;
        RECT 205.330 1191.810 217.650 1226.940 ;
        RECT 281.970 1212.950 316.720 1226.480 ;
        RECT 1063.110 1212.630 1067.320 1227.100 ;
        RECT 1213.610 1212.630 1217.820 1227.100 ;
        RECT 1364.910 1212.630 1366.570 1227.100 ;
        RECT 1515.840 1212.630 1517.300 1227.100 ;
        RECT 1665.110 1212.630 1669.320 1227.100 ;
        RECT 1815.610 1212.630 1819.820 1227.100 ;
        RECT 1966.050 1212.630 1969.000 1227.100 ;
        RECT 221.270 1172.660 233.590 1206.790 ;
        RECT 282.120 1193.120 316.720 1206.650 ;
        RECT 988.160 1192.670 991.610 1207.010 ;
        RECT 1138.660 1192.670 1142.110 1207.010 ;
        RECT 1289.160 1192.670 1292.610 1207.010 ;
        RECT 1440.340 1192.670 1442.830 1207.010 ;
        RECT 1591.130 1192.670 1592.870 1207.010 ;
        RECT 1740.660 1192.670 1744.110 1207.010 ;
        RECT 1890.660 1192.670 1894.110 1207.010 ;
        RECT 2042.050 1192.670 2043.670 1207.010 ;
        RECT 239.900 1172.940 253.390 1186.830 ;
        RECT 282.120 1172.970 315.610 1186.860 ;
        RECT 1054.790 1172.700 1058.610 1186.930 ;
        RECT 1205.290 1172.700 1209.110 1186.930 ;
        RECT 1356.720 1172.700 1359.610 1186.930 ;
        RECT 1507.570 1172.700 1510.110 1186.450 ;
        RECT 1657.070 1172.700 1660.610 1186.930 ;
        RECT 1807.290 1172.700 1811.110 1186.930 ;
        RECT 1959.170 1172.700 1961.110 1186.930 ;
        RECT 282.030 1153.030 315.090 1166.700 ;
        RECT 449.500 1156.990 469.840 1161.290 ;
        RECT 849.320 1156.960 869.660 1161.260 ;
        RECT 980.290 1152.690 982.780 1166.950 ;
        RECT 1130.790 1152.690 1133.280 1166.950 ;
        RECT 1281.290 1152.690 1283.780 1166.950 ;
        RECT 1431.790 1152.690 1434.280 1166.950 ;
        RECT 1582.290 1152.690 1584.780 1166.950 ;
        RECT 1732.790 1152.690 1735.280 1166.950 ;
        RECT 1882.790 1152.690 1885.280 1166.950 ;
        RECT 2033.300 1152.690 2035.280 1166.950 ;
        RECT 2149.550 1157.550 2169.890 1161.850 ;
        RECT 30.580 1058.030 34.440 1059.420 ;
        RECT 30.600 1041.200 34.480 1042.590 ;
        RECT 36.590 1066.440 40.460 1067.930 ;
        RECT 36.600 1049.590 40.460 1050.980 ;
        RECT 36.580 1032.640 40.450 1034.130 ;
        RECT 89.450 1085.280 93.230 1086.690 ;
        RECT 89.430 1061.230 93.290 1062.670 ;
        RECT 89.400 1044.320 93.260 1045.760 ;
        RECT 89.410 1027.410 93.270 1028.850 ;
        RECT 95.450 1081.760 99.230 1083.170 ;
        RECT 95.410 1052.780 99.270 1054.220 ;
        RECT 95.430 1035.880 99.290 1037.320 ;
        RECT 30.610 1024.200 34.480 1025.690 ;
        RECT 95.430 1018.980 99.290 1020.420 ;
        RECT 3377.040 1144.240 3382.450 1149.730 ;
        RECT 3358.510 1136.150 3363.920 1141.640 ;
        RECT 3495.950 1128.280 3499.730 1129.690 ;
        RECT 3489.950 1124.760 3493.730 1126.170 ;
        RECT 271.230 1101.240 276.640 1106.730 ;
        RECT 263.260 1093.150 268.670 1098.640 ;
        RECT 3489.910 1095.780 3493.770 1097.220 ;
        RECT 3489.890 1078.880 3493.750 1080.320 ;
        RECT 3495.890 1104.230 3499.750 1105.670 ;
        RECT 3495.920 1087.320 3499.780 1088.760 ;
        RECT 3548.730 1109.500 3552.560 1110.850 ;
        RECT 3548.740 1092.580 3552.570 1093.930 ;
        RECT 3548.730 1075.640 3552.600 1077.130 ;
        RECT 3554.740 1101.020 3558.570 1102.370 ;
        RECT 3554.710 1084.220 3558.540 1085.570 ;
        RECT 3495.910 1070.410 3499.770 1071.850 ;
        RECT 3554.700 1067.200 3558.570 1068.690 ;
        RECT 2992.990 1048.700 3005.490 1061.630 ;
        RECT 3037.260 1048.700 3049.760 1061.630 ;
        RECT 3205.760 1048.200 3210.050 1061.760 ;
        RECT 3489.890 1061.980 3493.750 1063.420 ;
        RECT 2981.660 1039.630 2988.320 1042.210 ;
        RECT 3012.280 1039.670 3026.630 1042.170 ;
        RECT 257.100 984.670 261.410 987.270 ;
        RECT 2993.420 985.540 3005.190 988.890 ;
        RECT 3030.080 986.190 3034.680 987.460 ;
        RECT 2980.580 919.510 2984.240 922.210 ;
        RECT 3012.280 919.590 3026.630 922.090 ;
        RECT 3377.040 919.240 3382.450 924.730 ;
        RECT 3358.510 911.150 3363.920 916.640 ;
        RECT 3495.950 903.280 3499.730 904.690 ;
        RECT 3489.950 899.760 3493.730 901.170 ;
        RECT 210.010 866.420 228.040 883.050 ;
        RECT 3489.910 870.780 3493.770 872.220 ;
        RECT 214.140 854.540 228.410 857.220 ;
        RECT 256.560 854.600 260.870 857.200 ;
        RECT 3489.890 853.880 3493.750 855.320 ;
        RECT 3495.890 879.230 3499.750 880.670 ;
        RECT 3495.920 862.320 3499.780 863.760 ;
        RECT 3548.730 884.500 3552.560 885.850 ;
        RECT 3548.740 867.580 3552.570 868.930 ;
        RECT 3548.730 850.640 3552.600 852.130 ;
        RECT 3554.740 876.020 3558.570 877.370 ;
        RECT 3554.710 859.220 3558.540 860.570 ;
        RECT 3495.910 845.410 3499.770 846.850 ;
        RECT 3554.700 842.200 3558.570 843.690 ;
        RECT 3489.890 836.980 3493.750 838.420 ;
        RECT 2993.420 832.340 3005.190 835.690 ;
        RECT 3029.930 833.040 3034.660 834.330 ;
        RECT 2970.570 789.530 2984.230 792.230 ;
        RECT 3012.150 789.650 3026.500 792.150 ;
        RECT 214.210 724.570 228.480 727.250 ;
        RECT 256.230 724.560 260.540 727.160 ;
        RECT 3377.040 693.240 3382.450 698.730 ;
        RECT 3358.510 685.150 3363.920 690.640 ;
        RECT 2993.420 679.140 3005.190 682.490 ;
        RECT 3029.860 679.820 3034.630 681.150 ;
        RECT 3495.950 677.280 3499.730 678.690 ;
        RECT 3489.950 673.760 3493.730 675.170 ;
        RECT 2970.620 659.500 2984.280 662.200 ;
        RECT 3012.280 659.570 3026.630 662.070 ;
        RECT 3489.910 644.780 3493.770 646.220 ;
        RECT 3489.890 627.880 3493.750 629.320 ;
        RECT 3495.890 653.230 3499.750 654.670 ;
        RECT 3495.920 636.320 3499.780 637.760 ;
        RECT 3548.730 658.500 3552.560 659.850 ;
        RECT 3548.740 641.580 3552.570 642.930 ;
        RECT 3548.730 624.640 3552.600 626.130 ;
        RECT 3554.740 650.020 3558.570 651.370 ;
        RECT 3554.710 633.220 3558.540 634.570 ;
        RECT 3495.910 619.410 3499.770 620.850 ;
        RECT 3554.700 616.200 3558.570 617.690 ;
        RECT 3489.890 610.980 3493.750 612.420 ;
        RECT 214.160 594.550 228.430 597.230 ;
        RECT 256.210 594.590 260.520 597.190 ;
        RECT 2970.630 529.530 2984.290 532.230 ;
        RECT 3012.300 529.630 3026.650 532.130 ;
        RECT 2993.420 524.540 3005.190 527.890 ;
        RECT 3029.900 526.630 3034.710 527.970 ;
        RECT 3127.780 480.370 3133.720 493.280 ;
        RECT 3181.080 482.920 3184.290 493.110 ;
        RECT 3282.110 480.710 3287.500 493.560 ;
        RECT 214.140 464.540 228.410 467.220 ;
        RECT 256.230 464.570 260.540 467.170 ;
        RECT 209.730 391.210 228.360 413.530 ;
        RECT 2970.600 399.580 2984.260 402.280 ;
        RECT 3012.270 399.690 3026.620 402.190 ;
        RECT 3161.000 391.630 3164.320 403.880 ;
        RECT 3201.050 391.280 3204.050 404.500 ;
        RECT 3124.030 383.130 3125.340 387.660 ;
        RECT 3131.790 376.120 3133.100 380.650 ;
        RECT 3139.590 383.200 3140.900 387.730 ;
        RECT 3147.260 376.140 3148.570 380.670 ;
        RECT 3155.040 383.180 3156.350 387.710 ;
        RECT 3162.800 376.160 3164.110 380.690 ;
        RECT 3170.510 383.180 3171.820 387.710 ;
        RECT 3178.320 376.120 3179.630 380.650 ;
        RECT 3186.050 383.240 3187.360 387.770 ;
        RECT 3193.830 376.250 3195.140 380.780 ;
        RECT 209.610 341.690 228.240 364.010 ;
        RECT 209.680 334.510 228.450 337.190 ;
        RECT 257.220 334.580 261.530 337.180 ;
        RECT 210.030 242.020 227.950 259.940 ;
        RECT 272.630 241.850 291.050 259.770 ;
        RECT 716.950 250.020 723.260 253.120 ;
        RECT 707.210 221.030 714.050 226.530 ;
        RECT 1208.700 214.210 1229.930 233.080 ;
        RECT 1256.960 214.280 1278.190 233.150 ;
        RECT 3240.830 233.300 3248.040 235.620 ;
        RECT 3332.300 235.150 3346.900 236.410 ;
      LAYER met5 ;
        RECT 2878.200 4973.980 3333.100 4986.980 ;
        RECT 89.230 4100.780 93.425 4100.895 ;
        RECT 71.550 4099.180 93.425 4100.780 ;
        RECT 89.230 4099.090 93.425 4099.180 ;
        RECT 95.260 4097.280 99.455 4097.350 ;
        RECT 71.550 4095.680 99.610 4097.280 ;
        RECT 95.260 4095.545 99.455 4095.680 ;
        RECT 36.395 4081.990 40.590 4082.095 ;
        RECT 36.300 4080.390 42.910 4081.990 ;
        RECT 36.395 4080.290 40.590 4080.390 ;
        RECT 89.245 4076.750 93.455 4076.840 ;
        RECT 87.120 4075.150 93.540 4076.750 ;
        RECT 89.245 4075.040 93.455 4075.150 ;
        RECT 30.440 4073.540 34.635 4073.700 ;
        RECT 30.240 4071.940 42.910 4073.540 ;
        RECT 30.440 4071.895 34.635 4071.940 ;
        RECT 95.280 4068.300 99.490 4068.365 ;
        RECT 87.120 4066.700 99.500 4068.300 ;
        RECT 95.280 4066.620 99.490 4066.700 ;
        RECT 36.485 4065.090 40.680 4065.205 ;
        RECT 36.330 4063.490 42.910 4065.090 ;
        RECT 36.485 4063.400 40.680 4063.490 ;
        RECT 89.285 4059.850 93.495 4059.890 ;
        RECT 87.120 4058.250 93.495 4059.850 ;
        RECT 89.285 4058.145 93.495 4058.250 ;
        RECT 30.170 4056.640 34.645 4056.770 ;
        RECT 30.170 4055.040 42.910 4056.640 ;
        RECT 30.170 4055.030 34.645 4055.040 ;
        RECT 95.265 4051.400 99.475 4051.475 ;
        RECT 87.120 4049.800 99.500 4051.400 ;
        RECT 95.265 4049.730 99.475 4049.800 ;
        RECT 36.385 4048.190 40.860 4048.265 ;
        RECT 36.385 4046.590 43.070 4048.190 ;
        RECT 36.385 4046.510 40.860 4046.590 ;
        RECT 89.265 4042.950 93.475 4043.025 ;
        RECT 87.120 4041.350 93.510 4042.950 ;
        RECT 89.265 4041.280 93.475 4041.350 ;
        RECT 30.425 4039.740 34.900 4039.850 ;
        RECT 30.425 4038.140 43.070 4039.740 ;
        RECT 30.425 4038.040 34.900 4038.140 ;
        RECT 95.310 4034.500 99.520 4034.575 ;
        RECT 87.120 4032.900 99.520 4034.500 ;
        RECT 95.310 4032.830 99.520 4032.900 ;
        RECT 89.230 3884.780 93.425 3884.895 ;
        RECT 71.550 3883.180 93.425 3884.780 ;
        RECT 89.230 3883.090 93.425 3883.180 ;
        RECT 95.260 3881.280 99.455 3881.350 ;
        RECT 71.550 3879.680 99.610 3881.280 ;
        RECT 95.260 3879.545 99.455 3879.680 ;
        RECT 36.395 3865.990 40.590 3866.095 ;
        RECT 36.300 3864.390 42.910 3865.990 ;
        RECT 36.395 3864.290 40.590 3864.390 ;
        RECT 89.245 3860.750 93.455 3860.840 ;
        RECT 87.120 3859.150 93.540 3860.750 ;
        RECT 89.245 3859.040 93.455 3859.150 ;
        RECT 30.440 3857.540 34.635 3857.700 ;
        RECT 30.240 3855.940 42.910 3857.540 ;
        RECT 30.440 3855.895 34.635 3855.940 ;
        RECT 95.280 3852.300 99.490 3852.365 ;
        RECT 87.120 3850.700 99.500 3852.300 ;
        RECT 95.280 3850.620 99.490 3850.700 ;
        RECT 36.485 3849.090 40.680 3849.205 ;
        RECT 36.330 3847.490 42.910 3849.090 ;
        RECT 36.485 3847.400 40.680 3847.490 ;
        RECT 89.285 3843.850 93.495 3843.890 ;
        RECT 87.120 3842.250 93.495 3843.850 ;
        RECT 89.285 3842.145 93.495 3842.250 ;
        RECT 30.170 3840.640 34.645 3840.770 ;
        RECT 30.170 3839.040 42.910 3840.640 ;
        RECT 30.170 3839.030 34.645 3839.040 ;
        RECT 95.265 3835.400 99.475 3835.475 ;
        RECT 87.120 3833.800 99.500 3835.400 ;
        RECT 95.265 3833.730 99.475 3833.800 ;
        RECT 36.385 3832.190 40.860 3832.265 ;
        RECT 36.385 3830.590 43.070 3832.190 ;
        RECT 36.385 3830.510 40.860 3830.590 ;
        RECT 89.265 3826.950 93.475 3827.025 ;
        RECT 87.120 3825.350 93.510 3826.950 ;
        RECT 89.265 3825.280 93.475 3825.350 ;
        RECT 30.425 3823.740 34.900 3823.850 ;
        RECT 30.425 3822.140 43.070 3823.740 ;
        RECT 30.425 3822.040 34.900 3822.140 ;
        RECT 95.310 3818.500 99.520 3818.575 ;
        RECT 87.120 3816.900 99.520 3818.500 ;
        RECT 95.310 3816.830 99.520 3816.900 ;
        RECT 89.230 3668.780 93.425 3668.895 ;
        RECT 71.550 3667.180 93.425 3668.780 ;
        RECT 89.230 3667.090 93.425 3667.180 ;
        RECT 95.260 3665.280 99.455 3665.350 ;
        RECT 71.550 3663.680 99.610 3665.280 ;
        RECT 95.260 3663.545 99.455 3663.680 ;
        RECT 36.395 3649.990 40.590 3650.095 ;
        RECT 36.300 3648.390 42.910 3649.990 ;
        RECT 36.395 3648.290 40.590 3648.390 ;
        RECT 89.245 3644.750 93.455 3644.840 ;
        RECT 87.120 3643.150 93.540 3644.750 ;
        RECT 89.245 3643.040 93.455 3643.150 ;
        RECT 30.440 3641.540 34.635 3641.700 ;
        RECT 30.240 3639.940 42.910 3641.540 ;
        RECT 30.440 3639.895 34.635 3639.940 ;
        RECT 95.280 3636.300 99.490 3636.365 ;
        RECT 87.120 3634.700 99.500 3636.300 ;
        RECT 95.280 3634.620 99.490 3634.700 ;
        RECT 36.485 3633.090 40.680 3633.205 ;
        RECT 36.330 3631.490 42.910 3633.090 ;
        RECT 36.485 3631.400 40.680 3631.490 ;
        RECT 89.285 3627.850 93.495 3627.890 ;
        RECT 87.120 3626.250 93.495 3627.850 ;
        RECT 89.285 3626.145 93.495 3626.250 ;
        RECT 30.170 3624.640 34.645 3624.770 ;
        RECT 30.170 3623.040 42.910 3624.640 ;
        RECT 30.170 3623.030 34.645 3623.040 ;
        RECT 95.265 3619.400 99.475 3619.475 ;
        RECT 87.120 3617.800 99.500 3619.400 ;
        RECT 95.265 3617.730 99.475 3617.800 ;
        RECT 36.385 3616.190 40.860 3616.265 ;
        RECT 36.385 3614.590 43.070 3616.190 ;
        RECT 36.385 3614.510 40.860 3614.590 ;
        RECT 89.265 3610.950 93.475 3611.025 ;
        RECT 87.120 3609.350 93.510 3610.950 ;
        RECT 89.265 3609.280 93.475 3609.350 ;
        RECT 30.425 3607.740 34.900 3607.850 ;
        RECT 30.425 3606.140 43.070 3607.740 ;
        RECT 30.425 3606.040 34.900 3606.140 ;
        RECT 95.310 3602.500 99.520 3602.575 ;
        RECT 87.120 3600.900 99.520 3602.500 ;
        RECT 95.310 3600.830 99.520 3600.900 ;
        RECT 89.230 3452.780 93.425 3452.895 ;
        RECT 71.550 3451.180 93.425 3452.780 ;
        RECT 89.230 3451.090 93.425 3451.180 ;
        RECT 95.260 3449.280 99.455 3449.350 ;
        RECT 71.550 3447.680 99.610 3449.280 ;
        RECT 95.260 3447.545 99.455 3447.680 ;
        RECT 36.395 3433.990 40.590 3434.095 ;
        RECT 36.300 3432.390 42.910 3433.990 ;
        RECT 36.395 3432.290 40.590 3432.390 ;
        RECT 89.245 3428.750 93.455 3428.840 ;
        RECT 87.120 3427.150 93.540 3428.750 ;
        RECT 89.245 3427.040 93.455 3427.150 ;
        RECT 30.440 3425.540 34.635 3425.700 ;
        RECT 30.240 3423.940 42.910 3425.540 ;
        RECT 30.440 3423.895 34.635 3423.940 ;
        RECT 95.280 3420.300 99.490 3420.365 ;
        RECT 87.120 3418.700 99.500 3420.300 ;
        RECT 95.280 3418.620 99.490 3418.700 ;
        RECT 36.485 3417.090 40.680 3417.205 ;
        RECT 36.330 3415.490 42.910 3417.090 ;
        RECT 36.485 3415.400 40.680 3415.490 ;
        RECT 89.285 3411.850 93.495 3411.890 ;
        RECT 87.120 3410.250 93.495 3411.850 ;
        RECT 89.285 3410.145 93.495 3410.250 ;
        RECT 30.170 3408.640 34.645 3408.770 ;
        RECT 30.170 3407.040 42.910 3408.640 ;
        RECT 30.170 3407.030 34.645 3407.040 ;
        RECT 95.265 3403.400 99.475 3403.475 ;
        RECT 87.120 3401.800 99.500 3403.400 ;
        RECT 95.265 3401.730 99.475 3401.800 ;
        RECT 36.385 3400.190 40.860 3400.265 ;
        RECT 36.385 3398.590 43.070 3400.190 ;
        RECT 36.385 3398.510 40.860 3398.590 ;
        RECT 89.265 3394.950 93.475 3395.025 ;
        RECT 87.120 3393.350 93.510 3394.950 ;
        RECT 89.265 3393.280 93.475 3393.350 ;
        RECT 30.425 3391.740 34.900 3391.850 ;
        RECT 30.425 3390.140 43.070 3391.740 ;
        RECT 30.425 3390.040 34.900 3390.140 ;
        RECT 95.310 3386.500 99.520 3386.575 ;
        RECT 87.120 3384.900 99.520 3386.500 ;
        RECT 95.310 3384.830 99.520 3384.900 ;
        RECT 89.230 3236.780 93.425 3236.895 ;
        RECT 71.550 3235.180 93.425 3236.780 ;
        RECT 89.230 3235.090 93.425 3235.180 ;
        RECT 95.260 3233.280 99.455 3233.350 ;
        RECT 71.550 3231.680 99.610 3233.280 ;
        RECT 95.260 3231.545 99.455 3231.680 ;
        RECT 36.395 3217.990 40.590 3218.095 ;
        RECT 36.300 3216.390 42.910 3217.990 ;
        RECT 36.395 3216.290 40.590 3216.390 ;
        RECT 89.245 3212.750 93.455 3212.840 ;
        RECT 87.120 3211.150 93.540 3212.750 ;
        RECT 89.245 3211.040 93.455 3211.150 ;
        RECT 30.440 3209.540 34.635 3209.700 ;
        RECT 30.240 3207.940 42.910 3209.540 ;
        RECT 30.440 3207.895 34.635 3207.940 ;
        RECT 95.280 3204.300 99.490 3204.365 ;
        RECT 87.120 3202.700 99.500 3204.300 ;
        RECT 95.280 3202.620 99.490 3202.700 ;
        RECT 36.485 3201.090 40.680 3201.205 ;
        RECT 36.330 3199.490 42.910 3201.090 ;
        RECT 36.485 3199.400 40.680 3199.490 ;
        RECT 89.285 3195.850 93.495 3195.890 ;
        RECT 87.120 3194.250 93.495 3195.850 ;
        RECT 89.285 3194.145 93.495 3194.250 ;
        RECT 30.170 3192.640 34.645 3192.770 ;
        RECT 30.170 3191.040 42.910 3192.640 ;
        RECT 30.170 3191.030 34.645 3191.040 ;
        RECT 95.265 3187.400 99.475 3187.475 ;
        RECT 87.120 3185.800 99.500 3187.400 ;
        RECT 95.265 3185.730 99.475 3185.800 ;
        RECT 36.385 3184.190 40.860 3184.265 ;
        RECT 36.385 3182.590 43.070 3184.190 ;
        RECT 36.385 3182.510 40.860 3182.590 ;
        RECT 89.265 3178.950 93.475 3179.025 ;
        RECT 87.120 3177.350 93.510 3178.950 ;
        RECT 89.265 3177.280 93.475 3177.350 ;
        RECT 30.425 3175.740 34.900 3175.850 ;
        RECT 30.425 3174.140 43.070 3175.740 ;
        RECT 30.425 3174.040 34.900 3174.140 ;
        RECT 95.310 3170.500 99.520 3170.575 ;
        RECT 87.120 3168.900 99.520 3170.500 ;
        RECT 95.310 3168.830 99.520 3168.900 ;
        RECT 89.230 3020.780 93.425 3020.895 ;
        RECT 71.550 3019.180 93.425 3020.780 ;
        RECT 89.230 3019.090 93.425 3019.180 ;
        RECT 95.260 3017.280 99.455 3017.350 ;
        RECT 71.550 3015.680 99.610 3017.280 ;
        RECT 95.260 3015.545 99.455 3015.680 ;
        RECT 36.395 3001.990 40.590 3002.095 ;
        RECT 36.300 3000.390 42.910 3001.990 ;
        RECT 36.395 3000.290 40.590 3000.390 ;
        RECT 89.245 2996.750 93.455 2996.840 ;
        RECT 87.120 2995.150 93.540 2996.750 ;
        RECT 89.245 2995.040 93.455 2995.150 ;
        RECT 30.440 2993.540 34.635 2993.700 ;
        RECT 30.240 2991.940 42.910 2993.540 ;
        RECT 30.440 2991.895 34.635 2991.940 ;
        RECT 95.280 2988.300 99.490 2988.365 ;
        RECT 87.120 2986.700 99.500 2988.300 ;
        RECT 95.280 2986.620 99.490 2986.700 ;
        RECT 36.485 2985.090 40.680 2985.205 ;
        RECT 36.330 2983.490 42.910 2985.090 ;
        RECT 36.485 2983.400 40.680 2983.490 ;
        RECT 89.285 2979.850 93.495 2979.890 ;
        RECT 87.120 2978.250 93.495 2979.850 ;
        RECT 89.285 2978.145 93.495 2978.250 ;
        RECT 30.170 2976.640 34.645 2976.770 ;
        RECT 30.170 2975.040 42.910 2976.640 ;
        RECT 30.170 2975.030 34.645 2975.040 ;
        RECT 95.265 2971.400 99.475 2971.475 ;
        RECT 87.120 2969.800 99.500 2971.400 ;
        RECT 95.265 2969.730 99.475 2969.800 ;
        RECT 36.385 2968.190 40.860 2968.265 ;
        RECT 36.385 2966.590 43.070 2968.190 ;
        RECT 36.385 2966.510 40.860 2966.590 ;
        RECT 89.265 2962.950 93.475 2963.025 ;
        RECT 87.120 2961.350 93.510 2962.950 ;
        RECT 89.265 2961.280 93.475 2961.350 ;
        RECT 30.425 2959.740 34.900 2959.850 ;
        RECT 30.425 2958.140 43.070 2959.740 ;
        RECT 30.425 2958.040 34.900 2958.140 ;
        RECT 95.310 2954.500 99.520 2954.575 ;
        RECT 87.120 2952.900 99.520 2954.500 ;
        RECT 95.310 2952.830 99.520 2952.900 ;
        RECT 89.230 2804.780 93.425 2804.895 ;
        RECT 71.550 2803.180 93.425 2804.780 ;
        RECT 89.230 2803.090 93.425 2803.180 ;
        RECT 95.260 2801.280 99.455 2801.350 ;
        RECT 71.550 2799.680 99.610 2801.280 ;
        RECT 95.260 2799.545 99.455 2799.680 ;
        RECT 36.395 2785.990 40.590 2786.095 ;
        RECT 36.300 2784.390 42.910 2785.990 ;
        RECT 36.395 2784.290 40.590 2784.390 ;
        RECT 89.245 2780.750 93.455 2780.840 ;
        RECT 87.120 2779.150 93.540 2780.750 ;
        RECT 89.245 2779.040 93.455 2779.150 ;
        RECT 30.440 2777.540 34.635 2777.700 ;
        RECT 30.240 2775.940 42.910 2777.540 ;
        RECT 30.440 2775.895 34.635 2775.940 ;
        RECT 95.280 2772.300 99.490 2772.365 ;
        RECT 87.120 2770.700 99.500 2772.300 ;
        RECT 95.280 2770.620 99.490 2770.700 ;
        RECT 36.485 2769.090 40.680 2769.205 ;
        RECT 36.330 2767.490 42.910 2769.090 ;
        RECT 36.485 2767.400 40.680 2767.490 ;
        RECT 89.285 2763.850 93.495 2763.890 ;
        RECT 87.120 2762.250 93.495 2763.850 ;
        RECT 89.285 2762.145 93.495 2762.250 ;
        RECT 30.170 2760.640 34.645 2760.770 ;
        RECT 30.170 2759.040 42.910 2760.640 ;
        RECT 30.170 2759.030 34.645 2759.040 ;
        RECT 95.265 2755.400 99.475 2755.475 ;
        RECT 87.120 2753.800 99.500 2755.400 ;
        RECT 95.265 2753.730 99.475 2753.800 ;
        RECT 36.385 2752.190 40.860 2752.265 ;
        RECT 36.385 2750.590 43.070 2752.190 ;
        RECT 36.385 2750.510 40.860 2750.590 ;
        RECT 89.265 2746.950 93.475 2747.025 ;
        RECT 87.120 2745.350 93.510 2746.950 ;
        RECT 89.265 2745.280 93.475 2745.350 ;
        RECT 30.425 2743.740 34.900 2743.850 ;
        RECT 30.425 2742.140 43.070 2743.740 ;
        RECT 30.425 2742.040 34.900 2742.140 ;
        RECT 95.310 2738.500 99.520 2738.575 ;
        RECT 87.120 2736.900 99.520 2738.500 ;
        RECT 95.310 2736.830 99.520 2736.900 ;
        RECT 89.230 2166.780 93.425 2166.895 ;
        RECT 71.550 2165.180 93.425 2166.780 ;
        RECT 89.230 2165.090 93.425 2165.180 ;
        RECT 95.260 2163.280 99.455 2163.350 ;
        RECT 71.550 2161.680 99.610 2163.280 ;
        RECT 95.260 2161.545 99.455 2161.680 ;
        RECT 36.395 2147.990 40.590 2148.095 ;
        RECT 36.300 2146.390 42.910 2147.990 ;
        RECT 36.395 2146.290 40.590 2146.390 ;
        RECT 89.245 2142.750 93.455 2142.840 ;
        RECT 87.120 2141.150 93.540 2142.750 ;
        RECT 89.245 2141.040 93.455 2141.150 ;
        RECT 30.440 2139.540 34.635 2139.700 ;
        RECT 30.240 2137.940 42.910 2139.540 ;
        RECT 30.440 2137.895 34.635 2137.940 ;
        RECT 95.280 2134.300 99.490 2134.365 ;
        RECT 87.120 2132.700 99.500 2134.300 ;
        RECT 95.280 2132.620 99.490 2132.700 ;
        RECT 36.485 2131.090 40.680 2131.205 ;
        RECT 36.330 2129.490 42.910 2131.090 ;
        RECT 36.485 2129.400 40.680 2129.490 ;
        RECT 89.285 2125.850 93.495 2125.890 ;
        RECT 87.120 2124.250 93.495 2125.850 ;
        RECT 89.285 2124.145 93.495 2124.250 ;
        RECT 30.170 2122.640 34.645 2122.770 ;
        RECT 30.170 2121.040 42.910 2122.640 ;
        RECT 30.170 2121.030 34.645 2121.040 ;
        RECT 95.265 2117.400 99.475 2117.475 ;
        RECT 87.120 2115.800 99.500 2117.400 ;
        RECT 95.265 2115.730 99.475 2115.800 ;
        RECT 36.385 2114.190 40.860 2114.265 ;
        RECT 36.385 2112.590 43.070 2114.190 ;
        RECT 36.385 2112.510 40.860 2112.590 ;
        RECT 89.265 2108.950 93.475 2109.025 ;
        RECT 87.120 2107.350 93.510 2108.950 ;
        RECT 89.265 2107.280 93.475 2107.350 ;
        RECT 30.425 2105.740 34.900 2105.850 ;
        RECT 30.425 2104.140 43.070 2105.740 ;
        RECT 30.425 2104.040 34.900 2104.140 ;
        RECT 95.310 2100.500 99.520 2100.575 ;
        RECT 87.120 2098.900 99.520 2100.500 ;
        RECT 95.310 2098.830 99.520 2098.900 ;
        RECT 89.230 1950.780 93.425 1950.895 ;
        RECT 71.550 1949.180 93.425 1950.780 ;
        RECT 89.230 1949.090 93.425 1949.180 ;
        RECT 95.260 1947.280 99.455 1947.350 ;
        RECT 71.550 1945.680 99.610 1947.280 ;
        RECT 95.260 1945.545 99.455 1945.680 ;
        RECT 36.395 1931.990 40.590 1932.095 ;
        RECT 36.300 1930.390 42.910 1931.990 ;
        RECT 36.395 1930.290 40.590 1930.390 ;
        RECT 89.245 1926.750 93.455 1926.840 ;
        RECT 87.120 1925.150 93.540 1926.750 ;
        RECT 89.245 1925.040 93.455 1925.150 ;
        RECT 30.440 1923.540 34.635 1923.700 ;
        RECT 30.240 1921.940 42.910 1923.540 ;
        RECT 30.440 1921.895 34.635 1921.940 ;
        RECT 95.280 1918.300 99.490 1918.365 ;
        RECT 87.120 1916.700 99.500 1918.300 ;
        RECT 95.280 1916.620 99.490 1916.700 ;
        RECT 36.485 1915.090 40.680 1915.205 ;
        RECT 36.330 1913.490 42.910 1915.090 ;
        RECT 36.485 1913.400 40.680 1913.490 ;
        RECT 89.285 1909.850 93.495 1909.890 ;
        RECT 87.120 1908.250 93.495 1909.850 ;
        RECT 89.285 1908.145 93.495 1908.250 ;
        RECT 30.170 1906.640 34.645 1906.770 ;
        RECT 30.170 1905.040 42.910 1906.640 ;
        RECT 30.170 1905.030 34.645 1905.040 ;
        RECT 95.265 1901.400 99.475 1901.475 ;
        RECT 87.120 1899.800 99.500 1901.400 ;
        RECT 95.265 1899.730 99.475 1899.800 ;
        RECT 36.385 1898.190 40.860 1898.265 ;
        RECT 36.385 1896.590 43.070 1898.190 ;
        RECT 36.385 1896.510 40.860 1896.590 ;
        RECT 89.265 1892.950 93.475 1893.025 ;
        RECT 87.120 1891.350 93.510 1892.950 ;
        RECT 89.265 1891.280 93.475 1891.350 ;
        RECT 30.425 1889.740 34.900 1889.850 ;
        RECT 30.425 1888.140 43.070 1889.740 ;
        RECT 30.425 1888.040 34.900 1888.140 ;
        RECT 95.310 1884.500 99.520 1884.575 ;
        RECT 87.120 1882.900 99.520 1884.500 ;
        RECT 95.310 1882.830 99.520 1882.900 ;
        RECT 89.230 1734.780 93.425 1734.895 ;
        RECT 71.550 1733.180 93.425 1734.780 ;
        RECT 89.230 1733.090 93.425 1733.180 ;
        RECT 95.260 1731.280 99.455 1731.350 ;
        RECT 71.550 1729.680 99.610 1731.280 ;
        RECT 95.260 1729.545 99.455 1729.680 ;
        RECT 36.395 1715.990 40.590 1716.095 ;
        RECT 36.300 1714.390 42.910 1715.990 ;
        RECT 36.395 1714.290 40.590 1714.390 ;
        RECT 89.245 1710.750 93.455 1710.840 ;
        RECT 87.120 1709.150 93.540 1710.750 ;
        RECT 89.245 1709.040 93.455 1709.150 ;
        RECT 30.440 1707.540 34.635 1707.700 ;
        RECT 30.240 1705.940 42.910 1707.540 ;
        RECT 30.440 1705.895 34.635 1705.940 ;
        RECT 95.280 1702.300 99.490 1702.365 ;
        RECT 87.120 1700.700 99.500 1702.300 ;
        RECT 95.280 1700.620 99.490 1700.700 ;
        RECT 36.485 1699.090 40.680 1699.205 ;
        RECT 36.330 1697.490 42.910 1699.090 ;
        RECT 36.485 1697.400 40.680 1697.490 ;
        RECT 89.285 1693.850 93.495 1693.890 ;
        RECT 87.120 1692.250 93.495 1693.850 ;
        RECT 89.285 1692.145 93.495 1692.250 ;
        RECT 30.170 1690.640 34.645 1690.770 ;
        RECT 30.170 1689.040 42.910 1690.640 ;
        RECT 30.170 1689.030 34.645 1689.040 ;
        RECT 95.265 1685.400 99.475 1685.475 ;
        RECT 87.120 1683.800 99.500 1685.400 ;
        RECT 95.265 1683.730 99.475 1683.800 ;
        RECT 36.385 1682.190 40.860 1682.265 ;
        RECT 36.385 1680.590 43.070 1682.190 ;
        RECT 36.385 1680.510 40.860 1680.590 ;
        RECT 89.265 1676.950 93.475 1677.025 ;
        RECT 87.120 1675.350 93.510 1676.950 ;
        RECT 89.265 1675.280 93.475 1675.350 ;
        RECT 30.425 1673.740 34.900 1673.850 ;
        RECT 30.425 1672.140 43.070 1673.740 ;
        RECT 30.425 1672.040 34.900 1672.140 ;
        RECT 95.310 1668.500 99.520 1668.575 ;
        RECT 87.120 1666.900 99.520 1668.500 ;
        RECT 95.310 1666.830 99.520 1666.900 ;
        RECT 89.230 1518.780 93.425 1518.895 ;
        RECT 71.550 1517.180 93.425 1518.780 ;
        RECT 89.230 1517.090 93.425 1517.180 ;
        RECT 95.260 1515.280 99.455 1515.350 ;
        RECT 71.550 1513.680 99.610 1515.280 ;
        RECT 95.260 1513.545 99.455 1513.680 ;
        RECT 36.395 1499.990 40.590 1500.095 ;
        RECT 36.300 1498.390 42.910 1499.990 ;
        RECT 36.395 1498.290 40.590 1498.390 ;
        RECT 89.245 1494.750 93.455 1494.840 ;
        RECT 87.120 1493.150 93.540 1494.750 ;
        RECT 89.245 1493.040 93.455 1493.150 ;
        RECT 30.440 1491.540 34.635 1491.700 ;
        RECT 30.240 1489.940 42.910 1491.540 ;
        RECT 30.440 1489.895 34.635 1489.940 ;
        RECT 95.280 1486.300 99.490 1486.365 ;
        RECT 87.120 1484.700 99.500 1486.300 ;
        RECT 95.280 1484.620 99.490 1484.700 ;
        RECT 36.485 1483.090 40.680 1483.205 ;
        RECT 36.330 1481.490 42.910 1483.090 ;
        RECT 36.485 1481.400 40.680 1481.490 ;
        RECT 89.285 1477.850 93.495 1477.890 ;
        RECT 87.120 1476.250 93.495 1477.850 ;
        RECT 89.285 1476.145 93.495 1476.250 ;
        RECT 30.170 1474.640 34.645 1474.770 ;
        RECT 30.170 1473.040 42.910 1474.640 ;
        RECT 30.170 1473.030 34.645 1473.040 ;
        RECT 95.265 1469.400 99.475 1469.475 ;
        RECT 87.120 1467.800 99.500 1469.400 ;
        RECT 95.265 1467.730 99.475 1467.800 ;
        RECT 36.385 1466.190 40.860 1466.265 ;
        RECT 36.385 1464.590 43.070 1466.190 ;
        RECT 36.385 1464.510 40.860 1464.590 ;
        RECT 89.265 1460.950 93.475 1461.025 ;
        RECT 87.120 1459.350 93.510 1460.950 ;
        RECT 89.265 1459.280 93.475 1459.350 ;
        RECT 30.425 1457.740 34.900 1457.850 ;
        RECT 30.425 1456.140 43.070 1457.740 ;
        RECT 30.425 1456.040 34.900 1456.140 ;
        RECT 95.310 1452.500 99.520 1452.575 ;
        RECT 87.120 1450.900 99.520 1452.500 ;
        RECT 95.310 1450.830 99.520 1450.900 ;
        RECT 89.230 1302.780 93.425 1302.895 ;
        RECT 71.550 1301.180 93.425 1302.780 ;
        RECT 89.230 1301.090 93.425 1301.180 ;
        RECT 95.260 1299.280 99.455 1299.350 ;
        RECT 71.550 1297.680 99.610 1299.280 ;
        RECT 95.260 1297.545 99.455 1297.680 ;
        RECT 238.990 1292.420 248.990 4212.800 ;
        RECT 36.395 1283.990 40.590 1284.095 ;
        RECT 36.300 1282.390 42.910 1283.990 ;
        RECT 36.395 1282.290 40.590 1282.390 ;
        RECT 89.245 1278.750 93.455 1278.840 ;
        RECT 87.120 1277.150 93.540 1278.750 ;
        RECT 89.245 1277.040 93.455 1277.150 ;
        RECT 30.440 1275.540 34.635 1275.700 ;
        RECT 30.240 1273.940 42.910 1275.540 ;
        RECT 30.440 1273.895 34.635 1273.940 ;
        RECT 250.990 1272.490 260.990 2489.960 ;
        RECT 95.280 1270.300 99.490 1270.365 ;
        RECT 87.120 1268.700 99.500 1270.300 ;
        RECT 95.280 1268.620 99.490 1268.700 ;
        RECT 36.485 1267.090 40.680 1267.205 ;
        RECT 36.330 1265.490 42.910 1267.090 ;
        RECT 36.485 1265.400 40.680 1265.490 ;
        RECT 89.285 1261.850 93.495 1261.890 ;
        RECT 87.120 1260.250 93.495 1261.850 ;
        RECT 89.285 1260.145 93.495 1260.250 ;
        RECT 30.170 1258.640 34.645 1258.770 ;
        RECT 30.170 1257.040 42.910 1258.640 ;
        RECT 30.170 1257.030 34.645 1257.040 ;
        RECT 95.265 1253.400 99.475 1253.475 ;
        RECT 87.120 1251.800 99.500 1253.400 ;
        RECT 95.265 1251.730 99.475 1251.800 ;
        RECT 36.385 1250.190 40.860 1250.265 ;
        RECT 36.385 1248.590 43.070 1250.190 ;
        RECT 36.385 1248.510 40.860 1248.590 ;
        RECT 89.265 1244.950 93.475 1245.025 ;
        RECT 87.120 1243.350 93.510 1244.950 ;
        RECT 89.265 1243.280 93.475 1243.350 ;
        RECT 30.425 1241.740 34.900 1241.850 ;
        RECT 30.425 1240.140 43.070 1241.740 ;
        RECT 30.425 1240.040 34.900 1240.140 ;
        RECT 95.310 1236.500 99.520 1236.575 ;
        RECT 87.120 1234.900 99.520 1236.500 ;
        RECT 95.310 1234.830 99.520 1234.900 ;
        RECT 205.330 1191.810 217.650 1226.940 ;
        RECT 221.270 1172.660 233.590 1206.790 ;
        RECT 89.230 1086.780 93.425 1086.895 ;
        RECT 71.550 1085.180 93.425 1086.780 ;
        RECT 89.230 1085.090 93.425 1085.180 ;
        RECT 95.260 1083.280 99.455 1083.350 ;
        RECT 71.550 1081.680 99.610 1083.280 ;
        RECT 95.260 1081.545 99.455 1081.680 ;
        RECT 36.395 1067.990 40.590 1068.095 ;
        RECT 36.300 1066.390 42.910 1067.990 ;
        RECT 36.395 1066.290 40.590 1066.390 ;
        RECT 89.245 1062.750 93.455 1062.840 ;
        RECT 87.120 1061.150 93.540 1062.750 ;
        RECT 89.245 1061.040 93.455 1061.150 ;
        RECT 30.440 1059.540 34.635 1059.700 ;
        RECT 30.240 1057.940 42.910 1059.540 ;
        RECT 30.440 1057.895 34.635 1057.940 ;
        RECT 95.280 1054.300 99.490 1054.365 ;
        RECT 87.120 1052.700 99.500 1054.300 ;
        RECT 95.280 1052.620 99.490 1052.700 ;
        RECT 239.180 1052.490 254.180 1188.060 ;
        RECT 262.990 1088.710 268.990 4113.290 ;
        RECT 270.990 1247.330 276.990 4121.450 ;
        RECT 3320.100 1347.330 3333.100 4973.980 ;
        RECT 3376.990 4512.240 3382.400 4517.730 ;
        RECT 3358.460 4504.150 3363.870 4509.640 ;
        RECT 3495.740 4497.780 3499.870 4497.840 ;
        RECT 3495.740 4496.180 3517.580 4497.780 ;
        RECT 3495.740 4496.125 3499.870 4496.180 ;
        RECT 3489.685 4494.280 3493.815 4494.355 ;
        RECT 3489.520 4492.680 3517.580 4494.280 ;
        RECT 3489.685 4492.640 3493.815 4492.680 ;
        RECT 3548.530 4478.990 3552.715 4479.075 ;
        RECT 3546.220 4477.390 3552.830 4478.990 ;
        RECT 3548.530 4477.300 3552.715 4477.390 ;
        RECT 3495.580 4473.750 3499.905 4473.850 ;
        RECT 3495.580 4472.150 3502.010 4473.750 ;
        RECT 3495.580 4472.080 3499.905 4472.150 ;
        RECT 3554.535 4470.540 3558.720 4470.620 ;
        RECT 3546.220 4468.940 3558.890 4470.540 ;
        RECT 3554.535 4468.845 3558.720 4468.940 ;
        RECT 3489.595 4465.300 3493.920 4465.360 ;
        RECT 3489.595 4463.700 3502.010 4465.300 ;
        RECT 3489.595 4463.590 3493.920 4463.700 ;
        RECT 3548.505 4462.090 3552.690 4462.205 ;
        RECT 3546.220 4460.490 3552.800 4462.090 ;
        RECT 3548.505 4460.430 3552.690 4460.490 ;
        RECT 3495.695 4456.850 3500.020 4456.935 ;
        RECT 3495.695 4455.250 3502.010 4456.850 ;
        RECT 3495.695 4455.165 3500.020 4455.250 ;
        RECT 3554.480 4453.640 3558.890 4453.750 ;
        RECT 3546.220 4452.140 3558.890 4453.640 ;
        RECT 3546.220 4452.060 3558.885 4452.140 ;
        RECT 3546.220 4452.040 3558.880 4452.060 ;
        RECT 3489.600 4448.400 3493.925 4448.460 ;
        RECT 3489.600 4446.800 3502.010 4448.400 ;
        RECT 3489.600 4446.690 3493.925 4446.800 ;
        RECT 3548.510 4445.190 3552.690 4445.280 ;
        RECT 3546.060 4443.590 3552.690 4445.190 ;
        RECT 3548.510 4443.480 3552.690 4443.590 ;
        RECT 3495.600 4439.950 3499.925 4440.055 ;
        RECT 3495.600 4438.350 3502.010 4439.950 ;
        RECT 3495.600 4438.285 3499.925 4438.350 ;
        RECT 3554.475 4436.740 3558.660 4436.820 ;
        RECT 3546.060 4435.140 3558.660 4436.740 ;
        RECT 3554.475 4435.045 3558.660 4435.140 ;
        RECT 3489.630 4431.500 3493.955 4431.600 ;
        RECT 3489.630 4429.900 3502.010 4431.500 ;
        RECT 3489.630 4429.830 3493.955 4429.900 ;
        RECT 291.110 1332.330 3333.100 1347.330 ;
        RECT 3336.100 1327.330 3349.100 4167.370 ;
        RECT 3377.040 3609.240 3382.450 3614.730 ;
        RECT 3358.510 3601.150 3363.920 3606.640 ;
        RECT 3495.790 3594.780 3499.920 3594.840 ;
        RECT 3495.790 3593.180 3517.630 3594.780 ;
        RECT 3495.790 3593.125 3499.920 3593.180 ;
        RECT 3489.735 3591.280 3493.865 3591.355 ;
        RECT 3489.570 3589.680 3517.630 3591.280 ;
        RECT 3489.735 3589.640 3493.865 3589.680 ;
        RECT 3548.580 3575.990 3552.765 3576.075 ;
        RECT 3546.270 3574.390 3552.880 3575.990 ;
        RECT 3548.580 3574.300 3552.765 3574.390 ;
        RECT 3495.630 3570.750 3499.955 3570.850 ;
        RECT 3495.630 3569.150 3502.060 3570.750 ;
        RECT 3495.630 3569.080 3499.955 3569.150 ;
        RECT 3554.585 3567.540 3558.770 3567.620 ;
        RECT 3546.270 3565.940 3558.940 3567.540 ;
        RECT 3554.585 3565.845 3558.770 3565.940 ;
        RECT 3489.645 3562.300 3493.970 3562.360 ;
        RECT 3489.645 3560.700 3502.060 3562.300 ;
        RECT 3489.645 3560.590 3493.970 3560.700 ;
        RECT 3548.555 3559.090 3552.740 3559.205 ;
        RECT 3546.270 3557.490 3552.850 3559.090 ;
        RECT 3548.555 3557.430 3552.740 3557.490 ;
        RECT 3495.745 3553.850 3500.070 3553.935 ;
        RECT 3495.745 3552.250 3502.060 3553.850 ;
        RECT 3495.745 3552.165 3500.070 3552.250 ;
        RECT 3554.530 3550.640 3558.940 3550.750 ;
        RECT 3546.270 3549.140 3558.940 3550.640 ;
        RECT 3546.270 3549.060 3558.935 3549.140 ;
        RECT 3546.270 3549.040 3558.930 3549.060 ;
        RECT 3489.650 3545.400 3493.975 3545.460 ;
        RECT 3489.650 3543.800 3502.060 3545.400 ;
        RECT 3489.650 3543.690 3493.975 3543.800 ;
        RECT 3548.560 3542.190 3552.740 3542.280 ;
        RECT 3546.110 3540.590 3552.740 3542.190 ;
        RECT 3548.560 3540.480 3552.740 3540.590 ;
        RECT 3495.650 3536.950 3499.975 3537.055 ;
        RECT 3495.650 3535.350 3502.060 3536.950 ;
        RECT 3495.650 3535.285 3499.975 3535.350 ;
        RECT 3554.525 3533.740 3558.710 3533.820 ;
        RECT 3546.110 3532.140 3558.710 3533.740 ;
        RECT 3554.525 3532.045 3558.710 3532.140 ;
        RECT 3489.680 3528.500 3494.005 3528.600 ;
        RECT 3489.680 3526.900 3502.060 3528.500 ;
        RECT 3489.680 3526.830 3494.005 3526.900 ;
        RECT 3377.040 3383.240 3382.450 3388.730 ;
        RECT 3358.510 3375.150 3363.920 3380.640 ;
        RECT 3495.790 3368.780 3499.920 3368.840 ;
        RECT 3495.790 3367.180 3517.630 3368.780 ;
        RECT 3495.790 3367.125 3499.920 3367.180 ;
        RECT 3489.735 3365.280 3493.865 3365.355 ;
        RECT 3489.570 3363.680 3517.630 3365.280 ;
        RECT 3489.735 3363.640 3493.865 3363.680 ;
        RECT 3548.580 3349.990 3552.765 3350.075 ;
        RECT 3546.270 3348.390 3552.880 3349.990 ;
        RECT 3548.580 3348.300 3552.765 3348.390 ;
        RECT 3495.630 3344.750 3499.955 3344.850 ;
        RECT 3495.630 3343.150 3502.060 3344.750 ;
        RECT 3495.630 3343.080 3499.955 3343.150 ;
        RECT 3554.585 3341.540 3558.770 3341.620 ;
        RECT 3546.270 3339.940 3558.940 3341.540 ;
        RECT 3554.585 3339.845 3558.770 3339.940 ;
        RECT 3489.645 3336.300 3493.970 3336.360 ;
        RECT 3489.645 3334.700 3502.060 3336.300 ;
        RECT 3489.645 3334.590 3493.970 3334.700 ;
        RECT 3548.555 3333.090 3552.740 3333.205 ;
        RECT 3546.270 3331.490 3552.850 3333.090 ;
        RECT 3548.555 3331.430 3552.740 3331.490 ;
        RECT 3495.745 3327.850 3500.070 3327.935 ;
        RECT 3495.745 3326.250 3502.060 3327.850 ;
        RECT 3495.745 3326.165 3500.070 3326.250 ;
        RECT 3554.530 3324.640 3558.940 3324.750 ;
        RECT 3546.270 3323.140 3558.940 3324.640 ;
        RECT 3546.270 3323.060 3558.935 3323.140 ;
        RECT 3546.270 3323.040 3558.930 3323.060 ;
        RECT 3489.650 3319.400 3493.975 3319.460 ;
        RECT 3489.650 3317.800 3502.060 3319.400 ;
        RECT 3489.650 3317.690 3493.975 3317.800 ;
        RECT 3548.560 3316.190 3552.740 3316.280 ;
        RECT 3546.110 3314.590 3552.740 3316.190 ;
        RECT 3548.560 3314.480 3552.740 3314.590 ;
        RECT 3495.650 3310.950 3499.975 3311.055 ;
        RECT 3495.650 3309.350 3502.060 3310.950 ;
        RECT 3495.650 3309.285 3499.975 3309.350 ;
        RECT 3554.525 3307.740 3558.710 3307.820 ;
        RECT 3546.110 3306.140 3558.710 3307.740 ;
        RECT 3554.525 3306.045 3558.710 3306.140 ;
        RECT 3489.680 3302.500 3494.005 3302.600 ;
        RECT 3489.680 3300.900 3502.060 3302.500 ;
        RECT 3489.680 3300.830 3494.005 3300.900 ;
        RECT 3377.040 3158.240 3382.450 3163.730 ;
        RECT 3358.510 3150.150 3363.920 3155.640 ;
        RECT 3495.790 3143.780 3499.920 3143.840 ;
        RECT 3495.790 3142.180 3517.630 3143.780 ;
        RECT 3495.790 3142.125 3499.920 3142.180 ;
        RECT 3489.735 3140.280 3493.865 3140.355 ;
        RECT 3489.570 3138.680 3517.630 3140.280 ;
        RECT 3489.735 3138.640 3493.865 3138.680 ;
        RECT 3548.580 3124.990 3552.765 3125.075 ;
        RECT 3546.270 3123.390 3552.880 3124.990 ;
        RECT 3548.580 3123.300 3552.765 3123.390 ;
        RECT 3495.630 3119.750 3499.955 3119.850 ;
        RECT 3495.630 3118.150 3502.060 3119.750 ;
        RECT 3495.630 3118.080 3499.955 3118.150 ;
        RECT 3554.585 3116.540 3558.770 3116.620 ;
        RECT 3546.270 3114.940 3558.940 3116.540 ;
        RECT 3554.585 3114.845 3558.770 3114.940 ;
        RECT 3489.645 3111.300 3493.970 3111.360 ;
        RECT 3489.645 3109.700 3502.060 3111.300 ;
        RECT 3489.645 3109.590 3493.970 3109.700 ;
        RECT 3548.555 3108.090 3552.740 3108.205 ;
        RECT 3546.270 3106.490 3552.850 3108.090 ;
        RECT 3548.555 3106.430 3552.740 3106.490 ;
        RECT 3495.745 3102.850 3500.070 3102.935 ;
        RECT 3495.745 3101.250 3502.060 3102.850 ;
        RECT 3495.745 3101.165 3500.070 3101.250 ;
        RECT 3554.530 3099.640 3558.940 3099.750 ;
        RECT 3546.270 3098.140 3558.940 3099.640 ;
        RECT 3546.270 3098.060 3558.935 3098.140 ;
        RECT 3546.270 3098.040 3558.930 3098.060 ;
        RECT 3489.650 3094.400 3493.975 3094.460 ;
        RECT 3489.650 3092.800 3502.060 3094.400 ;
        RECT 3489.650 3092.690 3493.975 3092.800 ;
        RECT 3548.560 3091.190 3552.740 3091.280 ;
        RECT 3546.110 3089.590 3552.740 3091.190 ;
        RECT 3548.560 3089.480 3552.740 3089.590 ;
        RECT 3495.650 3085.950 3499.975 3086.055 ;
        RECT 3495.650 3084.350 3502.060 3085.950 ;
        RECT 3495.650 3084.285 3499.975 3084.350 ;
        RECT 3554.525 3082.740 3558.710 3082.820 ;
        RECT 3546.110 3081.140 3558.710 3082.740 ;
        RECT 3554.525 3081.045 3558.710 3081.140 ;
        RECT 3489.680 3077.500 3494.005 3077.600 ;
        RECT 3489.680 3075.900 3502.060 3077.500 ;
        RECT 3489.680 3075.830 3494.005 3075.900 ;
        RECT 3377.040 2932.240 3382.450 2937.730 ;
        RECT 3358.510 2924.150 3363.920 2929.640 ;
        RECT 3495.790 2917.780 3499.920 2917.840 ;
        RECT 3495.790 2916.180 3517.630 2917.780 ;
        RECT 3495.790 2916.125 3499.920 2916.180 ;
        RECT 3489.735 2914.280 3493.865 2914.355 ;
        RECT 3489.570 2912.680 3517.630 2914.280 ;
        RECT 3489.735 2912.640 3493.865 2912.680 ;
        RECT 3548.580 2898.990 3552.765 2899.075 ;
        RECT 3546.270 2897.390 3552.880 2898.990 ;
        RECT 3548.580 2897.300 3552.765 2897.390 ;
        RECT 3495.630 2893.750 3499.955 2893.850 ;
        RECT 3495.630 2892.150 3502.060 2893.750 ;
        RECT 3495.630 2892.080 3499.955 2892.150 ;
        RECT 3554.585 2890.540 3558.770 2890.620 ;
        RECT 3546.270 2888.940 3558.940 2890.540 ;
        RECT 3554.585 2888.845 3558.770 2888.940 ;
        RECT 3489.645 2885.300 3493.970 2885.360 ;
        RECT 3489.645 2883.700 3502.060 2885.300 ;
        RECT 3489.645 2883.590 3493.970 2883.700 ;
        RECT 3548.555 2882.090 3552.740 2882.205 ;
        RECT 3546.270 2880.490 3552.850 2882.090 ;
        RECT 3548.555 2880.430 3552.740 2880.490 ;
        RECT 3495.745 2876.850 3500.070 2876.935 ;
        RECT 3495.745 2875.250 3502.060 2876.850 ;
        RECT 3495.745 2875.165 3500.070 2875.250 ;
        RECT 3554.530 2873.640 3558.940 2873.750 ;
        RECT 3546.270 2872.140 3558.940 2873.640 ;
        RECT 3546.270 2872.060 3558.935 2872.140 ;
        RECT 3546.270 2872.040 3558.930 2872.060 ;
        RECT 3489.650 2868.400 3493.975 2868.460 ;
        RECT 3489.650 2866.800 3502.060 2868.400 ;
        RECT 3489.650 2866.690 3493.975 2866.800 ;
        RECT 3548.560 2865.190 3552.740 2865.280 ;
        RECT 3546.110 2863.590 3552.740 2865.190 ;
        RECT 3548.560 2863.480 3552.740 2863.590 ;
        RECT 3495.650 2859.950 3499.975 2860.055 ;
        RECT 3495.650 2858.350 3502.060 2859.950 ;
        RECT 3495.650 2858.285 3499.975 2858.350 ;
        RECT 3554.525 2856.740 3558.710 2856.820 ;
        RECT 3546.110 2855.140 3558.710 2856.740 ;
        RECT 3554.525 2855.045 3558.710 2855.140 ;
        RECT 3489.680 2851.500 3494.005 2851.600 ;
        RECT 3489.680 2849.900 3502.060 2851.500 ;
        RECT 3489.680 2849.830 3494.005 2849.900 ;
        RECT 3377.040 2707.240 3382.450 2712.730 ;
        RECT 3358.510 2699.150 3363.920 2704.640 ;
        RECT 3495.790 2692.780 3499.920 2692.840 ;
        RECT 3495.790 2691.180 3517.630 2692.780 ;
        RECT 3495.790 2691.125 3499.920 2691.180 ;
        RECT 3489.735 2689.280 3493.865 2689.355 ;
        RECT 3489.570 2687.680 3517.630 2689.280 ;
        RECT 3489.735 2687.640 3493.865 2687.680 ;
        RECT 3548.580 2673.990 3552.765 2674.075 ;
        RECT 3546.270 2672.390 3552.880 2673.990 ;
        RECT 3548.580 2672.300 3552.765 2672.390 ;
        RECT 3495.630 2668.750 3499.955 2668.850 ;
        RECT 3495.630 2667.150 3502.060 2668.750 ;
        RECT 3495.630 2667.080 3499.955 2667.150 ;
        RECT 3554.585 2665.540 3558.770 2665.620 ;
        RECT 3546.270 2663.940 3558.940 2665.540 ;
        RECT 3554.585 2663.845 3558.770 2663.940 ;
        RECT 3489.645 2660.300 3493.970 2660.360 ;
        RECT 3489.645 2658.700 3502.060 2660.300 ;
        RECT 3489.645 2658.590 3493.970 2658.700 ;
        RECT 3548.555 2657.090 3552.740 2657.205 ;
        RECT 3546.270 2655.490 3552.850 2657.090 ;
        RECT 3548.555 2655.430 3552.740 2655.490 ;
        RECT 3495.745 2651.850 3500.070 2651.935 ;
        RECT 3495.745 2650.250 3502.060 2651.850 ;
        RECT 3495.745 2650.165 3500.070 2650.250 ;
        RECT 3554.530 2648.640 3558.940 2648.750 ;
        RECT 3546.270 2647.140 3558.940 2648.640 ;
        RECT 3546.270 2647.060 3558.935 2647.140 ;
        RECT 3546.270 2647.040 3558.930 2647.060 ;
        RECT 3489.650 2643.400 3493.975 2643.460 ;
        RECT 3489.650 2641.800 3502.060 2643.400 ;
        RECT 3489.650 2641.690 3493.975 2641.800 ;
        RECT 3548.560 2640.190 3552.740 2640.280 ;
        RECT 3546.110 2638.590 3552.740 2640.190 ;
        RECT 3548.560 2638.480 3552.740 2638.590 ;
        RECT 3495.650 2634.950 3499.975 2635.055 ;
        RECT 3495.650 2633.350 3502.060 2634.950 ;
        RECT 3495.650 2633.285 3499.975 2633.350 ;
        RECT 3554.525 2631.740 3558.710 2631.820 ;
        RECT 3546.110 2630.140 3558.710 2631.740 ;
        RECT 3554.525 2630.045 3558.710 2630.140 ;
        RECT 3489.680 2626.500 3494.005 2626.600 ;
        RECT 3489.680 2624.900 3502.060 2626.500 ;
        RECT 3489.680 2624.830 3494.005 2624.900 ;
        RECT 3377.040 2487.240 3382.450 2492.730 ;
        RECT 3358.510 2479.150 3363.920 2484.640 ;
        RECT 3495.790 2472.780 3499.920 2472.840 ;
        RECT 3495.790 2471.180 3517.630 2472.780 ;
        RECT 3495.790 2471.125 3499.920 2471.180 ;
        RECT 3489.735 2469.280 3493.865 2469.355 ;
        RECT 3489.570 2467.680 3517.630 2469.280 ;
        RECT 3489.735 2467.640 3493.865 2467.680 ;
        RECT 3548.580 2453.990 3552.765 2454.075 ;
        RECT 3546.270 2452.390 3552.880 2453.990 ;
        RECT 3548.580 2452.300 3552.765 2452.390 ;
        RECT 3495.630 2448.750 3499.955 2448.850 ;
        RECT 3495.630 2447.150 3502.060 2448.750 ;
        RECT 3495.630 2447.080 3499.955 2447.150 ;
        RECT 3554.585 2445.540 3558.770 2445.620 ;
        RECT 3546.270 2443.940 3558.940 2445.540 ;
        RECT 3554.585 2443.845 3558.770 2443.940 ;
        RECT 3489.645 2440.300 3493.970 2440.360 ;
        RECT 3489.645 2438.700 3502.060 2440.300 ;
        RECT 3489.645 2438.590 3493.970 2438.700 ;
        RECT 3548.555 2437.090 3552.740 2437.205 ;
        RECT 3546.270 2435.490 3552.850 2437.090 ;
        RECT 3548.555 2435.430 3552.740 2435.490 ;
        RECT 3495.745 2431.850 3500.070 2431.935 ;
        RECT 3495.745 2430.250 3502.060 2431.850 ;
        RECT 3495.745 2430.165 3500.070 2430.250 ;
        RECT 3554.530 2428.640 3558.940 2428.750 ;
        RECT 3546.270 2427.140 3558.940 2428.640 ;
        RECT 3546.270 2427.060 3558.935 2427.140 ;
        RECT 3546.270 2427.040 3558.930 2427.060 ;
        RECT 3489.650 2423.400 3493.975 2423.460 ;
        RECT 3489.650 2421.800 3502.060 2423.400 ;
        RECT 3489.650 2421.690 3493.975 2421.800 ;
        RECT 3548.560 2420.190 3552.740 2420.280 ;
        RECT 3546.110 2418.590 3552.740 2420.190 ;
        RECT 3548.560 2418.480 3552.740 2418.590 ;
        RECT 3495.650 2414.950 3499.975 2415.055 ;
        RECT 3495.650 2413.350 3502.060 2414.950 ;
        RECT 3495.650 2413.285 3499.975 2413.350 ;
        RECT 3554.525 2411.740 3558.710 2411.820 ;
        RECT 3546.110 2410.140 3558.710 2411.740 ;
        RECT 3554.525 2410.045 3558.710 2410.140 ;
        RECT 3489.680 2406.500 3494.005 2406.600 ;
        RECT 3489.680 2404.900 3502.060 2406.500 ;
        RECT 3489.680 2404.830 3494.005 2404.900 ;
        RECT 3377.040 2046.240 3382.450 2051.730 ;
        RECT 3358.510 2038.150 3363.920 2043.640 ;
        RECT 3495.790 2031.780 3499.920 2031.840 ;
        RECT 3495.790 2030.180 3517.630 2031.780 ;
        RECT 3495.790 2030.125 3499.920 2030.180 ;
        RECT 3489.735 2028.280 3493.865 2028.355 ;
        RECT 3489.570 2026.680 3517.630 2028.280 ;
        RECT 3489.735 2026.640 3493.865 2026.680 ;
        RECT 3548.580 2012.990 3552.765 2013.075 ;
        RECT 3546.270 2011.390 3552.880 2012.990 ;
        RECT 3548.580 2011.300 3552.765 2011.390 ;
        RECT 3495.630 2007.750 3499.955 2007.850 ;
        RECT 3495.630 2006.150 3502.060 2007.750 ;
        RECT 3495.630 2006.080 3499.955 2006.150 ;
        RECT 3554.585 2004.540 3558.770 2004.620 ;
        RECT 3546.270 2002.940 3558.940 2004.540 ;
        RECT 3554.585 2002.845 3558.770 2002.940 ;
        RECT 3489.645 1999.300 3493.970 1999.360 ;
        RECT 3489.645 1997.700 3502.060 1999.300 ;
        RECT 3489.645 1997.590 3493.970 1997.700 ;
        RECT 3548.555 1996.090 3552.740 1996.205 ;
        RECT 3546.270 1994.490 3552.850 1996.090 ;
        RECT 3548.555 1994.430 3552.740 1994.490 ;
        RECT 3495.745 1990.850 3500.070 1990.935 ;
        RECT 3495.745 1989.250 3502.060 1990.850 ;
        RECT 3495.745 1989.165 3500.070 1989.250 ;
        RECT 3554.530 1987.640 3558.940 1987.750 ;
        RECT 3546.270 1986.140 3558.940 1987.640 ;
        RECT 3546.270 1986.060 3558.935 1986.140 ;
        RECT 3546.270 1986.040 3558.930 1986.060 ;
        RECT 3489.650 1982.400 3493.975 1982.460 ;
        RECT 3489.650 1980.800 3502.060 1982.400 ;
        RECT 3489.650 1980.690 3493.975 1980.800 ;
        RECT 3548.560 1979.190 3552.740 1979.280 ;
        RECT 3546.110 1977.590 3552.740 1979.190 ;
        RECT 3548.560 1977.480 3552.740 1977.590 ;
        RECT 3495.650 1973.950 3499.975 1974.055 ;
        RECT 3495.650 1972.350 3502.060 1973.950 ;
        RECT 3495.650 1972.285 3499.975 1972.350 ;
        RECT 3554.525 1970.740 3558.710 1970.820 ;
        RECT 3546.110 1969.140 3558.710 1970.740 ;
        RECT 3554.525 1969.045 3558.710 1969.140 ;
        RECT 3489.680 1965.500 3494.005 1965.600 ;
        RECT 3489.680 1963.900 3502.060 1965.500 ;
        RECT 3489.680 1963.830 3494.005 1963.900 ;
        RECT 3377.040 1820.240 3382.450 1825.730 ;
        RECT 3358.510 1812.150 3363.920 1817.640 ;
        RECT 3495.790 1805.780 3499.920 1805.840 ;
        RECT 3495.790 1804.180 3517.630 1805.780 ;
        RECT 3495.790 1804.125 3499.920 1804.180 ;
        RECT 3489.735 1802.280 3493.865 1802.355 ;
        RECT 3489.570 1800.680 3517.630 1802.280 ;
        RECT 3489.735 1800.640 3493.865 1800.680 ;
        RECT 3548.580 1786.990 3552.765 1787.075 ;
        RECT 3546.270 1785.390 3552.880 1786.990 ;
        RECT 3548.580 1785.300 3552.765 1785.390 ;
        RECT 3495.630 1781.750 3499.955 1781.850 ;
        RECT 3495.630 1780.150 3502.060 1781.750 ;
        RECT 3495.630 1780.080 3499.955 1780.150 ;
        RECT 3554.585 1778.540 3558.770 1778.620 ;
        RECT 3546.270 1776.940 3558.940 1778.540 ;
        RECT 3554.585 1776.845 3558.770 1776.940 ;
        RECT 3489.645 1773.300 3493.970 1773.360 ;
        RECT 3489.645 1771.700 3502.060 1773.300 ;
        RECT 3489.645 1771.590 3493.970 1771.700 ;
        RECT 3548.555 1770.090 3552.740 1770.205 ;
        RECT 3546.270 1768.490 3552.850 1770.090 ;
        RECT 3548.555 1768.430 3552.740 1768.490 ;
        RECT 3495.745 1764.850 3500.070 1764.935 ;
        RECT 3495.745 1763.250 3502.060 1764.850 ;
        RECT 3495.745 1763.165 3500.070 1763.250 ;
        RECT 3554.530 1761.640 3558.940 1761.750 ;
        RECT 3546.270 1760.140 3558.940 1761.640 ;
        RECT 3546.270 1760.060 3558.935 1760.140 ;
        RECT 3546.270 1760.040 3558.930 1760.060 ;
        RECT 3489.650 1756.400 3493.975 1756.460 ;
        RECT 3489.650 1754.800 3502.060 1756.400 ;
        RECT 3489.650 1754.690 3493.975 1754.800 ;
        RECT 3548.560 1753.190 3552.740 1753.280 ;
        RECT 3546.110 1751.590 3552.740 1753.190 ;
        RECT 3548.560 1751.480 3552.740 1751.590 ;
        RECT 3495.650 1747.950 3499.975 1748.055 ;
        RECT 3495.650 1746.350 3502.060 1747.950 ;
        RECT 3495.650 1746.285 3499.975 1746.350 ;
        RECT 3554.525 1744.740 3558.710 1744.820 ;
        RECT 3546.110 1743.140 3558.710 1744.740 ;
        RECT 3554.525 1743.045 3558.710 1743.140 ;
        RECT 3489.680 1739.500 3494.005 1739.600 ;
        RECT 3489.680 1737.900 3502.060 1739.500 ;
        RECT 3489.680 1737.830 3494.005 1737.900 ;
        RECT 3377.040 1595.240 3382.450 1600.730 ;
        RECT 3358.510 1587.150 3363.920 1592.640 ;
        RECT 3495.790 1580.780 3499.920 1580.840 ;
        RECT 3495.790 1579.180 3517.630 1580.780 ;
        RECT 3495.790 1579.125 3499.920 1579.180 ;
        RECT 3489.735 1577.280 3493.865 1577.355 ;
        RECT 3489.570 1575.680 3517.630 1577.280 ;
        RECT 3489.735 1575.640 3493.865 1575.680 ;
        RECT 3548.580 1561.990 3552.765 1562.075 ;
        RECT 3546.270 1560.390 3552.880 1561.990 ;
        RECT 3548.580 1560.300 3552.765 1560.390 ;
        RECT 3495.630 1556.750 3499.955 1556.850 ;
        RECT 3495.630 1555.150 3502.060 1556.750 ;
        RECT 3495.630 1555.080 3499.955 1555.150 ;
        RECT 3554.585 1553.540 3558.770 1553.620 ;
        RECT 3546.270 1551.940 3558.940 1553.540 ;
        RECT 3554.585 1551.845 3558.770 1551.940 ;
        RECT 3489.645 1548.300 3493.970 1548.360 ;
        RECT 3489.645 1546.700 3502.060 1548.300 ;
        RECT 3489.645 1546.590 3493.970 1546.700 ;
        RECT 3548.555 1545.090 3552.740 1545.205 ;
        RECT 3546.270 1543.490 3552.850 1545.090 ;
        RECT 3548.555 1543.430 3552.740 1543.490 ;
        RECT 3495.745 1539.850 3500.070 1539.935 ;
        RECT 3495.745 1538.250 3502.060 1539.850 ;
        RECT 3495.745 1538.165 3500.070 1538.250 ;
        RECT 3554.530 1536.640 3558.940 1536.750 ;
        RECT 3546.270 1535.140 3558.940 1536.640 ;
        RECT 3546.270 1535.060 3558.935 1535.140 ;
        RECT 3546.270 1535.040 3558.930 1535.060 ;
        RECT 3489.650 1531.400 3493.975 1531.460 ;
        RECT 3489.650 1529.800 3502.060 1531.400 ;
        RECT 3489.650 1529.690 3493.975 1529.800 ;
        RECT 3548.560 1528.190 3552.740 1528.280 ;
        RECT 3546.110 1526.590 3552.740 1528.190 ;
        RECT 3548.560 1526.480 3552.740 1526.590 ;
        RECT 3495.650 1522.950 3499.975 1523.055 ;
        RECT 3495.650 1521.350 3502.060 1522.950 ;
        RECT 3495.650 1521.285 3499.975 1521.350 ;
        RECT 3554.525 1519.740 3558.710 1519.820 ;
        RECT 3546.110 1518.140 3558.710 1519.740 ;
        RECT 3554.525 1518.045 3558.710 1518.140 ;
        RECT 3489.680 1514.500 3494.005 1514.600 ;
        RECT 3489.680 1512.900 3502.060 1514.500 ;
        RECT 3489.680 1512.830 3494.005 1512.900 ;
        RECT 3377.040 1370.240 3382.450 1375.730 ;
        RECT 3358.510 1362.150 3363.920 1367.640 ;
        RECT 3495.790 1355.780 3499.920 1355.840 ;
        RECT 3495.790 1354.180 3517.630 1355.780 ;
        RECT 3495.790 1354.125 3499.920 1354.180 ;
        RECT 3489.735 1352.280 3493.865 1352.355 ;
        RECT 3489.570 1350.680 3517.630 1352.280 ;
        RECT 3489.735 1350.640 3493.865 1350.680 ;
        RECT 3548.580 1336.990 3552.765 1337.075 ;
        RECT 3546.270 1335.390 3552.880 1336.990 ;
        RECT 3548.580 1335.300 3552.765 1335.390 ;
        RECT 3495.630 1331.750 3499.955 1331.850 ;
        RECT 3495.630 1330.150 3502.060 1331.750 ;
        RECT 3495.630 1330.080 3499.955 1330.150 ;
        RECT 3554.585 1328.540 3558.770 1328.620 ;
        RECT 291.110 1312.330 3349.100 1327.330 ;
        RECT 3546.270 1326.940 3558.940 1328.540 ;
        RECT 3554.585 1326.845 3558.770 1326.940 ;
        RECT 3489.645 1323.300 3493.970 1323.360 ;
        RECT 3489.645 1321.700 3502.060 1323.300 ;
        RECT 3489.645 1321.590 3493.970 1321.700 ;
        RECT 3548.555 1320.090 3552.740 1320.205 ;
        RECT 3546.270 1318.490 3552.850 1320.090 ;
        RECT 3548.555 1318.430 3552.740 1318.490 ;
        RECT 3495.745 1314.850 3500.070 1314.935 ;
        RECT 3495.745 1313.250 3502.060 1314.850 ;
        RECT 3495.745 1313.165 3500.070 1313.250 ;
        RECT 3554.530 1311.640 3558.940 1311.750 ;
        RECT 3546.270 1310.140 3558.940 1311.640 ;
        RECT 3546.270 1310.060 3558.935 1310.140 ;
        RECT 3546.270 1310.040 3558.930 1310.060 ;
        RECT 281.850 1292.330 3255.870 1307.330 ;
        RECT 3489.650 1306.400 3493.975 1306.460 ;
        RECT 3489.650 1304.800 3502.060 1306.400 ;
        RECT 3489.650 1304.690 3493.975 1304.800 ;
        RECT 3548.560 1303.190 3552.740 1303.280 ;
        RECT 3546.110 1301.590 3552.740 1303.190 ;
        RECT 3548.560 1301.480 3552.740 1301.590 ;
        RECT 3495.650 1297.950 3499.975 1298.055 ;
        RECT 3495.650 1296.350 3502.060 1297.950 ;
        RECT 3495.650 1296.285 3499.975 1296.350 ;
        RECT 3554.525 1294.740 3558.710 1294.820 ;
        RECT 3546.110 1293.140 3558.710 1294.740 ;
        RECT 3554.525 1293.045 3558.710 1293.140 ;
        RECT 3489.680 1289.500 3494.005 1289.600 ;
        RECT 3489.680 1287.900 3502.060 1289.500 ;
        RECT 3489.680 1287.830 3494.005 1287.900 ;
        RECT 281.850 1272.330 3255.870 1287.330 ;
        RECT 280.630 1252.330 3354.930 1267.330 ;
        RECT 270.990 1232.330 3349.450 1247.330 ;
        RECT 3370.780 1233.080 3382.260 1246.480 ;
        RECT 270.990 1096.710 276.990 1232.330 ;
        RECT 281.390 1212.330 3254.730 1227.330 ;
        RECT 281.390 1192.330 3254.730 1207.330 ;
        RECT 281.440 1172.330 3026.950 1187.330 ;
        RECT 281.480 1152.330 3006.870 1167.330 ;
        RECT 36.485 1051.090 40.680 1051.205 ;
        RECT 36.330 1049.490 42.910 1051.090 ;
        RECT 36.485 1049.400 40.680 1049.490 ;
        RECT 239.180 1049.290 266.160 1052.490 ;
        RECT 2873.230 1049.290 2984.550 1052.490 ;
        RECT 89.285 1045.850 93.495 1045.890 ;
        RECT 87.120 1044.250 93.495 1045.850 ;
        RECT 89.285 1044.145 93.495 1044.250 ;
        RECT 30.170 1042.640 34.645 1042.770 ;
        RECT 30.170 1041.040 42.910 1042.640 ;
        RECT 30.170 1041.030 34.645 1041.040 ;
        RECT 95.265 1037.400 99.475 1037.475 ;
        RECT 87.120 1035.800 99.500 1037.400 ;
        RECT 95.265 1035.730 99.475 1035.800 ;
        RECT 36.385 1034.190 40.860 1034.265 ;
        RECT 36.385 1032.590 43.070 1034.190 ;
        RECT 36.385 1032.510 40.860 1032.590 ;
        RECT 89.265 1028.950 93.475 1029.025 ;
        RECT 87.120 1027.350 93.510 1028.950 ;
        RECT 89.265 1027.280 93.475 1027.350 ;
        RECT 30.425 1025.740 34.900 1025.850 ;
        RECT 30.425 1024.140 43.070 1025.740 ;
        RECT 30.425 1024.040 34.900 1024.140 ;
        RECT 95.310 1020.500 99.520 1020.575 ;
        RECT 87.120 1018.900 99.520 1020.500 ;
        RECT 95.310 1018.830 99.520 1018.900 ;
        RECT 239.180 922.490 254.180 1049.290 ;
        RECT 2981.350 1042.510 2984.550 1049.290 ;
        RECT 2981.350 1039.310 2988.710 1042.510 ;
        RECT 2991.870 987.490 3006.870 1152.330 ;
        RECT 256.720 984.290 266.080 987.490 ;
        RECT 2873.230 984.290 3006.870 987.490 ;
        RECT 239.180 919.290 266.060 922.490 ;
        RECT 2873.230 919.290 2984.550 922.490 ;
        RECT 208.840 240.370 228.840 884.370 ;
        RECT 239.180 833.940 254.180 919.290 ;
        RECT 2991.870 857.490 3006.870 984.290 ;
        RECT 256.230 854.290 266.200 857.490 ;
        RECT 2873.230 854.290 3006.870 857.490 ;
        RECT 234.180 792.490 254.180 833.940 ;
        RECT 234.180 789.290 266.100 792.490 ;
        RECT 2873.230 789.290 2984.550 792.490 ;
        RECT 234.180 662.490 254.180 789.290 ;
        RECT 2991.870 727.490 3006.870 854.290 ;
        RECT 255.890 724.290 266.330 727.490 ;
        RECT 2873.230 724.290 3006.870 727.490 ;
        RECT 234.180 659.290 266.030 662.490 ;
        RECT 2873.230 659.290 2984.550 662.490 ;
        RECT 234.180 532.490 254.180 659.290 ;
        RECT 2991.870 597.490 3006.870 724.290 ;
        RECT 255.890 594.290 266.330 597.490 ;
        RECT 2873.230 594.290 3006.870 597.490 ;
        RECT 234.180 529.290 266.110 532.490 ;
        RECT 2873.230 529.290 2984.550 532.490 ;
        RECT 234.180 402.490 254.180 529.290 ;
        RECT 2991.870 467.490 3006.870 594.290 ;
        RECT 255.890 464.290 266.330 467.490 ;
        RECT 2873.230 464.290 3006.870 467.490 ;
        RECT 234.180 399.290 265.840 402.490 ;
        RECT 2873.230 399.290 2984.550 402.490 ;
        RECT 234.180 233.940 254.180 399.290 ;
        RECT 2991.870 337.490 3006.870 464.290 ;
        RECT 256.810 334.290 265.860 337.490 ;
        RECT 2873.770 334.290 3006.870 337.490 ;
        RECT 2991.870 261.110 3006.870 334.290 ;
        RECT 271.870 241.110 3006.870 261.110 ;
        RECT 3011.950 1122.680 3026.950 1172.330 ;
        RECT 3377.040 1144.240 3382.450 1149.730 ;
        RECT 3358.510 1136.150 3363.920 1141.640 ;
        RECT 3243.330 1129.360 3255.950 1130.960 ;
        RECT 3011.950 1120.960 3205.220 1122.680 ;
        RECT 3011.950 1119.360 3209.950 1120.960 ;
        RECT 3011.950 1116.680 3205.220 1119.360 ;
        RECT 3011.950 911.050 3026.950 1116.680 ;
        RECT 3249.950 1110.960 3255.950 1129.360 ;
        RECT 3495.790 1129.780 3499.920 1129.840 ;
        RECT 3495.790 1128.180 3517.630 1129.780 ;
        RECT 3495.790 1128.125 3499.920 1128.180 ;
        RECT 3489.735 1126.280 3493.865 1126.355 ;
        RECT 3489.570 1124.680 3517.630 1126.280 ;
        RECT 3489.735 1124.640 3493.865 1124.680 ;
        RECT 3548.580 1110.990 3552.765 1111.075 ;
        RECT 3243.310 1109.360 3255.950 1110.960 ;
        RECT 3546.270 1109.390 3552.880 1110.990 ;
        RECT 3249.950 1062.520 3255.950 1109.360 ;
        RECT 3548.580 1109.300 3552.765 1109.390 ;
        RECT 3495.630 1105.750 3499.955 1105.850 ;
        RECT 3495.630 1104.150 3502.060 1105.750 ;
        RECT 3495.630 1104.080 3499.955 1104.150 ;
        RECT 3554.585 1102.540 3558.770 1102.620 ;
        RECT 3546.270 1100.940 3558.940 1102.540 ;
        RECT 3554.585 1100.845 3558.770 1100.940 ;
        RECT 3489.645 1097.300 3493.970 1097.360 ;
        RECT 3489.645 1095.700 3502.060 1097.300 ;
        RECT 3489.645 1095.590 3493.970 1095.700 ;
        RECT 3548.555 1094.090 3552.740 1094.205 ;
        RECT 3546.270 1092.490 3552.850 1094.090 ;
        RECT 3548.555 1092.430 3552.740 1092.490 ;
        RECT 3495.745 1088.850 3500.070 1088.935 ;
        RECT 3495.745 1087.250 3502.060 1088.850 ;
        RECT 3495.745 1087.165 3500.070 1087.250 ;
        RECT 3554.530 1085.640 3558.940 1085.750 ;
        RECT 3546.270 1084.140 3558.940 1085.640 ;
        RECT 3546.270 1084.060 3558.935 1084.140 ;
        RECT 3546.270 1084.040 3558.930 1084.060 ;
        RECT 3489.650 1080.400 3493.975 1080.460 ;
        RECT 3489.650 1078.800 3502.060 1080.400 ;
        RECT 3489.650 1078.690 3493.975 1078.800 ;
        RECT 3548.560 1077.190 3552.740 1077.280 ;
        RECT 3546.110 1075.590 3552.740 1077.190 ;
        RECT 3548.560 1075.480 3552.740 1075.590 ;
        RECT 3495.650 1071.950 3499.975 1072.055 ;
        RECT 3495.650 1070.350 3502.060 1071.950 ;
        RECT 3495.650 1070.285 3499.975 1070.350 ;
        RECT 3554.525 1068.740 3558.710 1068.820 ;
        RECT 3546.110 1067.140 3558.710 1068.740 ;
        RECT 3554.525 1067.045 3558.710 1067.140 ;
        RECT 3489.680 1063.500 3494.005 1063.600 ;
        RECT 3036.260 1047.520 3347.130 1062.520 ;
        RECT 3489.680 1061.900 3502.060 1063.500 ;
        RECT 3489.680 1061.830 3494.005 1061.900 ;
        RECT 3332.130 987.640 3347.130 1047.520 ;
        RECT 3029.880 986.040 3037.970 987.640 ;
        RECT 3326.190 986.040 3347.130 987.640 ;
        RECT 3011.950 909.450 3037.970 911.050 ;
        RECT 3011.950 757.870 3026.950 909.450 ;
        RECT 3332.130 834.460 3347.130 986.040 ;
        RECT 3377.040 919.240 3382.450 924.730 ;
        RECT 3358.510 911.150 3363.920 916.640 ;
        RECT 3495.790 904.780 3499.920 904.840 ;
        RECT 3495.790 903.180 3517.630 904.780 ;
        RECT 3495.790 903.125 3499.920 903.180 ;
        RECT 3489.735 901.280 3493.865 901.355 ;
        RECT 3489.570 899.680 3517.630 901.280 ;
        RECT 3489.735 899.640 3493.865 899.680 ;
        RECT 3548.580 885.990 3552.765 886.075 ;
        RECT 3546.270 884.390 3552.880 885.990 ;
        RECT 3548.580 884.300 3552.765 884.390 ;
        RECT 3495.630 880.750 3499.955 880.850 ;
        RECT 3495.630 879.150 3502.060 880.750 ;
        RECT 3495.630 879.080 3499.955 879.150 ;
        RECT 3554.585 877.540 3558.770 877.620 ;
        RECT 3546.270 875.940 3558.940 877.540 ;
        RECT 3554.585 875.845 3558.770 875.940 ;
        RECT 3489.645 872.300 3493.970 872.360 ;
        RECT 3489.645 870.700 3502.060 872.300 ;
        RECT 3489.645 870.590 3493.970 870.700 ;
        RECT 3548.555 869.090 3552.740 869.205 ;
        RECT 3546.270 867.490 3552.850 869.090 ;
        RECT 3548.555 867.430 3552.740 867.490 ;
        RECT 3495.745 863.850 3500.070 863.935 ;
        RECT 3495.745 862.250 3502.060 863.850 ;
        RECT 3495.745 862.165 3500.070 862.250 ;
        RECT 3554.530 860.640 3558.940 860.750 ;
        RECT 3546.270 859.140 3558.940 860.640 ;
        RECT 3546.270 859.060 3558.935 859.140 ;
        RECT 3546.270 859.040 3558.930 859.060 ;
        RECT 3489.650 855.400 3493.975 855.460 ;
        RECT 3489.650 853.800 3502.060 855.400 ;
        RECT 3489.650 853.690 3493.975 853.800 ;
        RECT 3548.560 852.190 3552.740 852.280 ;
        RECT 3546.110 850.590 3552.740 852.190 ;
        RECT 3548.560 850.480 3552.740 850.590 ;
        RECT 3495.650 846.950 3499.975 847.055 ;
        RECT 3495.650 845.350 3502.060 846.950 ;
        RECT 3495.650 845.285 3499.975 845.350 ;
        RECT 3554.525 843.740 3558.710 843.820 ;
        RECT 3546.110 842.140 3558.710 843.740 ;
        RECT 3554.525 842.045 3558.710 842.140 ;
        RECT 3489.680 838.500 3494.005 838.600 ;
        RECT 3489.680 836.900 3502.060 838.500 ;
        RECT 3489.680 836.830 3494.005 836.900 ;
        RECT 3029.760 832.860 3037.970 834.460 ;
        RECT 3326.030 832.860 3347.130 834.460 ;
        RECT 3011.950 756.270 3037.970 757.870 ;
        RECT 3011.950 604.690 3026.950 756.270 ;
        RECT 3332.130 681.280 3347.130 832.860 ;
        RECT 3377.040 693.240 3382.450 698.730 ;
        RECT 3358.510 685.150 3363.920 690.640 ;
        RECT 3029.700 679.680 3037.970 681.280 ;
        RECT 3325.820 679.680 3347.130 681.280 ;
        RECT 3011.950 603.090 3038.050 604.690 ;
        RECT 3011.950 494.780 3026.950 603.090 ;
        RECT 3332.130 528.100 3347.130 679.680 ;
        RECT 3495.790 678.780 3499.920 678.840 ;
        RECT 3495.790 677.180 3517.630 678.780 ;
        RECT 3495.790 677.125 3499.920 677.180 ;
        RECT 3489.735 675.280 3493.865 675.355 ;
        RECT 3489.570 673.680 3517.630 675.280 ;
        RECT 3489.735 673.640 3493.865 673.680 ;
        RECT 3548.580 659.990 3552.765 660.075 ;
        RECT 3546.270 658.390 3552.880 659.990 ;
        RECT 3548.580 658.300 3552.765 658.390 ;
        RECT 3495.630 654.750 3499.955 654.850 ;
        RECT 3495.630 653.150 3502.060 654.750 ;
        RECT 3495.630 653.080 3499.955 653.150 ;
        RECT 3554.585 651.540 3558.770 651.620 ;
        RECT 3546.270 649.940 3558.940 651.540 ;
        RECT 3554.585 649.845 3558.770 649.940 ;
        RECT 3489.645 646.300 3493.970 646.360 ;
        RECT 3489.645 644.700 3502.060 646.300 ;
        RECT 3489.645 644.590 3493.970 644.700 ;
        RECT 3548.555 643.090 3552.740 643.205 ;
        RECT 3546.270 641.490 3552.850 643.090 ;
        RECT 3548.555 641.430 3552.740 641.490 ;
        RECT 3495.745 637.850 3500.070 637.935 ;
        RECT 3495.745 636.250 3502.060 637.850 ;
        RECT 3495.745 636.165 3500.070 636.250 ;
        RECT 3554.530 634.640 3558.940 634.750 ;
        RECT 3546.270 633.140 3558.940 634.640 ;
        RECT 3546.270 633.060 3558.935 633.140 ;
        RECT 3546.270 633.040 3558.930 633.060 ;
        RECT 3489.650 629.400 3493.975 629.460 ;
        RECT 3489.650 627.800 3502.060 629.400 ;
        RECT 3489.650 627.690 3493.975 627.800 ;
        RECT 3548.560 626.190 3552.740 626.280 ;
        RECT 3546.110 624.590 3552.740 626.190 ;
        RECT 3548.560 624.480 3552.740 624.590 ;
        RECT 3495.650 620.950 3499.975 621.055 ;
        RECT 3495.650 619.350 3502.060 620.950 ;
        RECT 3495.650 619.285 3499.975 619.350 ;
        RECT 3554.525 617.740 3558.710 617.820 ;
        RECT 3546.110 616.140 3558.710 617.740 ;
        RECT 3554.525 616.045 3558.710 616.140 ;
        RECT 3489.680 612.500 3494.005 612.600 ;
        RECT 3489.680 610.900 3502.060 612.500 ;
        RECT 3489.680 610.830 3494.005 610.900 ;
        RECT 3029.700 526.500 3037.970 528.100 ;
        RECT 3325.880 526.500 3347.130 528.100 ;
        RECT 3011.950 479.780 3288.640 494.780 ;
        RECT 3011.950 235.940 3026.950 479.780 ;
        RECT 3124.120 453.700 3139.120 479.780 ;
        RECT 3217.720 467.370 3232.720 467.940 ;
        RECT 3209.530 465.770 3232.720 467.370 ;
        RECT 3115.380 447.370 3139.120 453.700 ;
        RECT 3115.380 445.770 3146.810 447.370 ;
        RECT 3115.380 445.060 3139.120 445.770 ;
        RECT 3115.380 380.960 3121.040 445.060 ;
        RECT 3217.720 427.370 3232.720 465.770 ;
        RECT 3254.970 462.950 3269.970 479.780 ;
        RECT 3332.130 467.030 3347.130 526.500 ;
        RECT 3312.610 465.430 3347.130 467.030 ;
        RECT 3254.970 461.350 3288.770 462.950 ;
        RECT 3254.970 454.790 3269.970 461.350 ;
        RECT 3332.130 458.870 3347.130 465.430 ;
        RECT 3312.420 457.270 3347.130 458.870 ;
        RECT 3254.970 453.190 3288.920 454.790 ;
        RECT 3254.970 452.610 3269.970 453.190 ;
        RECT 3332.130 450.710 3347.130 457.270 ;
        RECT 3312.520 449.110 3347.130 450.710 ;
        RECT 3209.840 425.770 3232.720 427.370 ;
        RECT 3217.720 405.410 3232.720 425.770 ;
        RECT 3332.130 405.410 3347.130 449.110 ;
        RECT 3160.010 390.410 3347.130 405.410 ;
        RECT 3210.450 387.960 3219.300 390.410 ;
        RECT 3122.800 382.960 3219.300 387.960 ;
        RECT 3102.590 375.960 3195.950 380.960 ;
        RECT 3102.590 360.600 3106.590 375.960 ;
        RECT 3205.920 369.050 3209.920 382.960 ;
        RECT 3202.180 367.450 3209.920 369.050 ;
        RECT 3102.590 359.000 3109.340 360.600 ;
        RECT 3102.590 343.700 3106.590 359.000 ;
        RECT 3205.920 352.150 3209.920 367.450 ;
        RECT 3202.010 350.550 3209.920 352.150 ;
        RECT 3102.590 342.100 3108.730 343.700 ;
        RECT 3102.590 331.080 3106.590 342.100 ;
        RECT 3205.920 335.250 3209.920 350.550 ;
        RECT 3202.620 333.650 3209.920 335.250 ;
        RECT 3205.920 329.790 3209.920 333.650 ;
        RECT 3011.950 233.940 3248.340 235.940 ;
        RECT 3332.130 234.890 3347.130 390.410 ;
        RECT 234.180 232.940 3248.340 233.940 ;
        RECT 234.180 228.940 3026.950 232.940 ;
        RECT 234.180 213.940 3026.980 228.940 ;
  END
END caravan_power_routing
END LIBRARY

