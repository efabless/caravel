module copyright_block ();
endmodule
