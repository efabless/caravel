VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_clocking
  CLASS BLOCK ;
  FOREIGN caravel_clocking ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.500 2.480 17.100 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.000 2.480 32.600 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.500 2.480 48.100 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.000 2.480 63.600 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 77.500 2.480 79.100 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.000 2.480 94.600 92.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 16.100 94.600 17.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 33.000 94.600 34.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 49.900 94.600 51.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 66.800 94.600 68.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 83.700 94.600 85.300 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 7.750 2.480 9.350 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.250 2.480 24.850 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.750 2.480 40.350 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.250 2.480 55.850 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.750 2.480 71.350 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.250 2.480 86.850 92.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 7.650 94.540 9.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 24.550 94.540 26.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 41.450 94.540 43.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 58.350 94.540 59.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 75.250 94.540 76.850 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 96.000 35.790 100.000 ;
    END
  END core_clk
  PIN ext_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 96.000 21.530 100.000 ;
    END
  END ext_clk
  PIN ext_clk_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END ext_clk_sel
  PIN ext_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 92.520 100.000 93.120 ;
    END
  END ext_reset
  PIN pll_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 96.000 78.570 100.000 ;
    END
  END pll_clk
  PIN pll_clk90
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 96.000 92.830 100.000 ;
    END
  END pll_clk90
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 96.000 7.270 100.000 ;
    END
  END resetb
  PIN resetb_sync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 96.000 64.310 100.000 ;
    END
  END resetb_sync
  PIN sel2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.800 100.000 56.400 ;
    END
  END sel2[0]
  PIN sel2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END sel2[1]
  PIN sel2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 80.280 100.000 80.880 ;
    END
  END sel2[2]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 19.080 100.000 19.680 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 31.320 100.000 31.920 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 43.560 100.000 44.160 ;
    END
  END sel[2]
  PIN user_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 96.000 50.050 100.000 ;
    END
  END user_clk
  OBS
      LAYER li1 ;
        RECT 0.920 2.635 94.300 92.565 ;
      LAYER met1 ;
        RECT 0.920 2.480 95.610 92.720 ;
      LAYER met2 ;
        RECT 2.860 95.720 6.710 96.290 ;
        RECT 7.550 95.720 20.970 96.290 ;
        RECT 21.810 95.720 35.230 96.290 ;
        RECT 36.070 95.720 49.490 96.290 ;
        RECT 50.330 95.720 63.750 96.290 ;
        RECT 64.590 95.720 78.010 96.290 ;
        RECT 78.850 95.720 92.270 96.290 ;
        RECT 93.110 95.720 95.590 96.290 ;
        RECT 2.860 2.535 95.590 95.720 ;
      LAYER met3 ;
        RECT 7.760 92.120 95.600 92.985 ;
        RECT 7.760 81.280 96.000 92.120 ;
        RECT 7.760 79.880 95.600 81.280 ;
        RECT 7.760 69.040 96.000 79.880 ;
        RECT 7.760 67.640 95.600 69.040 ;
        RECT 7.760 56.800 96.000 67.640 ;
        RECT 7.760 55.400 95.600 56.800 ;
        RECT 7.760 44.560 96.000 55.400 ;
        RECT 7.760 43.160 95.600 44.560 ;
        RECT 7.760 32.320 96.000 43.160 ;
        RECT 7.760 30.920 95.600 32.320 ;
        RECT 7.760 20.080 96.000 30.920 ;
        RECT 7.760 18.680 95.600 20.080 ;
        RECT 7.760 7.840 96.000 18.680 ;
        RECT 7.760 6.440 95.600 7.840 ;
        RECT 7.760 2.555 96.000 6.440 ;
  END
END caravel_clocking
END LIBRARY

