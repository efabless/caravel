* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_39_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6914_ _7081_/CLK _6914_/D fanout478/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6845_ _6951_/CLK _6845_/D fanout474/X VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6776_ _6777_/CLK _6776_/D fanout483/X VGND VGND VPWR VPWR _7195_/A sky130_fd_sc_hd__dfrtp_1
X_3988_ hold151/X hold99/X _3989_/S VGND VGND VPWR VPWR _3988_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5727_ _6909_/Q _5814_/B1 _5724_/X _5726_/X VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__a211o_1
XFILLER_148_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5658_ _5664_/A _5658_/B _5666_/B VGND VGND VPWR VPWR _5658_/X sky130_fd_sc_hd__and3b_4
XFILLER_191_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4609_ _4607_/A _4753_/B VGND VGND VPWR VPWR _4609_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5589_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5979_/A sky130_fd_sc_hd__and2b_4
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold340 _4055_/X VGND VGND VPWR VPWR _6491_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold351 _6463_/Q VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _4236_/X VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _6718_/Q VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _4108_/X VGND VGND VPWR VPWR _6523_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _7196_/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1040 _4061_/X VGND VGND VPWR VPWR _6494_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 hold1577/X VGND VGND VPWR VPWR _5172_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _5383_/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1073 _6611_/Q VGND VGND VPWR VPWR _4211_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1084 _5485_/X VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_202 _5652_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _6516_/Q VGND VGND VPWR VPWR _4099_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4960_ _4947_/C _4959_/Y _5018_/A _4775_/B VGND VGND VPWR VPWR _5088_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3911_ _3164_/Y _7158_/Q _3868_/S _3911_/B1 VGND VGND VPWR VPWR _3911_/X sky130_fd_sc_hd__a31o_1
XFILLER_17_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4891_ _4810_/A _4947_/C _4902_/B _4490_/B _4878_/C VGND VGND VPWR VPWR _5029_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6630_ _6632_/CLK _6630_/D fanout454/X VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3842_ _3866_/S VGND VGND VPWR VPWR _3851_/C sky130_fd_sc_hd__inv_2
XFILLER_20_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6561_ _6653_/CLK _6561_/D fanout452/X VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfrtp_2
X_3773_ _3773_/A _3773_/B _3773_/C VGND VGND VPWR VPWR _3794_/A sky130_fd_sc_hd__nor3_1
XFILLER_192_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5512_ hold145/X hold99/X _5513_/S VGND VGND VPWR VPWR _5512_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6492_ _6527_/CLK hold90/X fanout484/X VGND VGND VPWR VPWR _7183_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5443_ hold928/X _5548_/A1 _5444_/S VGND VGND VPWR VPWR _5443_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5374_ _5374_/A0 _5524_/A1 _5381_/S VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7113_ _7113_/CLK _7113_/D fanout459/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_2
X_4325_ hold431/X _5544_/A1 _4327_/S VGND VGND VPWR VPWR _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7044_ _7069_/CLK hold78/X fanout482/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_1
X_4256_ _4256_/A _4322_/B VGND VGND VPWR VPWR _4261_/S sky130_fd_sc_hd__and2_2
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3207_ _6917_/Q VGND VGND VPWR VPWR _3207_/Y sky130_fd_sc_hd__inv_2
X_4187_ _6638_/Q _6307_/B VGND VGND VPWR VPWR _4195_/S sky130_fd_sc_hd__nand2_8
XFILLER_95_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6828_ _6908_/CLK _6828_/D fanout475/X VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_1
X_6759_ _6953_/CLK _6759_/D fanout459/X VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold170 _7174_/A VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold181 _5297_/X VGND VGND VPWR VPWR _6862_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold192 _6559_/Q VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4110_ _4110_/A0 _5473_/A1 hold38/X VGND VGND VPWR VPWR _4110_/X sky130_fd_sc_hd__mux2_1
X_5090_ _4672_/B _4496_/Y _4542_/B VGND VGND VPWR VPWR _5090_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4041_ hold968/X _6355_/A1 _4043_/S VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5992_ _6818_/Q _5953_/X _5960_/X _7071_/Q _5991_/X VGND VGND VPWR VPWR _5992_/X
+ sky130_fd_sc_hd__a221o_1
X_4943_ _4673_/A _4619_/Y _4995_/B _4941_/X _5071_/A VGND VGND VPWR VPWR _4944_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4874_ _4542_/A _4947_/B _4652_/Y _4694_/Y _4873_/X VGND VGND VPWR VPWR _4875_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6613_ _6654_/CLK _6613_/D fanout454/X VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3825_ _6874_/Q _5310_/A _5229_/A _6802_/Q _3824_/X VGND VGND VPWR VPWR _3826_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6544_ _6709_/CLK _6544_/D fanout445/X VGND VGND VPWR VPWR _6544_/Q sky130_fd_sc_hd__dfstp_2
X_3756_ _7064_/Q _5523_/A _4286_/A _6681_/Q VGND VGND VPWR VPWR _3756_/X sky130_fd_sc_hd__a22o_2
XFILLER_9_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_6475_ _6707_/CLK _6475_/D fanout445/X VGND VGND VPWR VPWR _6475_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3687_ _6662_/Q _4262_/A _3684_/X _3686_/X VGND VGND VPWR VPWR _3688_/C sky130_fd_sc_hd__a211o_1
XFILLER_133_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5426_ hold700/X _5513_/A1 _5426_/S VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__mux2_1
Xoutput220 _7183_/X VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput231 _7193_/X VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput242 _7175_/X VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput253 _3948_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
Xoutput264 _6739_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
X_5357_ hold305/X _5465_/A1 _5363_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput275 _6431_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
Xoutput286 _6425_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xoutput297 _6751_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
X_4308_ hold748/X _6356_/A1 _4309_/S VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5288_ hold459/X _5528_/A1 _5291_/S VGND VGND VPWR VPWR _5288_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7027_ _7085_/CLK _7027_/D fanout477/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfstp_2
X_4239_ _4239_/A0 _6353_/A1 _4243_/S VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire347 _3437_/Y VGND VGND VPWR VPWR _3447_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_139_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire358 _3392_/Y VGND VGND VPWR VPWR _3410_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout480 fanout485/X VGND VGND VPWR VPWR fanout480/X sky130_fd_sc_hd__buf_4
XFILLER_93_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3610_ _6909_/Q _5346_/A _4102_/A input64/X _3609_/X VGND VGND VPWR VPWR _3611_/D
+ sky130_fd_sc_hd__a221o_1
X_4590_ _4591_/A _4664_/B VGND VGND VPWR VPWR _4747_/A sky130_fd_sc_hd__and2_1
X_3541_ _6854_/Q _5283_/A _5319_/A _6886_/Q _3540_/X VGND VGND VPWR VPWR _3552_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_183_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold906 _6976_/Q VGND VGND VPWR VPWR hold906/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold917 _5296_/X VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 _6992_/Q VGND VGND VPWR VPWR hold928/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6260_ _6633_/Q _5946_/X _5955_/X _6553_/Q VGND VGND VPWR VPWR _6260_/X sky130_fd_sc_hd__a22o_1
Xhold939 _5530_/X VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3472_ _3472_/A _3472_/B _3472_/C VGND VGND VPWR VPWR _3485_/A sky130_fd_sc_hd__nor3_1
XFILLER_143_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5211_ _5211_/A hold17/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__and2_4
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6191_ _6650_/Q _5973_/A _5948_/X _6695_/Q _6190_/X VGND VGND VPWR VPWR _6191_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5142_ _5142_/A _5142_/B _5142_/C _5142_/D VGND VGND VPWR VPWR _5142_/Y sky130_fd_sc_hd__nand4_1
XFILLER_96_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5073_ _5073_/A _5073_/B _5073_/C VGND VGND VPWR VPWR _5074_/C sky130_fd_sc_hd__and3_1
XFILLER_56_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4024_ hold351/X _5494_/A1 _4025_/S VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5975_ _5975_/A _5975_/B _5975_/C _5975_/D VGND VGND VPWR VPWR _5975_/Y sky130_fd_sc_hd__nor4_1
X_4926_ _4992_/A _4926_/B VGND VGND VPWR VPWR _5068_/C sky130_fd_sc_hd__nand2_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4857_ _4810_/A _4496_/Y _4856_/Y _4887_/A VGND VGND VPWR VPWR _4878_/C sky130_fd_sc_hd__o22a_1
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3808_ _6938_/Q _5382_/A _4304_/A _6695_/Q VGND VGND VPWR VPWR _3808_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4788_ _4689_/A _4616_/Y _4658_/C VGND VGND VPWR VPWR _5106_/A sky130_fd_sc_hd__o21a_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6527_ _6527_/CLK _6527_/D fanout484/X VGND VGND VPWR VPWR _6527_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ input15/X _3381_/Y _5148_/A _6738_/Q _3738_/X VGND VGND VPWR VPWR _3742_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_180_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6458_ _6747_/CLK _6458_/D fanout448/X VGND VGND VPWR VPWR _6458_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5409_ _5409_/A hold17/X VGND VGND VPWR VPWR _5417_/S sky130_fd_sc_hd__and2_4
XFILLER_0_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6389_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6389_/X sky130_fd_sc_hd__and2_1
XFILLER_121_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5760_ _6991_/Q _5627_/X _5635_/X _6831_/Q VGND VGND VPWR VPWR _5760_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4711_ _4701_/Y _4710_/Y _4627_/A VGND VGND VPWR VPWR _4711_/X sky130_fd_sc_hd__o21a_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5691_ _5681_/Y _5690_/Y _6787_/Q _5652_/Y VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4642_ _4642_/A _4673_/B VGND VGND VPWR VPWR _4644_/B sky130_fd_sc_hd__nor2_4
XFILLER_162_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4573_ _4965_/B _4724_/A VGND VGND VPWR VPWR _5041_/B sky130_fd_sc_hd__nand2_1
Xhold703 _5289_/X VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6312_ _6312_/A0 _6312_/A1 _6315_/S VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__mux2_1
Xhold714 _6824_/Q VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__dlygate4sd3_1
X_3524_ _3562_/A _3546_/A VGND VGND VPWR VPWR _4202_/A sky130_fd_sc_hd__nor2_8
Xhold725 _4296_/X VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold736 _6568_/Q VGND VGND VPWR VPWR hold736/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold747 _5255_/X VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _6543_/Q VGND VGND VPWR VPWR hold758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 _6356_/X VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6243_ _6562_/Q _5953_/X _5960_/X _6672_/Q _6242_/X VGND VGND VPWR VPWR _6243_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ _3455_/A _3577_/B VGND VGND VPWR VPWR _4102_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6174_ _7062_/Q _5954_/X _5976_/D _6881_/Q _6156_/X VGND VGND VPWR VPWR _6175_/D
+ sky130_fd_sc_hd__a221o_1
X_3386_ _7017_/Q _5463_/A _3370_/Y _7009_/Q VGND VGND VPWR VPWR _3386_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5125_ _4413_/Y _4946_/X _5124_/X _4823_/X VGND VGND VPWR VPWR _5126_/C sky130_fd_sc_hd__o211a_1
Xhold1403 _6798_/Q VGND VGND VPWR VPWR _5225_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1414 _6572_/Q VGND VGND VPWR VPWR hold1414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 _6583_/Q VGND VGND VPWR VPWR hold1425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1436 _7138_/Q VGND VGND VPWR VPWR _6313_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 _6595_/Q VGND VGND VPWR VPWR _4192_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5056_ _5089_/B _5089_/C _5142_/A _5056_/D VGND VGND VPWR VPWR _5058_/D sky130_fd_sc_hd__and4_1
Xhold1458 _6729_/Q VGND VGND VPWR VPWR _3702_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _6573_/Q VGND VGND VPWR VPWR _4167_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4007_ hold744/X _5540_/A1 _4007_/S VGND VGND VPWR VPWR _4007_/X sky130_fd_sc_hd__mux2_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5958_ _5968_/A _5981_/A _5979_/C VGND VGND VPWR VPWR _5958_/X sky130_fd_sc_hd__and3_4
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4909_ _4969_/A _5051_/B VGND VGND VPWR VPWR _4909_/Y sky130_fd_sc_hd__nand2_1
X_5889_ _6458_/Q _5645_/X _5646_/X _6653_/Q _5888_/X VGND VGND VPWR VPWR _5896_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold53/X VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__buf_12
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__buf_12
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_5 _5310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3240_ _6415_/Q _3264_/B VGND VGND VPWR VPWR _3867_/B sky130_fd_sc_hd__nand2_2
XFILLER_140_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3171_ _6487_/Q VGND VGND VPWR VPWR _3837_/B sky130_fd_sc_hd__inv_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6930_ _7006_/CLK _6930_/D fanout457/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6861_ _6951_/CLK _6861_/D fanout474/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_6_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7036_/CLK sky130_fd_sc_hd__clkbuf_16
X_5812_ _7001_/Q _5643_/X _5664_/X _6929_/Q VGND VGND VPWR VPWR _5812_/X sky130_fd_sc_hd__a22o_2
X_6792_ _7054_/CLK _6792_/D fanout461/X VGND VGND VPWR VPWR _6792_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5743_ _6902_/Q _5621_/X _5658_/X _6886_/Q VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5674_ _6963_/Q _5642_/X _5928_/A2 _6835_/Q _5673_/X VGND VGND VPWR VPWR _5681_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4625_ _4625_/A _4625_/B VGND VGND VPWR VPWR _4969_/B sky130_fd_sc_hd__nor2_1
Xhold500 _4260_/X VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold511 _6807_/Q VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _4556_/A _4562_/A _4972_/A VGND VGND VPWR VPWR _4557_/A sky130_fd_sc_hd__and3_1
Xhold522 _5434_/X VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _6479_/Q VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3573_/A _3571_/B VGND VGND VPWR VPWR _4292_/A sky130_fd_sc_hd__nor2_2
Xhold544 _5525_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _6539_/Q VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold566 _7155_/Q VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _4561_/B _4993_/A VGND VGND VPWR VPWR _4582_/B sky130_fd_sc_hd__nor2_1
Xhold577 _5408_/X VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold588 _7027_/Q VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ _6221_/X _6226_/B _6226_/C _6226_/D VGND VGND VPWR VPWR _6226_/X sky130_fd_sc_hd__and4b_1
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3438_ _7069_/Q _5523_/A _5328_/A _6896_/Q VGND VGND VPWR VPWR _3438_/X sky130_fd_sc_hd__a22o_1
Xhold599 _5509_/X VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6929_/Q _5938_/X _5952_/X _6961_/Q VGND VGND VPWR VPWR _6157_/X sky130_fd_sc_hd__a22o_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _5410_/X VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3369_ _3373_/B hold75/X VGND VGND VPWR VPWR _5463_/A sky130_fd_sc_hd__nor2_8
Xhold1211 _7010_/Q VGND VGND VPWR VPWR _5464_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 _5437_/X VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5108_ _5108_/A _5108_/B _5108_/C VGND VGND VPWR VPWR _5135_/B sky130_fd_sc_hd__and3_1
Xhold1233 _7079_/Q VGND VGND VPWR VPWR _5542_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ _6982_/Q _5945_/X _5975_/C _6838_/Q _6087_/X VGND VGND VPWR VPWR _6089_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1244 _4257_/X VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 _6645_/Q VGND VGND VPWR VPWR _4245_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _4215_/X VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1277 _6742_/Q VGND VGND VPWR VPWR _5155_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5039_ _5039_/A _5039_/B _5039_/C _5039_/D VGND VGND VPWR VPWR _5122_/A sky130_fd_sc_hd__and4_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 _4009_/X VGND VGND VPWR VPWR _6450_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _6737_/Q VGND VGND VPWR VPWR _5149_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR _3900_/C sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_cyc_i VGND VGND VPWR VPWR _3899_/C sky130_fd_sc_hd__clkbuf_1
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6333_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6338_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4410_ _4498_/A _4459_/B VGND VGND VPWR VPWR _4948_/A sky130_fd_sc_hd__nand2_4
X_5390_ hold658/X _5513_/A1 _5390_/S VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__mux2_1
X_4341_ _4753_/A _4607_/A VGND VGND VPWR VPWR _4690_/A sky130_fd_sc_hd__nand2_8
XFILLER_160_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7060_ _7078_/CLK hold88/X fanout482/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_1
X_4272_ hold355/X _5494_/A1 _4273_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6011_ _6971_/Q _5947_/X _5965_/X _6795_/Q _6010_/X VGND VGND VPWR VPWR _6014_/B
+ sky130_fd_sc_hd__a221o_2
X_3223_ _6543_/Q VGND VGND VPWR VPWR _3223_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6913_ _6969_/CLK _6913_/D fanout475/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_1
X_6844_ _6884_/CLK _6844_/D fanout475/X VGND VGND VPWR VPWR _6844_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3987_ hold630/X _5469_/A1 _3989_/S VGND VGND VPWR VPWR _3987_/X sky130_fd_sc_hd__mux2_1
X_6775_ _6777_/CLK hold92/X fanout483/X VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__dfrtp_1
X_5726_ _6901_/Q _5621_/X _5648_/X _6853_/Q _5725_/X VGND VGND VPWR VPWR _5726_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5657_ _5664_/A _5657_/B _5660_/C VGND VGND VPWR VPWR _5657_/X sky130_fd_sc_hd__and3b_2
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4608_ _4607_/A _4753_/B VGND VGND VPWR VPWR _4608_/X sky130_fd_sc_hd__and2b_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ _6508_/Q _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5594_/A sky130_fd_sc_hd__and3_1
XFILLER_163_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold330 _5336_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold341 _6785_/Q VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _4591_/A _4552_/A _4549_/A VGND VGND VPWR VPWR _4959_/B sky130_fd_sc_hd__and3_2
XFILLER_190_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold352 _4024_/X VGND VGND VPWR VPWR _6463_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold363 _6948_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _4332_/X VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _6996_/Q VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold396 _5201_/X VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6209_ _6556_/Q _5971_/B _5949_/X _6676_/Q _6208_/X VGND VGND VPWR VPWR _6225_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7189_ _7189_/A VGND VGND VPWR VPWR _7189_/X sky130_fd_sc_hd__clkbuf_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1030 _4028_/X VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 _6780_/Q VGND VGND VPWR VPWR _5205_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1052 _5172_/X VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1063 _6893_/Q VGND VGND VPWR VPWR _5332_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 _4211_/X VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 _7021_/Q VGND VGND VPWR VPWR _5476_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1096 _4099_/X VGND VGND VPWR VPWR _6516_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_71_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6926_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3910_ _3910_/A _3910_/B VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__nand2_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4890_ _4542_/A _4496_/Y _4892_/B _4381_/Y _4697_/Y VGND VGND VPWR VPWR _4895_/B
+ sky130_fd_sc_hd__o221a_1
X_3841_ _3837_/B _3867_/B _3840_/X _3860_/B VGND VGND VPWR VPWR _3866_/S sky130_fd_sc_hd__o31a_4
XFILLER_32_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3772_ _6540_/Q _4127_/A _3769_/X _3771_/X VGND VGND VPWR VPWR _3773_/C sky130_fd_sc_hd__a211o_1
X_6560_ _6653_/CLK _6560_/D fanout452/X VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5511_ hold403/X _5538_/A1 _5513_/S VGND VGND VPWR VPWR _5511_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6491_ _6527_/CLK _6491_/D fanout484/X VGND VGND VPWR VPWR _7182_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_157_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5442_ hold379/X _5538_/A1 _5444_/S VGND VGND VPWR VPWR _5442_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5373_ _5373_/A hold17/X VGND VGND VPWR VPWR _5381_/S sky130_fd_sc_hd__and2_4
XFILLER_114_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7112_ _7131_/CLK _7112_/D fanout459/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4324_ hold265/X _5534_/A1 _4327_/S VGND VGND VPWR VPWR _4324_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7043_ _7079_/CLK _7043_/D fanout478/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfrtp_4
X_4255_ _4255_/A0 hold60/X _4255_/S VGND VGND VPWR VPWR _4255_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3206_ _6925_/Q VGND VGND VPWR VPWR _3206_/Y sky130_fd_sc_hd__inv_2
X_4186_ _3410_/Y _4186_/A1 _4186_/S VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk _6888_/CLK VGND VGND VPWR VPWR _6969_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6827_ _6884_/CLK _6827_/D fanout475/X VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_51_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6758_ _6953_/CLK _6758_/D fanout460/X VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5709_ _6948_/Q _5637_/X _5660_/X _6804_/Q VGND VGND VPWR VPWR _5709_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6689_ _6707_/CLK _6689_/D fanout448/X VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold160 _6863_/Q VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _4074_/X VGND VGND VPWR VPWR _6500_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _7043_/Q VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold193 _4150_/X VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4040_ hold796/X _6354_/A1 _4043_/S VGND VGND VPWR VPWR _4040_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5991_ _7010_/Q _5940_/X _5947_/X _6970_/Q _5990_/X VGND VGND VPWR VPWR _5991_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_91_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4942_ _4942_/A _4942_/B _4942_/C VGND VGND VPWR VPWR _5071_/A sky130_fd_sc_hd__and3_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4873_ _4542_/A _4496_/Y _4700_/Y _4627_/B _4872_/X VGND VGND VPWR VPWR _4873_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6612_ _6671_/CLK _6612_/D _6383_/A VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3824_ _6768_/Q _5190_/A _5190_/B _4274_/A _6670_/Q VGND VGND VPWR VPWR _3824_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6543_ _6735_/CLK _6543_/D fanout445/X VGND VGND VPWR VPWR _6543_/Q sky130_fd_sc_hd__dfstp_2
X_3755_ _6427_/Q _3981_/A _4220_/A _6620_/Q _3754_/X VGND VGND VPWR VPWR _3760_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6474_ _6735_/CLK _6474_/D _3946_/B VGND VGND VPWR VPWR _6474_/Q sky130_fd_sc_hd__dfrtp_4
X_3686_ _6996_/Q _5445_/A _5211_/A _6788_/Q _3685_/X VGND VGND VPWR VPWR _3686_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_145_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput210 _3216_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
X_5425_ hold906/X _5548_/A1 _5426_/S VGND VGND VPWR VPWR _5425_/X sky130_fd_sc_hd__mux2_1
Xoutput221 _7184_/X VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput232 _7194_/X VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput243 _7176_/X VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
Xoutput254 _7198_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_5356_ _5356_/A0 hold667/X _5363_/S VGND VGND VPWR VPWR _5356_/X sky130_fd_sc_hd__mux2_1
Xoutput265 _6740_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
Xoutput276 _6432_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_160_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput287 _6748_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
X_4307_ hold956/X _6355_/A1 _4309_/S VGND VGND VPWR VPWR _4307_/X sky130_fd_sc_hd__mux2_1
Xoutput298 _6752_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
XFILLER_101_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5287_ hold912/X _5509_/A1 _5291_/S VGND VGND VPWR VPWR _5287_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7026_ _7026_/CLK _7026_/D fanout465/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfstp_2
X_4238_ _4238_/A _4322_/B VGND VGND VPWR VPWR _4243_/S sky130_fd_sc_hd__and2_2
XFILLER_87_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4169_ _3486_/Y _4169_/A1 _4171_/S VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire348 _3826_/Y VGND VGND VPWR VPWR _3827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout470 _6390_/A VGND VGND VPWR VPWR fanout470/X sky130_fd_sc_hd__buf_8
XFILLER_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout481 fanout485/X VGND VGND VPWR VPWR fanout481/X sky130_fd_sc_hd__buf_8
XFILLER_93_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3540_ _6918_/Q _5355_/A _6352_/A _7155_/Q VGND VGND VPWR VPWR _3540_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold907 _5425_/X VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 _6880_/Q VGND VGND VPWR VPWR hold918/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3471_ _6943_/Q _5382_/A _5274_/A _6847_/Q _3457_/X VGND VGND VPWR VPWR _3472_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold929 _5443_/X VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5210_ hold341/X _5540_/A1 _5210_/S VGND VGND VPWR VPWR _5210_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6190_ _6645_/Q _5976_/C _5971_/D _6565_/Q VGND VGND VPWR VPWR _6190_/X sky130_fd_sc_hd__a22o_1
X_5141_ _4542_/A _4946_/X _5058_/C _5140_/X VGND VGND VPWR VPWR _5142_/D sky130_fd_sc_hd__o211a_1
XFILLER_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5072_ _4565_/X _4741_/A _4650_/Y _5088_/C VGND VGND VPWR VPWR _5073_/C sky130_fd_sc_hd__o211a_1
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4023_ _4023_/A0 _6355_/A1 _4025_/S VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5974_ _5946_/X _5970_/X _5974_/C _5974_/D VGND VGND VPWR VPWR _5977_/A sky130_fd_sc_hd__and4bb_1
XFILLER_40_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4925_ _5088_/A _4925_/B _5114_/A VGND VGND VPWR VPWR _5103_/A sky130_fd_sc_hd__and3_1
XFILLER_21_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4856_ _4856_/A _4911_/B VGND VGND VPWR VPWR _4856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3807_ _3807_/A _3807_/B _3807_/C _3807_/D VGND VGND VPWR VPWR _3827_/B sky130_fd_sc_hd__nor4_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4787_ _4644_/Y _4714_/X _4782_/Y VGND VGND VPWR VPWR _4791_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6526_ _6527_/CLK hold7/X fanout484/X VGND VGND VPWR VPWR _6526_/Q sky130_fd_sc_hd__dfrtp_1
X_3738_ _6651_/Q _4250_/A _4133_/A _6546_/Q VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__a22o_2
XFILLER_109_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6457_ _6747_/CLK _6457_/D fanout447/X VGND VGND VPWR VPWR _6457_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_118_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3669_ _6940_/Q _5382_/A _4172_/A _6580_/Q _3668_/X VGND VGND VPWR VPWR _3670_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5408_ hold576/X _5513_/A1 _5408_/S VGND VGND VPWR VPWR _5408_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6388_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6388_/X sky130_fd_sc_hd__and2_1
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5339_ hold618/X _5543_/A1 _5345_/S VGND VGND VPWR VPWR _5339_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7017_/CLK _7009_/D fanout461/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4710_/A _4969_/B VGND VGND VPWR VPWR _4710_/Y sky130_fd_sc_hd__nand2_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _5690_/A _5690_/B _5690_/C _5690_/D VGND VGND VPWR VPWR _5690_/Y sky130_fd_sc_hd__nor4_1
XFILLER_187_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4641_ _4739_/A _4661_/B VGND VGND VPWR VPWR _4673_/B sky130_fd_sc_hd__nand2_2
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4572_ _4672_/A _4947_/B VGND VGND VPWR VPWR _4574_/B sky130_fd_sc_hd__nor2_2
XFILLER_175_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold704 _6839_/Q VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__dlygate4sd3_1
X_6311_ _3640_/Y _6311_/A1 _6315_/S VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__mux2_1
X_3523_ _3523_/A _3523_/B _3523_/C _3523_/D VGND VGND VPWR VPWR _3582_/B sky130_fd_sc_hd__nor4_1
Xhold715 _5254_/X VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 _6999_/Q VGND VGND VPWR VPWR hold726/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold737 _4161_/X VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold748 _6698_/Q VGND VGND VPWR VPWR hold748/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold759 _4131_/X VGND VGND VPWR VPWR _6543_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6242_ _6652_/Q _5973_/A _5948_/X _6697_/Q _6241_/X VGND VGND VPWR VPWR _6242_/X
+ sky130_fd_sc_hd__a221o_1
X_3454_ _3454_/A _3454_/B VGND VGND VPWR VPWR _3577_/B sky130_fd_sc_hd__nand2_8
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3385_ _6945_/Q _5382_/A _5436_/A _6993_/Q VGND VGND VPWR VPWR _3385_/X sky130_fd_sc_hd__a22o_1
X_6173_ _6817_/Q _5971_/B _5949_/X _6937_/Q _6172_/X VGND VGND VPWR VPWR _6175_/C
+ sky130_fd_sc_hd__a221o_1
X_5124_ _4672_/B _4496_/Y _4810_/A VGND VGND VPWR VPWR _5124_/X sky130_fd_sc_hd__a21o_1
Xhold1404 _6469_/Q VGND VGND VPWR VPWR _4031_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1415 _6573_/Q VGND VGND VPWR VPWR hold1415/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1426 _6584_/Q VGND VGND VPWR VPWR hold1426/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 _6592_/Q VGND VGND VPWR VPWR _4189_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5055_ _4413_/Y _4496_/Y _5092_/B _5054_/X VGND VGND VPWR VPWR _5056_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1448 _7137_/Q VGND VGND VPWR VPWR _6312_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _6732_/Q VGND VGND VPWR VPWR _3488_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4006_ hold892/X _5548_/A1 _4007_/S VGND VGND VPWR VPWR _4006_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5957_ _5969_/A _5968_/A _5969_/C VGND VGND VPWR VPWR _5975_/A sky130_fd_sc_hd__and3_4
X_4908_ _4845_/X _4907_/X _4465_/B VGND VGND VPWR VPWR _4915_/B sky130_fd_sc_hd__o21ai_1
XFILLER_178_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5888_ _7154_/Q _5625_/X _5642_/X _6718_/Q VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4839_ _5068_/A _4964_/B _5039_/C _4838_/X _4541_/X VGND VGND VPWR VPWR _4839_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_166_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6509_ _7131_/CLK _6509_/D fanout460/X VGND VGND VPWR VPWR _6509_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3224__1 net399_2/A VGND VGND VPWR VPWR _7157_/CLK sky130_fd_sc_hd__inv_2
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__buf_8
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__buf_8
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_6 _5310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3170_ _6635_/Q VGND VGND VPWR VPWR _3170_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6860_ _7079_/CLK _6860_/D fanout478/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5811_ _6937_/Q _5654_/X _5808_/X _5809_/X _5810_/X VGND VGND VPWR VPWR _5811_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_179_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6791_ _6953_/CLK _6791_/D fanout459/X VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtp_4
X_5742_ _6870_/Q _5628_/X _5634_/X _6974_/Q _5741_/X VGND VGND VPWR VPWR _5748_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5673_ _6947_/Q _5637_/X _5638_/X _6955_/Q VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4624_ _4620_/Y _4645_/B VGND VGND VPWR VPWR _4942_/B sky130_fd_sc_hd__nand2b_1
XFILLER_163_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold501 _6602_/Q VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlygate4sd3_1
X_4555_ _4724_/A _4650_/A VGND VGND VPWR VPWR _5088_/C sky130_fd_sc_hd__nand2_2
Xhold512 _5235_/X VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _6441_/Q VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _4043_/X VGND VGND VPWR VPWR _6479_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _6747_/Q VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _3554_/A _3692_/A VGND VGND VPWR VPWR _4250_/A sky130_fd_sc_hd__nor2_8
Xhold556 _4126_/X VGND VGND VPWR VPWR _6539_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4486_ _4690_/B _4626_/B VGND VGND VPWR VPWR _4689_/A sky130_fd_sc_hd__nand2_8
Xhold567 _6357_/X VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _6699_/Q VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _6225_/A _6225_/B _6225_/C _6225_/D VGND VGND VPWR VPWR _6225_/Y sky130_fd_sc_hd__nor4_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold589 _5483_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3437_ _6912_/Q _5346_/A _3432_/X _3434_/X _3436_/X VGND VGND VPWR VPWR _3437_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_103_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3368_ _3543_/A hold85/X VGND VGND VPWR VPWR _5373_/A sky130_fd_sc_hd__nor2_8
X_6156_ _7086_/Q _5976_/B _5971_/C _7046_/Q VGND VGND VPWR VPWR _6156_/X sky130_fd_sc_hd__a22o_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _6786_/Q VGND VGND VPWR VPWR _5212_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _5464_/X VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 _6954_/Q VGND VGND VPWR VPWR _5401_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5107_ _4611_/Y _4644_/Y _4663_/Y _4969_/Y VGND VGND VPWR VPWR _5108_/C sky130_fd_sc_hd__o22a_1
XFILLER_57_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1234 _5542_/X VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6087_ _6926_/Q _5938_/X _5952_/X _6958_/Q VGND VGND VPWR VPWR _6087_/X sky130_fd_sc_hd__a22o_1
X_3299_ _3347_/A hold72/X VGND VGND VPWR VPWR _3311_/C sky130_fd_sc_hd__nor2_2
XFILLER_73_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1245 _6660_/Q VGND VGND VPWR VPWR _4263_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _4245_/X VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 _6890_/Q VGND VGND VPWR VPWR _5329_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _5155_/X VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5038_ _5114_/B _5115_/A _5038_/C VGND VGND VPWR VPWR _5038_/X sky130_fd_sc_hd__and3_1
XFILLER_73_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1289 _6675_/Q VGND VGND VPWR VPWR _4281_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6989_ _7082_/CLK _6989_/D fanout480/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4556_/A sky130_fd_sc_hd__buf_8
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4625_/A sky130_fd_sc_hd__clkbuf_2
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6323_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6327_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6329_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6316_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4340_ _4753_/A _4607_/A VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__and2_4
XFILLER_141_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4271_ _4271_/A0 _6355_/A1 _4273_/S VGND VGND VPWR VPWR _4271_/X sky130_fd_sc_hd__mux2_1
X_3222_ _6789_/Q VGND VGND VPWR VPWR _3222_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6010_ _6891_/Q _5946_/X _5955_/X _6803_/Q VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6912_ _6951_/CLK _6912_/D fanout474/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6843_ _7067_/CLK _6843_/D fanout477/X VGND VGND VPWR VPWR _6843_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6774_ _7082_/CLK _6774_/D fanout483/X VGND VGND VPWR VPWR _7193_/A sky130_fd_sc_hd__dfrtp_1
X_3986_ hold620/X _6357_/A1 _3989_/S VGND VGND VPWR VPWR _3986_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5725_ _6869_/Q _5628_/X _5658_/X _6885_/Q VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5656_ _6930_/Q _5654_/X _5655_/X _6794_/Q _5653_/X VGND VGND VPWR VPWR _5669_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4607_ _4607_/A _4970_/A VGND VGND VPWR VPWR _4673_/A sky130_fd_sc_hd__nand2_8
X_5587_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5968_/A sky130_fd_sc_hd__and2_2
XFILLER_117_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold320 _5521_/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _6905_/Q VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__dlygate4sd3_1
X_4538_ _4424_/Y _4500_/Y _4504_/X _4537_/Y _5023_/A VGND VGND VPWR VPWR _4538_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_116_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold342 _5210_/X VGND VGND VPWR VPWR _6785_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _7012_/Q VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold364 _5394_/X VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold375 _6515_/Q VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold386 _5448_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4469_ _4469_/A _4672_/A VGND VGND VPWR VPWR _4472_/A sky130_fd_sc_hd__nor2_1
Xhold397 _7078_/Q VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _7035_/Q _5601_/X _5959_/X _6716_/Q VGND VGND VPWR VPWR _6208_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7188_ _7188_/A VGND VGND VPWR VPWR _7188_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _6984_/Q _5945_/X _5975_/C _6840_/Q _6138_/X VGND VGND VPWR VPWR _6140_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 _4135_/X VGND VGND VPWR VPWR _6546_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 _6451_/Q VGND VGND VPWR VPWR _4010_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1042 _5205_/X VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 _6447_/Q VGND VGND VPWR VPWR _4005_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1064 _5332_/X VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1075 _6909_/Q VGND VGND VPWR VPWR _5350_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 _5476_/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_204 _5971_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _6949_/Q VGND VGND VPWR VPWR _5395_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6632_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3840_ _7167_/Q _3875_/C _6485_/Q VGND VGND VPWR VPWR _3840_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3771_ _6794_/Q _3326_/Y _4032_/A _6470_/Q _3770_/X VGND VGND VPWR VPWR _3771_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5510_ hold483/X _5528_/A1 _5513_/S VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6490_ _6527_/CLK _6490_/D fanout481/X VGND VGND VPWR VPWR _7181_/A sky130_fd_sc_hd__dfrtp_1
X_5441_ hold439/X _5528_/A1 _5444_/S VGND VGND VPWR VPWR _5441_/X sky130_fd_sc_hd__mux2_1
X_5372_ hold654/X _5513_/A1 _5372_/S VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__mux2_1
X_7111_ _7131_/CLK _7111_/D fanout459/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4323_ _4323_/A0 hold667/X _4327_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7042_ _7086_/CLK _7042_/D fanout483/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_4
X_4254_ hold389/X _5494_/A1 _4255_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3205_ _6933_/Q VGND VGND VPWR VPWR _3205_/Y sky130_fd_sc_hd__inv_2
X_4185_ _3447_/Y _4185_/A1 _4186_/S VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6826_ _6908_/CLK _6826_/D fanout475/X VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_168_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6757_ _6953_/CLK _6757_/D fanout460/X VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3969_ hold1/X hold4/X _3975_/S VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__mux2_8
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5708_ _6836_/Q _5928_/A2 _5697_/X _5707_/X VGND VGND VPWR VPWR _5711_/B sky130_fd_sc_hd__a211o_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6688_ _6707_/CLK _6688_/D fanout448/X VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5639_ _6946_/Q _5637_/X _5638_/X _6954_/Q _5636_/X VGND VGND VPWR VPWR _5639_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold150 _5389_/X VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold161 _5298_/X VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _7148_/Q VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold183 _5501_/X VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _6678_/Q VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5990_ _6938_/Q _5961_/X _5976_/D _6874_/Q VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4941_ _4996_/C _4941_/B _5073_/B _4941_/D VGND VGND VPWR VPWR _4941_/X sky130_fd_sc_hd__and4_1
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4872_ _4872_/A _4872_/B _4872_/C _4872_/D VGND VGND VPWR VPWR _4872_/X sky130_fd_sc_hd__and4_1
XFILLER_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6611_ _6668_/CLK _6611_/D fanout452/X VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfstp_2
X_3823_ _6655_/Q _4256_/A _4172_/A _6578_/Q _3822_/X VGND VGND VPWR VPWR _3826_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6542_ _6709_/CLK _6542_/D fanout445/X VGND VGND VPWR VPWR _6542_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3754_ _6811_/Q _5238_/A hold67/A _6466_/Q VGND VGND VPWR VPWR _3754_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6473_ _6704_/CLK _6473_/D fanout448/X VGND VGND VPWR VPWR _6473_/Q sky130_fd_sc_hd__dfrtp_1
X_3685_ _6852_/Q _5283_/A _4208_/A _6611_/Q VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5424_ hold882/X _5538_/A1 _5426_/S VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput200 _3191_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput211 _3215_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _3932_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput233 _7174_/X VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
Xoutput244 _7177_/X VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
X_5355_ _5355_/A _5541_/B VGND VGND VPWR VPWR _5363_/S sky130_fd_sc_hd__and2_4
XFILLER_160_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput255 _3950_/A VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
Xoutput266 _6741_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput277 _6433_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
X_4306_ hold818/X _6354_/A1 _4309_/S VGND VGND VPWR VPWR _4306_/X sky130_fd_sc_hd__mux2_1
Xoutput288 _6749_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
Xoutput299 _6753_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
XFILLER_102_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5286_ hold333/X _5526_/A1 _5291_/S VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7025_ _7086_/CLK hold31/X fanout484/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4237_ hold842/X _5546_/A1 _4237_/S VGND VGND VPWR VPWR _4237_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4168_ _6312_/A0 _4168_/A1 _4171_/S VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4099_ _4099_/A0 _4098_/X _4101_/S VGND VGND VPWR VPWR _4099_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6809_ _7078_/CLK _6809_/D fanout481/X VGND VGND VPWR VPWR _6809_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire349 _3670_/Y VGND VGND VPWR VPWR _3699_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7037_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout460 fanout462/X VGND VGND VPWR VPWR fanout460/X sky130_fd_sc_hd__buf_6
XFILLER_120_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout471 _6396_/A VGND VGND VPWR VPWR _6390_/A sky130_fd_sc_hd__buf_6
Xfanout482 fanout485/X VGND VGND VPWR VPWR fanout482/X sky130_fd_sc_hd__buf_8
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6884_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_csclk _6888_/CLK VGND VGND VPWR VPWR _7070_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold908 _6808_/Q VGND VGND VPWR VPWR hold908/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 _5317_/X VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3470_ _6839_/Q _5265_/A _5463_/A _7015_/Q _3458_/X VGND VGND VPWR VPWR _3472_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5140_ _4542_/D _4672_/B _4518_/C _4821_/X VGND VGND VPWR VPWR _5140_/X sky130_fd_sc_hd__o211a_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5071_ _5071_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _5077_/A sky130_fd_sc_hd__and3_1
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4022_ _4022_/A0 _5492_/A1 _4025_/S VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5973_ _5973_/A _5973_/B VGND VGND VPWR VPWR _5974_/D sky130_fd_sc_hd__nor2_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4924_ _4456_/Y _4562_/Y _4673_/A _4689_/B _4768_/C VGND VGND VPWR VPWR _4999_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4855_ _4782_/A _4630_/X _4515_/Y VGND VGND VPWR VPWR _4855_/Y sky130_fd_sc_hd__a21oi_1
X_3806_ _6680_/Q _4286_/A _3585_/Y input98/X _3805_/X VGND VGND VPWR VPWR _3807_/D
+ sky130_fd_sc_hd__a221o_1
X_4786_ _4673_/A _4689_/B _4781_/X _5108_/B _4785_/X VGND VGND VPWR VPWR _4791_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_165_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6525_ _6527_/CLK _6525_/D fanout484/X VGND VGND VPWR VPWR _6525_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3737_ _7048_/Q _5505_/A _5274_/A _6843_/Q _3736_/X VGND VGND VPWR VPWR _3742_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_180_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6456_ _6704_/CLK _6456_/D fanout447/X VGND VGND VPWR VPWR _6456_/Q sky130_fd_sc_hd__dfrtp_2
X_3668_ _6462_/Q _4020_/A _4328_/A _6717_/Q VGND VGND VPWR VPWR _3668_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5407_ hold137/X hold99/X _5408_/S VGND VGND VPWR VPWR _5407_/X sky130_fd_sc_hd__mux2_1
X_6387_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6387_/X sky130_fd_sc_hd__and2_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3599_ _6683_/Q _4286_/A _4268_/A _6668_/Q _3598_/X VGND VGND VPWR VPWR _3604_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5338_ _5338_/A0 hold667/X _5345_/S VGND VGND VPWR VPWR _5338_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5269_ hold223/X _5494_/A1 _5273_/S VGND VGND VPWR VPWR _5269_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7008_ _7033_/CLK _7008_/D fanout464/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4640_ _4673_/A _4626_/Y _4639_/Y VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__a21o_1
XFILLER_175_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4571_ _4496_/Y _4570_/Y _5099_/A _4559_/X _4548_/X VGND VGND VPWR VPWR _4589_/C
+ sky130_fd_sc_hd__o2111a_1
X_6310_ _3700_/Y _6310_/A1 _6315_/S VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__mux2_1
Xhold705 _5271_/X VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3522_ _6838_/Q _5265_/A _3381_/Y input30/X _3521_/X VGND VGND VPWR VPWR _3523_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold716 _6872_/Q VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 _5451_/X VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold738 _6873_/Q VGND VGND VPWR VPWR hold738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 _4308_/X VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6241_ _6647_/Q _5976_/C _5971_/D _6567_/Q VGND VGND VPWR VPWR _6241_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3453_ _3453_/A hold64/X _3454_/A VGND VGND VPWR VPWR _5164_/B sky130_fd_sc_hd__and3_4
XFILLER_131_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6172_ _6449_/Q _5601_/X _5959_/X _6969_/Q VGND VGND VPWR VPWR _6172_/X sky130_fd_sc_hd__a22o_1
X_3384_ _7033_/Q hold49/A _5505_/A _7054_/Q VGND VGND VPWR VPWR _3384_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5123_ _5123_/A VGND VGND VPWR VPWR _5123_/Y sky130_fd_sc_hd__inv_2
Xhold1405 _6963_/Q VGND VGND VPWR VPWR _5411_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _6575_/Q VGND VGND VPWR VPWR hold1416/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1427 _6588_/Q VGND VGND VPWR VPWR hold1427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 _6594_/Q VGND VGND VPWR VPWR _4191_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5054_ _4413_/Y _4672_/B _5057_/A _5057_/B VGND VGND VPWR VPWR _5054_/X sky130_fd_sc_hd__o211a_1
Xhold1449 _6722_/Q VGND VGND VPWR VPWR _4988_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_4005_ _4005_/A0 _5469_/A1 _4007_/S VGND VGND VPWR VPWR _4005_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5956_ _5978_/A _5964_/A _5969_/C VGND VGND VPWR VPWR _5976_/C sky130_fd_sc_hd__and3_4
X_4907_ _4887_/B _4907_/B VGND VGND VPWR VPWR _4907_/X sky130_fd_sc_hd__and2b_1
X_5887_ _5887_/A1 _6279_/S _5885_/X _5886_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__o22a_1
XFILLER_21_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4838_ _4453_/B _4570_/Y _4837_/X _4925_/B VGND VGND VPWR VPWR _4838_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4769_ _4769_/A _4999_/A _4769_/C _4769_/D VGND VGND VPWR VPWR _4770_/D sky130_fd_sc_hd__and4_1
XFILLER_147_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6508_ _7113_/CLK _6508_/D fanout460/X VGND VGND VPWR VPWR _6508_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6439_ _6747_/CLK _6439_/D fanout447/X VGND VGND VPWR VPWR _6439_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__buf_6
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_7 _5391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5810_ _6873_/Q _5628_/X _5658_/X _6889_/Q _5801_/X VGND VGND VPWR VPWR _5810_/X
+ sky130_fd_sc_hd__a221o_2
X_6790_ _7006_/CLK _6790_/D fanout457/X VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5741_ _6982_/Q _5624_/X _5654_/X _6934_/Q VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__a22o_1
X_5672_ _5672_/A1 _6103_/B1 _5670_/Y _5671_/X VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4623_ _4653_/B _4638_/A VGND VGND VPWR VPWR _4623_/Y sky130_fd_sc_hd__nand2_2
XFILLER_175_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4554_ _4574_/A _4554_/B VGND VGND VPWR VPWR _4559_/B sky130_fd_sc_hd__nand2_1
Xhold502 _4200_/X VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold513 _6871_/Q VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _3998_/X VGND VGND VPWR VPWR _6441_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ hold74/X _3562_/B VGND VGND VPWR VPWR _4044_/A sky130_fd_sc_hd__nor2_4
Xhold535 _6883_/Q VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _5160_/X VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4485_ _4690_/B _4626_/B VGND VGND VPWR VPWR _4911_/B sky130_fd_sc_hd__and2_4
Xhold557 hold557/A VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold568 _6926_/Q VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _4309_/X VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _6456_/Q _5944_/X _5975_/A _6600_/Q _6205_/X VGND VGND VPWR VPWR _6225_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3436_ _7000_/Q _5445_/A _3964_/A _6424_/Q _3435_/X VGND VGND VPWR VPWR _3436_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_131_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _7033_/Q _5944_/X _5975_/A _6849_/Q VGND VGND VPWR VPWR _6155_/X sky130_fd_sc_hd__a22o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3370_/A _3511_/A VGND VGND VPWR VPWR _3367_/Y sky130_fd_sc_hd__nor2_8
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1202 _5212_/X VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5106_/A _5106_/B _5106_/C _5106_/D VGND VGND VPWR VPWR _5109_/B sky130_fd_sc_hd__and4_1
Xhold1213 _6994_/Q VGND VGND VPWR VPWR _5446_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1224 _5401_/X VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6086_ _6974_/Q _5947_/X _5965_/X _6798_/Q _6085_/X VGND VGND VPWR VPWR _6089_/B
+ sky130_fd_sc_hd__a221o_1
X_3298_ _3975_/S hold71/X _3298_/B1 VGND VGND VPWR VPWR _3298_/Y sky130_fd_sc_hd__o21ai_2
Xhold1235 _6619_/Q VGND VGND VPWR VPWR _4221_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1246 _4263_/X VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 _6475_/Q VGND VGND VPWR VPWR _4039_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5037_ _5114_/C _5086_/C _5037_/C _5115_/B VGND VGND VPWR VPWR _5038_/C sky130_fd_sc_hd__nand4_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1268 _5329_/X VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _6460_/Q VGND VGND VPWR VPWR _4021_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6988_ _7049_/CLK _6988_/D fanout456/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5939_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5981_/C sky130_fd_sc_hd__nor2_4
XFILLER_179_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4566_/A sky130_fd_sc_hd__clkbuf_4
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6330_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6336_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6341_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6319_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ _4270_/A0 _5492_/A1 _4273_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3221_ _6797_/Q VGND VGND VPWR VPWR _3221_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6911_ _6967_/CLK _6911_/D fanout474/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6842_ _7026_/CLK _6842_/D fanout463/X VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6773_ _6777_/CLK _6773_/D fanout479/X VGND VGND VPWR VPWR _7192_/A sky130_fd_sc_hd__dfrtp_1
X_3985_ hold770/X _6356_/A1 _3989_/S VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5724_ _6997_/Q _5643_/X _5667_/X _6813_/Q VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5655_ _5638_/A _5667_/C _5666_/C VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__and3b_4
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4606_ _4607_/A _4970_/A VGND VGND VPWR VPWR _4975_/A sky130_fd_sc_hd__and2_2
XFILLER_175_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5586_ _5586_/A VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__inv_2
Xhold310 _4224_/X VGND VGND VPWR VPWR _6622_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _6964_/Q VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4537_ _5068_/A _4925_/B _4537_/C _4537_/D VGND VGND VPWR VPWR _4537_/Y sky130_fd_sc_hd__nand4_1
XFILLER_190_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold332 _5345_/X VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _7004_/Q VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold354 _5466_/X VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _7195_/A VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold376 _4097_/X VGND VGND VPWR VPWR _6515_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ _4817_/A _4965_/B VGND VGND VPWR VPWR _5041_/A sky130_fd_sc_hd__nand2_2
Xhold387 _6956_/Q VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold398 _5540_/X VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _7152_/Q _5958_/X _5978_/X _6481_/Q VGND VGND VPWR VPWR _6207_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3419_ _6808_/Q _5229_/A hold86/A _7061_/Q VGND VGND VPWR VPWR _3419_/X sky130_fd_sc_hd__a22o_2
X_7187_ _7187_/A VGND VGND VPWR VPWR _7187_/X sky130_fd_sc_hd__clkbuf_1
X_4399_ _4551_/A _4813_/A VGND VGND VPWR VPWR _4459_/A sky130_fd_sc_hd__and2_2
XFILLER_98_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6928_/Q _5938_/X _5952_/X _6960_/Q VGND VGND VPWR VPWR _6138_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1010 _4252_/X VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 _6600_/Q VGND VGND VPWR VPWR _4198_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _4010_/X VGND VGND VPWR VPWR _6451_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1043 _6499_/Q VGND VGND VPWR VPWR _4072_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1054 _4005_/X VGND VGND VPWR VPWR _6447_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6069_ _6821_/Q _5953_/X _5960_/X _7074_/Q _6068_/X VGND VGND VPWR VPWR _6069_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1065 _7013_/Q VGND VGND VPWR VPWR _5467_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1076 _5350_/X VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _6989_/Q VGND VGND VPWR VPWR _5440_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_205 _3251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1098 _5395_/X VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3770_ _7010_/Q _5463_/A _4316_/A _6705_/Q VGND VGND VPWR VPWR _3770_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5440_ _5440_/A0 _5545_/A1 _5444_/S VGND VGND VPWR VPWR _5440_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5371_ hold114/X hold99/X _5372_/S VGND VGND VPWR VPWR _5371_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7110_ _7131_/CLK _7110_/D fanout456/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfrtp_1
X_4322_ _4322_/A _4322_/B VGND VGND VPWR VPWR _4327_/S sky130_fd_sc_hd__and2_2
XFILLER_99_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7041_ _7051_/CLK hold3/X fanout477/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_1
X_4253_ hold888/X _5493_/A1 _4255_/S VGND VGND VPWR VPWR _4253_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3204_ _6941_/Q VGND VGND VPWR VPWR _3204_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_79_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4184_ _3486_/Y _4184_/A1 _4186_/S VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _3937_/A1 sky130_fd_sc_hd__clkbuf_8
X_6825_ _7070_/CLK _6825_/D fanout473/X VGND VGND VPWR VPWR _6825_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3968_ hold247/X _5465_/A1 _3980_/S VGND VGND VPWR VPWR _3968_/X sky130_fd_sc_hd__mux2_1
X_6756_ _6769_/CLK _6756_/D fanout469/X VGND VGND VPWR VPWR _7173_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_149_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5707_ _6844_/Q _5902_/A2 _5905_/A2 _6796_/Q _5695_/X VGND VGND VPWR VPWR _5707_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6687_ _6707_/CLK _6687_/D fanout448/X VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_176_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3899_ input123/X input122/X _3899_/C _3899_/D VGND VGND VPWR VPWR _3901_/C sky130_fd_sc_hd__and4bb_1
XFILLER_109_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5638_ _5638_/A _5657_/B _5666_/C VGND VGND VPWR VPWR _5638_/X sky130_fd_sc_hd__and3_4
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5569_ _6508_/Q _5567_/Y _7092_/Q VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold140 _5218_/X VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _6958_/Q VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _3979_/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold184 _6902_/Q VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _4284_/X VGND VGND VPWR VPWR _6678_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4940_ _4948_/B _4562_/Y _4673_/A _4644_/Y _4738_/Y VGND VGND VPWR VPWR _4941_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4871_ _4947_/B _4456_/Y _4694_/Y _4627_/B VGND VGND VPWR VPWR _4872_/D sky130_fd_sc_hd__o22a_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6610_ _6668_/CLK _6610_/D _6400_/A VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_2
X_3822_ _6604_/Q _4202_/A _4262_/A _6660_/Q VGND VGND VPWR VPWR _3822_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6541_ _6709_/CLK _6541_/D fanout445/X VGND VGND VPWR VPWR _6541_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _6915_/Q _5355_/A hold49/A _7027_/Q _3752_/X VGND VGND VPWR VPWR _3760_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6472_ _6735_/CLK _6472_/D _3946_/B VGND VGND VPWR VPWR _6472_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3684_ input54/X _5193_/A _5229_/A _6804_/Q VGND VGND VPWR VPWR _3684_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5423_ hold437/X _5528_/A1 _5426_/S VGND VGND VPWR VPWR _5423_/X sky130_fd_sc_hd__mux2_1
Xoutput201 _3190_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 _3214_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
XFILLER_160_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput223 _7185_/X VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
Xoutput234 _7195_/X VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
X_5354_ hold675/X _5540_/A1 _5354_/S VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__mux2_1
Xoutput245 _3929_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
Xoutput256 _3950_/Y VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
Xoutput267 _6735_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
X_4305_ _4305_/A0 _5491_/A1 _4309_/S VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__mux2_1
Xoutput278 _6418_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
X_5285_ hold293/X _5465_/A1 _5291_/S VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__mux2_1
Xoutput289 _6436_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7024_ _7085_/CLK _7024_/D fanout482/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_2
X_4236_ hold361/X _5518_/A1 _4237_/S VGND VGND VPWR VPWR _4236_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4167_ _3640_/Y _4167_/A1 _4171_/S VGND VGND VPWR VPWR _6573_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4098_ hold291/X _5548_/A1 _5202_/B VGND VGND VPWR VPWR _4098_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_csclk clkbuf_leaf_4_csclk/A VGND VGND VPWR VPWR _6654_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6808_ _7085_/CLK _6808_/D fanout482/X VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6739_ _6739_/CLK _6739_/D _3946_/B VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout450 fanout486/X VGND VGND VPWR VPWR fanout450/X sky130_fd_sc_hd__buf_8
Xfanout461 fanout462/X VGND VGND VPWR VPWR fanout461/X sky130_fd_sc_hd__buf_8
XFILLER_59_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout472 fanout486/X VGND VGND VPWR VPWR _6396_/A sky130_fd_sc_hd__buf_6
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout483 fanout484/X VGND VGND VPWR VPWR fanout483/X sky130_fd_sc_hd__buf_8
XFILLER_171_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold909 _5236_/X VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5070_ _4542_/B _4428_/Y _4846_/B _4619_/Y _4771_/C VGND VGND VPWR VPWR _5071_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4021_ _4021_/A0 _6353_/A1 _4025_/S VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5972_ _5600_/A _5978_/A _5981_/B _5934_/X _5967_/X VGND VGND VPWR VPWR _5973_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4923_ _4921_/A _5043_/A _4747_/A _4747_/B _4740_/B VGND VGND VPWR VPWR _4923_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_178_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4854_ _4542_/B _4947_/B _4902_/B _4616_/Y VGND VGND VPWR VPWR _4877_/B sky130_fd_sc_hd__o22a_1
XFILLER_60_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3805_ _6834_/Q _5265_/A _4328_/A _6715_/Q VGND VGND VPWR VPWR _3805_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4785_ _4902_/B _4689_/B _4784_/X _4967_/A VGND VGND VPWR VPWR _4785_/X sky130_fd_sc_hd__o211a_1
X_3736_ _6676_/Q _4280_/A _4139_/A _6551_/Q VGND VGND VPWR VPWR _3736_/X sky130_fd_sc_hd__a22o_2
XFILLER_118_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6524_ _6527_/CLK _6524_/D fanout484/X VGND VGND VPWR VPWR _6524_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3667_ _7012_/Q _5463_/A _5182_/S _6759_/Q _3666_/X VGND VGND VPWR VPWR _3670_/C
+ sky130_fd_sc_hd__a221o_1
X_6455_ _6747_/CLK _6455_/D fanout447/X VGND VGND VPWR VPWR _6455_/Q sky130_fd_sc_hd__dfrtp_4
X_5406_ hold710/X _5469_/A1 _5408_/S VGND VGND VPWR VPWR _5406_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6386_ _6401_/A _6400_/B VGND VGND VPWR VPWR _6386_/X sky130_fd_sc_hd__and2_1
XFILLER_133_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3598_ input46/X hold37/A _5523_/A _7066_/Q VGND VGND VPWR VPWR _3598_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5337_ _5337_/A _5541_/B VGND VGND VPWR VPWR _5345_/S sky130_fd_sc_hd__and2_4
XFILLER_88_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5268_ hold369/X _5526_/A1 _5273_/S VGND VGND VPWR VPWR _5268_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7007_ _7017_/CLK _7007_/D fanout461/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_2
X_4219_ hold982/X _5546_/A1 _4219_/S VGND VGND VPWR VPWR _4219_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5199_ hold91/X hold42/X _5201_/S VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__mux2_1
XFILLER_56_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4570_ _4570_/A _4959_/B VGND VGND VPWR VPWR _4570_/Y sky130_fd_sc_hd__nand2_1
X_3521_ _7083_/Q _5541_/A _4172_/A _6582_/Q VGND VGND VPWR VPWR _3521_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold706 _6927_/Q VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 _5308_/X VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 _6740_/Q VGND VGND VPWR VPWR hold728/X sky130_fd_sc_hd__dlygate4sd3_1
X_6240_ _6240_/A _6240_/B _6240_/C VGND VGND VPWR VPWR _6240_/Y sky130_fd_sc_hd__nor3_1
X_3452_ _3714_/B _3562_/B VGND VGND VPWR VPWR _5154_/A sky130_fd_sc_hd__nor2_8
Xhold739 _5309_/X VGND VGND VPWR VPWR _6873_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6171_ _7025_/Q _5937_/X _5975_/D _6889_/Q _6155_/X VGND VGND VPWR VPWR _6175_/B
+ sky130_fd_sc_hd__a221o_1
X_3383_ _7025_/Q hold29/A _5409_/A _6969_/Q VGND VGND VPWR VPWR _3383_/X sky130_fd_sc_hd__a22o_2
XFILLER_130_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5122_ _5122_/A _5122_/B _5122_/C VGND VGND VPWR VPWR _5123_/A sky130_fd_sc_hd__and3_1
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1406 _5411_/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5053_ _4948_/A _4672_/B _4523_/Y _4824_/X _4953_/Y VGND VGND VPWR VPWR _5092_/B
+ sky130_fd_sc_hd__o2111a_1
Xhold1417 _7160_/Q VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1428 _6589_/Q VGND VGND VPWR VPWR hold1428/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 _6593_/Q VGND VGND VPWR VPWR _4190_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4004_ hold79/X _5519_/A1 _4007_/S VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__mux2_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5955_ _5978_/A _5981_/B _5969_/C VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__and3_4
X_4906_ _4381_/Y _4900_/Y _4869_/B VGND VGND VPWR VPWR _4906_/Y sky130_fd_sc_hd__o21ai_1
X_5886_ _5552_/B _7115_/Q _6103_/B1 VGND VGND VPWR VPWR _5886_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4837_ _5114_/A _5089_/A _5018_/A _4837_/D VGND VGND VPWR VPWR _4837_/X sky130_fd_sc_hd__and4_1
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4768_ _4768_/A _4768_/B _4768_/C _4768_/D VGND VGND VPWR VPWR _4769_/D sky130_fd_sc_hd__and4_1
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6507_ _7131_/CLK _6507_/D fanout460/X VGND VGND VPWR VPWR _6507_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3719_ _6443_/Q _3999_/A _5145_/A _6736_/Q _3718_/X VGND VGND VPWR VPWR _3720_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4699_ _4460_/A _4611_/B _4628_/Y _4967_/B _4625_/A VGND VGND VPWR VPWR _4706_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_134_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6438_ _6747_/CLK _6438_/D fanout447/X VGND VGND VPWR VPWR _6438_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_161_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6369_ _6383_/A _6396_/B VGND VGND VPWR VPWR _6369_/X sky130_fd_sc_hd__and2_1
XFILLER_96_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _6882_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__buf_6
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__buf_8
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7078_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 hold29/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5740_ _6990_/Q _5627_/X _5635_/X _6830_/Q VGND VGND VPWR VPWR _5740_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5671_ _6786_/Q _5652_/Y _5610_/Y VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__o21a_1
XFILLER_175_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4622_ _4653_/B _4638_/A VGND VGND VPWR VPWR _4645_/B sky130_fd_sc_hd__and2_2
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4553_ _4947_/C _4553_/B VGND VGND VPWR VPWR _4554_/B sky130_fd_sc_hd__nor2_1
XFILLER_144_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold503 _7030_/Q VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold514 _5307_/X VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _6649_/Q VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ _3504_/A _3504_/B _3504_/C _3504_/D VGND VGND VPWR VPWR _3504_/Y sky130_fd_sc_hd__nor4_1
XFILLER_116_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold536 _5321_/X VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _4562_/A _4972_/A VGND VGND VPWR VPWR _4484_/Y sky130_fd_sc_hd__nand2_1
Xhold547 _7190_/A VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold558 _7048_/Q VGND VGND VPWR VPWR hold558/X sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _6984_/Q _5427_/A _3381_/Y input32/X VGND VGND VPWR VPWR _3435_/X sky130_fd_sc_hd__a22o_1
Xhold569 _5369_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6681_/Q _5934_/X _5975_/B _6615_/Q _6222_/X VGND VGND VPWR VPWR _6225_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6178_/A0 _6153_/X _6304_/S VGND VGND VPWR VPWR _6154_/X sky130_fd_sc_hd__mux2_1
X_3366_ _3571_/A _3379_/A VGND VGND VPWR VPWR _5274_/A sky130_fd_sc_hd__nor2_8
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _6930_/Q VGND VGND VPWR VPWR _5374_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5105_ _4616_/Y _4970_/Y _5010_/Y _4613_/Y VGND VGND VPWR VPWR _5106_/D sky130_fd_sc_hd__o22a_1
Xhold1214 _5446_/X VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6085_ _6894_/Q _5946_/X _5955_/X _6806_/Q VGND VGND VPWR VPWR _6085_/X sky130_fd_sc_hd__a22o_1
Xhold1225 _6751_/Q VGND VGND VPWR VPWR _5167_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3297_ hold1003/X _3975_/S VGND VGND VPWR VPWR _3297_/Y sky130_fd_sc_hd__nand2b_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 _4221_/X VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 _6970_/Q VGND VGND VPWR VPWR _5419_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5036_ _4500_/A _4902_/B _4494_/Y _4882_/C _4909_/Y VGND VGND VPWR VPWR _5115_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_38_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1258 _4039_/X VGND VGND VPWR VPWR _6475_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1269 _6630_/Q VGND VGND VPWR VPWR _4239_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6987_ _7085_/CLK _6987_/D fanout477/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_41_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5938_ _5979_/A _5981_/A _5981_/B VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__and3_4
XFILLER_179_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5869_ _6697_/Q _5637_/X _5645_/X _6457_/Q VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4337_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4702_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__clkbuf_1
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6332_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6339_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6344_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6318_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3220_ _6805_/Q VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6910_ _7081_/CLK _6910_/D fanout478/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6841_ _6865_/CLK _6841_/D fanout464/X VGND VGND VPWR VPWR _6841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6772_ _7082_/CLK _6772_/D fanout479/X VGND VGND VPWR VPWR _7191_/A sky130_fd_sc_hd__dfrtp_1
X_3984_ hold993/X _6355_/A1 _3989_/S VGND VGND VPWR VPWR _3984_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5723_ _6981_/Q _5624_/X _5654_/X _6933_/Q _5717_/Y VGND VGND VPWR VPWR _5723_/X
+ sky130_fd_sc_hd__a221o_1
X_5654_ _5664_/A _5667_/C _5660_/C VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__and3_4
X_4605_ _4753_/A _4753_/B VGND VGND VPWR VPWR _4625_/B sky130_fd_sc_hd__nand2b_2
X_5585_ _5567_/Y _6508_/Q _7097_/Q VGND VGND VPWR VPWR _5586_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold300 _5429_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold311 _7046_/Q VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4536_ _5010_/A _4969_/A _4881_/B VGND VGND VPWR VPWR _4537_/D sky130_fd_sc_hd__o21ai_1
Xhold322 _5412_/X VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold333 _6852_/Q VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold344 _5457_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _6668_/Q VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _5200_/X VGND VGND VPWR VPWR _6776_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4467_ _4498_/A _4531_/B _4579_/B VGND VGND VPWR VPWR _5027_/A sky130_fd_sc_hd__nand3_1
Xhold377 _6683_/Q VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _5403_/X VGND VGND VPWR VPWR _6956_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold399 _6940_/Q VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _6610_/Q _5943_/X _5981_/X _6656_/Q VGND VGND VPWR VPWR _6206_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3418_ _7053_/Q _5505_/A _3367_/Y input27/X VGND VGND VPWR VPWR _3418_/X sky130_fd_sc_hd__a22o_1
X_7186_ _7186_/A VGND VGND VPWR VPWR _7186_/X sky130_fd_sc_hd__clkbuf_1
X_4398_ _4415_/A _4415_/B VGND VGND VPWR VPWR _4813_/A sky130_fd_sc_hd__and2b_1
Xhold1000 _4173_/X VGND VGND VPWR VPWR _6578_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6137_ _6976_/Q _5947_/X _5965_/X _6800_/Q _6136_/X VGND VGND VPWR VPWR _6140_/B
+ sky130_fd_sc_hd__a221o_1
X_3349_ hold75/A hold28/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__nor2_8
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _6610_/Q VGND VGND VPWR VPWR _4210_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1022 _4198_/X VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 _6615_/Q VGND VGND VPWR VPWR _4216_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _4072_/X VGND VGND VPWR VPWR _6499_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6068_ _6909_/Q _5973_/A _5948_/X _6949_/Q _6067_/X VGND VGND VPWR VPWR _6068_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1055 _7026_/Q VGND VGND VPWR VPWR _5482_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1066 _5467_/X VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 _6842_/Q VGND VGND VPWR VPWR _5275_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5019_ _5041_/B _4681_/Y _4710_/Y _4627_/A VGND VGND VPWR VPWR _5021_/D sky130_fd_sc_hd__a31o_1
Xhold1088 _5440_/X VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 _6802_/Q VGND VGND VPWR VPWR _5230_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_206 _5490_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5370_ hold706/X _5469_/A1 _5372_/S VGND VGND VPWR VPWR _5370_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4321_ hold580/X _6357_/A1 _4321_/S VGND VGND VPWR VPWR _4321_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4252_ _4252_/A0 _5492_/A1 _4255_/S VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7040_ _7081_/CLK _7040_/D fanout477/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_101_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3203_ _6949_/Q VGND VGND VPWR VPWR _3203_/Y sky130_fd_sc_hd__inv_2
X_4183_ _4192_/A0 _4183_/A1 _4186_/S VGND VGND VPWR VPWR _6587_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6824_ _6920_/CLK _6824_/D fanout473/X VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6755_ _6755_/CLK _6755_/D _6360_/A VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfrtp_1
X_3967_ hold8/X hold11/X _3975_/S VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__mux2_8
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5706_ _5706_/A _5706_/B _5706_/C _5706_/D VGND VGND VPWR VPWR _5706_/Y sky130_fd_sc_hd__nor4_4
XFILLER_176_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6686_ _6707_/CLK _6686_/D fanout448/X VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfrtp_4
X_3898_ _4334_/B _4334_/C VGND VGND VPWR VPWR _4702_/C sky130_fd_sc_hd__nor2_2
XFILLER_191_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5637_ _5664_/A _5658_/B _5657_/B VGND VGND VPWR VPWR _5637_/X sky130_fd_sc_hd__and3_4
XFILLER_164_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5568_ _6506_/Q _5610_/B VGND VGND VPWR VPWR _5568_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold130 _5180_/X VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold141 _6856_/Q VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ _4886_/B _4953_/A VGND VGND VPWR VPWR _4522_/B sky130_fd_sc_hd__nand2_1
Xhold152 _6998_/Q VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _5405_/X VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _5499_/A0 hold6/X hold77/A VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__mux2_1
Xhold174 hold21/X VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _5342_/X VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _6814_/Q VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7169_ _3945_/A1 _7169_/D _6399_/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4870_ _4870_/A _5027_/B _4870_/C VGND VGND VPWR VPWR _4872_/C sky130_fd_sc_hd__and3_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3821_ _6810_/Q _5238_/A _4208_/A _6609_/Q _3820_/X VGND VGND VPWR VPWR _3826_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6540_ _6735_/CLK _6540_/D fanout445/X VGND VGND VPWR VPWR _6540_/Q sky130_fd_sc_hd__dfrtp_2
X_3752_ _6995_/Q _5445_/A _5373_/A _6931_/Q VGND VGND VPWR VPWR _3752_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6471_ _6739_/CLK _6471_/D _3946_/B VGND VGND VPWR VPWR _6471_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3683_ _6482_/Q _4044_/A _4268_/A _6667_/Q _3682_/X VGND VGND VPWR VPWR _3688_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_173_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5422_ _5422_/A0 _5545_/A1 _5426_/S VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput202 _3189_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 _3933_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
XFILLER_173_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput224 _7186_/X VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
X_5353_ hold673/X _5521_/A1 _5354_/S VGND VGND VPWR VPWR _5353_/X sky130_fd_sc_hd__mux2_1
Xoutput235 _7196_/X VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
Xoutput246 _7178_/X VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
Xoutput257 _6745_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
X_4304_ _4304_/A _6352_/B VGND VGND VPWR VPWR _4309_/S sky130_fd_sc_hd__and2_2
Xoutput268 _6742_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
Xoutput279 _6419_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5284_ _5284_/A0 _5524_/A1 _5291_/S VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7023_ _7086_/CLK hold57/X fanout482/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__dfrtp_4
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4235_ hold461/X _5544_/A1 _4237_/S VGND VGND VPWR VPWR _4235_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4166_ _3700_/Y _4166_/A1 _4171_/S VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4097_ hold375/X _4096_/X _4101_/S VGND VGND VPWR VPWR _4097_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6807_ _7078_/CLK _6807_/D fanout481/X VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4999_ _4999_/A _4999_/B _4999_/C VGND VGND VPWR VPWR _5001_/B sky130_fd_sc_hd__and3_1
X_6738_ _6739_/CLK _6738_/D _3946_/B VGND VGND VPWR VPWR _6738_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6669_ _6677_/CLK _6669_/D fanout452/X VGND VGND VPWR VPWR _6669_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout440 _6396_/B VGND VGND VPWR VPWR _6400_/B sky130_fd_sc_hd__buf_6
Xfanout451 fanout452/X VGND VGND VPWR VPWR _6400_/A sky130_fd_sc_hd__buf_4
Xfanout462 fanout466/X VGND VGND VPWR VPWR fanout462/X sky130_fd_sc_hd__clkbuf_8
XFILLER_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout473 fanout474/X VGND VGND VPWR VPWR fanout473/X sky130_fd_sc_hd__buf_8
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout484 fanout485/X VGND VGND VPWR VPWR fanout484/X sky130_fd_sc_hd__buf_6
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4020_ _4020_/A _5490_/B VGND VGND VPWR VPWR _4025_/S sky130_fd_sc_hd__and2_2
XFILLER_77_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5971_ _5971_/A _5971_/B _5971_/C _5971_/D VGND VGND VPWR VPWR _5974_/C sky130_fd_sc_hd__nor4_1
XFILLER_18_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4922_ _4582_/B _4576_/B _4737_/A _4965_/B VGND VGND VPWR VPWR _4922_/X sky130_fd_sc_hd__o211a_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4853_ _4947_/B _4948_/C _4902_/B _4689_/B VGND VGND VPWR VPWR _4872_/A sky130_fd_sc_hd__o22a_1
XFILLER_178_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3804_ _7055_/Q hold86/A _4157_/A _6565_/Q _3803_/X VGND VGND VPWR VPWR _3807_/C
+ sky130_fd_sc_hd__a221o_2
X_4784_ _4625_/B _4702_/Y _4703_/Y _4716_/Y _4646_/Y VGND VGND VPWR VPWR _4784_/X
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_opt_2_0_csclk _6601_/CLK VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X sky130_fd_sc_hd__clkbuf_16
X_6523_ _6990_/CLK _6523_/D fanout478/X VGND VGND VPWR VPWR _6523_/Q sky130_fd_sc_hd__dfrtp_1
X_3735_ _6787_/Q _5211_/A _4151_/A _6561_/Q _3734_/X VGND VGND VPWR VPWR _3742_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6454_ _6655_/CLK _6454_/D _6383_/A VGND VGND VPWR VPWR _6454_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_174_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3666_ _6472_/Q _4032_/A _4322_/A _6712_/Q VGND VGND VPWR VPWR _3666_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5405_ hold162/X hold60/X _5408_/S VGND VGND VPWR VPWR _5405_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6385_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6385_/X sky130_fd_sc_hd__and2_1
X_3597_ _6869_/Q _5301_/A _4250_/A _6653_/Q _3596_/X VGND VGND VPWR VPWR _3597_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5336_ hold329/X _5540_/A1 _5336_/S VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5267_ hold297/X _5465_/A1 _5273_/S VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__mux2_1
X_7006_ _7006_/CLK _7006_/D fanout458/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4218_ hold495/X _5518_/A1 _4219_/S VGND VGND VPWR VPWR _4218_/X sky130_fd_sc_hd__mux2_1
X_5198_ hold443/X _5528_/A1 _5201_/S VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4149_ hold317/X _5518_/A1 _4150_/S VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3520_ _3562_/A _3577_/B VGND VGND VPWR VPWR _4172_/A sky130_fd_sc_hd__nor2_8
XFILLER_7_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold707 _5370_/X VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 _6920_/Q VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _5152_/X VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3451_ _3454_/A hold84/X VGND VGND VPWR VPWR _3562_/B sky130_fd_sc_hd__nand2_8
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3382_ _6857_/Q _5283_/A _5427_/A _6985_/Q VGND VGND VPWR VPWR _3382_/X sky130_fd_sc_hd__a22o_1
X_6170_ _7070_/Q _5934_/X _5975_/B _6873_/Q _6169_/X VGND VGND VPWR VPWR _6175_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6653_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5121_ _5087_/D _5118_/X _5120_/X _5116_/Y VGND VGND VPWR VPWR _5129_/B sky130_fd_sc_hd__a31o_1
XFILLER_57_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1407 _7150_/Q VGND VGND VPWR VPWR _3963_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1418 _6597_/Q VGND VGND VPWR VPWR hold1418/X sky130_fd_sc_hd__dlygate4sd3_1
X_5052_ _4551_/A _5041_/Y _4957_/Y VGND VGND VPWR VPWR _5142_/A sky130_fd_sc_hd__a21oi_1
XFILLER_97_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1429 _6571_/Q VGND VGND VPWR VPWR hold1429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4003_ hold646/X _5509_/A1 _4007_/S VGND VGND VPWR VPWR _4003_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5954_ _5978_/A _5966_/A _5981_/B VGND VGND VPWR VPWR _5954_/X sky130_fd_sc_hd__and3_4
XFILLER_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4905_ _5080_/A _4905_/B _5131_/A VGND VGND VPWR VPWR _4916_/B sky130_fd_sc_hd__and3_1
X_5885_ _6542_/Q _5652_/Y _5875_/X _5884_/X _6303_/S VGND VGND VPWR VPWR _5885_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4836_ _4810_/A _4810_/B _4834_/X _4835_/Y _5088_/B VGND VGND VPWR VPWR _4837_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4767_ _4764_/X _4767_/B _4767_/C _4996_/B VGND VGND VPWR VPWR _4768_/D sky130_fd_sc_hd__and4b_1
X_6506_ _7131_/CLK _6506_/D fanout459/X VGND VGND VPWR VPWR _6506_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_181_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3718_ _6875_/Q _5310_/A _5463_/A _7011_/Q VGND VGND VPWR VPWR _3718_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4698_ _4984_/A _4970_/A _4698_/C VGND VGND VPWR VPWR _4967_/B sky130_fd_sc_hd__nand3_1
XFILLER_107_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6437_ _7155_/CLK _6437_/D fanout449/X VGND VGND VPWR VPWR _6437_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3649_ _7081_/Q _5541_/A _3999_/A _6444_/Q VGND VGND VPWR VPWR _3649_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6368_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6368_/X sky130_fd_sc_hd__and2_1
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5319_ _5319_/A _5541_/B VGND VGND VPWR VPWR _5327_/S sky130_fd_sc_hd__and2_4
XFILLER_130_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6299_ _6694_/Q _5954_/X _5976_/D _6623_/Q _6280_/X VGND VGND VPWR VPWR _6300_/D
+ sky130_fd_sc_hd__a221o_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _5328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5670_/A _5670_/B VGND VGND VPWR VPWR _5670_/Y sky130_fd_sc_hd__nand2_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4621_ _4846_/B _4616_/Y _4619_/Y _4673_/A VGND VGND VPWR VPWR _4621_/X sky130_fd_sc_hd__o22a_1
XFILLER_129_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4552_ _4552_/A _4664_/A VGND VGND VPWR VPWR _4574_/A sky130_fd_sc_hd__nor2_2
XFILLER_156_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold504 _5486_/X VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _6862_/Q _5292_/A _5418_/A _6974_/Q _3502_/X VGND VGND VPWR VPWR _3504_/D
+ sky130_fd_sc_hd__a221o_1
Xhold515 _6879_/Q VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold526 _4249_/X VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4483_ _4984_/A _4636_/A VGND VGND VPWR VPWR _4483_/Y sky130_fd_sc_hd__nand2_2
XFILLER_116_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold537 _6803_/Q VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _5195_/X VGND VGND VPWR VPWR _6771_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ _6701_/Q _5971_/A _5979_/X _6471_/Q VGND VGND VPWR VPWR _6222_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold559 _5507_/X VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3434_ _6960_/Q _5400_/A _3999_/A _6448_/Q _3433_/X VGND VGND VPWR VPWR _3434_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _7124_/Q _6152_/X _6303_/S VGND VGND VPWR VPWR _6153_/X sky130_fd_sc_hd__mux2_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _3373_/B _3511_/A VGND VGND VPWR VPWR _3365_/Y sky130_fd_sc_hd__nor2_8
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5004_/A _5077_/A _5099_/X _5138_/B _5103_/Y VGND VGND VPWR VPWR _5129_/D
+ sky130_fd_sc_hd__a41o_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _5374_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6084_ _6942_/Q _5961_/X _6080_/X _6083_/X VGND VGND VPWR VPWR _6089_/A sky130_fd_sc_hd__a211o_1
Xhold1215 _6978_/Q VGND VGND VPWR VPWR _5428_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3296_ _3292_/A hold70/X _6488_/Q VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__mux2_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _5167_/X VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1237 _6690_/Q VGND VGND VPWR VPWR _4299_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _5419_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5035_ _4899_/B _5118_/B _5083_/C _5035_/D VGND VGND VPWR VPWR _5037_/C sky130_fd_sc_hd__and4b_1
Xhold1259 _6510_/Q VGND VGND VPWR VPWR _4087_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6986_ _7049_/CLK _6986_/D fanout457/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5937_ _5979_/A _5964_/A _5981_/A VGND VGND VPWR VPWR _5937_/X sky130_fd_sc_hd__and3_4
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5868_ _6687_/Q _5632_/X _5638_/X _6707_/Q VGND VGND VPWR VPWR _5868_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4819_ _4413_/Y _4902_/A _4562_/Y _4542_/B VGND VGND VPWR VPWR _5057_/A sky130_fd_sc_hd__o22a_1
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5799_ _6507_/Q _7111_/Q _6103_/B1 VGND VGND VPWR VPWR _5799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4336_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _4334_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4753_/A sky130_fd_sc_hd__clkbuf_16
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6335_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6342_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6333_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6320_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6840_ _6997_/CLK _6840_/D fanout463/X VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6771_ _7082_/CLK _6771_/D fanout479/X VGND VGND VPWR VPWR _7190_/A sky130_fd_sc_hd__dfrtp_1
X_3983_ hold828/X _6354_/A1 _3989_/S VGND VGND VPWR VPWR _3983_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5722_ _7013_/Q _5630_/X _5719_/X _5720_/X _5721_/X VGND VGND VPWR VPWR _5722_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6683_/CLK sky130_fd_sc_hd__clkbuf_16
X_5653_ _6850_/Q _5648_/X _5652_/B _6914_/Q _5651_/Y VGND VGND VPWR VPWR _5653_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4604_ _4753_/A _4753_/B VGND VGND VPWR VPWR _4970_/A sky130_fd_sc_hd__and2b_2
X_5584_ _5584_/A VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7076_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold301 _6939_/Q VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlygate4sd3_1
X_4535_ _4535_/A _4535_/B _4535_/C _4535_/D VGND VGND VPWR VPWR _4537_/C sky130_fd_sc_hd__and4_1
XFILLER_116_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold312 _5504_/X VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _7058_/Q VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _5286_/X VGND VGND VPWR VPWR _6852_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold345 _6693_/Q VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _4272_/X VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4466_ _4493_/B VGND VGND VPWR VPWR _4846_/A sky130_fd_sc_hd__inv_2
Xhold367 _6753_/Q VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold378 _4290_/X VGND VGND VPWR VPWR _6683_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6205_ _6466_/Q _5937_/X _5975_/D _6626_/Q VGND VGND VPWR VPWR _6205_/X sky130_fd_sc_hd__a22o_1
Xhold389 _6653_/Q VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3417_ _7131_/Q _6761_/Q _6762_/Q VGND VGND VPWR VPWR _3417_/X sky130_fd_sc_hd__mux2_2
X_7185_ _7185_/A VGND VGND VPWR VPWR _7185_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4397_ _4739_/A _4396_/A _4400_/B VGND VGND VPWR VPWR _4415_/B sky130_fd_sc_hd__o21a_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6896_/Q _5946_/X _5955_/X _6808_/Q VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__a22o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3348_ _3586_/A _3714_/B VGND VGND VPWR VPWR _5211_/A sky130_fd_sc_hd__nor2_8
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _6666_/Q VGND VGND VPWR VPWR _4270_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 _4210_/X VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _6676_/Q VGND VGND VPWR VPWR _4282_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1034 _4216_/X VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ _6901_/Q _5976_/C _5971_/D _6829_/Q VGND VGND VPWR VPWR _6067_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3279_ hold62/X hold81/A _6488_/Q VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__mux2_2
Xhold1045 _6820_/Q VGND VGND VPWR VPWR _5250_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 _5482_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1067 _6834_/Q VGND VGND VPWR VPWR _5266_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5018_ _5018_/A _5112_/C _5018_/C _5018_/D VGND VGND VPWR VPWR _5021_/C sky130_fd_sc_hd__and4_1
Xhold1078 _5275_/X VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _6805_/Q VGND VGND VPWR VPWR _5233_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_207 _5171_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _6969_/CLK _6969_/D fanout474/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold890 _6738_/Q VGND VGND VPWR VPWR hold890/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1590 _7181_/A VGND VGND VPWR VPWR hold1590/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4320_ hold740/X _6356_/A1 _4321_/S VGND VGND VPWR VPWR _4320_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4251_ _4251_/A0 _6353_/A1 _4255_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3202_ _6957_/Q VGND VGND VPWR VPWR _3202_/Y sky130_fd_sc_hd__inv_2
X_4182_ _3640_/Y _4182_/A1 _4186_/S VGND VGND VPWR VPWR _6586_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6823_ _6951_/CLK _6823_/D fanout474/X VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_2
X_6754_ _7011_/CLK _6754_/D fanout456/X VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfrtp_4
X_3966_ _3966_/A0 _5491_/A1 _3980_/S VGND VGND VPWR VPWR _3966_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5705_ _6820_/Q _5818_/A2 _5814_/B1 _6908_/Q _5704_/X VGND VGND VPWR VPWR _5706_/D
+ sky130_fd_sc_hd__a221o_1
X_6685_ _6707_/CLK _6685_/D fanout448/X VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_2
X_3897_ _4702_/A _4566_/A VGND VGND VPWR VPWR _4374_/A sky130_fd_sc_hd__and2_1
X_5636_ _6970_/Q _5634_/X _5635_/X _6826_/Q VGND VGND VPWR VPWR _5636_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5567_ _6506_/Q _6508_/Q VGND VGND VPWR VPWR _5567_/Y sky130_fd_sc_hd__nor2_1
Xhold120 _6412_/Q VGND VGND VPWR VPWR _3292_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _7014_/Q VGND VGND VPWR VPWR hold131/X sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _4515_/Y _4518_/B _4518_/C _4518_/D VGND VGND VPWR VPWR _4522_/A sky130_fd_sc_hd__and4b_1
Xhold142 _5290_/X VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold153 _5450_/X VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5498_ hold602/X _5543_/A1 hold77/X VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold164 _7008_/Q VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _5318_/X VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _4551_/A _4813_/A _4579_/B VGND VGND VPWR VPWR _4948_/B sky130_fd_sc_hd__nand3_4
Xhold186 _6684_/Q VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _5243_/X VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7168_ _3945_/A1 _7168_/D _6398_/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6119_ _7052_/Q _5971_/A _5979_/X _6991_/Q _6105_/X VGND VGND VPWR VPWR _6125_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_19_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7113_/CLK _7099_/D fanout464/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_85_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ _7071_/Q _5532_/A _4139_/A _6550_/Q VGND VGND VPWR VPWR _3820_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3751_ _3751_/A _3751_/B _3751_/C _3751_/D VGND VGND VPWR VPWR _3761_/C sky130_fd_sc_hd__nor4_1
XFILLER_186_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6470_ _6735_/CLK _6470_/D _3946_/B VGND VGND VPWR VPWR _6470_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3682_ _6567_/Q _4157_/A _4250_/A _6652_/Q VGND VGND VPWR VPWR _3682_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5421_ hold880/X _5484_/A1 _5426_/S VGND VGND VPWR VPWR _5421_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput203 _3922_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
XFILLER_114_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5352_ hold449/X _5538_/A1 _5354_/S VGND VGND VPWR VPWR _5352_/X sky130_fd_sc_hd__mux2_1
Xoutput214 _3926_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
Xoutput225 _7187_/X VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
XFILLER_99_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput236 _3923_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
Xoutput247 _3928_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput258 _6746_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
X_4303_ hold838/X _5546_/A1 _4303_/S VGND VGND VPWR VPWR _4303_/X sky130_fd_sc_hd__mux2_1
X_5283_ _5283_/A hold17/X VGND VGND VPWR VPWR _5291_/S sky130_fd_sc_hd__and2_4
Xoutput269 _6743_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
XFILLER_141_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7022_ _7051_/CLK _7022_/D fanout476/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfrtp_4
X_4234_ hold413/X _5534_/A1 _4237_/S VGND VGND VPWR VPWR _4234_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4165_ _3762_/Y _4165_/A1 _4171_/S VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4096_ hold168/X hold42/X _5202_/B VGND VGND VPWR VPWR _4096_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6806_ _7051_/CLK _6806_/D fanout476/X VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4998_ _5068_/C _5069_/C _4998_/C VGND VGND VPWR VPWR _5001_/A sky130_fd_sc_hd__and3_1
XFILLER_11_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3949_ _6403_/Q _3949_/B VGND VGND VPWR VPWR _3950_/A sky130_fd_sc_hd__nor2_2
X_6737_ _6739_/CLK _6737_/D _3946_/B VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6668_ _6668_/CLK _6668_/D fanout452/X VGND VGND VPWR VPWR _6668_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5619_ _5664_/A _5666_/B _5666_/C VGND VGND VPWR VPWR _5619_/X sky130_fd_sc_hd__and3_4
XFILLER_191_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6599_ _6654_/CLK _6599_/D fanout454/X VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout430 hold16/X VGND VGND VPWR VPWR _4322_/B sky130_fd_sc_hd__buf_6
Xfanout441 _6396_/B VGND VGND VPWR VPWR _6401_/B sky130_fd_sc_hd__clkbuf_4
Xfanout452 fanout455/X VGND VGND VPWR VPWR fanout452/X sky130_fd_sc_hd__buf_6
Xfanout463 fanout465/X VGND VGND VPWR VPWR fanout463/X sky130_fd_sc_hd__buf_8
XFILLER_58_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout474 fanout475/X VGND VGND VPWR VPWR fanout474/X sky130_fd_sc_hd__clkbuf_16
Xfanout485 fanout486/X VGND VGND VPWR VPWR fanout485/X sky130_fd_sc_hd__buf_8
XFILLER_74_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5970_ _5600_/A _5969_/A _5981_/C _5943_/X _5965_/X VGND VGND VPWR VPWR _5970_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4921_ _4921_/A _5043_/A VGND VGND VPWR VPWR _4921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4852_ _4947_/B _4456_/Y _4902_/B _4628_/Y VGND VGND VPWR VPWR _4852_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3803_ input43/X _4058_/S _4102_/A input61/X VGND VGND VPWR VPWR _3803_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4783_ _4846_/B _4644_/Y _4663_/Y _4782_/Y VGND VGND VPWR VPWR _5108_/B sky130_fd_sc_hd__o22a_1
X_6522_ _6990_/CLK _6522_/D fanout478/X VGND VGND VPWR VPWR _6522_/Q sky130_fd_sc_hd__dfrtp_1
X_3734_ _6656_/Q _4256_/A _4298_/A _6691_/Q VGND VGND VPWR VPWR _3734_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6453_ _6655_/CLK _6453_/D _6383_/A VGND VGND VPWR VPWR _6453_/Q sky130_fd_sc_hd__dfrtp_4
X_3665_ _6436_/Q _3372_/Y _4280_/A _6677_/Q _3664_/X VGND VGND VPWR VPWR _3670_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5404_ hold221/X _5494_/A1 _5408_/S VGND VGND VPWR VPWR _5404_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6384_ _6401_/A _6400_/B VGND VGND VPWR VPWR _6384_/X sky130_fd_sc_hd__and2_1
X_3596_ _6861_/Q _5292_/A _3593_/X _3595_/X VGND VGND VPWR VPWR _3596_/X sky130_fd_sc_hd__a211o_1
XFILLER_127_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5335_ hold940/X _5548_/A1 _5336_/S VGND VGND VPWR VPWR _5335_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5266_ _5266_/A0 hold666/X _5273_/S VGND VGND VPWR VPWR _5266_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7005_ _7017_/CLK _7005_/D fanout466/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfrtp_4
X_4217_ hold662/X _5544_/A1 _4219_/S VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
X_5197_ _5197_/A0 _5545_/A1 _5201_/S VGND VGND VPWR VPWR _5197_/X sky130_fd_sc_hd__mux2_1
X_4148_ hold453/X _5544_/A1 _4150_/S VGND VGND VPWR VPWR _4148_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4079_ hold742/X hold42/X _4083_/S VGND VGND VPWR VPWR _4079_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold708 _6919_/Q VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold719 _5362_/X VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3450_ _7118_/Q _6760_/Q _6762_/Q VGND VGND VPWR VPWR _3450_/X sky130_fd_sc_hd__mux2_2
X_3381_ _3511_/A hold66/A VGND VGND VPWR VPWR _3381_/Y sky130_fd_sc_hd__nor2_8
X_5120_ _4906_/Y _5120_/B _5120_/C VGND VGND VPWR VPWR _5120_/X sky130_fd_sc_hd__and3b_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5051_ _5051_/A _5051_/B VGND VGND VPWR VPWR _5089_/C sky130_fd_sc_hd__nand2_1
Xhold1408 _7005_/Q VGND VGND VPWR VPWR _5458_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 _6586_/Q VGND VGND VPWR VPWR hold1419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4002_ hold886/X _5484_/A1 _4007_/S VGND VGND VPWR VPWR _4002_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5953_ _5969_/A _5969_/C _5981_/C VGND VGND VPWR VPWR _5953_/X sky130_fd_sc_hd__and3_4
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4904_ _4359_/Y _4900_/Y _4850_/Y VGND VGND VPWR VPWR _5131_/A sky130_fd_sc_hd__o21a_1
XFILLER_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5884_ _6547_/Q _5655_/X _5879_/X _5881_/X _5883_/X VGND VGND VPWR VPWR _5884_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4835_ _4551_/B _4554_/B _4574_/A VGND VGND VPWR VPWR _4835_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4766_ _4627_/A _4626_/Y _4643_/Y _4948_/C _4672_/B VGND VGND VPWR VPWR _4767_/C
+ sky130_fd_sc_hd__o32a_1
X_6505_ _6537_/CLK _6505_/D fanout464/X VGND VGND VPWR VPWR _7178_/A sky130_fd_sc_hd__dfrtp_1
X_3717_ hold28/X _3717_/B VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__nor2_4
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4697_ _4911_/B _4703_/B VGND VGND VPWR VPWR _4697_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6436_ _6747_/CLK _6436_/D fanout447/X VGND VGND VPWR VPWR _6436_/Q sky130_fd_sc_hd__dfstp_2
X_3648_ _3957_/A _4102_/A _3585_/Y input97/X _3647_/X VGND VGND VPWR VPWR _3651_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6367_ _6383_/A _6367_/B VGND VGND VPWR VPWR _6367_/X sky130_fd_sc_hd__and2_1
XFILLER_88_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3579_ _6870_/Q _5301_/A _4014_/A _6459_/Q _3578_/X VGND VGND VPWR VPWR _3580_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5318_ _5318_/A0 hold22/X _5318_/S VGND VGND VPWR VPWR _5318_/X sky130_fd_sc_hd__mux2_1
X_6298_ _6559_/Q _5971_/B _5949_/X _6679_/Q _6297_/X VGND VGND VPWR VPWR _6300_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold13 hold9/X VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__buf_6
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ hold287/X _5534_/A1 _5255_/S VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4620_ _4716_/A _4975_/A VGND VGND VPWR VPWR _4620_/Y sky130_fd_sc_hd__nand2_2
XFILLER_187_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4551_ _4551_/A _4551_/B VGND VGND VPWR VPWR _5088_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3502_ hold79/A _3999_/A _4256_/A _6659_/Q VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__a22o_1
Xhold505 _6553_/Q VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _5316_/X VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4482_/A _4482_/B VGND VGND VPWR VPWR _4972_/A sky130_fd_sc_hd__nor2_2
XFILLER_171_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold527 _6425_/Q VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _5231_/X VGND VGND VPWR VPWR _6803_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6561_/Q _5953_/X _5960_/X _6671_/Q _6220_/X VGND VGND VPWR VPWR _6221_/X
+ sky130_fd_sc_hd__a221o_1
X_3433_ _7032_/Q hold49/A _5463_/A _7016_/Q VGND VGND VPWR VPWR _3433_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold549 _6891_/Q VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6140_/Y _6151_/X _6792_/Q _6226_/B VGND VGND VPWR VPWR _6152_/X sky130_fd_sc_hd__o2bb2a_1
X_3364_ _3714_/A hold74/X VGND VGND VPWR VPWR _5436_/A sky130_fd_sc_hd__nor2_8
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5103_/A _5103_/B _5103_/C VGND VGND VPWR VPWR _5103_/Y sky130_fd_sc_hd__nand3_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6862_/Q _5943_/X _5981_/X _6918_/Q _6079_/X VGND VGND VPWR VPWR _6083_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _7002_/Q VGND VGND VPWR VPWR _5455_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3295_ _3295_/A _3323_/B VGND VGND VPWR VPWR _3295_/Y sky130_fd_sc_hd__nor2_4
Xhold1216 _5428_/X VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A _5034_/B _5085_/B _5034_/D VGND VGND VPWR VPWR _5035_/D sky130_fd_sc_hd__and4_1
Xhold1227 _6898_/Q VGND VGND VPWR VPWR _5338_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 _4299_/X VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _7063_/Q VGND VGND VPWR VPWR _5524_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6985_ _7033_/CLK _6985_/D fanout464/X VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5936_ _5968_/A _5981_/B _5969_/C VGND VGND VPWR VPWR _5971_/B sky130_fd_sc_hd__and3_4
XFILLER_179_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5867_ _7153_/Q _5625_/X _5661_/X _6621_/Q VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4818_ _4902_/A _4456_/Y _4562_/Y _4948_/C VGND VGND VPWR VPWR _4818_/X sky130_fd_sc_hd__o22a_1
XFILLER_166_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5798_ _3227_/Y _5651_/Y _5787_/Y _5797_/Y _5552_/B VGND VGND VPWR VPWR _5798_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _4413_/Y _4581_/B _4611_/Y _4616_/Y VGND VGND VPWR VPWR _5099_/C sky130_fd_sc_hd__o22a_1
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6419_ _7049_/CLK _6419_/D fanout457/X VGND VGND VPWR VPWR _6419_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_103_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4336_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _4334_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _4642_/A sky130_fd_sc_hd__clkbuf_8
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6338_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6345_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6336_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_stb_i VGND VGND VPWR VPWR _3899_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_57_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6668_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3982_ _3982_/A0 _6353_/A1 _3989_/S VGND VGND VPWR VPWR _3982_/X sky130_fd_sc_hd__mux2_1
X_6770_ _7080_/CLK _6770_/D fanout479/X VGND VGND VPWR VPWR _7189_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5721_ _6949_/Q _5637_/X _5645_/X _7029_/Q VGND VGND VPWR VPWR _5721_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5652_ _5899_/B _5652_/B VGND VGND VPWR VPWR _5652_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_175_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4603_ _4607_/A _4993_/B VGND VGND VPWR VPWR _4682_/A sky130_fd_sc_hd__nand2_1
X_5583_ _5582_/Y _5664_/A _5583_/S VGND VGND VPWR VPWR _5584_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4534_ _4782_/A _4881_/B _5088_/A VGND VGND VPWR VPWR _4535_/D sky130_fd_sc_hd__a21boi_1
Xhold302 _5384_/X VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold313 _7062_/Q VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _5518_/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _7049_/Q VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _4302_/X VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _4489_/A _4465_/B VGND VGND VPWR VPWR _4493_/B sky130_fd_sc_hd__and2_1
Xhold357 _6980_/Q VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _5169_/X VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ _3714_/B _3571_/B VGND VGND VPWR VPWR _5182_/S sky130_fd_sc_hd__nor2_8
X_6204_ _6204_/A0 _6203_/X _6279_/S VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold379 _6991_/Q VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlygate4sd3_1
X_7184_ _7184_/A VGND VGND VPWR VPWR _7184_/X sky130_fd_sc_hd__clkbuf_1
X_4396_ _4396_/A _4396_/B VGND VGND VPWR VPWR _4415_/A sky130_fd_sc_hd__nor2_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _6944_/Q _5961_/X _6131_/X _6134_/X VGND VGND VPWR VPWR _6140_/A sky130_fd_sc_hd__a211o_1
X_3347_ _3347_/A _3356_/B VGND VGND VPWR VPWR _3714_/B sky130_fd_sc_hd__nand2_8
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _4270_/X VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _6519_/Q VGND VGND VPWR VPWR _4104_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1024 _4282_/X VGND VGND VPWR VPWR _6676_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6066_ _6066_/A _6066_/B _6066_/C VGND VGND VPWR VPWR _6075_/C sky130_fd_sc_hd__nor3_2
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1035 _6551_/Q VGND VGND VPWR VPWR _4141_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3278_ hold83/X VGND VGND VPWR VPWR _3453_/A sky130_fd_sc_hd__clkinv_2
Xhold1046 _5250_/X VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 _6973_/Q VGND VGND VPWR VPWR _5422_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ _5106_/B _5064_/B _5062_/D VGND VGND VPWR VPWR _5018_/D sky130_fd_sc_hd__and3_1
Xhold1068 _5266_/X VGND VGND VPWR VPWR _6834_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1079 _6813_/Q VGND VGND VPWR VPWR _5242_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6968_ _7069_/CLK _6968_/D fanout482/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_2
X_5919_ _7038_/Q _5614_/X _5917_/X _5918_/X VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__a211o_1
X_6899_ _7080_/CLK _6899_/D fanout479/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_139_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold880 _6972_/Q VGND VGND VPWR VPWR hold880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 _5150_/X VGND VGND VPWR VPWR _6738_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1580 _7100_/Q VGND VGND VPWR VPWR _5596_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1591 _6528_/Q VGND VGND VPWR VPWR hold812/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4250_ _4250_/A _5490_/B VGND VGND VPWR VPWR _4255_/S sky130_fd_sc_hd__and2_2
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3201_ _6965_/Q VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__inv_2
X_4181_ _3700_/Y _4181_/A1 _4186_/S VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6822_ _6884_/CLK _6822_/D fanout475/X VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6753_ _7011_/CLK _6753_/D fanout459/X VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfrtp_4
X_3965_ _3251_/A hold664/X _3975_/S VGND VGND VPWR VPWR _3965_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5704_ _6996_/Q _5643_/X _5652_/B _6916_/Q _5651_/Y VGND VGND VPWR VPWR _5704_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3896_ _5552_/B _3887_/Y _5959_/A _5966_/A _3895_/X VGND VGND VPWR VPWR _6509_/D
+ sky130_fd_sc_hd__a41o_1
X_6684_ _6714_/CLK _6684_/D fanout470/X VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_2
X_5635_ _5638_/A _5657_/B _5666_/C VGND VGND VPWR VPWR _5635_/X sky130_fd_sc_hd__and3b_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5566_ _3176_/Y _5564_/B _5565_/X VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__a21boi_1
Xhold110 _7006_/Q VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _3292_/X VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold132 _5468_/X VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ _4953_/A _5042_/B VGND VGND VPWR VPWR _4518_/C sky130_fd_sc_hd__nand2_1
X_5497_ _5497_/A0 hold667/X hold77/A VGND VGND VPWR VPWR _5497_/X sky130_fd_sc_hd__mux2_1
Xhold143 _6985_/Q VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold154 _7144_/Q VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _5461_/X VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold176 _7070_/Q VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _4408_/B _4448_/B VGND VGND VPWR VPWR _4579_/B sky130_fd_sc_hd__and2b_4
Xhold187 _4291_/X VGND VGND VPWR VPWR _6684_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _7037_/Q VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7167_ _3945_/A1 _7167_/D _6397_/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_1
X_4379_ _4360_/B _4379_/B VGND VGND VPWR VPWR _4384_/A sky130_fd_sc_hd__nand2b_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6118_ _6823_/Q _5953_/X _5960_/X _7076_/Q _6117_/X VGND VGND VPWR VPWR _6118_/X
+ sky130_fd_sc_hd__a221o_1
X_7098_ _7113_/CLK _7098_/D fanout462/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfstp_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6049_ _6049_/A _6049_/B _6049_/C _6049_/D VGND VGND VPWR VPWR _6049_/Y sky130_fd_sc_hd__nor4_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6714_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6527_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ input12/X _3358_/Y _4208_/A _6610_/Q _3749_/X VGND VGND VPWR VPWR _3751_/D
+ sky130_fd_sc_hd__a221o_1
X_3681_ _6836_/Q _5265_/A _5319_/A _6884_/Q _3680_/X VGND VGND VPWR VPWR _3688_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5420_ hold634/X _5543_/A1 _5426_/S VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5351_ hold485/X _5528_/A1 _5354_/S VGND VGND VPWR VPWR _5351_/X sky130_fd_sc_hd__mux2_1
Xoutput204 _3921_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
Xoutput215 _7179_/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput226 _7188_/X VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput237 _3924_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
Xoutput248 _3946_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
X_4302_ hold345/X _5518_/A1 _4303_/S VGND VGND VPWR VPWR _4302_/X sky130_fd_sc_hd__mux2_1
Xoutput259 _6747_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
X_5282_ hold624/X _5513_/A1 _5282_/S VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4233_ _4233_/A0 hold667/X _4237_/S VGND VGND VPWR VPWR _4233_/X sky130_fd_sc_hd__mux2_1
X_7021_ _7082_/CLK _7021_/D fanout483/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4164_ _3828_/Y _4164_/A1 _4171_/S VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4095_ hold393/X _4094_/X _4101_/S VGND VGND VPWR VPWR _4095_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6805_ _7085_/CLK _6805_/D fanout477/X VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4997_ _5073_/A _5103_/A _4997_/C _4997_/D VGND VGND VPWR VPWR _4998_/C sky130_fd_sc_hd__and4_1
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6736_ _6739_/CLK _6736_/D _3946_/B VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfstp_2
X_3948_ _3948_/A VGND VGND VPWR VPWR _3948_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6667_ _6668_/CLK _6667_/D fanout452/X VGND VGND VPWR VPWR _6667_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_164_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3879_ _6642_/Q _3962_/B _3879_/B1 VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__a21o_1
XFILLER_176_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5618_ _7093_/Q _7092_/Q VGND VGND VPWR VPWR _5666_/C sky130_fd_sc_hd__and2b_2
XFILLER_192_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6598_ _7137_/CLK _6598_/D VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5549_ _5549_/A0 hold22/X _5549_/S VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__mux2_1
XFILLER_117_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout420 hold13/X VGND VGND VPWR VPWR _5534_/A1 sky130_fd_sc_hd__buf_12
Xfanout431 _5505_/B VGND VGND VPWR VPWR _5541_/B sky130_fd_sc_hd__buf_6
Xfanout442 _3268_/Y VGND VGND VPWR VPWR _6396_/B sky130_fd_sc_hd__clkbuf_16
Xfanout453 fanout454/X VGND VGND VPWR VPWR _6401_/A sky130_fd_sc_hd__clkbuf_8
Xfanout464 fanout465/X VGND VGND VPWR VPWR fanout464/X sky130_fd_sc_hd__buf_8
Xfanout475 fanout486/X VGND VGND VPWR VPWR fanout475/X sky130_fd_sc_hd__buf_8
Xfanout486 input75/X VGND VGND VPWR VPWR fanout486/X sky130_fd_sc_hd__buf_12
XFILLER_101_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _7150_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4920_ _5023_/B _4920_/B _4964_/C VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__and3_1
XFILLER_80_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4851_ _4413_/Y _4496_/Y _4616_/Y _4689_/A VGND VGND VPWR VPWR _4877_/A sky130_fd_sc_hd__o22a_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3802_ input4/X _3381_/Y _4044_/A _6480_/Q _3801_/X VGND VGND VPWR VPWR _3807_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4782_ _4782_/A _4975_/A VGND VGND VPWR VPWR _4782_/Y sky130_fd_sc_hd__nor2_1
X_6521_ _6755_/CLK _6521_/D _6360_/A VGND VGND VPWR VPWR _6521_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3733_ _6979_/Q _5427_/A _3414_/Y _3732_/X VGND VGND VPWR VPWR _3733_/X sky130_fd_sc_hd__a211o_1
XFILLER_118_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6452_ _6677_/CLK _6452_/D fanout452/X VGND VGND VPWR VPWR _6452_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_118_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3664_ _6988_/Q _5436_/A _4139_/A _6552_/Q VGND VGND VPWR VPWR _3664_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5403_ hold387/X _5526_/A1 _5408_/S VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__mux2_1
X_6383_ _6383_/A _6401_/B VGND VGND VPWR VPWR _6383_/X sky130_fd_sc_hd__and2_1
X_3595_ input38/X _3331_/Y _4298_/A _6693_/Q _3594_/X VGND VGND VPWR VPWR _3595_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5334_ hold417/X _5538_/A1 _5336_/S VGND VGND VPWR VPWR _5334_/X sky130_fd_sc_hd__mux2_1
X_5265_ _5265_/A hold17/X VGND VGND VPWR VPWR _5273_/S sky130_fd_sc_hd__and2_4
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7004_ _7012_/CLK _7004_/D fanout466/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_141_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4216_ _4216_/A0 _5492_/A1 _4219_/S VGND VGND VPWR VPWR _4216_/X sky130_fd_sc_hd__mux2_1
X_5196_ hold858/X _5484_/A1 _5201_/S VGND VGND VPWR VPWR _5196_/X sky130_fd_sc_hd__mux2_1
X_4147_ hold281/X _5534_/A1 _4150_/S VGND VGND VPWR VPWR _4147_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4078_ hold349/X _4077_/X _4084_/S VGND VGND VPWR VPWR _4078_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6719_ _7038_/CLK _6719_/D fanout455/X VGND VGND VPWR VPWR _6719_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold709 _5361_/X VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap439 _4434_/B VGND VGND VPWR VPWR _4591_/A sky130_fd_sc_hd__buf_2
XFILLER_109_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3380_ hold65/X _3415_/B VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__nand2_8
XFILLER_170_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5050_ _4456_/Y _4946_/X _5049_/X _4820_/X VGND VGND VPWR VPWR _5058_/C sky130_fd_sc_hd__o211a_1
XFILLER_69_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1409 _6750_/Q VGND VGND VPWR VPWR _5165_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4001_ hold263/X _5465_/A1 _4007_/S VGND VGND VPWR VPWR _4001_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5952_ _5969_/A _5979_/A _5981_/A VGND VGND VPWR VPWR _5952_/X sky130_fd_sc_hd__and3_4
XFILLER_46_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4903_ _4493_/B _5024_/B _4841_/X VGND VGND VPWR VPWR _4905_/B sky130_fd_sc_hd__a21oi_1
X_5883_ _6580_/Q _5928_/A2 _5913_/B1 _6552_/Q _5882_/X VGND VGND VPWR VPWR _5883_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4834_ _4413_/Y _4810_/B _4823_/X _4833_/X VGND VGND VPWR VPWR _4834_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4765_ _4921_/A _4992_/B _4588_/Y VGND VGND VPWR VPWR _4767_/B sky130_fd_sc_hd__a21oi_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6504_ _6755_/CLK _6504_/D _6360_/A VGND VGND VPWR VPWR _6504_/Q sky130_fd_sc_hd__dfrtp_1
X_3716_ _6605_/Q _4202_/A _3714_/Y _6749_/Q _3715_/X VGND VGND VPWR VPWR _3720_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4696_ _4694_/Y _4695_/Y _4482_/B VGND VGND VPWR VPWR _4706_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _6746_/CLK _6435_/D fanout447/X VGND VGND VPWR VPWR _6435_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_161_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3647_ _7020_/Q hold29/A _4196_/A _6601_/Q VGND VGND VPWR VPWR _3647_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6366_ _6383_/A _6401_/B VGND VGND VPWR VPWR _6366_/X sky130_fd_sc_hd__and2_1
XFILLER_115_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3578_ _6806_/Q _5229_/A _4102_/A _7199_/A VGND VGND VPWR VPWR _3578_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5317_ hold918/X _5548_/A1 _5318_/S VGND VGND VPWR VPWR _5317_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6297_ _7038_/Q _5601_/X _5959_/X _6719_/Q VGND VGND VPWR VPWR _6297_/X sky130_fd_sc_hd__a22o_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5248_ _5248_/A0 _5473_/A1 _5255_/S VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__mux2_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__buf_6
XFILLER_102_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ hold696/X _5469_/A1 _5181_/S VGND VGND VPWR VPWR _5179_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4550_ _4947_/B _4553_/B VGND VGND VPWR VPWR _4551_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3501_ _3555_/A _3546_/A VGND VGND VPWR VPWR _4256_/A sky130_fd_sc_hd__nor2_4
XFILLER_144_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold506 _4143_/X VGND VGND VPWR VPWR _6553_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4481_ _4615_/B _4653_/C VGND VGND VPWR VPWR _4482_/B sky130_fd_sc_hd__nand2_4
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold517 _7068_/Q VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 _3980_/X VGND VGND VPWR VPWR _6425_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold539 _6484_/Q VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ _6651_/Q _5973_/A _5948_/X _6696_/Q _6219_/X VGND VGND VPWR VPWR _6220_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_144_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3432_ _6880_/Q _5310_/A _5238_/A _6816_/Q VGND VGND VPWR VPWR _3432_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3363_ _3814_/A _3714_/A VGND VGND VPWR VPWR _5505_/A sky130_fd_sc_hd__nor2_8
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _6143_/X _6145_/X _6151_/C _6226_/B VGND VGND VPWR VPWR _6151_/X sky130_fd_sc_hd__and4bb_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _4626_/Y _4663_/Y _4933_/C _5101_/X VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__o211a_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3294_ hold32/X _3975_/S hold121/X _3293_/Y VGND VGND VPWR VPWR _3294_/X sky130_fd_sc_hd__o31a_2
X_6082_ _7083_/Q _5976_/B _5971_/C _7043_/Q VGND VGND VPWR VPWR _6099_/B sky130_fd_sc_hd__a22o_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _5455_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _6946_/Q VGND VGND VPWR VPWR _5392_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5033_ _5033_/A _5080_/B _5033_/C _5120_/B VGND VGND VPWR VPWR _5034_/D sky130_fd_sc_hd__and4_1
Xhold1228 _5338_/X VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 _7055_/Q VGND VGND VPWR VPWR _5515_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6984_ _7001_/CLK _6984_/D fanout461/X VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5935_ _7101_/Q _7102_/Q VGND VGND VPWR VPWR _5969_/C sky130_fd_sc_hd__nor2_8
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5866_ _3185_/Y _5899_/B _5651_/B VGND VGND VPWR VPWR _5866_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4817_ _4817_/A _4972_/A VGND VGND VPWR VPWR _5018_/A sky130_fd_sc_hd__nand2_2
X_5797_ _5797_/A _5797_/B _5797_/C _5797_/D VGND VGND VPWR VPWR _5797_/Y sky130_fd_sc_hd__nor4_4
XFILLER_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4748_ _4921_/A _4926_/B VGND VGND VPWR VPWR _5074_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4679_ _4925_/B _4679_/B _4679_/C _4679_/D VGND VGND VPWR VPWR _4682_/C sky130_fd_sc_hd__and4_1
XFILLER_107_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6418_ _6749_/CLK _6418_/D fanout449/X VGND VGND VPWR VPWR _6418_/Q sky130_fd_sc_hd__dfstp_1
X_6349_ _6643_/Q _6319_/B _6348_/X VGND VGND VPWR VPWR _6349_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3904_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_102_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR _4739_/A sky130_fd_sc_hd__buf_6
XFILLER_76_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6341_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6324_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6339_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3981_ _3981_/A _6352_/B VGND VGND VPWR VPWR _3989_/S sky130_fd_sc_hd__and2_2
X_5720_ _6941_/Q _5632_/X _5638_/X _6957_/Q VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5651_ _5899_/B _5651_/B VGND VGND VPWR VPWR _5651_/Y sky130_fd_sc_hd__nor2_8
X_4602_ _4993_/B VGND VGND VPWR VPWR _4602_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5582_ _5664_/A _5602_/A VGND VGND VPWR VPWR _5582_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4533_ _4490_/Y _5083_/A _4912_/A _4533_/D VGND VGND VPWR VPWR _4535_/C sky130_fd_sc_hd__and4b_1
XFILLER_190_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold303 _6713_/Q VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _5522_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 _6924_/Q VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _5508_/X VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4464_ _5051_/B VGND VGND VPWR VPWR _4464_/Y sky130_fd_sc_hd__inv_2
Xhold347 _6663_/Q VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _5430_/X VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6203_ _6203_/A0 _6202_/X _6303_/S VGND VGND VPWR VPWR _6203_/X sky130_fd_sc_hd__mux2_1
Xhold369 _6836_/Q VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3415_ hold84/X _3415_/B VGND VGND VPWR VPWR _3571_/B sky130_fd_sc_hd__nand2_8
X_7183_ _7183_/A VGND VGND VPWR VPWR _7183_/X sky130_fd_sc_hd__clkbuf_1
X_4395_ _4642_/A _4441_/B VGND VGND VPWR VPWR _4396_/B sky130_fd_sc_hd__nor2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _7016_/Q _5940_/X _5967_/X _6856_/Q _6130_/X VGND VGND VPWR VPWR _6134_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _3347_/A _3355_/B hold72/X VGND VGND VPWR VPWR _5190_/B sky130_fd_sc_hd__and3_2
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1003 _6725_/Q VGND VGND VPWR VPWR hold1003/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _4104_/X VGND VGND VPWR VPWR _6519_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6065_ _6981_/Q _5945_/X _5975_/C _6837_/Q _6064_/X VGND VGND VPWR VPWR _6066_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 _6561_/Q VGND VGND VPWR VPWR _4153_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3277_ hold82/X _4988_/B2 _3975_/S VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__mux2_2
Xhold1036 _4141_/X VGND VGND VPWR VPWR _6551_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1047 _6884_/Q VGND VGND VPWR VPWR _5322_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 _5422_/X VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5016_ _4644_/Y _4975_/Y _4991_/X _5011_/X VGND VGND VPWR VPWR _5062_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1069 _6933_/Q VGND VGND VPWR VPWR _5377_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _6967_/CLK _6967_/D fanout474/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5918_ _6484_/Q _5643_/X _5664_/X _6669_/Q VGND VGND VPWR VPWR _5918_/X sky130_fd_sc_hd__a22o_1
X_6898_ _7083_/CLK _6898_/D fanout476/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5849_ _7035_/Q _5614_/X _5643_/X _6481_/Q VGND VGND VPWR VPWR _5849_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold870 _6467_/Q VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold881 _5421_/X VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _6448_/Q VGND VGND VPWR VPWR hold892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1570 _7158_/Q VGND VGND VPWR VPWR _3868_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1581 _6760_/Q VGND VGND VPWR VPWR hold696/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1592 _7101_/Q VGND VGND VPWR VPWR _5598_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3200_ _6973_/Q VGND VGND VPWR VPWR _3200_/Y sky130_fd_sc_hd__inv_2
X_4180_ _3762_/Y _4180_/A1 _4186_/S VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6821_ _7076_/CLK _6821_/D fanout481/X VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6752_ _7011_/CLK _6752_/D fanout456/X VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_4
X_3964_ _3964_/A _6352_/B VGND VGND VPWR VPWR _3980_/S sky130_fd_sc_hd__and2_2
X_5703_ _6444_/Q _5614_/X _5664_/X _6924_/Q _5702_/X VGND VGND VPWR VPWR _5706_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6683_ _6683_/CLK _6683_/D _6390_/A VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfrtp_1
X_3895_ _7088_/Q _3886_/B _7090_/Q _7091_/Q _6509_/Q VGND VGND VPWR VPWR _3895_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_176_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5634_ _5638_/A _5667_/B _5657_/B VGND VGND VPWR VPWR _5634_/X sky130_fd_sc_hd__and3_4
XFILLER_176_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5565_ _3176_/Y _5564_/B _5564_/A VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__o21a_1
XFILLER_163_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 _4125_/X VGND VGND VPWR VPWR _6538_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _5459_/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4531_/B _4953_/A VGND VGND VPWR VPWR _4518_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold122 _3294_/X VGND VGND VPWR VPWR _3323_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _6757_/Q VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5496_ hold76/X _5541_/B VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__and2_4
Xhold144 _5435_/X VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold155 _3971_/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _6838_/Q VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _4454_/A _4611_/B VGND VGND VPWR VPWR _4902_/A sky130_fd_sc_hd__nand2_8
XFILLER_171_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold177 _5531_/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold188 _6822_/Q VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _5494_/X VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7166_ net399_2/A _7166_/D _6396_/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dfrtp_1
X_4378_ _4360_/B _4379_/B VGND VGND VPWR VPWR _4900_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_1_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6677_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6911_/Q _5973_/A _5948_/X _6951_/Q _6116_/X VGND VGND VPWR VPWR _6117_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3329_ hold47/X hold65/X VGND VGND VPWR VPWR _3373_/B sky130_fd_sc_hd__nand2_8
X_7097_ _7113_/CLK _7097_/D fanout462/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfstp_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6048_ _6812_/Q _5971_/B _5949_/X _6932_/Q _6047_/X VGND VGND VPWR VPWR _6049_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3680_ _6812_/Q _5238_/A hold76/A _7041_/Q VGND VGND VPWR VPWR _3680_/X sky130_fd_sc_hd__a22o_1
X_5350_ _5350_/A0 _5545_/A1 _5354_/S VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput205 _3920_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
Xoutput216 _7180_/X VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
XFILLER_160_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput227 _7189_/X VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
XFILLER_114_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4301_ hold457/X _5544_/A1 _4303_/S VGND VGND VPWR VPWR _4301_/X sky130_fd_sc_hd__mux2_1
Xoutput238 _7197_/X VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
Xoutput249 _3943_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
X_5281_ hold922/X _5548_/A1 _5282_/S VGND VGND VPWR VPWR _5281_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7020_ _7051_/CLK _7020_/D fanout476/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_4
X_4232_ _4232_/A _4322_/B VGND VGND VPWR VPWR _4237_/S sky130_fd_sc_hd__and2_2
X_4163_ _6639_/Q _6307_/B VGND VGND VPWR VPWR _4171_/S sky130_fd_sc_hd__nand2_4
XFILLER_68_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4094_ hold766/X _5519_/A1 _5202_/B VGND VGND VPWR VPWR _4094_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6804_ _7067_/CLK _6804_/D fanout477/X VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4996_ _5021_/A _4996_/B _4996_/C _4996_/D VGND VGND VPWR VPWR _4997_/D sky130_fd_sc_hd__and4_1
X_6735_ _6735_/CLK _6735_/D _3946_/B VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3947_ _6404_/Q _3947_/B VGND VGND VPWR VPWR _3948_/A sky130_fd_sc_hd__nand2b_1
X_6666_ _6668_/CLK _6666_/D fanout452/X VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3878_ hold15/A _6402_/Q _6396_/B VGND VGND VPWR VPWR _3961_/B sky130_fd_sc_hd__o21ai_1
XFILLER_136_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5617_ _6442_/Q _5614_/X _5616_/X _6842_/Q VGND VGND VPWR VPWR _5617_/X sky130_fd_sc_hd__a22o_1
X_6597_ _7137_/CLK _6597_/D VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5548_ hold926/X _5548_/A1 _5549_/S VGND VGND VPWR VPWR _5548_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5479_ hold315/X _5521_/A1 hold30/X VGND VGND VPWR VPWR _5479_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout410 hold156/X VGND VGND VPWR VPWR _5518_/A1 sky130_fd_sc_hd__buf_6
Xfanout421 _6353_/A1 VGND VGND VPWR VPWR _5491_/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout432 hold16/X VGND VGND VPWR VPWR _5505_/B sky130_fd_sc_hd__buf_4
Xfanout454 fanout455/X VGND VGND VPWR VPWR fanout454/X sky130_fd_sc_hd__buf_6
X_7149_ _3937_/A1 _7149_/D fanout487/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout465 fanout466/X VGND VGND VPWR VPWR fanout465/X sky130_fd_sc_hd__buf_8
Xfanout476 fanout485/X VGND VGND VPWR VPWR fanout476/X sky130_fd_sc_hd__buf_8
Xfanout487 _6307_/B VGND VGND VPWR VPWR fanout487/X sky130_fd_sc_hd__buf_8
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4850_ _4456_/A _4843_/B _4689_/Y VGND VGND VPWR VPWR _4850_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3801_ _6978_/Q _5427_/A _3714_/Y _6748_/Q VGND VGND VPWR VPWR _3801_/X sky130_fd_sc_hd__a22o_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _4846_/B _4689_/B _4780_/Y _4627_/A VGND VGND VPWR VPWR _4781_/X sky130_fd_sc_hd__o22a_1
X_6520_ _6777_/CLK _6520_/D fanout484/X VGND VGND VPWR VPWR _7197_/A sky130_fd_sc_hd__dfrtp_1
X_3732_ _6626_/Q _4232_/A _3692_/Y _6766_/Q _3731_/X VGND VGND VPWR VPWR _3732_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6451_ _6677_/CLK _6451_/D fanout452/X VGND VGND VPWR VPWR _6451_/Q sky130_fd_sc_hd__dfrtp_2
X_3663_ _6964_/Q _5409_/A _3381_/Y input26/X _3662_/X VGND VGND VPWR VPWR _3670_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5402_ hold249/X _5465_/A1 _5408_/S VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__mux2_1
X_6382_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6382_/X sky130_fd_sc_hd__and2_1
X_3594_ _6612_/Q _4208_/A _4196_/A _6602_/Q VGND VGND VPWR VPWR _3594_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5333_ hold479/X _5528_/A1 _5336_/S VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5264_ hold679/X _5540_/A1 _5264_/S VGND VGND VPWR VPWR _5264_/X sky130_fd_sc_hd__mux2_1
X_7003_ _7012_/CLK _7003_/D fanout458/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfstp_1
X_4215_ _4215_/A0 _6353_/A1 _4219_/S VGND VGND VPWR VPWR _4215_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5195_ hold547/X _5543_/A1 _5201_/S VGND VGND VPWR VPWR _5195_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4146_ _4146_/A0 hold667/X _4150_/S VGND VGND VPWR VPWR _4146_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4077_ hold158/X hold60/X _4083_/S VGND VGND VPWR VPWR _4077_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4979_ _4626_/Y _4644_/Y _4663_/Y _4782_/Y _4978_/X VGND VGND VPWR VPWR _4981_/C
+ sky130_fd_sc_hd__o221a_1
X_6718_ _7038_/CLK _6718_/D fanout455/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6649_ _6654_/CLK _6649_/D _6383_/A VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6777_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_csclk _7001_/CLK VGND VGND VPWR VPWR _7033_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4000_ _4000_/A0 _5524_/A1 _4007_/S VGND VGND VPWR VPWR _4000_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5951_ _5969_/A _5966_/A _5979_/A VGND VGND VPWR VPWR _5976_/B sky130_fd_sc_hd__and3_4
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _4902_/A _4902_/B VGND VGND VPWR VPWR _5024_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5882_ _6467_/Q _5619_/X _5663_/X _6611_/Q VGND VGND VPWR VPWR _5882_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4833_ _4542_/B _4810_/B _5057_/A _4832_/X VGND VGND VPWR VPWR _4833_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4764_ _4737_/A _4608_/X _4686_/B _4738_/A _4763_/X VGND VGND VPWR VPWR _4764_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_193_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6503_ _6537_/CLK _6503_/D fanout464/X VGND VGND VPWR VPWR _7177_/A sky130_fd_sc_hd__dfrtp_1
X_3715_ _6955_/Q _5400_/A _4157_/A _6566_/Q VGND VGND VPWR VPWR _3715_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4695_ _4716_/A _4969_/A VGND VGND VPWR VPWR _4695_/Y sky130_fd_sc_hd__nand2_4
XFILLER_119_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6434_ _6746_/CLK _6434_/D fanout447/X VGND VGND VPWR VPWR _6434_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_174_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3646_ _6682_/Q _4286_/A _4145_/A _6557_/Q _3645_/X VGND VGND VPWR VPWR _3651_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6365_ _6383_/A _6401_/B VGND VGND VPWR VPWR _6365_/X sky130_fd_sc_hd__and2_1
X_3577_ hold74/X _3577_/B VGND VGND VPWR VPWR _4014_/A sky130_fd_sc_hd__nor2_4
XFILLER_115_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5316_ hold515/X _5538_/A1 _5318_/S VGND VGND VPWR VPWR _5316_/X sky130_fd_sc_hd__mux2_1
X_6296_ _6459_/Q _5944_/X _5975_/A _6603_/Q _6295_/X VGND VGND VPWR VPWR _6300_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5247_ _5247_/A _5541_/B VGND VGND VPWR VPWR _5255_/S sky130_fd_sc_hd__and2_4
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__buf_8
X_5178_ hold359/X _5526_/A1 _5181_/S VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__mux2_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4129_ hold808/X _6354_/A1 _4132_/S VGND VGND VPWR VPWR _4129_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3500_ input7/X _3365_/Y _4280_/A _6679_/Q _3498_/X VGND VGND VPWR VPWR _3504_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4480_ _4615_/B _4653_/C VGND VGND VPWR VPWR _4636_/A sky130_fd_sc_hd__and2_2
Xhold507 _6453_/Q VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _5529_/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 _6608_/Q VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3431_ _3431_/A _3431_/B VGND VGND VPWR VPWR _3447_/A sky130_fd_sc_hd__nor2_2
XFILLER_171_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6150_ _6150_/A _6150_/B _6150_/C _6150_/D VGND VGND VPWR VPWR _6151_/C sky130_fd_sc_hd__nor4_1
X_3362_ _3714_/A _3573_/A VGND VGND VPWR VPWR _5364_/A sky130_fd_sc_hd__nor2_8
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5101_ _4846_/B _4644_/Y _4997_/D _5100_/Y VGND VGND VPWR VPWR _5101_/X sky130_fd_sc_hd__o211a_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6081_ _7059_/Q _5954_/X _5976_/D _6878_/Q VGND VGND VPWR VPWR _6099_/A sky130_fd_sc_hd__a22o_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _6726_/Q _3975_/S VGND VGND VPWR VPWR _3293_/Y sky130_fd_sc_hd__nand2b_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _6426_/Q VGND VGND VPWR VPWR _3982_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _4662_/Y _4695_/Y _4847_/Y _4905_/B _4508_/D VGND VGND VPWR VPWR _5120_/B
+ sky130_fd_sc_hd__o2111a_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _5392_/X VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1229 _7039_/Q VGND VGND VPWR VPWR _5497_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6983_ _6997_/CLK _6983_/D fanout465/X VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5934_ _5966_/A _5968_/A _5981_/B VGND VGND VPWR VPWR _5934_/X sky130_fd_sc_hd__and3_4
XFILLER_179_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5865_ _5864_/Y _5863_/X _6279_/S _5865_/B2 VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_178_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4816_ _4947_/B _4947_/C _4553_/B VGND VGND VPWR VPWR _4816_/Y sky130_fd_sc_hd__a21oi_1
X_5796_ _6880_/Q _5661_/X _5663_/X _6864_/Q _5795_/X VGND VGND VPWR VPWR _5797_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4747_ _4747_/A _4747_/B _4747_/C VGND VGND VPWR VPWR _4926_/B sky130_fd_sc_hd__and3_1
XFILLER_119_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4678_ _4741_/A wire380/X _4660_/X _4648_/X _4942_/B VGND VGND VPWR VPWR _4679_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_162_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6417_ _3945_/A1 _6417_/D _6373_/X VGND VGND VPWR VPWR _6417_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3629_ _7005_/Q _3370_/Y _5490_/A _7037_/Q VGND VGND VPWR VPWR _3629_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6348_ _6644_/Q _6320_/A _6318_/B _6642_/Q VGND VGND VPWR VPWR _6348_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6279_ _6279_/A0 _6278_/X _6279_/S VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__mux2_1
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4336_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_130_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR _3906_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4631_/D sky130_fd_sc_hd__clkbuf_8
XFILLER_102_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6344_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6327_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980_ hold527/X _5513_/A1 _3980_/S VGND VGND VPWR VPWR _3980_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5650_ _5658_/B _5667_/C VGND VGND VPWR VPWR _5651_/B sky130_fd_sc_hd__nand2_8
XFILLER_31_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4601_ _4601_/A _4601_/B VGND VGND VPWR VPWR _4993_/B sky130_fd_sc_hd__nor2_1
X_5581_ _5583_/S _5580_/X _5574_/Y VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__o21a_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4810_/A _4453_/B _4530_/X _4823_/A VGND VGND VPWR VPWR _4533_/D sky130_fd_sc_hd__o211a_1
XFILLER_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold304 _4326_/X VGND VGND VPWR VPWR _6713_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _7024_/Q VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _5367_/X VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ _4911_/A _4856_/A VGND VGND VPWR VPWR _5051_/B sky130_fd_sc_hd__and2_2
Xhold337 _6988_/Q VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _4266_/X VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6189_/Y _6201_/X _6540_/Q _6226_/B VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__o2bb2a_1
Xhold359 _6759_/Q VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ hold85/A _3511_/A VGND VGND VPWR VPWR _3414_/Y sky130_fd_sc_hd__nor2_2
X_7182_ _7182_/A VGND VGND VPWR VPWR _7182_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4394_ _4393_/A _4393_/B _4568_/B VGND VGND VPWR VPWR _4551_/A sky130_fd_sc_hd__o21a_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _7085_/Q _5976_/B _5971_/C _7045_/Q VGND VGND VPWR VPWR _6150_/B sky130_fd_sc_hd__a22o_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3355_/B hold72/X VGND VGND VPWR VPWR _3356_/B sky130_fd_sc_hd__and2_2
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6925_/Q _5938_/X _5952_/X _6957_/Q VGND VGND VPWR VPWR _6064_/X sky130_fd_sc_hd__a22o_1
Xhold1004 _3297_/Y VGND VGND VPWR VPWR _3298_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 _6461_/Q VGND VGND VPWR VPWR _4022_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3276_ hold81/X hold24/X _6488_/Q VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__mux2_1
Xhold1026 _4153_/X VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1037 _6716_/Q VGND VGND VPWR VPWR _4330_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5015_ _4653_/Y _4970_/Y _5010_/Y _4645_/Y _4807_/X VGND VGND VPWR VPWR _5064_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1048 _5322_/X VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 _6901_/Q VGND VGND VPWR VPWR _5341_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6966_ _7083_/CLK _6966_/D fanout476/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5917_ _6564_/Q _5631_/X _5646_/X _6654_/Q VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__a22o_1
X_6897_ _7076_/CLK _6897_/D fanout481/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5848_ _6476_/Q _5630_/X _5634_/X _6451_/Q VGND VGND VPWR VPWR _5848_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5779_ _6960_/Q _5638_/X _5648_/X _6856_/Q VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold860 _6876_/Q VGND VGND VPWR VPWR hold860/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 _4029_/X VGND VGND VPWR VPWR _6467_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 _6975_/Q VGND VGND VPWR VPWR hold882/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold893 _4006_/X VGND VGND VPWR VPWR _6448_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1560 hold70/A VGND VGND VPWR VPWR _3855_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1571 _7170_/Q VGND VGND VPWR VPWR _3235_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1582 _6533_/Q VGND VGND VPWR VPWR hold824/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1593 _6498_/Q VGND VGND VPWR VPWR hold1593/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6820_ _6884_/CLK _6820_/D fanout475/X VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6751_ _7011_/CLK _6751_/D fanout459/X VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_4
X_3963_ hold15/X _3963_/A1 _3963_/S VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__mux2_8
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_5702_ _6964_/Q _5642_/X _5667_/X _6812_/Q VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__a22o_1
X_6682_ _6683_/CLK _6682_/D _6390_/A VGND VGND VPWR VPWR _6682_/Q sky130_fd_sc_hd__dfstp_1
X_3894_ _5552_/B _3887_/Y _3893_/Y _6763_/Q _3894_/B2 VGND VGND VPWR VPWR _6508_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5633_ _6818_/Q _5631_/X _5632_/X _6938_/Q VGND VGND VPWR VPWR _5633_/X sky130_fd_sc_hd__a22o_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5564_ _5564_/A _5564_/B _5564_/C VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__and3_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4515_ _4542_/A _4947_/B VGND VGND VPWR VPWR _4515_/Y sky130_fd_sc_hd__nor2_1
Xhold101 _6724_/Q VGND VGND VPWR VPWR hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _7000_/Q VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ hold235/X hold60/X _5495_/S VGND VGND VPWR VPWR _5495_/X sky130_fd_sc_hd__mux2_1
Xhold123 _3295_/Y VGND VGND VPWR VPWR _3355_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _5176_/X VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _7053_/Q VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold94/X VGND VGND VPWR VPWR hold156/X sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4495_/A _4993_/A VGND VGND VPWR VPWR _4531_/B sky130_fd_sc_hd__nor2_2
Xhold167 _5270_/X VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold178 _7059_/Q VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _5252_/X VGND VGND VPWR VPWR _6822_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7165_ net399_2/A _7165_/D _6395_/X VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__dfrtp_1
X_4377_ _4471_/B _4568_/B VGND VGND VPWR VPWR _4887_/A sky130_fd_sc_hd__nand2_2
XFILLER_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6903_/Q _5976_/C _5971_/D _6831_/Q VGND VGND VPWR VPWR _6116_/X sky130_fd_sc_hd__a22o_1
X_3328_ _3571_/A hold85/X VGND VGND VPWR VPWR _5229_/A sky130_fd_sc_hd__nor2_8
X_7096_ _7113_/CLK _7096_/D fanout462/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfstp_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6444_/Q _5601_/X _5959_/X _6964_/Q VGND VGND VPWR VPWR _6047_/X sky130_fd_sc_hd__a22o_1
X_3259_ _3260_/A1 _3259_/A1 _3260_/S VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__mux2_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6949_ _7085_/CLK _6949_/D fanout477/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold690 _7033_/Q VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1390 _5214_/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput206 _3173_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput217 _3938_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
X_4300_ hold277/X _5534_/A1 _4303_/S VGND VGND VPWR VPWR _4300_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput228 _7190_/X VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5280_ hold780/X _5538_/A1 _5282_/S VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput239 _3925_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4231_ _6624_/Q _3170_/Y _4228_/Y _5006_/A _3168_/A VGND VGND VPWR VPWR _4231_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4162_ hold233/X hold60/X _4162_/S VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4093_ _4093_/A0 _4092_/X _4101_/S VGND VGND VPWR VPWR _4093_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6803_ _7067_/CLK _6803_/D fanout477/X VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4995_ _4995_/A _4995_/B _4995_/C VGND VGND VPWR VPWR _5004_/A sky130_fd_sc_hd__and3_1
XFILLER_168_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6734_ _3945_/A1 _6734_/D _6386_/X VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfrtn_1
X_3946_ _6403_/Q _3946_/B VGND VGND VPWR VPWR _3946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6665_ _6755_/CLK _6665_/D _6360_/A VGND VGND VPWR VPWR _6665_/Q sky130_fd_sc_hd__dfrtp_2
X_3877_ hold15/A _6402_/Q _6396_/B VGND VGND VPWR VPWR _3962_/B sky130_fd_sc_hd__o21a_1
XFILLER_177_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5616_ _5638_/A _5667_/B _5657_/B VGND VGND VPWR VPWR _5616_/X sky130_fd_sc_hd__and3b_4
XFILLER_136_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6596_ _7137_/CLK _6596_/D VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfxtp_1
X_5547_ _5547_/A0 hold42/X _5549_/S VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__mux2_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5478_ hold56/X hold42/X hold30/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__mux2_1
XFILLER_132_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4429_ _4685_/A _4992_/A VGND VGND VPWR VPWR _5068_/A sky130_fd_sc_hd__nand2_2
Xfanout400 hold54/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__buf_8
Xfanout411 _5526_/A1 VGND VGND VPWR VPWR _6355_/A1 sky130_fd_sc_hd__buf_6
Xfanout422 hold666/X VGND VGND VPWR VPWR _6353_/A1 sky130_fd_sc_hd__buf_8
XFILLER_160_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout433 _3178_/Y VGND VGND VPWR VPWR _6303_/S sky130_fd_sc_hd__buf_8
XFILLER_58_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout444 fanout486/X VGND VGND VPWR VPWR _3946_/B sky130_fd_sc_hd__buf_8
X_7148_ _3937_/A1 _7148_/D _6307_/B VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout455 fanout486/X VGND VGND VPWR VPWR fanout455/X sky130_fd_sc_hd__buf_8
Xfanout466 fanout486/X VGND VGND VPWR VPWR fanout466/X sky130_fd_sc_hd__buf_6
Xfanout477 fanout485/X VGND VGND VPWR VPWR fanout477/X sky130_fd_sc_hd__buf_8
Xfanout488 input164/X VGND VGND VPWR VPWR _6307_/B sky130_fd_sc_hd__clkbuf_16
X_7079_ _7079_/CLK _7079_/D fanout478/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ _6614_/Q _4214_/A _4133_/A _6545_/Q _3799_/X VGND VGND VPWR VPWR _3807_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4780_ _4782_/A _4707_/C _4574_/B VGND VGND VPWR VPWR _4780_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _6803_/Q _5229_/A _4172_/A _6579_/Q VGND VGND VPWR VPWR _3731_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_0_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6709_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3662_ _6687_/Q _4292_/A hold67/A _6467_/Q VGND VGND VPWR VPWR _3662_/X sky130_fd_sc_hd__a22o_1
X_6450_ _6677_/CLK _6450_/D fanout452/X VGND VGND VPWR VPWR _6450_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5401_ _5401_/A0 _5524_/A1 _5408_/S VGND VGND VPWR VPWR _5401_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6381_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6381_/X sky130_fd_sc_hd__and2_1
X_3593_ _6901_/Q _5337_/A _5274_/A _6845_/Q _3592_/X VGND VGND VPWR VPWR _3593_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5332_ _5332_/A0 _5545_/A1 _5336_/S VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5263_ hold671/X _5521_/A1 _5264_/S VGND VGND VPWR VPWR _5263_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7002_ _7006_/CLK _7002_/D fanout458/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfstp_1
X_4214_ _4214_/A _4322_/B VGND VGND VPWR VPWR _4219_/S sky130_fd_sc_hd__and2_2
X_5194_ _5194_/A0 _5473_/A1 _5201_/S VGND VGND VPWR VPWR _5194_/X sky130_fd_sc_hd__mux2_1
X_4145_ _4145_/A _4322_/B VGND VGND VPWR VPWR _4150_/S sky130_fd_sc_hd__and2_2
X_4076_ _4076_/A0 hold95/X _4084_/S VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__mux2_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4978_ _4639_/Y _4692_/Y _4969_/Y _4663_/Y VGND VGND VPWR VPWR _4978_/X sky130_fd_sc_hd__o22a_1
X_6717_ _7038_/CLK _6717_/D fanout455/X VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfstp_1
X_3929_ _6504_/Q input77/X _3956_/B VGND VGND VPWR VPWR _3929_/X sky130_fd_sc_hd__mux2_4
XFILLER_20_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6648_ _6671_/CLK _6648_/D fanout468/X VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6579_ _6677_/CLK _6579_/D fanout452/X VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5950_ _6946_/Q _5948_/X _5949_/X _6930_/Q VGND VGND VPWR VPWR _5950_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4901_ _4491_/Y _4900_/Y _4707_/Y _4498_/Y VGND VGND VPWR VPWR _5080_/A sky130_fd_sc_hd__o211a_1
X_5881_ _6601_/Q _5616_/X _5880_/X VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4832_ _4948_/A _4810_/B _5092_/A _4831_/X VGND VGND VPWR VPWR _4832_/X sky130_fd_sc_hd__o211a_1
XANTENNA_190 _5513_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4763_ _4921_/A _4737_/A _4668_/C _4671_/A VGND VGND VPWR VPWR _4763_/X sky130_fd_sc_hd__a31o_1
XFILLER_159_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6502_ _6539_/CLK _6502_/D fanout461/X VGND VGND VPWR VPWR _7176_/A sky130_fd_sc_hd__dfrtp_1
X_3714_ _3714_/A _3714_/B VGND VGND VPWR VPWR _3714_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4694_ _4716_/A _4782_/A VGND VGND VPWR VPWR _4694_/Y sky130_fd_sc_hd__nand2_4
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6433_ _6749_/CLK _6433_/D fanout449/X VGND VGND VPWR VPWR _6433_/Q sky130_fd_sc_hd__dfstp_4
X_3645_ input37/X _3331_/Y _4202_/A _6606_/Q VGND VGND VPWR VPWR _3645_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3576_ _6982_/Q _5427_/A _5490_/A _7038_/Q _3574_/X VGND VGND VPWR VPWR _3580_/C
+ sky130_fd_sc_hd__a221o_1
X_6364_ _6383_/A _6401_/B VGND VGND VPWR VPWR _6364_/X sky130_fd_sc_hd__and2_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5315_ hold465/X _5528_/A1 _5318_/S VGND VGND VPWR VPWR _5315_/X sky130_fd_sc_hd__mux2_1
X_6295_ _6469_/Q _5937_/X _5975_/D _6629_/Q VGND VGND VPWR VPWR _6295_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5246_ hold762/X _5540_/A1 _5246_/S VGND VGND VPWR VPWR _5246_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__buf_6
XFILLER_130_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5177_ hold209/X _5494_/A1 _5181_/S VGND VGND VPWR VPWR _5177_/X sky130_fd_sc_hd__mux2_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4128_ _4128_/A0 _5491_/A1 _4132_/S VGND VGND VPWR VPWR _4128_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4059_ hold997/X _4058_/X _4067_/S VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6755_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold508 _4012_/X VGND VGND VPWR VPWR _6453_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3430_ _5182_/S _3417_/X _3426_/X _3428_/X _3429_/X VGND VGND VPWR VPWR _3431_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold519 _6682_/Q VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3361_ _3562_/A hold48/X VGND VGND VPWR VPWR _5265_/A sky130_fd_sc_hd__nor2_8
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _4992_/A _4737_/A _4735_/X _4588_/Y VGND VGND VPWR VPWR _5100_/Y sky130_fd_sc_hd__a31oi_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6080_ _7006_/Q _5958_/X _5978_/X _6998_/Q VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__a22o_1
X_3292_ _3292_/A _6488_/Q VGND VGND VPWR VPWR _3292_/X sky130_fd_sc_hd__and2_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _4542_/A _4902_/A _4695_/Y _4627_/B _4872_/D VGND VGND VPWR VPWR _5033_/C
+ sky130_fd_sc_hd__o221a_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _3982_/X VGND VGND VPWR VPWR _6426_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1219 _7047_/Q VGND VGND VPWR VPWR _5506_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6982_ _7065_/CLK _6982_/D fanout465/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfrtp_2
X_5933_ _5966_/A _5979_/A _5981_/B VGND VGND VPWR VPWR _5971_/A sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7086_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5864_ _5552_/B _7114_/Q _6103_/B1 VGND VGND VPWR VPWR _5864_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_178_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4815_ _4947_/C _4553_/B _5041_/A VGND VGND VPWR VPWR _4815_/Y sky130_fd_sc_hd__o21ai_1
X_5795_ _7024_/Q _5619_/X _5666_/X _6896_/Q VGND VGND VPWR VPWR _5795_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_csclk _7001_/CLK VGND VGND VPWR VPWR _6981_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4746_ _4948_/A _4581_/B _4611_/Y _4645_/Y VGND VGND VPWR VPWR _4942_/C sky130_fd_sc_hd__o22a_1
XFILLER_193_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4677_ _4500_/A _4902_/B _4535_/A _5021_/A VGND VGND VPWR VPWR _4679_/C sky130_fd_sc_hd__o211a_1
XFILLER_162_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6416_ _3927_/A1 _6416_/D _6372_/X VGND VGND VPWR VPWR _6416_/Q sky130_fd_sc_hd__dfrtp_2
X_3628_ _3628_/A _3628_/B _3628_/C _3628_/D VGND VGND VPWR VPWR _3639_/B sky130_fd_sc_hd__nor4_1
XFILLER_162_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6347_ _6347_/A1 _4228_/Y _4229_/X _3910_/A VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__o211a_2
X_3559_ _3714_/B _3814_/B VGND VGND VPWR VPWR _4133_/A sky130_fd_sc_hd__nor2_8
XFILLER_163_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6278_ _6278_/A0 _6277_/X _6303_/S VGND VGND VPWR VPWR _6278_/X sky130_fd_sc_hd__mux2_1
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4335_/B sky130_fd_sc_hd__clkbuf_1
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR _3900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4633_/B sky130_fd_sc_hd__buf_4
XFILLER_88_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5229_ _5229_/A _5541_/B VGND VGND VPWR VPWR _5237_/S sky130_fd_sc_hd__and2_4
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6323_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _6558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_79_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4600_ _4739_/A _4600_/B _4747_/B _4739_/B VGND VGND VPWR VPWR _4601_/B sky130_fd_sc_hd__nand4b_1
X_5580_ _7094_/Q _5576_/B _7095_/Q VGND VGND VPWR VPWR _5580_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4531_ _4810_/A _4531_/B VGND VGND VPWR VPWR _4823_/A sky130_fd_sc_hd__nand2b_1
XFILLER_184_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold305 _6915_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 _5479_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4462_ _4896_/A _4462_/B VGND VGND VPWR VPWR _4856_/A sky130_fd_sc_hd__and2_1
Xhold327 _6857_/Q VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _5439_/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 hold349/A VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _6192_/X _6201_/B _6226_/B VGND VGND VPWR VPWR _6201_/X sky130_fd_sc_hd__and3b_1
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3413_ _3412_/X _3413_/A1 _3829_/B VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7181_ _7181_/A VGND VGND VPWR VPWR _7181_/X sky130_fd_sc_hd__clkbuf_1
X_4393_ _4393_/A _4393_/B VGND VGND VPWR VPWR _4552_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3374_/A hold48/X VGND VGND VPWR VPWR _5337_/A sky130_fd_sc_hd__nor2_8
X_6132_ _7061_/Q _5954_/X _5976_/D _6880_/Q VGND VGND VPWR VPWR _6150_/A sky130_fd_sc_hd__a22o_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6063_ _6973_/Q _5947_/X _5965_/X _6797_/Q _6062_/X VGND VGND VPWR VPWR _6066_/B
+ sky130_fd_sc_hd__a221o_1
X_3275_ hold46/X hold26/X VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__and2b_4
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _3298_/Y VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 _4022_/X VGND VGND VPWR VPWR _6461_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1027 _6601_/Q VGND VGND VPWR VPWR _4199_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 _4330_/X VGND VGND VPWR VPWR _6716_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5014_ _4628_/Y _5010_/Y _4982_/X _4796_/A VGND VGND VPWR VPWR _5018_/C sky130_fd_sc_hd__o211a_1
Xhold1049 _6844_/Q VGND VGND VPWR VPWR _5277_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7080_/CLK _6965_/D fanout479/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfrtp_4
X_5916_ _6719_/Q _5642_/X _5666_/X _6634_/Q VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__a22o_1
X_6896_ _7069_/CLK _6896_/D fanout482/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _6600_/Q _5616_/X _5648_/X _6605_/Q _5846_/X VGND VGND VPWR VPWR _5852_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5778_ _5778_/A1 _6279_/S _5776_/X _5777_/X VGND VGND VPWR VPWR _5778_/X sky130_fd_sc_hd__o22a_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4729_ _4964_/A _4725_/Y _4728_/X _4229_/X VGND VGND VPWR VPWR _4729_/X sky130_fd_sc_hd__a211o_1
XFILLER_108_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold850 _6804_/Q VGND VGND VPWR VPWR hold850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _5313_/X VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold872 _7020_/Q VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _5424_/X VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 _7032_/Q VGND VGND VPWR VPWR hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1550 _6641_/Q VGND VGND VPWR VPWR _3168_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1561 _7159_/Q VGND VGND VPWR VPWR _3912_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1572 _7116_/Q VGND VGND VPWR VPWR _5887_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1583 _6412_/Q VGND VGND VPWR VPWR _3852_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1594 _7176_/A VGND VGND VPWR VPWR hold349/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6750_ _7006_/CLK _6750_/D fanout457/X VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfstp_1
X_3962_ _3962_/A _3962_/B VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__nor2_1
X_5701_ _6852_/Q _5648_/X _5666_/X _6892_/Q _5700_/X VGND VGND VPWR VPWR _5706_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6681_ _6714_/CLK _6681_/D fanout470/X VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_4
X_3893_ _5959_/A _5966_/A VGND VGND VPWR VPWR _3893_/Y sky130_fd_sc_hd__nand2_1
X_5632_ _5638_/A _5667_/B _5667_/C VGND VGND VPWR VPWR _5632_/X sky130_fd_sc_hd__and3_4
XFILLER_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5563_ _7088_/Q _7089_/Q _5562_/D _7090_/Q VGND VGND VPWR VPWR _5564_/C sky130_fd_sc_hd__a31o_1
XFILLER_129_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4514_ _4514_/A _4514_/B _4514_/C VGND VGND VPWR VPWR _4518_/D sky130_fd_sc_hd__and3_1
Xhold102 _3287_/Y VGND VGND VPWR VPWR _3356_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _5452_/X VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ hold198/X _5494_/A1 _5495_/S VGND VGND VPWR VPWR _5494_/X sky130_fd_sc_hd__mux2_1
Xhold124 _3300_/Y VGND VGND VPWR VPWR _3571_/A sky130_fd_sc_hd__buf_12
Xhold135 _6840_/Q VGND VGND VPWR VPWR hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold146 _5512_/X VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4556_/A _4611_/B VGND VGND VPWR VPWR _5051_/A sky130_fd_sc_hd__and2_2
Xhold157 _4030_/X VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _6783_/Q VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _5519_/X VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_113_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7164_ net399_2/A _7164_/D _6394_/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfrtp_1
X_4376_ _4376_/A _4376_/B _4568_/B VGND VGND VPWR VPWR _4465_/B sky130_fd_sc_hd__and3_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6115_ _6115_/A _6115_/B _6115_/C VGND VGND VPWR VPWR _6126_/C sky130_fd_sc_hd__nor3_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3327_ hold47/X hold84/X VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__nand2_8
X_7095_ _7113_/CLK _7095_/D fanout462/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6046_ _7020_/Q _5937_/X _5975_/D _6884_/Q _6029_/X VGND VGND VPWR VPWR _6049_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3258_ _3259_/A1 hold93/A _3260_/S VGND VGND VPWR VPWR _3258_/X sky130_fd_sc_hd__mux2_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _7058_/Q VGND VGND VPWR VPWR _3189_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6948_ _7065_/CLK _6948_/D fanout463/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6879_ _7078_/CLK _6879_/D fanout481/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold680 _5264_/X VGND VGND VPWR VPWR _6833_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _5489_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1380 _6531_/Q VGND VGND VPWR VPWR _4117_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1391 _6654_/Q VGND VGND VPWR VPWR _4255_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3219_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
Xoutput218 _7181_/X VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
Xoutput229 _7191_/X VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
XFILLER_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ _6640_/Q _4230_/B VGND VGND VPWR VPWR _5006_/A sky130_fd_sc_hd__nand2b_2
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4161_ hold736/X _6356_/A1 _4162_/S VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4092_ hold904/X _5509_/A1 _5202_/B VGND VGND VPWR VPWR _4092_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6802_ _7051_/CLK _6802_/D fanout476/X VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_36_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4994_ _4413_/Y _4428_/Y _4621_/X VGND VGND VPWR VPWR _4995_/C sky130_fd_sc_hd__o21a_1
X_6733_ _3927_/A1 _6733_/D _6385_/X VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfrtn_1
X_3945_ input83/X _3945_/A1 _6403_/Q VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__mux2_1
X_6664_ _6712_/CLK _6664_/D _6396_/A VGND VGND VPWR VPWR _6664_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3876_ _6485_/Q _3867_/B _3875_/X _6487_/Q VGND VGND VPWR VPWR _6485_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5615_ _7095_/Q _7094_/Q VGND VGND VPWR VPWR _5657_/B sky130_fd_sc_hd__and2b_2
XFILLER_137_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6595_ _7137_/CLK _6595_/D VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5546_ hold816/X _5546_/A1 _5549_/S VGND VGND VPWR VPWR _5546_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5477_ hold455/X _5528_/A1 hold30/X VGND VGND VPWR VPWR _5477_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4428_ _4753_/A _4607_/A _4600_/B VGND VGND VPWR VPWR _4428_/Y sky130_fd_sc_hd__nand3b_4
Xfanout401 hold60/X VGND VGND VPWR VPWR _6357_/A1 sky130_fd_sc_hd__buf_8
Xfanout412 _5526_/A1 VGND VGND VPWR VPWR _5493_/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR net399_2/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout423 hold666/X VGND VGND VPWR VPWR _5524_/A1 sky130_fd_sc_hd__buf_6
Xfanout434 _5638_/A VGND VGND VPWR VPWR _5664_/A sky130_fd_sc_hd__buf_4
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7147_ _3937_/A1 _7147_/D _6307_/B VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout445 _6360_/A VGND VGND VPWR VPWR fanout445/X sky130_fd_sc_hd__buf_8
X_4359_ _4382_/B _4359_/B VGND VGND VPWR VPWR _4359_/Y sky130_fd_sc_hd__nand2_2
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout456 fanout466/X VGND VGND VPWR VPWR fanout456/X sky130_fd_sc_hd__buf_8
Xfanout467 fanout469/X VGND VGND VPWR VPWR _6383_/A sky130_fd_sc_hd__buf_6
Xfanout478 fanout480/X VGND VGND VPWR VPWR fanout478/X sky130_fd_sc_hd__buf_8
X_7078_ _7078_/CLK _7078_/D fanout485/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout489 _4625_/A VGND VGND VPWR VPWR _4607_/A sky130_fd_sc_hd__buf_12
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6029_ _7028_/Q _5944_/X _5975_/A _6844_/Q VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _3730_/A _3730_/B _3730_/C VGND VGND VPWR VPWR _3762_/A sky130_fd_sc_hd__and3_1
XFILLER_158_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3661_ _3661_/A _3661_/B _3661_/C _3661_/D VGND VGND VPWR VPWR _3661_/Y sky130_fd_sc_hd__nor4_1
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5400_ _5400_/A hold17/X VGND VGND VPWR VPWR _5408_/S sky130_fd_sc_hd__and2_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6380_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6380_/X sky130_fd_sc_hd__and2_1
X_3592_ _6877_/Q _5310_/A _5319_/A _6885_/Q VGND VGND VPWR VPWR _3592_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ hold868/X _5484_/A1 _5336_/S VGND VGND VPWR VPWR _5331_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5262_ hold790/X _5538_/A1 _5264_/S VGND VGND VPWR VPWR _5262_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7001_ _7001_/CLK _7001_/D fanout464/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4213_ hold447/X _6357_/A1 _4213_/S VGND VGND VPWR VPWR _4213_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5193_ _5193_/A _5541_/B VGND VGND VPWR VPWR _5201_/S sky130_fd_sc_hd__and2_2
X_4144_ hold944/X _5546_/A1 _4144_/S VGND VGND VPWR VPWR _4144_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4075_ _6535_/Q hold94/X _4083_/S VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__mux2_1
XFILLER_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_4_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _6601_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4977_ _4631_/Y _4689_/B _4970_/Y VGND VGND VPWR VPWR _4981_/B sky130_fd_sc_hd__a21o_1
X_6716_ _7038_/CLK _6716_/D fanout455/X VGND VGND VPWR VPWR _6716_/Q sky130_fd_sc_hd__dfrtp_4
X_3928_ _6510_/Q _3268_/C _6406_/Q VGND VGND VPWR VPWR _3928_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6647_ _6671_/CLK _6647_/D _6383_/A VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_20_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3859_ hold44/A _6488_/Q _3851_/C hold24/A VGND VGND VPWR VPWR _3861_/A sky130_fd_sc_hd__o211a_1
XFILLER_137_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6578_ _6709_/CLK _6578_/D fanout445/X VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5529_ hold517/X _5538_/A1 _5531_/S VGND VGND VPWR VPWR _5529_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4900_ _4900_/A _4900_/B VGND VGND VPWR VPWR _4900_/Y sky130_fd_sc_hd__nand2_1
X_5880_ _6472_/Q _5627_/X _5635_/X _6567_/Q VGND VGND VPWR VPWR _5880_/X sky130_fd_sc_hd__a22o_1
X_4831_ _4542_/D _4810_/B _4824_/X _4830_/X VGND VGND VPWR VPWR _4831_/X sky130_fd_sc_hd__o211a_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_180 _6542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 _5494_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4762_ _4627_/A _4627_/B _4611_/Y _4581_/B _4542_/A VGND VGND VPWR VPWR _4769_/C
+ sky130_fd_sc_hd__o32a_1
X_6501_ _6539_/CLK hold96/X fanout459/X VGND VGND VPWR VPWR _7175_/A sky130_fd_sc_hd__dfrtp_1
X_3713_ input62/X _4102_/A _4244_/A _6646_/Q _3712_/X VGND VGND VPWR VPWR _3720_/B
+ sky130_fd_sc_hd__a221o_2
X_4693_ _4881_/A _4630_/X _4753_/C _4975_/B _4689_/Y VGND VGND VPWR VPWR _4693_/X
+ sky130_fd_sc_hd__a221o_1
X_6432_ _6749_/CLK _6432_/D fanout449/X VGND VGND VPWR VPWR _6432_/Q sky130_fd_sc_hd__dfstp_2
X_3644_ _6876_/Q _5310_/A _3964_/A _6420_/Q _3643_/X VGND VGND VPWR VPWR _3651_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6363_ _6383_/A _6401_/B VGND VGND VPWR VPWR _6363_/X sky130_fd_sc_hd__and2_1
X_3575_ hold75/X _3692_/A VGND VGND VPWR VPWR _5490_/A sky130_fd_sc_hd__nor2_4
X_5314_ hold628/X _5509_/A1 _5318_/S VGND VGND VPWR VPWR _5314_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6294_ _6684_/Q _5934_/X _5975_/B _6618_/Q _6293_/X VGND VGND VPWR VPWR _6300_/A
+ sky130_fd_sc_hd__a221o_1
X_5245_ hold920/X _5548_/A1 _5246_/S VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__buf_8
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__buf_12
X_5176_ hold133/X hold60/X _5181_/S VGND VGND VPWR VPWR _5176_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4127_ _4127_/A _6352_/B VGND VGND VPWR VPWR _4132_/S sky130_fd_sc_hd__and2_2
XFILLER_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4058_ hold692/X _5509_/A1 _4058_/S VGND VGND VPWR VPWR _4058_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold509 _6633_/Q VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__dlygate4sd3_1
X_3360_ hold48/X hold75/A VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__nor2_8
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3291_ hold34/X VGND VGND VPWR VPWR _3295_/A sky130_fd_sc_hd__inv_2
XFILLER_151_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _4542_/A _4902_/A _4628_/Y _4691_/A _4852_/X VGND VGND VPWR VPWR _5131_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1209 _6794_/Q VGND VGND VPWR VPWR _5221_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6981_ _6981_/CLK _6981_/D fanout463/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5932_ _7100_/Q _7099_/Q VGND VGND VPWR VPWR _5981_/B sky130_fd_sc_hd__nor2_4
XFILLER_34_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5863_ _3184_/Y _5651_/Y _5852_/Y _5862_/Y _5552_/B VGND VGND VPWR VPWR _5863_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4814_ _4886_/B _4958_/B VGND VGND VPWR VPWR _5089_/A sky130_fd_sc_hd__nand2_1
X_5794_ _6968_/Q _5642_/X _5905_/A2 _6800_/Q _5793_/X VGND VGND VPWR VPWR _5797_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4745_ _4456_/Y _4672_/B _4626_/Y _4639_/Y VGND VGND VPWR VPWR _4768_/A sky130_fd_sc_hd__o22a_1
XFILLER_193_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4676_ _4737_/A _4676_/B VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6415_ _3945_/A1 _6415_/D _6371_/X VGND VGND VPWR VPWR _6415_/Q sky130_fd_sc_hd__dfrtp_2
X_3627_ input6/X _3365_/Y _3381_/Y input29/X _3626_/X VGND VGND VPWR VPWR _3628_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6346_ _6345_/X _6346_/A1 _6346_/S VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__mux2_1
X_3558_ hold35/X _3573_/B VGND VGND VPWR VPWR _4274_/A sky130_fd_sc_hd__nor2_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6277_ _6543_/Q _6226_/B _6276_/X VGND VGND VPWR VPWR _6277_/X sky130_fd_sc_hd__o21ba_1
XFILLER_88_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3489_ _3554_/A _3573_/B VGND VGND VPWR VPWR _4232_/A sky130_fd_sc_hd__nor2_4
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4335_/A sky130_fd_sc_hd__clkbuf_1
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__clkbuf_1
X_5228_ hold687/X _5513_/A1 _5228_/S VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__mux2_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4337_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5159_ hold553/X _6357_/A1 _5160_/S VGND VGND VPWR VPWR _5159_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_80 _6869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _6558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4530_ _4413_/Y _4453_/B _4528_/X _4529_/Y VGND VGND VPWR VPWR _4530_/X sky130_fd_sc_hd__o211a_1
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold306 _5357_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _4690_/B _4611_/B VGND VGND VPWR VPWR _4902_/B sky130_fd_sc_hd__nand2_8
Xhold317 _6558_/Q VGND VGND VPWR VPWR hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold328 _5291_/X VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6200_ _6200_/A _6200_/B _6200_/C _6200_/D VGND VGND VPWR VPWR _6200_/Y sky130_fd_sc_hd__nor4_1
Xhold339 _7182_/A VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ _3410_/Y _3449_/A1 _3829_/A VGND VGND VPWR VPWR _3412_/X sky130_fd_sc_hd__mux2_1
X_7180_ _7180_/A VGND VGND VPWR VPWR _7180_/X sky130_fd_sc_hd__clkbuf_2
X_4392_ _4566_/A _4564_/A _4392_/C VGND VGND VPWR VPWR _4393_/B sky130_fd_sc_hd__and3_1
XFILLER_131_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _7008_/Q _5958_/X _5978_/X _7000_/Q VGND VGND VPWR VPWR _6131_/X sky130_fd_sc_hd__a22o_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3573_/A hold28/X VGND VGND VPWR VPWR _5400_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6893_/Q _5946_/X _5955_/X _6805_/Q VGND VGND VPWR VPWR _6062_/X sky130_fd_sc_hd__a22o_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3274_ hold45/X _6720_/Q _3975_/S VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__mux2_2
XFILLER_39_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _3355_/X VGND VGND VPWR VPWR _5171_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1017 _6579_/Q VGND VGND VPWR VPWR _4174_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _4619_/Y _4970_/Y _5010_/Y _4616_/Y _4796_/C VGND VGND VPWR VPWR _5106_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1028 _4199_/X VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 hold1598/X VGND VGND VPWR VPWR _4061_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6964_ _7006_/CLK _6964_/D fanout458/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5915_ _6469_/Q _5619_/X _5663_/X _6613_/Q _5914_/X VGND VGND VPWR VPWR _5915_/X
+ sky130_fd_sc_hd__a221o_1
X_6895_ _7076_/CLK _6895_/D fanout481/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_4
X_5846_ _6466_/Q _5619_/X _5663_/X _6610_/Q VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5777_ _6507_/Q _7110_/Q _6103_/B1 VGND VGND VPWR VPWR _5777_/X sky130_fd_sc_hd__a21o_1
X_4728_ _5039_/A _4964_/A _4727_/X VGND VGND VPWR VPWR _4728_/X sky130_fd_sc_hd__o21ba_1
XFILLER_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4659_ _4846_/B _4644_/Y _4646_/Y _4657_/X _4658_/X VGND VGND VPWR VPWR _4660_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold840 _7035_/Q VGND VGND VPWR VPWR hold840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 _5232_/X VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold862 _6900_/Q VGND VGND VPWR VPWR hold862/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _5475_/X VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 _6736_/Q VGND VGND VPWR VPWR hold884/X sky130_fd_sc_hd__dlygate4sd3_1
X_6329_ _6642_/Q _6329_/A2 _6329_/B1 _4230_/B VGND VGND VPWR VPWR _6329_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold895 _5488_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1540 _6351_/X VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 _4231_/X VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1562 _7113_/Q VGND VGND VPWR VPWR _5821_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1573 _6761_/Q VGND VGND VPWR VPWR hold129/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1584 _7197_/A VGND VGND VPWR VPWR hold237/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1595 _6725_/Q VGND VGND VPWR VPWR _5113_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7069_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_47_csclk _7001_/CLK VGND VGND VPWR VPWR _6997_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ _6644_/Q _3961_/B VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__and2_1
XFILLER_16_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5700_ _6900_/Q _5621_/X _5658_/X _6884_/Q VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__a22o_1
XFILLER_189_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6680_ _6683_/CLK _6680_/D _6390_/A VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfrtp_4
X_3892_ _5600_/A _7102_/Q VGND VGND VPWR VPWR _5966_/A sky130_fd_sc_hd__and2_2
X_5631_ _5664_/A _5658_/B _5657_/B VGND VGND VPWR VPWR _5631_/X sky130_fd_sc_hd__and3b_4
X_5562_ _7088_/Q _7089_/Q _7090_/Q _5562_/D VGND VGND VPWR VPWR _5564_/B sky130_fd_sc_hd__nand4_1
XFILLER_191_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4513_ _4902_/A _4453_/B _4542_/A VGND VGND VPWR VPWR _4514_/C sky130_fd_sc_hd__a21o_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5493_ _5493_/A0 _5493_/A1 _5495_/S VGND VGND VPWR VPWR _5493_/X sky130_fd_sc_hd__mux2_1
Xhold103 _3511_/A VGND VGND VPWR VPWR _3717_/B sky130_fd_sc_hd__buf_6
XFILLER_144_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold114 _6928_/Q VGND VGND VPWR VPWR hold114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 hold125/A VGND VGND VPWR VPWR _3562_/A sky130_fd_sc_hd__buf_12
XFILLER_144_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold136 _5272_/X VGND VGND VPWR VPWR _6840_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4444_ _4607_/A _4753_/A VGND VGND VPWR VPWR _4993_/A sky130_fd_sc_hd__nand2b_4
Xhold147 _6982_/Q VGND VGND VPWR VPWR hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 hold158/A VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _5208_/X VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ net399_2/A _7163_/D _6393_/X VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__dfrtp_1
X_4375_ _4334_/B _4334_/C _4374_/A _4372_/X VGND VGND VPWR VPWR _4568_/B sky130_fd_sc_hd__a31o_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6983_/Q _5945_/X _5975_/C _6839_/Q _6113_/X VGND VGND VPWR VPWR _6115_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3326_ _3562_/A _3714_/A VGND VGND VPWR VPWR _3326_/Y sky130_fd_sc_hd__nor2_8
X_7094_ _7113_/CLK _7094_/D fanout462/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _7065_/Q _5934_/X _5975_/B _6868_/Q _6044_/X VGND VGND VPWR VPWR _6045_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ hold93/A _3257_/A1 _3260_/S VGND VGND VPWR VPWR _3257_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3188_ _7066_/Q VGND VGND VPWR VPWR _3188_/Y sky130_fd_sc_hd__inv_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6947_ _7011_/CLK hold10/X fanout456/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfstp_4
X_6878_ _7051_/CLK _6878_/D fanout476/X VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5829_ _6460_/Q _5624_/X _5654_/X _6675_/Q _5822_/Y VGND VGND VPWR VPWR _5829_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold670 _5299_/X VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 _6889_/Q VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 hold692/A VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1370 hold1370/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
XFILLER_18_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1381 _6526_/Q VGND VGND VPWR VPWR _4112_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1392 _4255_/X VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput208 _3218_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XFILLER_153_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput219 _7182_/X VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ _4160_/A0 _5493_/A1 _4162_/S VGND VGND VPWR VPWR _4160_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4091_ _4091_/A0 _4090_/X _4101_/S VGND VGND VPWR VPWR _4091_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6801_ _7053_/CLK _6801_/D fanout459/X VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4993_ _4993_/A _4993_/B VGND VGND VPWR VPWR _5069_/C sky130_fd_sc_hd__nand2_1
X_3944_ _6404_/Q _3946_/B VGND VGND VPWR VPWR _3944_/Y sky130_fd_sc_hd__nor2_1
X_6732_ _3945_/A1 _6732_/D _6384_/X VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_177_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6663_ _7058_/CLK _6663_/D _6396_/A VGND VGND VPWR VPWR _6663_/Q sky130_fd_sc_hd__dfstp_2
X_3875_ _7167_/Q _3875_/B _3875_/C VGND VGND VPWR VPWR _3875_/X sky130_fd_sc_hd__and3_1
XFILLER_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5614_ _5638_/A _5667_/B _5666_/B VGND VGND VPWR VPWR _5614_/X sky130_fd_sc_hd__and3_4
XFILLER_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6594_ _7130_/CLK _6594_/D VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5545_ _5545_/A0 _5545_/A1 _5549_/S VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_145_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5476_ _5476_/A0 _5545_/A1 hold30/X VGND VGND VPWR VPWR _5476_/X sky130_fd_sc_hd__mux2_1
X_4427_ _4561_/B _4632_/B VGND VGND VPWR VPWR _4992_/A sky130_fd_sc_hd__nor2_4
XFILLER_99_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout402 hold59/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__buf_12
Xfanout413 hold6/X VGND VGND VPWR VPWR _5526_/A1 sky130_fd_sc_hd__buf_8
X_7146_ _3937_/A1 _7146_/D _6307_/B VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfrtp_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout424 hold666/X VGND VGND VPWR VPWR hold667/A sky130_fd_sc_hd__buf_8
X_4358_ _4739_/A _4356_/B _4357_/B _4661_/A VGND VGND VPWR VPWR _4359_/B sky130_fd_sc_hd__a2bb2o_1
Xfanout435 _5899_/B VGND VGND VPWR VPWR _5638_/A sky130_fd_sc_hd__clkbuf_4
Xfanout446 fanout486/X VGND VGND VPWR VPWR _6360_/A sky130_fd_sc_hd__buf_6
XFILLER_101_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout457 fanout466/X VGND VGND VPWR VPWR fanout457/X sky130_fd_sc_hd__buf_8
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout468 fanout469/X VGND VGND VPWR VPWR fanout468/X sky130_fd_sc_hd__buf_4
X_3309_ hold27/X hold65/X VGND VGND VPWR VPWR _3370_/A sky130_fd_sc_hd__nand2_8
X_7077_ _7086_/CLK _7077_/D fanout483/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4289_ hold519/X _5544_/A1 _4291_/S VGND VGND VPWR VPWR _4289_/X sky130_fd_sc_hd__mux2_1
Xfanout479 fanout480/X VGND VGND VPWR VPWR fanout479/X sky130_fd_sc_hd__buf_8
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6028_ _6028_/A0 _6027_/X _6279_/S VGND VGND VPWR VPWR _6028_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3660_ _7073_/Q _5532_/A _5148_/A _6739_/Q _3659_/X VGND VGND VPWR VPWR _3661_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3591_ _6617_/Q _4214_/A _4238_/A _6633_/Q VGND VGND VPWR VPWR _3591_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5330_ hold549/X _5543_/A1 _5336_/S VGND VGND VPWR VPWR _5330_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5261_ hold190/X _5519_/A1 _5264_/S VGND VGND VPWR VPWR _5261_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7000_ _7017_/CLK _7000_/D fanout461/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4212_ hold493/X _5518_/A1 _4213_/S VGND VGND VPWR VPWR _4212_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5192_ hold423/X _5534_/A1 _5192_/S VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4143_ hold505/X _5518_/A1 _4144_/S VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4074_ hold170/X _4073_/X _4084_/S VGND VGND VPWR VPWR _4074_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4976_ _4576_/Y _4701_/Y _4975_/Y _4613_/Y VGND VGND VPWR VPWR _4981_/A sky130_fd_sc_hd__o22a_1
X_6715_ _7038_/CLK _6715_/D fanout455/X VGND VGND VPWR VPWR _6715_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3927_ _6511_/Q _3927_/A1 _6405_/Q VGND VGND VPWR VPWR _3927_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3858_ _3858_/A1 _3851_/C _3857_/X VGND VGND VPWR VPWR _6410_/D sky130_fd_sc_hd__o21a_1
X_6646_ _6671_/CLK _6646_/D fanout468/X VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3789_ _5186_/A _3355_/X _3788_/Y hold49/A _7026_/Q VGND VGND VPWR VPWR _3789_/X
+ sky130_fd_sc_hd__a32o_1
X_6577_ _7140_/CLK _6577_/D VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5528_ hold435/X _5528_/A1 _5531_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ hold110/X hold60/X _5461_/S VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7129_ _7130_/CLK _7129_/D fanout486/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4830_ _4542_/A _4810_/B _4821_/X _4828_/X _4829_/X VGND VGND VPWR VPWR _4830_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _4108_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_181 _6925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_192 _5544_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _4627_/A _4615_/Y _4626_/Y _4810_/A _4672_/B VGND VGND VPWR VPWR _4772_/C
+ sky130_fd_sc_hd__o32a_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6500_ _6539_/CLK _6500_/D fanout461/X VGND VGND VPWR VPWR _7174_/A sky130_fd_sc_hd__dfrtp_1
X_3712_ _7019_/Q hold29/A _5256_/A _6827_/Q VGND VGND VPWR VPWR _3712_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4692_ _4975_/B VGND VGND VPWR VPWR _4692_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6431_ _6749_/CLK _6431_/D fanout449/X VGND VGND VPWR VPWR _6431_/Q sky130_fd_sc_hd__dfstp_2
X_3643_ _6972_/Q _5418_/A _4058_/S input45/X VGND VGND VPWR VPWR _3643_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6362_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6362_/X sky130_fd_sc_hd__and2_1
X_3574_ _6990_/Q _5436_/A _4304_/A _6699_/Q VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__a22o_1
X_5313_ hold860/X _5484_/A1 _5318_/S VGND VGND VPWR VPWR _5313_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6293_ _6704_/Q _5971_/A _5979_/X _6474_/Q VGND VGND VPWR VPWR _6293_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5244_ hold764/X _5538_/A1 _5246_/S VGND VGND VPWR VPWR _5244_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5175_ _5182_/S hold17/X VGND VGND VPWR VPWR _5181_/S sky130_fd_sc_hd__and2_2
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4126_ hold555/X _5513_/A1 _4126_/S VGND VGND VPWR VPWR _4126_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4057_ hold89/X _4056_/X _4067_/S VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__mux2_1
XFILLER_37_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4959_ _4959_/A _4959_/B VGND VGND VPWR VPWR _4959_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6629_ _6629_/CLK _6629_/D _6390_/A VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3975_/S hold33/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__nand2b_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6980_ _7065_/CLK _6980_/D fanout465/X VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5931_ _7118_/Q _6279_/S _5929_/X _5930_/X VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__o22a_1
X_5862_ _5862_/A _5862_/B _5862_/C _5862_/D VGND VGND VPWR VPWR _5862_/Y sky130_fd_sc_hd__nor4_2
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4813_ _4813_/A _4959_/B VGND VGND VPWR VPWR _4958_/B sky130_fd_sc_hd__and2_1
XFILLER_179_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5793_ _6872_/Q _5628_/X _5643_/X _7000_/Q VGND VGND VPWR VPWR _5793_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4744_ _4542_/B _4581_/B _4611_/Y _4619_/Y VGND VGND VPWR VPWR _4771_/A sky130_fd_sc_hd__o22a_1
XFILLER_159_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4675_ _4565_/X _4741_/A _4609_/Y _4663_/Y _5002_/A VGND VGND VPWR VPWR _4682_/B
+ sky130_fd_sc_hd__o221a_1
X_3626_ _6688_/Q _4292_/A _4032_/A _6473_/Q VGND VGND VPWR VPWR _3626_/X sky130_fd_sc_hd__a22o_1
X_6414_ _3568_/A1 _6414_/D _6370_/X VGND VGND VPWR VPWR _6414_/Q sky130_fd_sc_hd__dfrtp_1
X_3557_ _6694_/Q _4298_/A _4268_/A _6669_/Q _3556_/X VGND VGND VPWR VPWR _3565_/A
+ sky130_fd_sc_hd__a221o_1
X_6345_ _6642_/Q _6345_/A2 _6345_/B1 _6350_/A2 _6344_/X VGND VGND VPWR VPWR _6345_/X
+ sky130_fd_sc_hd__a221o_1
X_6276_ _6267_/X _6301_/C _6276_/C _6276_/D VGND VGND VPWR VPWR _6276_/X sky130_fd_sc_hd__and4b_2
X_3488_ _3487_/X _3488_/A1 _3829_/B VGND VGND VPWR VPWR _3488_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5227_ hold722/X _5521_/A1 _5227_/S VGND VGND VPWR VPWR _5227_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4335_/D sky130_fd_sc_hd__clkbuf_1
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5158_ hold754/X _6356_/A1 _5160_/S VGND VGND VPWR VPWR _5158_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4109_ _6396_/B hold37/X _5505_/B VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__and3b_4
X_5089_ _5089_/A _5089_/B _5089_/C _5089_/D VGND VGND VPWR VPWR _5122_/C sky130_fd_sc_hd__and4_1
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_70 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 _6619_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_92 _6558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4460_ _4460_/A _4993_/A VGND VGND VPWR VPWR _4782_/A sky130_fd_sc_hd__nor2_8
XFILLER_171_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold307 _6937_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold318 _4149_/X VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _7170_/Q _6487_/Q VGND VGND VPWR VPWR _3829_/B sky130_fd_sc_hd__nand2_4
Xhold329 _6897_/Q VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4391_ _4564_/A _4392_/C _4566_/A VGND VGND VPWR VPWR _4393_/A sky130_fd_sc_hd__a21oi_1
X_6130_ _6864_/Q _5943_/X _5981_/X _6920_/Q VGND VGND VPWR VPWR _6130_/X sky130_fd_sc_hd__a22o_1
X_3342_ hold27/X _3454_/B VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__nand2_8
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6941_/Q _5961_/X _6055_/X _6060_/X VGND VGND VPWR VPWR _6066_/A sky130_fd_sc_hd__a211o_1
XFILLER_97_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3273_ hold44/X _3251_/A _6488_/Q VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__mux2_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1007 _5164_/X VGND VGND VPWR VPWR _5165_/S sky130_fd_sc_hd__dlygate4sd3_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5012_ _4689_/B _4970_/Y _5010_/Y _4628_/Y _4796_/A VGND VGND VPWR VPWR _5134_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _4174_/X VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 _6466_/Q VGND VGND VPWR VPWR _4028_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6963_ _6963_/CLK hold14/X fanout458/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5914_ _6549_/Q _5655_/X _5912_/X _5913_/X VGND VGND VPWR VPWR _5914_/X sky130_fd_sc_hd__a211o_1
X_6894_ _7051_/CLK _6894_/D fanout476/X VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5845_ _6646_/Q _5621_/X _5628_/X _6615_/Q _5844_/X VGND VGND VPWR VPWR _5852_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5776_ _6791_/Q _5652_/Y _5769_/X _5775_/X _6303_/S VGND VGND VPWR VPWR _5776_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _4500_/A _4611_/Y _4964_/B _5039_/B VGND VGND VPWR VPWR _4727_/X sky130_fd_sc_hd__o211a_1
XFILLER_175_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4658_ _5088_/A _5099_/B _4658_/C VGND VGND VPWR VPWR _4658_/X sky130_fd_sc_hd__and3_1
XFILLER_174_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3609_ _6622_/Q _4220_/A _4151_/A _6563_/Q VGND VGND VPWR VPWR _3609_/X sky130_fd_sc_hd__a22o_1
Xhold830 _6664_/Q VGND VGND VPWR VPWR hold830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 _5492_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold852 _6749_/Q VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4589_ _4589_/A _4589_/B _4589_/C _4589_/D VGND VGND VPWR VPWR _4589_/Y sky130_fd_sc_hd__nand4_2
XFILLER_103_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold863 _5340_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 _6916_/Q VGND VGND VPWR VPWR hold874/X sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ _6327_/X _6328_/A1 _6346_/S VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__mux2_1
Xhold885 _5147_/X VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _6885_/Q VGND VGND VPWR VPWR hold896/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6259_ _6688_/Q _5961_/X _6257_/X _6258_/X VGND VGND VPWR VPWR _6264_/A sky130_fd_sc_hd__a211o_2
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1530 _7104_/Q VGND VGND VPWR VPWR _5607_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1541 _6723_/Q VGND VGND VPWR VPWR _5061_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 _7117_/Q VGND VGND VPWR VPWR _5909_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1563 _7091_/Q VGND VGND VPWR VPWR _3176_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1574 _7168_/Q VGND VGND VPWR VPWR _3249_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1585 _6527_/Q VGND VGND VPWR VPWR hold692/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1596 _6536_/Q VGND VGND VPWR VPWR hold158/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3960_ _6769_/Q _3960_/B VGND VGND VPWR VPWR _3960_/X sky130_fd_sc_hd__and2_4
XFILLER_73_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3891_ _5978_/A _5969_/A VGND VGND VPWR VPWR _5959_/A sky130_fd_sc_hd__and2_1
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5630_ _5664_/A _5658_/B _5666_/B VGND VGND VPWR VPWR _5630_/X sky130_fd_sc_hd__and3_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5561_ _5561_/A1 _5554_/Y _5604_/B _5560_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4512_ _4947_/B _4947_/C _4456_/Y VGND VGND VPWR VPWR _4514_/B sky130_fd_sc_hd__a21o_1
X_5492_ hold840/X _5492_/A1 _5495_/S VGND VGND VPWR VPWR _5492_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold104 _3372_/Y VGND VGND VPWR VPWR _3990_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 _5371_/X VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold126 _3326_/Y VGND VGND VPWR VPWR _5220_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4443_ _4607_/A _4753_/A VGND VGND VPWR VPWR _4611_/B sky130_fd_sc_hd__and2b_4
Xhold137 _6960_/Q VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _5432_/X VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold159 _4123_/X VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7162_ net399_2/A _7162_/D _6392_/X VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__dfrtp_1
X_4374_ _4374_/A _4374_/B VGND VGND VPWR VPWR _4471_/C sky130_fd_sc_hd__nor2_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6927_/Q _5938_/X _5952_/X _6959_/Q VGND VGND VPWR VPWR _6113_/X sky130_fd_sc_hd__a22o_1
X_3325_ _3379_/A _3543_/A VGND VGND VPWR VPWR _5418_/A sky130_fd_sc_hd__nor2_8
X_7093_ _7113_/CLK _7093_/D fanout462/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfstp_2
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _7049_/Q _5971_/A _5979_/X _6988_/Q VGND VGND VPWR VPWR _6044_/X sky130_fd_sc_hd__a22o_1
X_3256_ _3257_/A1 _3256_/A1 _3260_/S VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__mux2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3187_ _7074_/Q VGND VGND VPWR VPWR _3187_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6946_ _7049_/CLK _6946_/D fanout457/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6877_ _7076_/CLK _6877_/D fanout481/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfrtp_4
X_5828_ _6475_/Q _5630_/X _5824_/X _5825_/X _5827_/X VGND VGND VPWR VPWR _5828_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5759_ _7007_/Q _5625_/X _5661_/X _6879_/Q VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold660 _6793_/Q VGND VGND VPWR VPWR hold660/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold671 _6832_/Q VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold682 _5327_/X VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold693 _4113_/X VGND VGND VPWR VPWR _6527_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1360 hold1360/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
Xhold1371 _4188_/A1 VGND VGND VPWR VPWR hold1371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1382 _4112_/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1393 _7041_/Q VGND VGND VPWR VPWR _5499_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput209 _3217_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XFILLER_5_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4090_ _5205_/A0 _5484_/A1 _5202_/B VGND VGND VPWR VPWR _4090_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6800_ _6920_/CLK _6800_/D fanout474/X VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4992_ _4992_/A _4992_/B VGND VGND VPWR VPWR _4996_/D sky130_fd_sc_hd__nand2_1
X_6731_ _3945_/A1 _6731_/D _6383_/X VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfrtn_1
X_3943_ input84/X _3268_/C _6404_/Q VGND VGND VPWR VPWR _3943_/X sky130_fd_sc_hd__mux2_2
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6662_ _7058_/CLK _6662_/D _6396_/A VGND VGND VPWR VPWR _6662_/Q sky130_fd_sc_hd__dfrtp_1
X_3874_ _7104_/Q _6757_/Q _6762_/Q VGND VGND VPWR VPWR _5606_/A sky130_fd_sc_hd__mux2_4
XFILLER_177_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5613_ _7095_/Q _7094_/Q VGND VGND VPWR VPWR _5666_/B sky130_fd_sc_hd__and2_2
X_6593_ _7130_/CLK _6593_/D VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5544_ hold215/X _5544_/A1 _5549_/S VGND VGND VPWR VPWR _5544_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ hold872/X _5484_/A1 hold30/X VGND VGND VPWR VPWR _5475_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4426_ _4753_/A _4607_/A VGND VGND VPWR VPWR _4632_/B sky130_fd_sc_hd__nand2b_4
XFILLER_160_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout403 _5519_/A1 VGND VGND VPWR VPWR _5546_/A1 sky130_fd_sc_hd__buf_6
XFILLER_160_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout414 _5544_/A1 VGND VGND VPWR VPWR _5484_/A1 sky130_fd_sc_hd__buf_6
X_7145_ _3937_/A1 _7145_/D _6307_/B VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout425 hold666/X VGND VGND VPWR VPWR _5473_/A1 sky130_fd_sc_hd__buf_6
X_4357_ _4642_/A _4357_/B VGND VGND VPWR VPWR _4382_/B sky130_fd_sc_hd__xnor2_1
Xfanout436 _7096_/Q VGND VGND VPWR VPWR _5899_/B sky130_fd_sc_hd__buf_8
Xfanout447 fanout450/X VGND VGND VPWR VPWR fanout447/X sky130_fd_sc_hd__buf_6
Xfanout458 fanout466/X VGND VGND VPWR VPWR fanout458/X sky130_fd_sc_hd__buf_8
X_3308_ _3453_/A hold64/X VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__nor2_8
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout469 fanout486/X VGND VGND VPWR VPWR fanout469/X sky130_fd_sc_hd__buf_6
XFILLER_100_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4288_ hold269/X _5534_/A1 _4291_/S VGND VGND VPWR VPWR _4288_/X sky130_fd_sc_hd__mux2_1
X_7076_ _7076_/CLK _7076_/D fanout481/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_171_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6027_ _7119_/Q _6026_/X _6303_/S VGND VGND VPWR VPWR _6027_/X sky130_fd_sc_hd__mux2_1
X_3239_ _3837_/A _3239_/B VGND VGND VPWR VPWR _3875_/B sky130_fd_sc_hd__nor2_2
XFILLER_100_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _7054_/CLK _6929_/D fanout461/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7085_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_csclk _7001_/CLK VGND VGND VPWR VPWR _7065_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold490 _5363_/X VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_104_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1190 _6353_/X VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3590_ _6837_/Q _5265_/A _4172_/A _6581_/Q VGND VGND VPWR VPWR _3590_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5260_ hold652/X _5509_/A1 _5264_/S VGND VGND VPWR VPWR _5260_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4211_ _4211_/A0 _5493_/A1 _4213_/S VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
X_5191_ _5191_/A0 hold667/X _5192_/S VGND VGND VPWR VPWR _5191_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4142_ _4142_/A0 _5493_/A1 _4144_/S VGND VGND VPWR VPWR _4142_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4073_ hold401/X hold6/X _4083_/S VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4975_ _4975_/A _4975_/B VGND VGND VPWR VPWR _4975_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6714_ _6714_/CLK _6714_/D fanout470/X VGND VGND VPWR VPWR _6714_/Q sky130_fd_sc_hd__dfrtp_1
X_3926_ _6512_/Q _3251_/A _6406_/Q VGND VGND VPWR VPWR _3926_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6645_ _6671_/CLK _6645_/D fanout468/X VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfrtp_4
X_3857_ hold81/A _6488_/Q _3850_/Y _3856_/X _3866_/S VGND VGND VPWR VPWR _3857_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6576_ _7140_/CLK _6576_/D VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3788_ _3788_/A VGND VGND VPWR VPWR _3788_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5527_ _5527_/A0 _5545_/A1 _5531_/S VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5458_ _5458_/A0 _5494_/A1 _5462_/S VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4409_ _4551_/A _4570_/A _4459_/B VGND VGND VPWR VPWR _4584_/A sky130_fd_sc_hd__and3_1
X_5389_ hold149/X hold99/X _5390_/S VGND VGND VPWR VPWR _5389_/X sky130_fd_sc_hd__mux2_1
X_7128_ _7130_/CLK _7128_/D fanout486/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7059_ _7083_/CLK _7059_/D _6396_/A VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 hold666/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_171 _5291_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _7066_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_193 _5465_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4948_/A _4672_/B _4626_/Y _4653_/Y VGND VGND VPWR VPWR _5003_/A sky130_fd_sc_hd__o22a_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3711_ _6435_/Q _3372_/Y _5319_/A _6883_/Q _3710_/X VGND VGND VPWR VPWR _3720_/A
+ sky130_fd_sc_hd__a221o_1
X_4691_ _4691_/A _4902_/B VGND VGND VPWR VPWR _4975_/B sky130_fd_sc_hd__nand2_2
X_6430_ _6749_/CLK _6430_/D fanout449/X VGND VGND VPWR VPWR _6430_/Q sky130_fd_sc_hd__dfrtp_2
X_3642_ _3641_/X _3642_/A1 _3829_/B VGND VGND VPWR VPWR _3642_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6361_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6361_/X sky130_fd_sc_hd__and2_1
XFILLER_127_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3573_ _3573_/A _3573_/B VGND VGND VPWR VPWR _4304_/A sky130_fd_sc_hd__nor2_4
XFILLER_114_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5312_ hold541/X _5543_/A1 _5318_/S VGND VGND VPWR VPWR _5312_/X sky130_fd_sc_hd__mux2_1
X_6292_ _6564_/Q _5953_/X _5960_/X _6674_/Q _6291_/X VGND VGND VPWR VPWR _6292_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5243_ hold196/X _5519_/A1 _5246_/S VGND VGND VPWR VPWR _5243_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ hold48/X _3717_/B hold667/X _5173_/X hold16/X VGND VGND VPWR VPWR _5174_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4125_ _4125_/A0 hold99/X _4126_/S VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4056_ _4112_/A0 hold6/X _4058_/S VGND VGND VPWR VPWR _4056_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4958_ _5042_/B _4958_/B VGND VGND VPWR VPWR _5046_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3909_ _3909_/A _3909_/B VGND VGND VPWR VPWR _3910_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4889_ _4689_/A _4645_/Y _4892_/B _4491_/Y _4523_/Y VGND VGND VPWR VPWR _5084_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6628_ _6683_/CLK _6628_/D _6390_/A VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6559_ _6629_/CLK _6559_/D _6390_/A VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5930_ _5552_/B _7117_/Q _6103_/B1 VGND VGND VPWR VPWR _5930_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5861_ _6471_/Q _5627_/X _5655_/X _6546_/Q _5860_/X VGND VGND VPWR VPWR _5862_/D
+ sky130_fd_sc_hd__a221o_1
X_4812_ _4562_/Y _4810_/B _4948_/D VGND VGND VPWR VPWR _4812_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5792_ _6984_/Q _5624_/X _5818_/A2 _6824_/Q _5791_/X VGND VGND VPWR VPWR _5797_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4743_ _4810_/A _4581_/B _4611_/Y _4613_/Y VGND VGND VPWR VPWR _4772_/A sky130_fd_sc_hd__o22a_1
XFILLER_187_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4674_ _4608_/X _4644_/B _4984_/B _4673_/Y _4472_/A VGND VGND VPWR VPWR _4674_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_6413_ _3568_/A1 _6413_/D _6369_/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfrtp_2
X_3625_ _6437_/Q _3372_/Y _3964_/A _6421_/Q _3624_/X VGND VGND VPWR VPWR _3628_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6344_ _6644_/Q _6344_/A2 _6344_/B1 _6643_/Q VGND VGND VPWR VPWR _6344_/X sky130_fd_sc_hd__a22o_1
X_3556_ _7022_/Q hold29/A _4238_/A _6634_/Q VGND VGND VPWR VPWR _3556_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6275_ _6275_/A _6275_/B _6275_/C _6275_/D VGND VGND VPWR VPWR _6276_/D sky130_fd_sc_hd__nor4_1
XFILLER_163_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3487_ _3486_/Y _6731_/Q _3829_/A VGND VGND VPWR VPWR _3487_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5226_ _5226_/A0 _5538_/A1 _5227_/S VGND VGND VPWR VPWR _5226_/X sky130_fd_sc_hd__mux2_1
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4335_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_69_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5157_ hold950/X _6355_/A1 _5160_/S VGND VGND VPWR VPWR _5157_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4108_ hold383/X _5538_/A1 _4108_/S VGND VGND VPWR VPWR _4108_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5088_ _5088_/A _5088_/B _5088_/C _5088_/D VGND VGND VPWR VPWR _5089_/D sky130_fd_sc_hd__and4_1
XFILLER_56_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4039_ _4039_/A0 _5491_/A1 _4043_/S VGND VGND VPWR VPWR _4039_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_60 _6025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _6898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_93 _6568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold308 _5381_/X VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold319 _7061_/Q VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_3410_ _3410_/A _3410_/B VGND VGND VPWR VPWR _3410_/Y sky130_fd_sc_hd__nand2_4
XFILLER_144_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4390_ _4631_/D _4633_/B _4661_/A _4441_/B VGND VGND VPWR VPWR _4392_/C sky130_fd_sc_hd__and4_1
XFILLER_125_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3341_ hold36/X hold85/X VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__nor2_8
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _7013_/Q _5940_/X _5967_/X _6853_/Q _6054_/X VGND VGND VPWR VPWR _6060_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ hold25/X _4885_/B2 _3975_/S VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__mux2_2
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1008 _5165_/X VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5011_ _4689_/A _4644_/Y _5010_/Y _4639_/Y VGND VGND VPWR VPWR _5011_/X sky130_fd_sc_hd__o22a_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1019 _6546_/Q VGND VGND VPWR VPWR _4135_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6962_ _7006_/CLK _6962_/D fanout457/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5913_ _6603_/Q _5616_/X _5913_/B1 _6554_/Q VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__a22o_1
X_6893_ _7076_/CLK _6893_/D fanout481/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5844_ _6456_/Q _5645_/X _5910_/B1 _6626_/Q VGND VGND VPWR VPWR _5844_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5775_ _6935_/Q _5654_/X _5770_/X _5772_/X _5774_/X VGND VGND VPWR VPWR _5775_/X
+ sky130_fd_sc_hd__a2111o_2
X_4726_ _4984_/A _4965_/B _4975_/A VGND VGND VPWR VPWR _5039_/B sky130_fd_sc_hd__nand3_1
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4657_ _4611_/Y _4639_/Y _4652_/Y _4620_/Y VGND VGND VPWR VPWR _4657_/X sky130_fd_sc_hd__o22a_1
XFILLER_175_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3608_ input55/X _5193_/A _4256_/A _6658_/Q _3589_/X VGND VGND VPWR VPWR _3611_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold820 _6623_/Q VGND VGND VPWR VPWR hold820/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_2
X_4588_ _4948_/B _4672_/B VGND VGND VPWR VPWR _4588_/Y sky130_fd_sc_hd__nor2_1
Xhold831 _4267_/X VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 _6629_/Q VGND VGND VPWR VPWR hold842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 _5163_/X VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold864 _6932_/Q VGND VGND VPWR VPWR hold864/X sky130_fd_sc_hd__dlygate4sd3_1
X_6327_ _6644_/Q _6327_/A2 _6327_/B1 _6350_/A2 _6326_/X VGND VGND VPWR VPWR _6327_/X
+ sky130_fd_sc_hd__a221o_1
X_3539_ hold74/X _3571_/B VGND VGND VPWR VPWR _6352_/A sky130_fd_sc_hd__nor2_4
Xmgmt_gpio_15_buff_inst _3936_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_8
Xhold875 _5358_/X VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold886 _6444_/Q VGND VGND VPWR VPWR hold886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 _5323_/X VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6258_ _6478_/Q _5940_/X _5967_/X _6607_/Q _6256_/X VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5209_ hold291/X _5521_/A1 _5210_/S VGND VGND VPWR VPWR _5209_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6189_ _6189_/A _6189_/B _6189_/C VGND VGND VPWR VPWR _6189_/Y sky130_fd_sc_hd__nor3_1
Xhold1520 _7110_/Q VGND VGND VPWR VPWR _5757_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 hold52/A VGND VGND VPWR VPWR _6340_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 _6640_/Q VGND VGND VPWR VPWR _3954_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1553 _7114_/Q VGND VGND VPWR VPWR _5843_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1564 _7126_/Q VGND VGND VPWR VPWR _6179_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1575 _7087_/Q VGND VGND VPWR VPWR _5551_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1586 _7098_/Q VGND VGND VPWR VPWR _5590_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1597 _6784_/Q VGND VGND VPWR VPWR hold291/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3890_ _7100_/Q _7099_/Q VGND VGND VPWR VPWR _5969_/A sky130_fd_sc_hd__and2b_4
XFILLER_149_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5560_ _7088_/Q _7089_/Q _6509_/Q _5552_/B _3885_/Y VGND VGND VPWR VPWR _5560_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_129_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4511_ _4453_/B _4948_/C _4508_/X _4510_/X VGND VGND VPWR VPWR _4514_/A sky130_fd_sc_hd__o211a_1
XFILLER_157_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5491_ _5491_/A0 _5491_/A1 _5495_/S VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__mux2_1
Xhold105 _3997_/X VGND VGND VPWR VPWR _6440_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold116 _6942_/Q VGND VGND VPWR VPWR hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4442_ _4465_/B _4900_/A _4896_/B _4724_/A VGND VGND VPWR VPWR _4442_/Y sky130_fd_sc_hd__nand4_1
Xhold127 _5227_/S VGND VGND VPWR VPWR _5228_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _5407_/X VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _6944_/Q VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7161_ net399_2/A _7161_/D _6391_/X VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4373_ _4702_/B _4434_/B VGND VGND VPWR VPWR _4627_/A sky130_fd_sc_hd__nand2_4
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6975_/Q _5947_/X _5965_/X _6799_/Q _6111_/X VGND VGND VPWR VPWR _6115_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3356_/A hold73/X VGND VGND VPWR VPWR _3543_/A sky130_fd_sc_hd__nand2_8
X_7092_ _7113_/CLK _7092_/D fanout462/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6820_/Q _5953_/X _5960_/X _7073_/Q _6042_/X VGND VGND VPWR VPWR _6043_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3256_/A1 _3255_/A1 _3260_/S VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__mux2_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3186_ _7082_/Q VGND VGND VPWR VPWR _3186_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _7054_/CLK _6945_/D fanout461/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6876_ _7067_/CLK _6876_/D fanout476/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5827_ _6578_/Q _5928_/A2 _5913_/B1 _6550_/Q _5826_/X VGND VGND VPWR VPWR _5827_/X
+ sky130_fd_sc_hd__a221o_1
X_5758_ _3226_/Y _5899_/B _5651_/B VGND VGND VPWR VPWR _5758_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_148_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4709_ _4691_/A _4902_/B _4619_/Y VGND VGND VPWR VPWR _5084_/C sky130_fd_sc_hd__a21o_1
XFILLER_135_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5689_ _6939_/Q _5632_/X _5663_/X _6859_/Q _5688_/X VGND VGND VPWR VPWR _5690_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold650 _7054_/Q VGND VGND VPWR VPWR hold650/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold661 _5219_/X VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold672 _5263_/X VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold683 _6791_/Q VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap391 _4230_/B VGND VGND VPWR VPWR _6350_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold694 _6935_/Q VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1350 hold1350/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1361 _6313_/A1 VGND VGND VPWR VPWR hold1361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1372 hold1372/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_85_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 hold1578/X VGND VGND VPWR VPWR _4125_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _5499_/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4991_ _4626_/Y _4644_/Y _4646_/Y VGND VGND VPWR VPWR _4991_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6730_ _3945_/A1 _6730_/D _6382_/X VGND VGND VPWR VPWR _6730_/Q sky130_fd_sc_hd__dfrtn_1
X_3942_ _3975_/S _3942_/A2 _6396_/B _3941_/Y VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__a22o_2
XFILLER_189_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ _6712_/CLK _6661_/D _6396_/A VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfrtp_4
X_3873_ _3264_/B _3838_/A _3872_/X _3832_/B _6402_/Q VGND VGND VPWR VPWR _6402_/D
+ sky130_fd_sc_hd__a32o_1
X_5612_ _5552_/B _5606_/A _5610_/Y VGND VGND VPWR VPWR _6304_/S sky130_fd_sc_hd__a21o_2
XFILLER_149_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6592_ _7130_/CLK _6592_/D VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfxtp_1
X_5543_ hold644/X _5543_/A1 _5549_/S VGND VGND VPWR VPWR _5543_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5474_ hold594/X _5543_/A1 hold30/X VGND VGND VPWR VPWR _5474_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4425_ _4685_/A _4921_/A VGND VGND VPWR VPWR _5023_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout404 _5519_/A1 VGND VGND VPWR VPWR _5528_/A1 sky130_fd_sc_hd__buf_6
X_7144_ _3937_/A1 _7144_/D fanout487/X VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfrtp_1
X_4356_ _4356_/A _4356_/B VGND VGND VPWR VPWR _4492_/D sky130_fd_sc_hd__nor2_2
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout415 hold6/X VGND VGND VPWR VPWR _5544_/A1 sky130_fd_sc_hd__buf_8
Xfanout426 hold665/X VGND VGND VPWR VPWR hold666/A sky130_fd_sc_hd__buf_8
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout437 _3963_/S VGND VGND VPWR VPWR _3975_/S sky130_fd_sc_hd__clkbuf_16
Xfanout448 fanout450/X VGND VGND VPWR VPWR fanout448/X sky130_fd_sc_hd__buf_4
XFILLER_100_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3307_ _3586_/A _3374_/A VGND VGND VPWR VPWR _5355_/A sky130_fd_sc_hd__nor2_8
Xfanout459 fanout462/X VGND VGND VPWR VPWR fanout459/X sky130_fd_sc_hd__buf_8
XFILLER_113_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7075_ _7083_/CLK _7075_/D _6396_/A VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4287_ _4287_/A0 hold667/X _4291_/S VGND VGND VPWR VPWR _4287_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6026_ _6014_/Y _6025_/X _6787_/Q _6226_/B VGND VGND VPWR VPWR _6026_/X sky130_fd_sc_hd__o2bb2a_1
X_3238_ _6416_/Q _3837_/A _6485_/Q _3829_/A _3239_/B VGND VGND VPWR VPWR _3249_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _6642_/Q VGND VGND VPWR VPWR _3962_/A sky130_fd_sc_hd__inv_2
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ _7017_/CLK _6928_/D fanout461/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6859_ _7011_/CLK _6859_/D fanout456/X VGND VGND VPWR VPWR _6859_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold480 _5333_/X VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _6648_/Q VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1180 _5293_/X VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 _6922_/Q VGND VGND VPWR VPWR _5365_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4210_ _4210_/A0 _5492_/A1 _4213_/S VGND VGND VPWR VPWR _4210_/X sky130_fd_sc_hd__mux2_1
X_5190_ _5190_/A _5190_/B hold16/X VGND VGND VPWR VPWR _5192_/S sky130_fd_sc_hd__and3_1
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4141_ _4141_/A0 _5492_/A1 _4144_/S VGND VGND VPWR VPWR _4141_/X sky130_fd_sc_hd__mux2_1
X_4072_ _4072_/A0 _4071_/X _4084_/S VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4974_ _5021_/B _4974_/B _5008_/C _4974_/D VGND VGND VPWR VPWR _4983_/B sky130_fd_sc_hd__and4_1
X_3925_ _6521_/Q input81/X _3957_/B VGND VGND VPWR VPWR _3925_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6713_ _7083_/CLK _6713_/D _6396_/A VGND VGND VPWR VPWR _6713_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6644_ _3937_/A1 _6644_/D fanout487/X VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfrtp_4
X_3856_ hold81/A hold24/A hold44/A hold62/A VGND VGND VPWR VPWR _3856_/X sky130_fd_sc_hd__a31o_1
XFILLER_177_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6575_ _7140_/CLK _6575_/D VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfxtp_1
X_3787_ _7159_/Q _6404_/Q _6755_/Q VGND VGND VPWR VPWR _3788_/A sky130_fd_sc_hd__nor3_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5526_ hold371/X _5526_/A1 _5531_/S VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5457_ hold343/X _5526_/A1 _5462_/S VGND VGND VPWR VPWR _5457_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4408_ _4633_/B _4408_/B VGND VGND VPWR VPWR _4459_/B sky130_fd_sc_hd__and2b_4
XFILLER_132_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5388_ hold712/X _5469_/A1 _5390_/S VGND VGND VPWR VPWR _5388_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7127_ _7130_/CLK _7127_/D fanout486/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_1
X_4339_ _4739_/A _4642_/A VGND VGND VPWR VPWR _4661_/A sky130_fd_sc_hd__and2_4
XFILLER_115_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7058_ _7058_/CLK _7058_/D _6396_/A VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6009_ _6939_/Q _5961_/X _6006_/X _6008_/X VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__a211o_1
XFILLER_74_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_161 hold666/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _5948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _6558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 _5473_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _6923_/Q _5364_/A _4044_/A _6481_/Q VGND VGND VPWR VPWR _3710_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4690_ _4690_/A _4690_/B VGND VGND VPWR VPWR _4690_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3641_ _3640_/Y _6729_/Q _3829_/A VGND VGND VPWR VPWR _3641_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6360_ _6360_/A _6400_/B VGND VGND VPWR VPWR _6360_/X sky130_fd_sc_hd__and2_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3572_ _6950_/Q _3781_/A2 _4145_/A _6559_/Q _3570_/X VGND VGND VPWR VPWR _3580_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5311_ _5311_/A0 _5473_/A1 _5318_/S VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__mux2_1
X_6291_ _6654_/Q _5973_/A _5948_/X _6699_/Q _6290_/X VGND VGND VPWR VPWR _6291_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5242_ _5242_/A0 _5545_/A1 _5246_/S VGND VGND VPWR VPWR _5242_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7082_/CLK sky130_fd_sc_hd__clkbuf_16
X_5173_ _3320_/X _3355_/X _5173_/B1 VGND VGND VPWR VPWR _5173_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4124_ hold742/X _5469_/A1 _4126_/S VGND VGND VPWR VPWR _4124_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_2
X_4055_ hold339/X _4054_/X _4067_/S VGND VGND VPWR VPWR _4055_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_csclk clkbuf_opt_4_0_csclk/X VGND VGND VPWR VPWR _6908_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4957_ _4574_/Y _4956_/Y _4575_/Y VGND VGND VPWR VPWR _4957_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3908_ _3909_/B VGND VGND VPWR VPWR _3908_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4888_ _4469_/A _4947_/C _4887_/A _4633_/B _4379_/B VGND VGND VPWR VPWR _4892_/B
+ sky130_fd_sc_hd__a2111o_2
X_3839_ _6488_/Q _3867_/A VGND VGND VPWR VPWR _3860_/B sky130_fd_sc_hd__nand2_2
X_6627_ _6629_/CLK _6627_/D _6390_/A VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_192_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6558_ _6712_/CLK _6558_/D _6390_/A VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5509_ hold598/X _5509_/A1 _5513_/S VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__mux2_1
X_6489_ _3927_/A1 _6489_/D _6378_/X VGND VGND VPWR VPWR _6489_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire443 _3268_/Y VGND VGND VPWR VPWR _6367_/B sky130_fd_sc_hd__buf_4
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5860_ _6461_/Q _5624_/X _5664_/X _6666_/Q VGND VGND VPWR VPWR _5860_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4811_ _4581_/B _4947_/C _4500_/A VGND VGND VPWR VPWR _5039_/C sky130_fd_sc_hd__a21o_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5791_ _6976_/Q _5634_/X _5652_/B _5790_/Y VGND VGND VPWR VPWR _5791_/X sky130_fd_sc_hd__a22o_1
X_4742_ _4472_/A _4574_/B _4737_/A VGND VGND VPWR VPWR _4996_/B sky130_fd_sc_hd__o21ai_1
XFILLER_193_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4673_ _4673_/A _4673_/B VGND VGND VPWR VPWR _4673_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6412_ _3568_/A1 _6412_/D _6368_/X VGND VGND VPWR VPWR _6412_/Q sky130_fd_sc_hd__dfrtp_1
X_3624_ _6933_/Q _5373_/A _4316_/A _6708_/Q VGND VGND VPWR VPWR _3624_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6343_ _6342_/X _6343_/A1 _6346_/S VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__mux2_1
X_3555_ _3555_/A hold66/X VGND VGND VPWR VPWR _4238_/A sky130_fd_sc_hd__nor2_4
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6274_ _6693_/Q _5954_/X _5976_/D _6622_/Q _6255_/X VGND VGND VPWR VPWR _6275_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3486_ _3486_/A _3486_/B VGND VGND VPWR VPWR _3486_/Y sky130_fd_sc_hd__nand2_4
XFILLER_88_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5225_ _5225_/A0 hold60/X _5228_/S VGND VGND VPWR VPWR _5225_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5156_ hold832/X _6354_/A1 _5160_/S VGND VGND VPWR VPWR _5156_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4107_ hold433/X _5528_/A1 _4108_/S VGND VGND VPWR VPWR _4107_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5087_ _5087_/A _5087_/B _5115_/C _5087_/D VGND VGND VPWR VPWR _5087_/Y sky130_fd_sc_hd__nand4_1
XFILLER_84_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4038_ _4038_/A _6352_/B VGND VGND VPWR VPWR _4043_/S sky130_fd_sc_hd__and2_2
XFILLER_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5989_ _5989_/A _5989_/B _5989_/C VGND VGND VPWR VPWR _6001_/C sky130_fd_sc_hd__nor3_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 _5654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _6025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_83 _6949_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 _6837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput190 _3200_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_121_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold309 _6622_/Q VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7137_/CLK sky130_fd_sc_hd__clkbuf_8
X_3340_ _3370_/A _3455_/A VGND VGND VPWR VPWR _5523_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ hold24/X hold44/A _6488_/Q VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__mux2_1
XFILLER_98_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/A _5010_/B VGND VGND VPWR VPWR _5010_/Y sky130_fd_sc_hd__nor2_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1009 _6651_/Q VGND VGND VPWR VPWR _4252_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7103__490 VGND VGND VPWR VPWR _7103_/D _7103__490/LO sky130_fd_sc_hd__conb_1
XFILLER_93_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6961_ _7017_/CLK _6961_/D fanout461/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5912_ _6474_/Q _5627_/X _5635_/X _6569_/Q VGND VGND VPWR VPWR _5912_/X sky130_fd_sc_hd__a22o_1
X_6892_ _7067_/CLK _6892_/D fanout477/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_2
X_5843_ _5843_/A1 _6279_/S _5842_/X VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__o21a_1
XFILLER_179_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5774_ _6839_/Q _5657_/X _5660_/X _6807_/Q _5773_/X VGND VGND VPWR VPWR _5774_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4725_ _5114_/A _4725_/B VGND VGND VPWR VPWR _4725_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4656_ _4632_/Y _4645_/Y _4654_/X _4655_/X VGND VGND VPWR VPWR _4660_/C sky130_fd_sc_hd__o211a_1
XFILLER_174_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _3959_/B sky130_fd_sc_hd__clkbuf_4
X_3607_ _6853_/Q _5283_/A _5256_/A _6829_/Q _3590_/X VGND VGND VPWR VPWR _3611_/B
+ sky130_fd_sc_hd__a221o_1
Xhold810 _6566_/Q VGND VGND VPWR VPWR hold810/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4587_ _4690_/A _4495_/A _4570_/Y _4580_/X _4586_/X VGND VGND VPWR VPWR _4589_/D
+ sky130_fd_sc_hd__o311a_1
Xhold821 _4225_/X VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 _6743_/Q VGND VGND VPWR VPWR hold832/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_2
Xhold843 _4237_/X VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3538_ _3538_/A _3538_/B _3538_/C _3538_/D VGND VGND VPWR VPWR _3538_/Y sky130_fd_sc_hd__nor4_1
Xhold854 _6812_/Q VGND VGND VPWR VPWR hold854/X sky130_fd_sc_hd__dlygate4sd3_1
X_6326_ _6642_/Q _6326_/A2 _6326_/B1 _6643_/Q VGND VGND VPWR VPWR _6326_/X sky130_fd_sc_hd__a22o_1
Xhold865 _5376_/X VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold876 _6471_/Q VGND VGND VPWR VPWR hold876/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold887 _4002_/X VGND VGND VPWR VPWR _6444_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold898 _7077_/Q VGND VGND VPWR VPWR hold898/X sky130_fd_sc_hd__dlygate4sd3_1
X_6257_ _7154_/Q _5958_/X _5978_/X _6483_/Q VGND VGND VPWR VPWR _6257_/X sky130_fd_sc_hd__a22o_1
X_3469_ _3956_/A _4083_/S _5337_/A _6903_/Q _3468_/X VGND VGND VPWR VPWR _3472_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5208_ hold168/X hold42/X _5210_/S VGND VGND VPWR VPWR _5208_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6188_ _6665_/Q _5938_/X _5952_/X _6705_/Q _6187_/X VGND VGND VPWR VPWR _6189_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1510 hold20/A VGND VGND VPWR VPWR _3254_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 _5757_/X VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5139_ _5001_/B _5077_/C _5138_/X _5103_/Y VGND VGND VPWR VPWR _5143_/B sky130_fd_sc_hd__a31o_1
Xhold1532 _7160_/Q VGND VGND VPWR VPWR _3260_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 _7169_/Q VGND VGND VPWR VPWR _3248_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1554 _6720_/Q VGND VGND VPWR VPWR _4731_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 hold44/A VGND VGND VPWR VPWR _3866_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1576 _6524_/Q VGND VGND VPWR VPWR hold1576/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1587 _6525_/Q VGND VGND VPWR VPWR hold622/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 _7185_/A VGND VGND VPWR VPWR hold1598/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ _4902_/A _4456_/Y _4509_/X VGND VGND VPWR VPWR _4510_/X sky130_fd_sc_hd__o21a_1
XFILLER_157_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5490_ _5490_/A _5490_/B VGND VGND VPWR VPWR _5495_/S sky130_fd_sc_hd__and2_2
XFILLER_171_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4441_ _4441_/A _4441_/B VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__nand2_8
Xhold106 _7147_/Q VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _5387_/X VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _5225_/X VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _6792_/Q VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7160_ net399_2/A _7160_/D _6390_/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4372_ _4702_/B _4591_/A VGND VGND VPWR VPWR _4372_/X sky130_fd_sc_hd__and2_1
XFILLER_171_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6895_/Q _5946_/X _5955_/X _6807_/Q VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3323_ hold34/X _3323_/B hold72/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__and3_4
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7113_/CLK _7091_/D fanout460/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6908_/Q _5973_/A _5948_/X _6948_/Q _6041_/X VGND VGND VPWR VPWR _6042_/X
+ sky130_fd_sc_hd__a221o_1
X_3254_ hold97/A _3254_/A1 _3260_/S VGND VGND VPWR VPWR _3254_/X sky130_fd_sc_hd__mux2_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _6657_/Q VGND VGND VPWR VPWR _3185_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6944_ _6981_/CLK _6944_/D fanout463/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtp_1
X_6875_ _7067_/CLK _6875_/D fanout477/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_179_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5826_ _6465_/Q _5619_/X _5663_/X _6609_/Q VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5757_ _5757_/A0 _5756_/X _6279_/S VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4708_ _4469_/A _4689_/B _4639_/Y _4690_/Y VGND VGND VPWR VPWR _5062_/B sky130_fd_sc_hd__o22a_1
XFILLER_175_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5688_ _6987_/Q _5627_/X _5661_/X _6875_/Q VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__a22o_1
X_4639_ _4716_/A _4707_/C VGND VGND VPWR VPWR _4639_/Y sky130_fd_sc_hd__nand2_8
Xhold640 _6422_/Q VGND VGND VPWR VPWR hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold651 _5513_/X VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold662 _6616_/Q VGND VGND VPWR VPWR hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap370 hold36/X VGND VGND VPWR VPWR _3814_/A sky130_fd_sc_hd__buf_12
Xhold673 _6912_/Q VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _5217_/X VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6309_ _3762_/Y _6309_/A1 _6315_/S VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold695 _5379_/X VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1340 hold1340/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1351 _4164_/A1 VGND VGND VPWR VPWR hold1351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 hold1362/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
Xhold1373 _6308_/A1 VGND VGND VPWR VPWR hold1373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 _7175_/A VGND VGND VPWR VPWR _4076_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1395 _7025_/Q VGND VGND VPWR VPWR _5480_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4990_ _4948_/A _4428_/Y _4846_/B _4645_/Y VGND VGND VPWR VPWR _5003_/C sky130_fd_sc_hd__o22a_1
XFILLER_63_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3941_ _3975_/S _3941_/B VGND VGND VPWR VPWR _3941_/Y sky130_fd_sc_hd__nor2_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3872_ _7170_/Q _6402_/Q _3867_/A VGND VGND VPWR VPWR _3872_/X sky130_fd_sc_hd__o21a_1
X_6660_ _7058_/CLK _6660_/D _6396_/A VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5611_ _5552_/B _5606_/A _5610_/Y VGND VGND VPWR VPWR _5611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6591_ _7130_/CLK _6591_/D VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfxtp_1
X_5542_ _5542_/A0 hold667/X _5549_/S VGND VGND VPWR VPWR _5542_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5473_ _5473_/A0 _5473_/A1 hold30/X VGND VGND VPWR VPWR _5473_/X sky130_fd_sc_hd__mux2_1
X_4424_ _4500_/A _4581_/B VGND VGND VPWR VPWR _4424_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4355_ _4556_/A _4563_/A _4753_/A _4607_/A _4642_/A VGND VGND VPWR VPWR _4356_/B
+ sky130_fd_sc_hd__o2111a_1
X_7143_ _7150_/CLK _7143_/D fanout487/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfrtp_1
XFILLER_113_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout405 hold59/X VGND VGND VPWR VPWR _5519_/A1 sky130_fd_sc_hd__buf_6
Xfanout416 _5465_/A1 VGND VGND VPWR VPWR _6354_/A1 sky130_fd_sc_hd__buf_6
Xfanout427 _5490_/B VGND VGND VPWR VPWR _6352_/B sky130_fd_sc_hd__buf_6
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3306_ _3554_/A _3379_/A VGND VGND VPWR VPWR _5346_/A sky130_fd_sc_hd__nor2_8
Xfanout438 _6507_/Q VGND VGND VPWR VPWR _5552_/B sky130_fd_sc_hd__buf_6
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7074_ _7085_/CLK _7074_/D fanout479/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout449 fanout450/X VGND VGND VPWR VPWR fanout449/X sky130_fd_sc_hd__buf_6
XFILLER_59_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4286_ _4286_/A _4322_/B VGND VGND VPWR VPWR _4291_/S sky130_fd_sc_hd__and2_2
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3237_ _6417_/Q _6416_/Q VGND VGND VPWR VPWR _3239_/B sky130_fd_sc_hd__nand2_1
X_6025_ _6017_/X _6025_/B _6226_/B VGND VGND VPWR VPWR _6025_/X sky130_fd_sc_hd__and3b_2
XFILLER_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3168_ _3168_/A VGND VGND VPWR VPWR _3910_/A sky130_fd_sc_hd__inv_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _7054_/CLK _6927_/D fanout460/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6858_ _6926_/CLK _6858_/D fanout457/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5809_ _6985_/Q _5624_/X _5634_/X _6977_/Q _5802_/Y VGND VGND VPWR VPWR _5809_/X
+ sky130_fd_sc_hd__a221o_1
X_6789_ _6963_/CLK _6789_/D fanout456/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold470 _5415_/X VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold481 _6673_/Q VGND VGND VPWR VPWR hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _4248_/X VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1170 _4070_/X VGND VGND VPWR VPWR _6498_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1181 _6764_/Q VGND VGND VPWR VPWR _5185_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1192 _5365_/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4140_ _4140_/A0 _6353_/A1 _4144_/S VGND VGND VPWR VPWR _4140_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4071_ hold824/X _6354_/A1 _4118_/B VGND VGND VPWR VPWR _4071_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4973_ _4616_/Y _4628_/Y _4970_/Y VGND VGND VPWR VPWR _4974_/D sky130_fd_sc_hd__a21o_1
X_6712_ _6712_/CLK _6712_/D fanout470/X VGND VGND VPWR VPWR _6712_/Q sky130_fd_sc_hd__dfstp_2
X_3924_ _6519_/Q input78/X _3957_/B VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6643_ _7150_/CLK _6643_/D fanout487/X VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfrtp_4
X_3855_ _3854_/X _3855_/A1 _3866_/S VGND VGND VPWR VPWR _6411_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3786_ _6866_/Q _5301_/A _4038_/A _6475_/Q _3785_/X VGND VGND VPWR VPWR _3793_/B
+ sky130_fd_sc_hd__a221o_1
X_6574_ _7137_/CLK _6574_/D VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5525_ hold543/X _5543_/A1 _5531_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5456_ hold253/X _5465_/A1 _5462_/S VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4407_ _4551_/A _4570_/A VGND VGND VPWR VPWR _4498_/A sky130_fd_sc_hd__and2_2
X_5387_ hold116/X hold60/X _5390_/S VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7126_ _7126_/CLK _7126_/D fanout459/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4338_ _4338_/A _4338_/B _4338_/C VGND VGND VPWR VPWR _4564_/A sky130_fd_sc_hd__and3_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4269_ _4269_/A0 _6353_/A1 _4273_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
X_7057_ _7079_/CLK _7057_/D fanout478/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6008_ _7011_/Q _5940_/X _5967_/X _6851_/Q _6005_/X VGND VGND VPWR VPWR _6008_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_101_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _6226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_151 _5473_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _5193_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _5953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _6853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _5490_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _3597_/X _3640_/B _3640_/C _3640_/D VGND VGND VPWR VPWR _3640_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3571_ _3571_/A _3571_/B VGND VGND VPWR VPWR _4145_/A sky130_fd_sc_hd__nor2_2
XFILLER_155_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5310_ _5310_/A _5541_/B VGND VGND VPWR VPWR _5318_/S sky130_fd_sc_hd__and2_4
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6290_ _6649_/Q _5976_/C _5971_/D _6569_/Q VGND VGND VPWR VPWR _6290_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5241_ hold854/X _5484_/A1 _5246_/S VGND VGND VPWR VPWR _5241_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5172_ _5172_/A0 _5491_/A1 _5172_/S VGND VGND VPWR VPWR _5172_/X sky130_fd_sc_hd__mux2_1
X_4123_ hold158/X hold60/X _4126_/S VGND VGND VPWR VPWR _4123_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
X_4054_ hold622/X _5534_/A1 _4058_/S VGND VGND VPWR VPWR _4054_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_opt_1_0_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR clkbuf_leaf_4_csclk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4956_ _4965_/B _5051_/A _4554_/B VGND VGND VPWR VPWR _4956_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3907_ _3907_/A _3907_/B _3907_/C _3907_/D VGND VGND VPWR VPWR _3909_/B sky130_fd_sc_hd__nand4_2
X_4887_ _4887_/A _4887_/B VGND VGND VPWR VPWR _4900_/B sky130_fd_sc_hd__nor2_1
X_6626_ _6769_/CLK _6626_/D fanout469/X VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfrtp_4
X_3838_ _3838_/A _3838_/B VGND VGND VPWR VPWR _6415_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6557_ _6629_/CLK _6557_/D _6390_/A VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfrtp_4
X_3769_ _6786_/Q _5211_/A _4280_/A _6675_/Q VGND VGND VPWR VPWR _3769_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5508_ hold335/X _5526_/A1 _5513_/S VGND VGND VPWR VPWR _5508_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6488_ _3927_/A1 _6488_/D _6377_/X VGND VGND VPWR VPWR _6488_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5439_ hold337/X _5526_/A1 _5444_/S VGND VGND VPWR VPWR _5439_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _7126_/CLK _7109_/D fanout456/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4810_ _4810_/A _4810_/B VGND VGND VPWR VPWR _4810_/Y sky130_fd_sc_hd__nor2_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _6920_/Q _5899_/B VGND VGND VPWR VPWR _5790_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_178_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4741_/A _4741_/B VGND VGND VPWR VPWR _4992_/B sky130_fd_sc_hd__nor2_1
X_4672_ _4672_/A _4672_/B VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__nor2_1
X_6411_ _3568_/A1 _6411_/D _6367_/X VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__dfrtp_1
X_3623_ _7021_/Q hold29/A _4127_/A _6543_/Q _3587_/X VGND VGND VPWR VPWR _3628_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6342_ _6642_/Q _6342_/A2 _6342_/B1 _6350_/A2 _6341_/X VGND VGND VPWR VPWR _6342_/X
+ sky130_fd_sc_hd__a221o_1
X_3554_ _3554_/A _3814_/B VGND VGND VPWR VPWR _4268_/A sky130_fd_sc_hd__nor2_4
XFILLER_142_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6273_ _6558_/Q _5971_/B _5949_/X _6678_/Q _6272_/X VGND VGND VPWR VPWR _6275_/C
+ sky130_fd_sc_hd__a221o_2
X_3485_ _3485_/A _3485_/B _3485_/C VGND VGND VPWR VPWR _3486_/B sky130_fd_sc_hd__and3_1
XFILLER_103_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5224_ hold200/X _5494_/A1 _5228_/S VGND VGND VPWR VPWR _5224_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5155_ _5155_/A0 _5491_/A1 _5160_/S VGND VGND VPWR VPWR _5155_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4106_ hold752/X _6356_/A1 _4108_/S VGND VGND VPWR VPWR _4106_/X sky130_fd_sc_hd__mux2_1
X_5086_ _5088_/A _5086_/B _5086_/C VGND VGND VPWR VPWR _5114_/D sky130_fd_sc_hd__and3_1
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4037_ hold582/X _6357_/A1 _4037_/S VGND VGND VPWR VPWR _4037_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _7047_/Q _5971_/A _5938_/X _6922_/Q _5980_/X VGND VGND VPWR VPWR _5989_/C
+ sky130_fd_sc_hd__a221o_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4939_ _4460_/A _4484_/Y _4967_/A _4563_/A _4923_/Y VGND VGND VPWR VPWR _5073_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA_40 _5300_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _5940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _6025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_73 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _6653_/CLK _6609_/D fanout454/X VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_84 _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_95 _6405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput180 _3209_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput191 _3199_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_csclk _6888_/CLK VGND VGND VPWR VPWR _7016_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _7171_/Q hold15/A _6487_/Q _3875_/B VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__o211a_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk _6447_/CLK VGND VGND VPWR VPWR _7053_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6960_ _6997_/CLK _6960_/D fanout465/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5911_ _3225_/Y _5899_/B _5651_/B VGND VGND VPWR VPWR _5911_/Y sky130_fd_sc_hd__a21oi_1
X_6891_ _7067_/CLK _6891_/D fanout477/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfstp_1
X_5842_ _5552_/B _7113_/Q _6103_/B1 _5841_/X VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5773_ hold56/A _5619_/X _5663_/X _6863_/Q VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4724_ _4724_/A _4972_/A VGND VGND VPWR VPWR _4775_/B sky130_fd_sc_hd__nand2_1
XFILLER_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4655_ _4626_/Y _4628_/Y _4653_/Y _4609_/Y VGND VGND VPWR VPWR _4655_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3606_ _6797_/Q _3326_/Y _4139_/A _6553_/Q _3605_/X VGND VGND VPWR VPWR _3611_/A
+ sky130_fd_sc_hd__a221o_1
Xhold800 _6823_/Q VGND VGND VPWR VPWR hold800/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_2
Xhold811 _4159_/X VGND VGND VPWR VPWR _6566_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4586_ _4563_/A _4951_/B _4942_/A _4583_/X VGND VGND VPWR VPWR _4586_/X sky130_fd_sc_hd__o211a_1
XFILLER_162_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold822 _6605_/Q VGND VGND VPWR VPWR hold822/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_4
Xhold833 _5156_/X VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 _6828_/Q VGND VGND VPWR VPWR hold844/X sky130_fd_sc_hd__dlygate4sd3_1
X_6325_ _6324_/X _6325_/A1 _6346_/S VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__mux2_1
X_3537_ _6926_/Q _5364_/A _3964_/A _6422_/Q _3536_/X VGND VGND VPWR VPWR _3538_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold855 _5241_/X VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 _6547_/Q VGND VGND VPWR VPWR hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold877 _4034_/X VGND VGND VPWR VPWR _6471_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _6652_/Q VGND VGND VPWR VPWR hold888/X sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ _6612_/Q _5943_/X _5981_/X _6658_/Q VGND VGND VPWR VPWR _6256_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold899 _5539_/X VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3468_ _7076_/Q _5532_/A _5319_/A _6887_/Q VGND VGND VPWR VPWR _3468_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5207_ hold766/X _5528_/A1 _5210_/S VGND VGND VPWR VPWR _5207_/X sky130_fd_sc_hd__mux2_1
X_6187_ _6460_/Q _5945_/X _5975_/C _6578_/Q VGND VGND VPWR VPWR _6187_/X sky130_fd_sc_hd__a22o_1
X_3399_ _6841_/Q _5265_/A hold76/A _7046_/Q _3398_/X VGND VGND VPWR VPWR _3409_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1500 hold4/A VGND VGND VPWR VPWR _6331_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1511 _3254_/X VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1522 hold11/A VGND VGND VPWR VPWR _6328_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5138_ _5138_/A _5138_/B _5138_/C VGND VGND VPWR VPWR _5138_/X sky130_fd_sc_hd__and3_1
Xhold1533 _7148_/Q VGND VGND VPWR VPWR _6346_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1544 _3248_/X VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 hold62/A VGND VGND VPWR VPWR _3858_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1566 _6637_/Q VGND VGND VPWR VPWR _3879_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 _6755_/Q VGND VGND VPWR VPWR hold1577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1588 _7177_/A VGND VGND VPWR VPWR hold405/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5069_ _5069_/A _5069_/B _5069_/C _5069_/D VGND VGND VPWR VPWR _5103_/B sky130_fd_sc_hd__and4_1
Xhold1599 _7089_/Q VGND VGND VPWR VPWR _5561_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4440_ _4690_/A _4495_/A VGND VGND VPWR VPWR _4724_/A sky130_fd_sc_hd__nor2_8
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold107 _3977_/X VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _6790_/Q VGND VGND VPWR VPWR hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold129 hold129/A VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4371_ _4702_/A _4566_/A VGND VGND VPWR VPWR _4374_/B sky130_fd_sc_hd__nor2_1
X_6110_ _6943_/Q _5961_/X _6108_/X _6109_/X VGND VGND VPWR VPWR _6115_/A sky130_fd_sc_hd__a211o_1
XFILLER_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3455_/A hold48/X VGND VGND VPWR VPWR _5193_/A sky130_fd_sc_hd__nor2_8
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _7113_/CLK _7090_/D fanout460/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6041_ _6900_/Q _5976_/C _5971_/D _6828_/Q VGND VGND VPWR VPWR _6041_/X sky130_fd_sc_hd__a22o_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3252_/Y _3253_/A1 _3253_/S VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__mux2_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _6541_/Q VGND VGND VPWR VPWR _3184_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6943_ _6999_/CLK _6943_/D fanout464/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6874_ _7051_/CLK _6874_/D fanout476/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_179_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5825_ _6695_/Q _5637_/X _5645_/X _6455_/Q VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5756_ _7109_/Q _5755_/X _6303_/S VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__mux2_1
X_4707_ _4716_/A _4911_/B _4707_/C VGND VGND VPWR VPWR _4707_/Y sky130_fd_sc_hd__nand3_2
X_5687_ _7011_/Q _5630_/X _5635_/X _6827_/Q _5686_/X VGND VGND VPWR VPWR _5690_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4638_ _4638_/A _4661_/B VGND VGND VPWR VPWR _4638_/Y sky130_fd_sc_hd__nand2_2
Xhold630 _6431_/Q VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold641 _3974_/X VGND VGND VPWR VPWR _6422_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _4636_/A _5043_/A _4737_/A VGND VGND VPWR VPWR _5099_/A sky130_fd_sc_hd__nand3_2
Xhold652 _6829_/Q VGND VGND VPWR VPWR hold652/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold663 _4217_/X VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap371 hold35/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__buf_12
XFILLER_162_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap382 _5660_/X VGND VGND VPWR VPWR _5913_/B1 sky130_fd_sc_hd__buf_6
X_6308_ _3828_/Y _6308_/A1 _6315_/S VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__mux2_1
Xhold674 _5353_/X VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 _6993_/Q VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 hold696/A VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6239_ _6462_/Q _5945_/X _5975_/C _6580_/Q _6238_/X VGND VGND VPWR VPWR _6240_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 hold1330/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
Xhold1341 hold1426/X VGND VGND VPWR VPWR hold1341/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1352 hold1352/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1363 _6309_/A1 VGND VGND VPWR VPWR hold1363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1374 hold1374/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _6529_/Q VGND VGND VPWR VPWR _4115_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 _7161_/Q VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3940_ _7105_/Q _6758_/Q _6762_/Q VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3871_ _3837_/B _3912_/B1 _3837_/C _6403_/Q VGND VGND VPWR VPWR _6403_/D sky130_fd_sc_hd__a31o_1
X_5610_ _6507_/Q _5610_/B VGND VGND VPWR VPWR _5610_/Y sky130_fd_sc_hd__nor2_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6590_ _7137_/CLK _6590_/D VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfxtp_1
X_5541_ _5541_/A _5541_/B VGND VGND VPWR VPWR _5549_/S sky130_fd_sc_hd__and2_4
XFILLER_191_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5472_ hold29/X _5541_/B VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__and2_4
XFILLER_144_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4423_ _4600_/B _4626_/B VGND VGND VPWR VPWR _4581_/B sky130_fd_sc_hd__nand2_8
XFILLER_132_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7142_ _3937_/A1 _7142_/D fanout487/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfrtp_1
X_4354_ _4642_/A _4357_/B VGND VGND VPWR VPWR _4356_/A sky130_fd_sc_hd__nor2_1
Xfanout406 _5494_/A1 VGND VGND VPWR VPWR _6356_/A1 sky130_fd_sc_hd__buf_6
Xfanout417 _5465_/A1 VGND VGND VPWR VPWR _5492_/A1 sky130_fd_sc_hd__buf_6
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout428 hold17/X VGND VGND VPWR VPWR _5490_/B sky130_fd_sc_hd__buf_4
X_3305_ _3313_/A hold27/X VGND VGND VPWR VPWR _3379_/A sky130_fd_sc_hd__nand2_8
X_7073_ _7083_/CLK _7073_/D _6390_/A VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_4
X_4285_ hold229/X hold60/X _4285_/S VGND VGND VPWR VPWR _4285_/X sky130_fd_sc_hd__mux2_1
X_6024_ _6024_/A _6024_/B _6024_/C _6024_/D VGND VGND VPWR VPWR _6025_/B sky130_fd_sc_hd__nor4_1
X_3236_ _6417_/Q _6416_/Q VGND VGND VPWR VPWR _3264_/B sky130_fd_sc_hd__and2_1
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3167_ hold44/A VGND VGND VPWR VPWR _3167_/Y sky130_fd_sc_hd__inv_2
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _6926_/CLK _6926_/D fanout457/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfrtp_4
X_6857_ _7086_/CLK _6857_/D fanout482/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5808_ _6945_/Q _5632_/X _5804_/X _5805_/X _5807_/X VGND VGND VPWR VPWR _5808_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6788_ _7012_/CLK hold19/X fanout458/X VGND VGND VPWR VPWR _6788_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5739_ _7022_/Q _5619_/X _5663_/X _6862_/Q VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold460 _5288_/X VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold471 _6662_/Q VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _4278_/X VGND VGND VPWR VPWR _6673_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold493 _6612_/Q VGND VGND VPWR VPWR hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1160 _5194_/X VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _6810_/Q VGND VGND VPWR VPWR _5239_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 _5185_/X VGND VGND VPWR VPWR _6764_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _6700_/Q VGND VGND VPWR VPWR _4311_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3568_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4070_ _4070_/A0 _4069_/X _4084_/S VGND VGND VPWR VPWR _4070_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4972_ _4972_/A _5010_/B VGND VGND VPWR VPWR _5008_/C sky130_fd_sc_hd__nand2_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6711_ _6714_/CLK _6711_/D fanout470/X VGND VGND VPWR VPWR _6711_/Q sky130_fd_sc_hd__dfrtp_1
X_3923_ _6518_/Q input80/X _3957_/B VGND VGND VPWR VPWR _3923_/X sky130_fd_sc_hd__mux2_8
XFILLER_189_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6642_ _7150_/CLK _6642_/D fanout487/X VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfrtp_4
X_3854_ _3284_/X _3283_/Y _3854_/S VGND VGND VPWR VPWR _3854_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6573_ _7140_/CLK _6573_/D VGND VGND VPWR VPWR _6573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3785_ _7039_/Q hold76/A _4322_/A _6710_/Q VGND VGND VPWR VPWR _3785_/X sky130_fd_sc_hd__a22o_2
XFILLER_164_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5524_ _5524_/A0 _5524_/A1 _5531_/S VGND VGND VPWR VPWR _5524_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5455_ _5455_/A0 _5524_/A1 _5462_/S VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4406_ _4739_/A _4415_/A VGND VGND VPWR VPWR _4570_/A sky130_fd_sc_hd__and2b_1
X_5386_ hold217/X _5494_/A1 _5390_/S VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7125_ _7126_/CLK _7125_/D fanout459/X VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4337_ _4337_/A _4337_/B _4337_/C _4337_/D VGND VGND VPWR VPWR _4338_/C sky130_fd_sc_hd__and4_1
XFILLER_59_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7056_ _7085_/CLK _7056_/D fanout485/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfstp_1
X_4268_ _4268_/A _5490_/B VGND VGND VPWR VPWR _4273_/S sky130_fd_sc_hd__and2_2
X_6007_ _7080_/Q _5976_/B _5954_/X _7056_/Q _6004_/X VGND VGND VPWR VPWR _6024_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3219_ _6821_/Q VGND VGND VPWR VPWR _3219_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4199_ _4199_/A0 _5544_/A1 _4201_/S VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6909_ _7076_/CLK _6909_/D fanout481/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold290 _5222_/X VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _3923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_141 _6226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_152 _5552_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_163 _5532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _5976_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _7173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 hold94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3570_ _7059_/Q hold86/A _4008_/A _6454_/Q VGND VGND VPWR VPWR _3570_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5240_ hold604/X _5543_/A1 _5246_/S VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5171_ _5186_/A _5171_/B _6352_/B VGND VGND VPWR VPWR _5172_/S sky130_fd_sc_hd__and3_1
XFILLER_96_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4122_ hold243/X _5494_/A1 _4126_/S VGND VGND VPWR VPWR _4122_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4053_ _4053_/A0 _4052_/X _4067_/S VGND VGND VPWR VPWR _4053_/X sky130_fd_sc_hd__mux2_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4955_ _5068_/A _4964_/B _5068_/B VGND VGND VPWR VPWR _5039_/D sky130_fd_sc_hd__and3_1
X_3906_ _3906_/A _3906_/B _3906_/C VGND VGND VPWR VPWR _3907_/D sky130_fd_sc_hd__and3_1
X_4886_ _5010_/A _4886_/B VGND VGND VPWR VPWR _4887_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6625_ _6629_/CLK _6625_/D _6390_/A VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfrtp_4
X_3837_ _3837_/A _3837_/B _3837_/C VGND VGND VPWR VPWR _3838_/B sky130_fd_sc_hd__and3_1
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6556_ _6629_/CLK _6556_/D _6390_/A VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfrtp_4
X_3768_ _6418_/Q _3964_/A _4014_/A _6455_/Q _3767_/X VGND VGND VPWR VPWR _3773_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5507_ hold558/X _5543_/A1 _5513_/S VGND VGND VPWR VPWR _5507_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6487_ _3945_/A1 _6487_/D _6376_/X VGND VGND VPWR VPWR _6487_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_173_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3699_ _3699_/A _3699_/B _3699_/C _3699_/D VGND VGND VPWR VPWR _3700_/C sky130_fd_sc_hd__and4_1
X_5438_ hold570/X _5543_/A1 _5444_/S VGND VGND VPWR VPWR _5438_/X sky130_fd_sc_hd__mux2_1
Xoutput340 hold1375/X VGND VGND VPWR VPWR hold1376/A sky130_fd_sc_hd__buf_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5369_ hold568/X _6357_/A1 _5372_/S VGND VGND VPWR VPWR _5369_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7108_ _7126_/CLK _7108_/D fanout456/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7039_ _7083_/CLK _7039_/D fanout470/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_75_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4740_/A _4740_/B VGND VGND VPWR VPWR _4741_/B sky130_fd_sc_hd__nand2_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4671_ _4671_/A VGND VGND VPWR VPWR _4679_/B sky130_fd_sc_hd__clkinv_2
X_6410_ _3568_/A1 _6410_/D _6366_/X VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__dfrtp_1
X_3622_ _6429_/Q _3981_/A _4304_/A _6698_/Q _3621_/X VGND VGND VPWR VPWR _3628_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6341_ _6644_/Q _6341_/A2 _6341_/B1 _6643_/Q VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__a22o_1
X_3553_ hold36/X _3562_/B VGND VGND VPWR VPWR _4298_/A sky130_fd_sc_hd__nor2_2
X_6272_ _7037_/Q _5601_/X _5959_/X _6718_/Q VGND VGND VPWR VPWR _6272_/X sky130_fd_sc_hd__a22o_1
X_3484_ _3484_/A _3484_/B _3484_/C _3484_/D VGND VGND VPWR VPWR _3485_/C sky130_fd_sc_hd__nor4_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5223_ hold381/X _5526_/A1 _5228_/S VGND VGND VPWR VPWR _5223_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5154_ _5154_/A _6352_/B VGND VGND VPWR VPWR _5160_/S sky130_fd_sc_hd__and2_2
XFILLER_111_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4105_ hold237/X _5544_/A1 _4108_/S VGND VGND VPWR VPWR _4105_/X sky130_fd_sc_hd__mux2_1
X_5085_ _5085_/A _5085_/B _5085_/C VGND VGND VPWR VPWR _5087_/D sky130_fd_sc_hd__and3_1
X_4036_ hold778/X _6356_/A1 _4037_/S VGND VGND VPWR VPWR _4036_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _6442_/Q _5601_/X _5981_/X _6914_/Q _5950_/X VGND VGND VPWR VPWR _5989_/B
+ sky130_fd_sc_hd__a221o_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4938_ _5068_/A _5046_/A _5068_/B _5103_/A VGND VGND VPWR VPWR _4941_/B sky130_fd_sc_hd__and4_1
XFILLER_178_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_30 _3612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4841_/X _4869_/B _4869_/C _4869_/D VGND VGND VPWR VPWR _4870_/C sky130_fd_sc_hd__and4b_1
XANTENNA_41 _5300_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 _5973_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_63 _6025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6608_ _6746_/CLK _6608_/D fanout448/X VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_119_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_74 _6268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _6467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _6406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6539_ _6539_/CLK _6539_/D fanout461/X VGND VGND VPWR VPWR _6539_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput181 _3208_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3198_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__1177_ clkbuf_0__1177_/X VGND VGND VPWR VPWR _6312_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5910_ _6618_/Q _5628_/X _5910_/B1 _6629_/Q VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__a22o_1
X_6890_ _6890_/CLK _6890_/D fanout476/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5841_ _6540_/Q _5652_/Y _5828_/X _5840_/X _6303_/S VGND VGND VPWR VPWR _5841_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5772_ _6903_/Q _5621_/X _5648_/X _6855_/Q _5771_/X VGND VGND VPWR VPWR _5772_/X
+ sky130_fd_sc_hd__a221o_1
X_4723_ _4984_/A _4723_/B VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__nand2_1
XFILLER_187_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4654_ _4619_/Y _4653_/Y _4846_/B VGND VGND VPWR VPWR _4654_/X sky130_fd_sc_hd__a21o_1
X_3605_ _6628_/Q _4232_/A _4244_/A _6648_/Q VGND VGND VPWR VPWR _3605_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_2
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold801 _5253_/X VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4585_ _5051_/A _4881_/B VGND VGND VPWR VPWR _4951_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold812 hold812/A VGND VGND VPWR VPWR hold812/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 _4204_/X VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_2
Xinput94 uart_enabled VGND VGND VPWR VPWR _3956_/B sky130_fd_sc_hd__clkbuf_1
Xhold834 _6701_/Q VGND VGND VPWR VPWR hold834/X sky130_fd_sc_hd__dlygate4sd3_1
X_6324_ _6644_/Q _6324_/A2 _6324_/B1 _6643_/Q _6323_/X VGND VGND VPWR VPWR _6324_/X
+ sky130_fd_sc_hd__a221o_1
X_3536_ _7075_/Q _5532_/A _4286_/A _6684_/Q VGND VGND VPWR VPWR _3536_/X sky130_fd_sc_hd__a22o_2
Xhold845 _5259_/X VGND VGND VPWR VPWR _6828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _6908_/Q VGND VGND VPWR VPWR hold856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 _4136_/X VGND VGND VPWR VPWR _6547_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold878 _7028_/Q VGND VGND VPWR VPWR hold878/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 _4253_/X VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ _6663_/Q _5976_/B _5971_/C _6713_/Q VGND VGND VPWR VPWR _6255_/X sky130_fd_sc_hd__a22o_1
X_3467_ _3467_/A _3467_/B _3467_/C _3467_/D VGND VGND VPWR VPWR _3467_/Y sky130_fd_sc_hd__nor4_1
X_5206_ hold904/X _5509_/A1 _5210_/S VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6186_ _6450_/Q _5947_/X _5965_/X _6545_/Q _6185_/X VGND VGND VPWR VPWR _6189_/B
+ sky130_fd_sc_hd__a221o_1
X_3398_ input28/X _3367_/Y _3964_/A _6425_/Q _3384_/X VGND VGND VPWR VPWR _3398_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1501 _7120_/Q VGND VGND VPWR VPWR _6028_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1512 _6598_/Q VGND VGND VPWR VPWR _4195_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5137_ _4428_/Y _4542_/D _4846_/B _4653_/Y _4769_/A VGND VGND VPWR VPWR _5138_/C
+ sky130_fd_sc_hd__o221a_1
Xhold1523 _7144_/Q VGND VGND VPWR VPWR _6334_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _7123_/Q VGND VGND VPWR VPWR _6104_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1545 _7183_/A VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 _6506_/Q VGND VGND VPWR VPWR _3894_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1567 _6417_/Q VGND VGND VPWR VPWR _3834_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_5068_ _5068_/A _5068_/B _5068_/C VGND VGND VPWR VPWR _5069_/D sky130_fd_sc_hd__and3_1
Xhold1578 _6538_/Q VGND VGND VPWR VPWR hold1578/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1589 _6532_/Q VGND VGND VPWR VPWR hold1589/X sky130_fd_sc_hd__dlygate4sd3_1
X_4019_ hold616/X _6357_/A1 _4019_/S VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold108 hold98/X VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold119 _5216_/X VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4370_ _4556_/A _4441_/A VGND VGND VPWR VPWR _4495_/A sky130_fd_sc_hd__nand2_4
XFILLER_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3321_ hold47/X _3454_/B VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__nand2_8
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6040_/B _6040_/C VGND VGND VPWR VPWR _6040_/Y sky130_fd_sc_hd__nor3_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _7167_/Q _6485_/Q _3262_/C VGND VGND VPWR VPWR _3252_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_79_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3183_ _6655_/Q VGND VGND VPWR VPWR _3183_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6942_ _7006_/CLK _6942_/D fanout457/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6873_ _7070_/CLK _6873_/D fanout473/X VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5824_ _6599_/Q _5616_/X _5655_/X _6545_/Q _5823_/X VGND VGND VPWR VPWR _5824_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5755_ wire367/X _5754_/Y _6790_/Q _5652_/Y VGND VGND VPWR VPWR _5755_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4706_ _4693_/X _4706_/B _4706_/C _4706_/D VGND VGND VPWR VPWR _4722_/B sky130_fd_sc_hd__and4b_1
X_5686_ _6851_/Q _5648_/X _5910_/B1 _6883_/Q VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4637_ _4638_/A _4661_/B VGND VGND VPWR VPWR _4707_/C sky130_fd_sc_hd__and2_2
XFILLER_147_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold620 _6430_/Q VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _3987_/X VGND VGND VPWR VPWR _6431_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _4664_/B _4568_/B VGND VGND VPWR VPWR _4741_/A sky130_fd_sc_hd__nand2b_2
Xhold642 _6657_/Q VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold653 _5260_/X VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap361 hold37/X VGND VGND VPWR VPWR _4058_/S sky130_fd_sc_hd__buf_6
X_3519_ _6910_/Q _5346_/A _4214_/A _6618_/Q _3518_/X VGND VGND VPWR VPWR _3523_/C
+ sky130_fd_sc_hd__a221o_1
X_6307_ _6636_/Q _6307_/B VGND VGND VPWR VPWR _6315_/S sky130_fd_sc_hd__nand2_4
Xhold664 _7141_/Q VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap383 _5658_/X VGND VGND VPWR VPWR _5910_/B1 sky130_fd_sc_hd__buf_8
Xhold675 _6913_/Q VGND VGND VPWR VPWR hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _5444_/X VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4499_ _5051_/B _4582_/B VGND VGND VPWR VPWR _4535_/A sky130_fd_sc_hd__nand2_1
Xhold697 _5179_/X VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6238_ _6667_/Q _5938_/X _5952_/X _6707_/Q VGND VGND VPWR VPWR _6238_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _7054_/Q _5971_/A _5979_/X _6993_/Q VGND VGND VPWR VPWR _6169_/X sky130_fd_sc_hd__a22o_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 hold1320/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
Xhold1331 hold1420/X VGND VGND VPWR VPWR hold1331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1342 hold1342/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1353 _4183_/A1 VGND VGND VPWR VPWR hold1353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 hold1364/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
XFILLER_45_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1375 _4192_/A1 VGND VGND VPWR VPWR hold1375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 _7044_/Q VGND VGND VPWR VPWR _5502_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1397 _7086_/Q VGND VGND VPWR VPWR _5549_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_43_csclk _6888_/CLK VGND VGND VPWR VPWR _6920_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_csclk _6447_/CLK VGND VGND VPWR VPWR _6953_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3870_ _6404_/Q _3912_/A1 _3870_/S VGND VGND VPWR VPWR _6404_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ hold397/X _5540_/A1 _5540_/S VGND VGND VPWR VPWR _5540_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5471_ hold626/X _5513_/A1 _5471_/S VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4422_ _4607_/A _4947_/A VGND VGND VPWR VPWR _4921_/A sky130_fd_sc_hd__nor2_4
X_7141_ _7150_/CLK _7141_/D fanout487/X VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4353_ _4379_/B _4360_/B VGND VGND VPWR VPWR _4896_/A sky130_fd_sc_hd__and2_1
Xfanout407 hold156/X VGND VGND VPWR VPWR _5494_/A1 sky130_fd_sc_hd__buf_12
Xfanout418 hold13/X VGND VGND VPWR VPWR _5465_/A1 sky130_fd_sc_hd__clkbuf_16
X_3304_ _3313_/A hold27/X VGND VGND VPWR VPWR _5190_/A sky130_fd_sc_hd__and2_4
X_7072_ _7083_/CLK _7072_/D fanout470/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfstp_4
X_4284_ hold194/X _5494_/A1 _4285_/S VGND VGND VPWR VPWR _4284_/X sky130_fd_sc_hd__mux2_1
Xfanout429 hold16/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__buf_8
XFILLER_98_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6023_ _6811_/Q _5971_/B _5949_/X _6931_/Q _6022_/X VGND VGND VPWR VPWR _6024_/D
+ sky130_fd_sc_hd__a221o_2
X_3235_ _3235_/A0 _3251_/A _3235_/S VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3166_ _6415_/Q VGND VGND VPWR VPWR _3837_/A sky130_fd_sc_hd__clkinv_2
XFILLER_27_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6925_/CLK _6925_/D fanout461/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6856_ _6981_/CLK _6856_/D fanout464/X VGND VGND VPWR VPWR _6856_/Q sky130_fd_sc_hd__dfrtp_1
X_5807_ _7017_/Q _5630_/X _5638_/X _6961_/Q _5806_/X VGND VGND VPWR VPWR _5807_/X
+ sky130_fd_sc_hd__a221o_1
X_6787_ _7012_/CLK _6787_/D fanout458/X VGND VGND VPWR VPWR _6787_/Q sky130_fd_sc_hd__dfstp_1
X_3999_ _3999_/A _5541_/B VGND VGND VPWR VPWR _4007_/S sky130_fd_sc_hd__and2_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5738_ _6966_/Q _5642_/X _5667_/X _6814_/Q VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5669_ _5669_/A _5669_/B _5669_/C _5669_/D VGND VGND VPWR VPWR _5670_/B sky130_fd_sc_hd__nor4_1
XFILLER_136_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold450 _5352_/X VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold461 _6627_/Q VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _4265_/X VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _7051_/Q VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _4212_/X VGND VGND VPWR VPWR _6612_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1150 _5347_/X VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1161 _7018_/Q VGND VGND VPWR VPWR _5473_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 _5239_/X VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1183 _6455_/Q VGND VGND VPWR VPWR _4015_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _4311_/X VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _4691_/A _4902_/B _4625_/B _4645_/Y VGND VGND VPWR VPWR _4974_/B sky130_fd_sc_hd__a31o_1
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6710_ _6714_/CLK _6710_/D fanout470/X VGND VGND VPWR VPWR _6710_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3922_ _3188_/Y input82/X _3957_/B VGND VGND VPWR VPWR _3922_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3853_ _3853_/A _3853_/B VGND VGND VPWR VPWR _6412_/D sky130_fd_sc_hd__xnor2_1
XFILLER_177_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6641_ _7150_/CLK _6641_/D fanout487/X VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfrtp_1
X_3784_ _6954_/Q _5400_/A _5154_/A _6742_/Q _3783_/X VGND VGND VPWR VPWR _3793_/A
+ sky130_fd_sc_hd__a221o_1
X_6572_ _7140_/CLK _6572_/D VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5523_ _5523_/A _5541_/B VGND VGND VPWR VPWR _5531_/S sky130_fd_sc_hd__and2_4
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5454_ _5454_/A hold17/X VGND VGND VPWR VPWR _5461_/S sky130_fd_sc_hd__and2_4
XFILLER_105_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4405_ _4459_/A _4549_/A VGND VGND VPWR VPWR _4810_/A sky130_fd_sc_hd__nand2_4
X_5385_ hold399/X _5526_/A1 _5390_/S VGND VGND VPWR VPWR _5385_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7124_ _7131_/CLK _7124_/D fanout459/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4336_ _4336_/A _4336_/B _4336_/C _4336_/D VGND VGND VPWR VPWR _4338_/B sky130_fd_sc_hd__and4_1
XFILLER_113_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7055_ _7079_/CLK _7055_/D _6396_/A VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4267_ hold830/X _5546_/A1 _4267_/S VGND VGND VPWR VPWR _4267_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6006_ _7003_/Q _5958_/X _5978_/X _6995_/Q VGND VGND VPWR VPWR _6006_/X sky130_fd_sc_hd__a22o_1
X_3218_ _6829_/Q VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__inv_2
X_4198_ _4198_/A0 _5492_/A1 _4201_/S VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ _6908_/CLK _6908_/D fanout475/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_1
X_6839_ _6865_/CLK _6839_/D fanout464/X VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold280 _5188_/X VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 hold291/A VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _3925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 _6279_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_153 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _4157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_175 _5975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_186 _7118_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_197 hold99/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5170_ hold211/X _5494_/A1 _5170_/S VGND VGND VPWR VPWR _5170_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4121_ hold401/X _5526_/A1 _4126_/S VGND VGND VPWR VPWR _4121_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4052_ _4110_/A0 _5473_/A1 _4058_/S VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__mux2_1
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4954_ _4413_/Y _4946_/X _5047_/A _5057_/B _4953_/Y VGND VGND VPWR VPWR _4962_/B
+ sky130_fd_sc_hd__o2111a_1
X_3905_ _4336_/C _4336_/D _4335_/A _4335_/B VGND VGND VPWR VPWR _3906_/C sky130_fd_sc_hd__nor4_1
X_4885_ _4884_/X _4839_/X _5006_/A _4885_/B2 VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6624_ _7150_/CLK _6624_/D fanout487/X VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_4
X_3836_ _3836_/A _3836_/B VGND VGND VPWR VPWR _6416_/D sky130_fd_sc_hd__nor2_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3767_ _7047_/Q _5505_/A _5166_/A _6751_/Q VGND VGND VPWR VPWR _3767_/X sky130_fd_sc_hd__a22o_1
X_6555_ _6712_/CLK _6555_/D fanout470/X VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5506_ _5506_/A0 _5524_/A1 _5513_/S VGND VGND VPWR VPWR _5506_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6486_ _3945_/A1 _6486_/D _6375_/X VGND VGND VPWR VPWR _6486_/Q sky130_fd_sc_hd__dfrtp_1
X_3698_ _3698_/A _3698_/B _3698_/C _3698_/D VGND VGND VPWR VPWR _3699_/D sky130_fd_sc_hd__nor4_1
X_5437_ _5437_/A0 _5524_/A1 _5444_/S VGND VGND VPWR VPWR _5437_/X sky130_fd_sc_hd__mux2_1
Xoutput330 hold1373/X VGND VGND VPWR VPWR hold1374/A sky130_fd_sc_hd__buf_12
XFILLER_160_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput341 hold1331/X VGND VGND VPWR VPWR hold1332/A sky130_fd_sc_hd__buf_12
XFILLER_160_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5368_ hold241/X _5494_/A1 _5372_/S VGND VGND VPWR VPWR _5368_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7107_ _7126_/CLK _7107_/D fanout456/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4319_ hold954/X _6355_/A1 _4321_/S VGND VGND VPWR VPWR _4319_/X sky130_fd_sc_hd__mux2_1
X_5299_ hold669/X _5521_/A1 _5300_/S VGND VGND VPWR VPWR _5299_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7038_ _7038_/CLK _7038_/D fanout455/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4670_ _4928_/A _4676_/B VGND VGND VPWR VPWR _4671_/A sky130_fd_sc_hd__and2_1
XFILLER_187_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3621_ _6981_/Q _5427_/A _4020_/A _6463_/Q VGND VGND VPWR VPWR _3621_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3552_ _3552_/A _3552_/B _3552_/C _3552_/D VGND VGND VPWR VPWR _3581_/B sky130_fd_sc_hd__nor4_1
X_6340_ _6339_/X _6340_/A1 _6346_/S VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6271_ _6458_/Q _5944_/X _5975_/A _6602_/Q _6270_/X VGND VGND VPWR VPWR _6275_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3483_ _6895_/Q _5328_/A _5256_/A _6831_/Q _3482_/X VGND VGND VPWR VPWR _3484_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5222_ hold289/X _5465_/A1 _5228_/S VGND VGND VPWR VPWR _5222_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5153_ hold564/X _6357_/A1 _5153_/S VGND VGND VPWR VPWR _5153_/X sky130_fd_sc_hd__mux2_1
X_4104_ _4104_/A0 _5492_/A1 _4108_/S VGND VGND VPWR VPWR _4104_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5084_ _5084_/A _5084_/B _5084_/C _5084_/D VGND VGND VPWR VPWR _5085_/C sky130_fd_sc_hd__and4_1
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4035_ hold948/X _6355_/A1 _4037_/S VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _7039_/Q _5971_/C _5982_/X _5985_/X VGND VGND VPWR VPWR _5989_/A sky130_fd_sc_hd__a211o_1
XFILLER_80_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4937_ _4921_/A _4737_/A _4668_/C _4671_/A _4922_/X VGND VGND VPWR VPWR _4996_/C
+ sky130_fd_sc_hd__a311oi_2
XANTENNA_20 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _3618_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4846_/A _4672_/B _4643_/Y _4694_/Y _4442_/Y VGND VGND VPWR VPWR _4869_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA_42 _5300_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _5948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_64 _6051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _6707_/CLK _6607_/D fanout447/X VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_75 _6276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ _6555_/Q _4145_/A _3692_/Y _6767_/Q _3818_/X VGND VGND VPWR VPWR _3826_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_86 _7021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _4483_/Y _4673_/A _5008_/A _4798_/X VGND VGND VPWR VPWR _4799_/X sky130_fd_sc_hd__o211a_1
XANTENNA_97 _6406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6538_ _6735_/CLK _6538_/D _6360_/A VGND VGND VPWR VPWR _6538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6469_ _6654_/CLK hold69/X fanout454/X VGND VGND VPWR VPWR _6469_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_121_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput171 _3958_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
XFILLER_161_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput182 _3207_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 _3197_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5840_ _6450_/Q _5634_/X _5829_/X _5833_/X _5839_/X VGND VGND VPWR VPWR _5840_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_62_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5771_ _6871_/Q _5628_/X _5658_/X _6887_/Q VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4722_ _4722_/A _4722_/B _4722_/C _4722_/D VGND VGND VPWR VPWR _4725_/B sky130_fd_sc_hd__and4_1
XFILLER_187_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4653_ _4716_/A _4653_/B _4653_/C VGND VGND VPWR VPWR _4653_/Y sky130_fd_sc_hd__nand3_4
XFILLER_147_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
X_3604_ _3604_/A _3604_/B _3604_/C _3604_/D VGND VGND VPWR VPWR _3604_/Y sky130_fd_sc_hd__nor4_1
XFILLER_162_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
X_4584_ _4584_/A _5043_/A VGND VGND VPWR VPWR _4942_/A sky130_fd_sc_hd__nand2_1
Xhold802 _6966_/Q VGND VGND VPWR VPWR hold802/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_2
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _3952_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_116_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_2
Xhold813 _4114_/X VGND VGND VPWR VPWR _6528_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_4
Xhold824 hold824/A VGND VGND VPWR VPWR hold824/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6323_ _6642_/Q _6323_/A2 _6323_/B1 _4230_/B VGND VGND VPWR VPWR _6323_/X sky130_fd_sc_hd__a22o_1
Xhold835 _4312_/X VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3535_ hold36/X _3571_/B VGND VGND VPWR VPWR _4286_/A sky130_fd_sc_hd__nor2_2
Xhold846 _6456_/Q VGND VGND VPWR VPWR hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 _5349_/X VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold868 _6892_/Q VGND VGND VPWR VPWR hold868/X sky130_fd_sc_hd__dlygate4sd3_1
X_6254_ _6278_/A0 _6253_/X _6279_/S VGND VGND VPWR VPWR _6254_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3466_ _6983_/Q _5427_/A _5247_/A _6823_/Q _3460_/X VGND VGND VPWR VPWR _3467_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold879 _5484_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5205_ _5205_/A0 _5484_/A1 _5210_/S VGND VGND VPWR VPWR _5205_/X sky130_fd_sc_hd__mux2_1
X_3397_ _3959_/B _4083_/S _5211_/A _6793_/Q _3396_/X VGND VGND VPWR VPWR _3409_/A
+ sky130_fd_sc_hd__a221o_1
X_6185_ _6630_/Q _5946_/X _5955_/X _6550_/Q VGND VGND VPWR VPWR _6185_/X sky130_fd_sc_hd__a22o_1
Xhold1502 _6028_/X VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _7119_/Q VGND VGND VPWR VPWR _6003_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5136_ _6726_/Q _4229_/X _5112_/X _5135_/Y VGND VGND VPWR VPWR _5136_/X sky130_fd_sc_hd__a22o_1
Xhold1524 _7109_/Q VGND VGND VPWR VPWR _5736_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1535 _6584_/Q VGND VGND VPWR VPWR _4180_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1546 _7115_/Q VGND VGND VPWR VPWR _5865_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 _7132_/Q VGND VGND VPWR VPWR hold1557/X sky130_fd_sc_hd__dlygate4sd3_1
X_5067_ _5134_/B _5066_/X _5006_/Y VGND VGND VPWR VPWR _5067_/Y sky130_fd_sc_hd__a21oi_1
Xhold1568 _7093_/Q VGND VGND VPWR VPWR _5575_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1579 _6416_/Q VGND VGND VPWR VPWR _3835_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4018_ hold756/X _6356_/A1 _4019_/S VGND VGND VPWR VPWR _4018_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5969_ _5969_/A _5979_/A _5969_/C VGND VGND VPWR VPWR _5971_/D sky130_fd_sc_hd__and3_4
XFILLER_185_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold109 _3978_/X VGND VGND VPWR VPWR _6424_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3320_ hold47/X _3453_/A hold64/X VGND VGND VPWR VPWR _3320_/X sky130_fd_sc_hd__and3_2
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3251_/A _6485_/Q VGND VGND VPWR VPWR _3262_/C sky130_fd_sc_hd__nand2_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3182_ _6489_/Q VGND VGND VPWR VPWR _3182_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6941_ _7054_/CLK _6941_/D fanout461/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6872_ _6920_/CLK _6872_/D fanout473/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5823_ _6470_/Q _5627_/X _5635_/X _6565_/Q VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__a22o_1
X_5754_ _5754_/A _5754_/B _5754_/C VGND VGND VPWR VPWR _5754_/Y sky130_fd_sc_hd__nor3_2
XFILLER_148_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4705_ _4689_/A _4644_/Y _4702_/Y _4673_/A _4704_/X VGND VGND VPWR VPWR _4706_/D
+ sky130_fd_sc_hd__o221a_1
X_5685_ _6979_/Q _5624_/X _5654_/X _6931_/Q _5684_/X VGND VGND VPWR VPWR _5690_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4636_ _4636_/A _4646_/A VGND VGND VPWR VPWR _4658_/C sky130_fd_sc_hd__nand2_1
XFILLER_147_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold610 _6511_/Q VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 _3986_/X VGND VGND VPWR VPWR _6430_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4567_ _4664_/B _4568_/B VGND VGND VPWR VPWR _4737_/A sky130_fd_sc_hd__and2b_2
Xhold632 _6841_/Q VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 _4259_/X VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold654 _6929_/Q VGND VGND VPWR VPWR hold654/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap362 _3331_/Y VGND VGND VPWR VPWR _5202_/B sky130_fd_sc_hd__buf_6
X_6306_ _6636_/Q _3910_/B _6305_/Y _6306_/B2 VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__a22o_1
X_3518_ _6474_/Q _4032_/A _4038_/A _6479_/Q VGND VGND VPWR VPWR _3518_/X sky130_fd_sc_hd__a22o_1
Xmax_cap373 _3555_/A VGND VGND VPWR VPWR _3554_/A sky130_fd_sc_hd__buf_12
Xhold665 hold665/A VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap384 _5657_/X VGND VGND VPWR VPWR _5928_/A2 sky130_fd_sc_hd__buf_8
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold676 _5354_/X VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _4498_/A _4843_/B VGND VGND VPWR VPWR _4498_/Y sky130_fd_sc_hd__nand2_1
Xhold687 _6801_/Q VGND VGND VPWR VPWR hold687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold698 _6983_/Q VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__dlygate4sd3_1
X_6237_ _6452_/Q _5947_/X _5965_/X _6547_/Q _6236_/X VGND VGND VPWR VPWR _6240_/B
+ sky130_fd_sc_hd__a221o_1
X_3449_ _3448_/X _3449_/A1 _3829_/B VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6825_/Q _5953_/X _5960_/X _7078_/Q _6167_/X VGND VGND VPWR VPWR _6168_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _4033_/X VGND VGND VPWR VPWR _6470_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1321 hold1415/X VGND VGND VPWR VPWR hold1321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 hold1332/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_85_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1343 hold1427/X VGND VGND VPWR VPWR hold1343/X sky130_fd_sc_hd__dlygate4sd3_1
X_5119_ _4465_/B _4644_/B _4975_/B _4450_/Y VGND VGND VPWR VPWR _5120_/C sky130_fd_sc_hd__a31oi_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1354 hold1354/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
X_6099_ _6099_/A _6099_/B _6099_/C _6099_/D VGND VGND VPWR VPWR _6100_/C sky130_fd_sc_hd__nor4_1
Xhold1365 _4189_/A1 VGND VGND VPWR VPWR hold1365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1376 hold1376/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_84_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1387 _7060_/Q VGND VGND VPWR VPWR _5520_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _7145_/Q VGND VGND VPWR VPWR _3973_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7113_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5470_ hold750/X _5521_/A1 _5471_/S VGND VGND VPWR VPWR _5470_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4421_ _4753_/A _4607_/A VGND VGND VPWR VPWR _4626_/B sky130_fd_sc_hd__nor2_8
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7140_ _7140_/CLK _7140_/D VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfxtp_1
X_4352_ _4633_/B _4352_/B VGND VGND VPWR VPWR _4360_/B sky130_fd_sc_hd__xor2_1
XFILLER_125_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3303_ hold26/X hold46/X VGND VGND VPWR VPWR _3303_/Y sky130_fd_sc_hd__nor2_8
Xfanout408 _5509_/A1 VGND VGND VPWR VPWR _5545_/A1 sky130_fd_sc_hd__buf_6
X_4283_ _4283_/A0 _5493_/A1 _4285_/S VGND VGND VPWR VPWR _4283_/X sky130_fd_sc_hd__mux2_1
X_7071_ _7083_/CLK _7071_/D fanout470/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfstp_2
Xfanout419 _5534_/A1 VGND VGND VPWR VPWR _5543_/A1 sky130_fd_sc_hd__buf_6
XFILLER_58_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6022_ _6443_/Q _5601_/X _5959_/X _6963_/Q VGND VGND VPWR VPWR _6022_/X sky130_fd_sc_hd__a22o_1
X_3234_ _6415_/Q _6485_/Q _3234_/C VGND VGND VPWR VPWR _3235_/S sky130_fd_sc_hd__and3_1
XFILLER_101_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3165_ _7158_/Q VGND VGND VPWR VPWR _3165_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6924_ _7006_/CLK _6924_/D fanout458/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6855_ _6865_/CLK _6855_/D fanout464/X VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5806_ _7009_/Q _5625_/X _5661_/X _6881_/Q VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__a22o_1
X_6786_ _7006_/CLK _6786_/D fanout456/X VGND VGND VPWR VPWR _6786_/Q sky130_fd_sc_hd__dfstp_1
X_3998_ hold523/X _5513_/A1 _3998_/S VGND VGND VPWR VPWR _3998_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5737_ _6958_/Q _5638_/X _5661_/X _6878_/Q VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5668_ _6890_/Q _5666_/X _5667_/X _6810_/Q _5665_/X VGND VGND VPWR VPWR _5669_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4619_ _4716_/A _4653_/B _4635_/B VGND VGND VPWR VPWR _4619_/Y sky130_fd_sc_hd__nand3_4
XFILLER_190_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5599_ _5597_/B _5598_/Y _5602_/B VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__a21oi_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold440 _5441_/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold451 _6806_/Q VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold462 _4235_/X VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold473 _6918_/Q VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold484 _5510_/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _6617_/Q VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1140 _5191_/X VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1151 _6866_/Q VGND VGND VPWR VPWR _5302_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _5473_/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 _6555_/Q VGND VGND VPWR VPWR _4146_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _4015_/X VGND VGND VPWR VPWR _6455_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1195 _6850_/Q VGND VGND VPWR VPWR _5284_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4970_ _4970_/A _4975_/B VGND VGND VPWR VPWR _4970_/Y sky130_fd_sc_hd__nor2_2
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3921_ _3187_/Y input90/X _3921_/S VGND VGND VPWR VPWR _3921_/X sky130_fd_sc_hd__mux2_2
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6640_ _7150_/CLK _6640_/D fanout487/X VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3852_ _3852_/A _3860_/B VGND VGND VPWR VPWR _3853_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6571_ _7137_/CLK _6571_/D VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfxtp_1
X_3783_ _6685_/Q _4292_/A _5490_/A _7034_/Q VGND VGND VPWR VPWR _3783_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5522_ hold313/X _5540_/A1 hold87/X VGND VGND VPWR VPWR _5522_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5453_ hold497/X hold22/X _5453_/S VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4404_ _4408_/B _4448_/B VGND VGND VPWR VPWR _4549_/A sky130_fd_sc_hd__nor2_4
X_5384_ hold301/X _5465_/A1 _5390_/S VGND VGND VPWR VPWR _5384_/X sky130_fd_sc_hd__mux2_1
X_7123_ _7131_/CLK _7123_/D fanout459/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_1
X_4335_ _4335_/A _4335_/B _4335_/C _4335_/D VGND VGND VPWR VPWR _4338_/A sky130_fd_sc_hd__and4_1
XFILLER_87_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7054_ _7054_/CLK _7054_/D fanout461/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfrtp_1
X_4266_ hold347/X _5518_/A1 _4267_/S VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_57_csclk _6447_/CLK VGND VGND VPWR VPWR _6925_/CLK sky130_fd_sc_hd__clkbuf_16
X_6005_ _6859_/Q _5943_/X _5981_/X _6915_/Q VGND VGND VPWR VPWR _6005_/X sky130_fd_sc_hd__a22o_1
X_3217_ _6837_/Q VGND VGND VPWR VPWR _3217_/Y sky130_fd_sc_hd__inv_2
X_4197_ hold976/X hold666/X _4201_/S VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6907_ _7082_/CLK _6907_/D fanout479/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfstp_1
X_6838_ _7026_/CLK _6838_/D fanout463/X VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6769_ _6769_/CLK _6769_/D fanout469/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold270 _4288_/X VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _6556_/Q VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _5209_/X VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _3956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_121 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_132 _6747_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _5902_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 hold6/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _4238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _5960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_187 _3957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _5171_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4120_ hold824/X _6354_/A1 _4126_/S VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4051_ _6396_/B _3692_/A hold37/X _4050_/X _4322_/B VGND VGND VPWR VPWR _4067_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_83_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4953_ _4953_/A _5043_/B VGND VGND VPWR VPWR _4953_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3904_ _4335_/C _4335_/D _3904_/C VGND VGND VPWR VPWR _3906_/B sky130_fd_sc_hd__nor3_1
X_4884_ _5006_/A _4884_/B _4884_/C _4884_/D VGND VGND VPWR VPWR _4884_/X sky130_fd_sc_hd__and4_1
X_6623_ _6712_/CLK _6623_/D _6390_/A VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfrtp_4
X_3835_ _3835_/A _3838_/A VGND VGND VPWR VPWR _3836_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6554_ _6674_/CLK _6554_/D _6383_/A VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3766_ input52/X _5193_/A _4220_/A _6619_/Q _3765_/X VGND VGND VPWR VPWR _3773_/A
+ sky130_fd_sc_hd__a221o_1
X_5505_ _5505_/A _5505_/B VGND VGND VPWR VPWR _5513_/S sky130_fd_sc_hd__and2_4
XFILLER_192_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6485_ _3927_/A1 _6485_/D _6374_/X VGND VGND VPWR VPWR _6485_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_146_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3697_ _6820_/Q _5247_/A _4298_/A _6692_/Q _3696_/X VGND VGND VPWR VPWR _3698_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5436_ _5436_/A _5505_/B VGND VGND VPWR VPWR _5444_/S sky130_fd_sc_hd__and2_4
Xoutput320 hold1339/X VGND VGND VPWR VPWR hold1340/A sky130_fd_sc_hd__buf_12
XFILLER_105_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput331 hold1363/X VGND VGND VPWR VPWR hold1364/A sky130_fd_sc_hd__buf_12
Xoutput342 hold1335/X VGND VGND VPWR VPWR hold1336/A sky130_fd_sc_hd__buf_12
XFILLER_161_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5367_ hold325/X _5526_/A1 _5372_/S VGND VGND VPWR VPWR _5367_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7106_ _7126_/CLK _7106_/D fanout456/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_1
X_4318_ hold814/X _6354_/A1 _4321_/S VGND VGND VPWR VPWR _4318_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5298_ hold160/X hold42/X _5300_/S VGND VGND VPWR VPWR _5298_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7037_ _7037_/CLK _7037_/D fanout450/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4249_ hold525/X _5546_/A1 _4249_/S VGND VGND VPWR VPWR _4249_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3620_ _3620_/A _3620_/B _3620_/C _3620_/D VGND VGND VPWR VPWR _3639_/A sky130_fd_sc_hd__nor4_1
XFILLER_147_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3551_ _6830_/Q _5256_/A _4196_/A _6603_/Q _3549_/X VGND VGND VPWR VPWR _3552_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6270_ _6468_/Q _5937_/X _5975_/D _6628_/Q VGND VGND VPWR VPWR _6270_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3482_ input57/X _5193_/A _5541_/A _7084_/Q VGND VGND VPWR VPWR _3482_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5221_ _5221_/A0 _5524_/A1 _5228_/S VGND VGND VPWR VPWR _5221_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5152_ hold728/X _6356_/A1 _5153_/S VGND VGND VPWR VPWR _5152_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4103_ _4103_/A0 _5491_/A1 _4108_/S VGND VGND VPWR VPWR _4103_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5083_ _5083_/A _5083_/B _5083_/C VGND VGND VPWR VPWR _5115_/C sky130_fd_sc_hd__and3_1
XFILLER_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4034_ hold876/X _6354_/A1 _4037_/S VGND VGND VPWR VPWR _4034_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5985_ _7018_/Q _5937_/X _5944_/X _7026_/Q _5984_/X VGND VGND VPWR VPWR _5985_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4936_ _4999_/B _5003_/B _5076_/A VGND VGND VPWR VPWR _4944_/B sky130_fd_sc_hd__and3_1
XANTENNA_10 _3355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _3504_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4902_/B _4639_/Y _4508_/C VGND VGND VPWR VPWR _5027_/B sky130_fd_sc_hd__o21a_1
XANTENNA_32 _3638_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_43 _5399_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _6746_/CLK _6606_/D fanout447/X VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_54 _5976_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3818_ _6898_/Q _5337_/A _4232_/A _6625_/Q VGND VGND VPWR VPWR _3818_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _6276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _4627_/B _4638_/Y _4673_/A _4627_/A VGND VGND VPWR VPWR _4798_/X sky130_fd_sc_hd__a211o_1
XANTENNA_87 _7040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 _7157_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ _6537_/CLK _6537_/D fanout464/X VGND VGND VPWR VPWR _6537_/Q sky130_fd_sc_hd__dfrtp_1
X_3749_ _6835_/Q _5265_/A _4008_/A _6451_/Q VGND VGND VPWR VPWR _3749_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6468_ _6654_/CLK _6468_/D _6401_/A VGND VGND VPWR VPWR _6468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5419_ _5419_/A0 _5524_/A1 _5426_/S VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__mux2_1
X_6399_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__and2_1
XFILLER_121_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput172 _7173_/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
Xoutput183 _3206_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 _3196_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5770_ _6983_/Q _5624_/X _5634_/X _6975_/Q _5758_/Y VGND VGND VPWR VPWR _5770_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4721_/A _4721_/B _4721_/C VGND VGND VPWR VPWR _4722_/D sky130_fd_sc_hd__and3_1
X_4652_ _4653_/B _4653_/C VGND VGND VPWR VPWR _4652_/Y sky130_fd_sc_hd__nand2_4
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__buf_2
XFILLER_147_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3603_ _6805_/Q _5229_/A _4145_/A _6558_/Q _3588_/X VGND VGND VPWR VPWR _3604_/D
+ sky130_fd_sc_hd__a221o_1
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4583_ _4581_/B _4582_/Y _4810_/A VGND VGND VPWR VPWR _4583_/X sky130_fd_sc_hd__a21o_1
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_4
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _3957_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_162_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold803 _5414_/X VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 _6706_/Q VGND VGND VPWR VPWR hold814/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _3953_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6322_ _6643_/Q _6319_/Y _6321_/X _6317_/Y VGND VGND VPWR VPWR _6346_/S sky130_fd_sc_hd__a211o_4
Xhold825 _4120_/X VGND VGND VPWR VPWR _6533_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3534_ _6741_/Q _5148_/A hold67/A _6469_/Q _3531_/X VGND VGND VPWR VPWR _3538_/C
+ sky130_fd_sc_hd__a221o_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_2
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold836 _7152_/Q VGND VGND VPWR VPWR hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _4016_/X VGND VGND VPWR VPWR _6456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _7191_/A VGND VGND VPWR VPWR hold858/X sky130_fd_sc_hd__dlygate4sd3_1
X_6253_ _7128_/Q _6252_/X _6303_/S VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__mux2_1
Xhold869 _5331_/X VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3465_ _6863_/Q _5292_/A _5154_/A _6747_/Q _3464_/X VGND VGND VPWR VPWR _3467_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5204_ hold257/X _5534_/A1 _5210_/S VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__mux2_1
X_6184_ _6685_/Q _5961_/X _6182_/X _6183_/X VGND VGND VPWR VPWR _6189_/A sky130_fd_sc_hd__a211o_1
X_3396_ _6441_/Q _3372_/Y _3393_/X _3395_/X VGND VGND VPWR VPWR _3396_/X sky130_fd_sc_hd__a211o_1
XFILLER_97_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1503 _7130_/Q VGND VGND VPWR VPWR _6279_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5135_ _5135_/A _5135_/B _5135_/C VGND VGND VPWR VPWR _5135_/Y sky130_fd_sc_hd__nand3_2
Xhold1514 _7147_/Q VGND VGND VPWR VPWR _6343_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 hold58/A VGND VGND VPWR VPWR _3257_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1536 hold40/A VGND VGND VPWR VPWR _3256_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 _6489_/Q VGND VGND VPWR VPWR _3912_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1558 hold32/A VGND VGND VPWR VPWR _3849_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5066_ _5066_/A _5112_/C _5106_/C _5066_/D VGND VGND VPWR VPWR _5066_/X sky130_fd_sc_hd__and4_1
XFILLER_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1569 _7167_/Q VGND VGND VPWR VPWR _3253_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4017_ hold960/X _6355_/A1 _4019_/S VGND VGND VPWR VPWR _4017_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5968_ _5968_/A _5969_/C _5979_/C VGND VGND VPWR VPWR _5976_/D sky130_fd_sc_hd__and3_4
XFILLER_52_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4919_ _5023_/A _5023_/B _5023_/C _4919_/D VGND VGND VPWR VPWR _4919_/X sky130_fd_sc_hd__and4_1
XFILLER_21_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5899_ _6658_/Q _5899_/B VGND VGND VPWR VPWR _5899_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3250_ _3250_/A _3250_/B VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__xnor2_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3181_ _4566_/A VGND VGND VPWR VPWR _4702_/B sky130_fd_sc_hd__clkinv_2
XFILLER_79_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6940_ _7063_/CLK _6940_/D fanout463/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ _7078_/CLK _6871_/D fanout482/X VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5822_ _3183_/Y _5899_/B _5651_/B VGND VGND VPWR VPWR _5822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5753_ _7006_/Q _5625_/X _5632_/X _6942_/Q _5737_/X VGND VGND VPWR VPWR _5754_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4704_ _4460_/A _4626_/B _4616_/Y _4703_/Y VGND VGND VPWR VPWR _4704_/X sky130_fd_sc_hd__o31a_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5684_ _6971_/Q _5634_/X _5652_/B _6915_/Q _5651_/Y VGND VGND VPWR VPWR _5684_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_187_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4635_ _4716_/A _4635_/B _4661_/B VGND VGND VPWR VPWR _4689_/B sky130_fd_sc_hd__nand3_4
XFILLER_147_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 _7056_/Q VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 _4089_/X VGND VGND VPWR VPWR _6511_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _4566_/A _4566_/B VGND VGND VPWR VPWR _4664_/B sky130_fd_sc_hd__xnor2_2
Xhold622 hold622/A VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _5273_/X VGND VGND VPWR VPWR _6841_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold644 _7080_/Q VGND VGND VPWR VPWR hold644/X sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ _6636_/Q _6641_/Q _6635_/Q _3910_/B VGND VGND VPWR VPWR _6305_/Y sky130_fd_sc_hd__o31ai_1
X_3517_ hold74/X _3573_/B VGND VGND VPWR VPWR _4038_/A sky130_fd_sc_hd__nor2_4
XFILLER_89_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap363 _4118_/B VGND VGND VPWR VPWR _4083_/S sky130_fd_sc_hd__buf_8
Xhold655 _5372_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap374 _3571_/A VGND VGND VPWR VPWR hold125/A sky130_fd_sc_hd__buf_12
X_4497_ _4579_/B _5042_/B VGND VGND VPWR VPWR _4843_/B sky130_fd_sc_hd__and2_1
Xhold666 hold666/A VGND VGND VPWR VPWR hold666/X sky130_fd_sc_hd__buf_8
Xmax_cap385 _5655_/X VGND VGND VPWR VPWR _5905_/A2 sky130_fd_sc_hd__buf_6
Xhold677 _6969_/Q VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 _5228_/X VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6236_ _6632_/Q _5946_/X _5955_/X _6552_/Q VGND VGND VPWR VPWR _6236_/X sky130_fd_sc_hd__a22o_1
Xhold699 _5433_/X VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3448_ _3447_/Y _3488_/A1 _3829_/A VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__mux2_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6913_/Q _5973_/A _5948_/X _6953_/Q _6166_/X VGND VGND VPWR VPWR _6167_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 _5149_/X VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3379_ _3379_/A hold75/X VGND VGND VPWR VPWR _3999_/A sky130_fd_sc_hd__nor2_8
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _6418_/Q VGND VGND VPWR VPWR _3966_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 hold1322/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5118_ _5118_/A _5118_/B _5118_/C VGND VGND VPWR VPWR _5118_/X sky130_fd_sc_hd__and3_1
Xhold1333 hold1419/X VGND VGND VPWR VPWR hold1333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1344 hold1344/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
Xclkbuf_0__1177_ _3582_/Y VGND VGND VPWR VPWR clkbuf_0__1177_/X sky130_fd_sc_hd__clkbuf_16
X_6098_ _6814_/Q _5971_/B _5949_/X _6934_/Q _6097_/X VGND VGND VPWR VPWR _6099_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1355 _6315_/A1 VGND VGND VPWR VPWR hold1355/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1366 hold1366/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1377 _6312_/A1 VGND VGND VPWR VPWR hold1377/X sky130_fd_sc_hd__dlygate4sd3_1
X_5049_ _4672_/B _4496_/Y _4542_/A VGND VGND VPWR VPWR _5049_/X sky130_fd_sc_hd__a21o_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1388 _7084_/Q VGND VGND VPWR VPWR _5547_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _3973_/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4420_ _4753_/A _4600_/B VGND VGND VPWR VPWR _4947_/A sky130_fd_sc_hd__nand2b_2
XFILLER_144_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4351_ _4352_/B _4351_/B VGND VGND VPWR VPWR _4379_/B sky130_fd_sc_hd__nand2_1
X_3302_ hold72/X _3355_/B _3347_/A VGND VGND VPWR VPWR _3555_/A sky130_fd_sc_hd__nand3b_4
X_7070_ _7070_/CLK _7070_/D fanout482/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout409 _5518_/A1 VGND VGND VPWR VPWR _5509_/A1 sky130_fd_sc_hd__buf_6
X_4282_ _4282_/A0 _5492_/A1 _4285_/S VGND VGND VPWR VPWR _4282_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6021_ _7027_/Q _5944_/X _5975_/A _6843_/Q _6020_/X VGND VGND VPWR VPWR _6024_/C
+ sky130_fd_sc_hd__a221o_1
X_3233_ _3233_/A0 _3251_/A _3233_/S VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_66_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3164_ _7159_/Q VGND VGND VPWR VPWR _3164_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6923_ _7006_/CLK _6923_/D fanout458/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_81_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6854_ _7081_/CLK _6854_/D fanout478/X VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfrtp_4
X_5805_ _6953_/Q _5637_/X _5645_/X _7033_/Q VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__a22o_1
X_6785_ _7076_/CLK _6785_/D fanout481/X VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtp_1
X_3997_ _3997_/A0 hold99/X _3998_/S VGND VGND VPWR VPWR _3997_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5736_ _5736_/A1 _6279_/S _5734_/X _5735_/X VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__o22a_1
XFILLER_148_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5667_ _5664_/A _5667_/B _5667_/C VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__and3b_4
XFILLER_135_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4618_ _4653_/B _4635_/B VGND VGND VPWR VPWR _4618_/Y sky130_fd_sc_hd__nand2_2
X_5598_ _5598_/A _5602_/A VGND VGND VPWR VPWR _5598_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold430 _5343_/X VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _4549_/A _4549_/B VGND VGND VPWR VPWR _4553_/B sky130_fd_sc_hd__nand2_1
Xhold441 _6765_/Q VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold452 _5234_/X VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _6563_/Q VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _5360_/X VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold485 _6910_/Q VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold496 _4218_/X VGND VGND VPWR VPWR _6617_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6219_ _6646_/Q _5976_/C _5971_/D _6566_/Q VGND VGND VPWR VPWR _6219_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7199_ _7199_/A VGND VGND VPWR VPWR _7199_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1130 _4160_/X VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1141 _6767_/Q VGND VGND VPWR VPWR _5189_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1152 _5302_/X VGND VGND VPWR VPWR _6866_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1163 _6465_/Q VGND VGND VPWR VPWR _4027_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 _4146_/X VGND VGND VPWR VPWR _6555_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 _6882_/Q VGND VGND VPWR VPWR _5320_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1196 _5284_/X VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3920_ _3186_/Y input92/X _3921_/S VGND VGND VPWR VPWR _3920_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3851_ _3850_/Y hold70/A _3851_/C VGND VGND VPWR VPWR _3853_/A sky130_fd_sc_hd__and3b_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6570_ _7137_/CLK _6570_/D VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfxtp_1
X_3782_ _3782_/A _3782_/B _3782_/C _3782_/D VGND VGND VPWR VPWR _3794_/B sky130_fd_sc_hd__nor4_1
XFILLER_164_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5521_ hold319/X _5521_/A1 hold87/X VGND VGND VPWR VPWR _5521_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5452_ hold112/X hold99/X _5453_/S VGND VGND VPWR VPWR _5452_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4403_ _4633_/B _4389_/Y _4653_/B _4563_/D VGND VGND VPWR VPWR _4448_/B sky130_fd_sc_hd__a22o_1
XFILLER_145_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5383_ _5383_/A0 hold666/X _5390_/S VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__mux2_1
X_7122_ _7131_/CLK _7122_/D fanout456/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4334_ _4702_/A _4334_/B _4334_/C VGND VGND VPWR VPWR _4434_/B sky130_fd_sc_hd__nor3_2
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7053_ _7053_/CLK _7053_/D fanout459/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4265_ hold471/X _5544_/A1 _4267_/S VGND VGND VPWR VPWR _4265_/X sky130_fd_sc_hd__mux2_1
X_6004_ _7040_/Q _5971_/C _5976_/D _6875_/Q VGND VGND VPWR VPWR _6004_/X sky130_fd_sc_hd__a22o_1
X_3216_ _6845_/Q VGND VGND VPWR VPWR _3216_/Y sky130_fd_sc_hd__inv_2
X_4196_ _4196_/A _4322_/B VGND VGND VPWR VPWR _4201_/S sky130_fd_sc_hd__and2_2
XFILLER_67_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6906_ _6908_/CLK _6906_/D fanout463/X VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6837_ _6865_/CLK _6837_/D fanout464/X VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_145_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6768_ _6769_/CLK _6768_/D fanout469/X VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5719_ _7005_/Q _5625_/X _5661_/X _6877_/Q VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6699_ _6709_/CLK _6699_/D _6360_/A VGND VGND VPWR VPWR _6699_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold260 _5447_/X VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _6752_/Q VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _4147_/X VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold293 _6851_/Q VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _7157_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _7199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 _6739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _5902_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 hold60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _5166_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _5975_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _5229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4050_ _6396_/B _5193_/A VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__and2b_2
XFILLER_49_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4952_ _4542_/B _5043_/B VGND VGND VPWR VPWR _5057_/B sky130_fd_sc_hd__nand2b_1
X_3903_ _4337_/C _4337_/D _4336_/A _4336_/B VGND VGND VPWR VPWR _3907_/C sky130_fd_sc_hd__nor4_1
X_4883_ _5023_/C _4882_/X _5023_/A VGND VGND VPWR VPWR _4884_/D sky130_fd_sc_hd__a21bo_1
XFILLER_20_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3834_ _3867_/B _3832_/B _3836_/A _3834_/B2 VGND VGND VPWR VPWR _6417_/D sky130_fd_sc_hd__o22a_1
X_6622_ _6629_/CLK _6622_/D _6390_/A VGND VGND VPWR VPWR _6622_/Q sky130_fd_sc_hd__dfrtp_2
X_6553_ _6659_/CLK _6553_/D fanout469/X VGND VGND VPWR VPWR _6553_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3765_ _7018_/Q hold29/A _5409_/A _6962_/Q VGND VGND VPWR VPWR _3765_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5504_ hold311/X _5540_/A1 hold77/X VGND VGND VPWR VPWR _5504_/X sky130_fd_sc_hd__mux2_1
X_6484_ _6707_/CLK _6484_/D fanout450/X VGND VGND VPWR VPWR _6484_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_106_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3696_ _6621_/Q _4220_/A _4244_/A _6647_/Q VGND VGND VPWR VPWR _3696_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpad_flashh_clk_buff_inst _3945_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_145_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5435_ hold143/X hold22/X _5435_/S VGND VGND VPWR VPWR _5435_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput310 _3953_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
Xoutput321 hold1351/X VGND VGND VPWR VPWR hold1352/A sky130_fd_sc_hd__buf_12
Xoutput332 hold1357/X VGND VGND VPWR VPWR hold1358/A sky130_fd_sc_hd__buf_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 hold1337/X VGND VGND VPWR VPWR hold1338/A sky130_fd_sc_hd__buf_12
X_5366_ hold245/X _5465_/A1 _5372_/S VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4317_ _4317_/A0 _5491_/A1 _4321_/S VGND VGND VPWR VPWR _4317_/X sky130_fd_sc_hd__mux2_1
X_7105_ _7113_/CLK _7105_/D fanout460/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_1
X_5297_ hold180/X _5519_/A1 _5300_/S VGND VGND VPWR VPWR _5297_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7036_ _7036_/CLK _7036_/D fanout455/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_59_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4248_ hold491/X _5518_/A1 _4249_/S VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4179_ _3828_/Y _4179_/A1 _4186_/S VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_csclk clkbuf_opt_3_0_csclk/X VGND VGND VPWR VPWR _6967_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_csclk _6447_/CLK VGND VGND VPWR VPWR _6539_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3550_ _3562_/A _3692_/A VGND VGND VPWR VPWR _4196_/A sky130_fd_sc_hd__nor2_4
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3481_ _6855_/Q _5283_/A _5202_/B input40/X _3480_/X VGND VGND VPWR VPWR _3484_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5220_ _5220_/A hold17/X VGND VGND VPWR VPWR _5227_/S sky130_fd_sc_hd__and2_4
XFILLER_115_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5151_ hold995/X _6355_/A1 _5153_/S VGND VGND VPWR VPWR _5151_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4102_ _4102_/A _5541_/B VGND VGND VPWR VPWR _4108_/S sky130_fd_sc_hd__and2_4
X_5082_ _5088_/A _5114_/A _5082_/C VGND VGND VPWR VPWR _5087_/B sky130_fd_sc_hd__and3_1
XFILLER_84_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4033_ _4033_/A0 _5491_/A1 _4037_/S VGND VGND VPWR VPWR _4033_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5984_ _6794_/Q _5965_/X _5971_/D _6826_/Q VGND VGND VPWR VPWR _5984_/X sky130_fd_sc_hd__a22o_1
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4935_ _4948_/C _4562_/Y _4620_/Y _4638_/Y _4768_/B VGND VGND VPWR VPWR _5076_/A
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_3_7_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 _5265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _4220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _4948_/C _4496_/Y _4639_/Y _4689_/A VGND VGND VPWR VPWR _4870_/A sky130_fd_sc_hd__o22a_1
XFILLER_177_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_33 _3688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ _6746_/CLK _6605_/D fanout447/X VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_44 _5471_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_55 _5958_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3817_ _3817_/A _3817_/B _3817_/C _3817_/D VGND VGND VPWR VPWR _3827_/C sky130_fd_sc_hd__nor4_1
XANTENNA_66 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4797_ _4673_/A _4611_/Y _4476_/Y VGND VGND VPWR VPWR _5008_/A sky130_fd_sc_hd__a21o_1
XANTENNA_77 _6276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _7040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 _7157_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _6539_/CLK _6536_/D fanout461/X VGND VGND VPWR VPWR _6536_/Q sky130_fd_sc_hd__dfrtp_1
X_3748_ _6661_/Q _4262_/A _4127_/A _6541_/Q _3747_/X VGND VGND VPWR VPWR _3751_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6467_ _6654_/CLK _6467_/D _6401_/A VGND VGND VPWR VPWR _6467_/Q sky130_fd_sc_hd__dfstp_2
X_3679_ _3679_/A _3679_/B _3679_/C _3679_/D VGND VGND VPWR VPWR _3699_/B sky130_fd_sc_hd__nor4_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5418_ _5418_/A _5541_/B VGND VGND VPWR VPWR _5426_/S sky130_fd_sc_hd__and2_4
X_6398_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__and2_1
Xoutput173 _3959_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
XFILLER_121_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5349_ hold856/X _5484_/A1 _5354_/S VGND VGND VPWR VPWR _5349_/X sky130_fd_sc_hd__mux2_1
Xoutput184 _3205_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput195 _3195_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_87_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7019_ _7085_/CLK _7019_/D fanout479/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4689_/A _4616_/Y _4626_/Y _4483_/Y _4719_/X VGND VGND VPWR VPWR _4721_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_187_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4651_ _4441_/A _4484_/Y _4609_/Y _4619_/Y _4650_/Y VGND VGND VPWR VPWR _4660_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_2
X_3602_ _6917_/Q _5355_/A _5247_/A _6821_/Q _3601_/X VGND VGND VPWR VPWR _3604_/C
+ sky130_fd_sc_hd__a221o_1
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
X_4582_ _4992_/A _4582_/B VGND VGND VPWR VPWR _4582_/Y sky130_fd_sc_hd__nor2_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_2
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_1
Xhold804 _6435_/Q VGND VGND VPWR VPWR hold804/X sky130_fd_sc_hd__dlygate4sd3_1
X_3533_ hold74/A hold66/X VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__nor2_8
X_6321_ _6642_/Q _6318_/Y _6320_/Y _6644_/Q _4229_/X VGND VGND VPWR VPWR _6321_/X
+ sky130_fd_sc_hd__a221o_1
Xhold815 _4318_/X VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _3947_/B sky130_fd_sc_hd__clkbuf_4
Xhold826 _6714_/Q VGND VGND VPWR VPWR hold826/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold837 _6354_/X VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold848 _6481_/Q VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6252_ _6240_/Y _6251_/X _6542_/Q _6226_/B VGND VGND VPWR VPWR _6252_/X sky130_fd_sc_hd__o2bb2a_1
X_3464_ _6911_/Q _5346_/A _5391_/A _6951_/Q VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold859 _5196_/X VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5203_ _5203_/A0 _5473_/A1 _5210_/S VGND VGND VPWR VPWR _5203_/X sky130_fd_sc_hd__mux2_1
X_6183_ _6475_/Q _5940_/X _5967_/X _6604_/Q _6181_/X VGND VGND VPWR VPWR _6183_/X
+ sky130_fd_sc_hd__a221o_1
X_3395_ _6865_/Q _5292_/A _5532_/A _7078_/Q _3394_/X VGND VGND VPWR VPWR _3395_/X
+ sky130_fd_sc_hd__a221o_4
X_5134_ _5134_/A _5134_/B _5134_/C VGND VGND VPWR VPWR _5135_/C sky130_fd_sc_hd__and3_1
XFILLER_97_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1504 _7124_/Q VGND VGND VPWR VPWR _6129_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1515 _7145_/Q VGND VGND VPWR VPWR _6337_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _3257_/X VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1537 _7112_/Q VGND VGND VPWR VPWR _5820_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5065_ _4483_/Y _4625_/B _4650_/Y _4716_/Y _5018_/A VGND VGND VPWR VPWR _5066_/D
+ sky130_fd_sc_hd__o2111a_1
Xhold1548 _3182_/Y VGND VGND VPWR VPWR _3869_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 _6635_/Q VGND VGND VPWR VPWR _3909_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4016_ hold846/X _6354_/A1 _4019_/S VGND VGND VPWR VPWR _4016_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5967_ _5969_/C _5981_/C _5979_/C VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__and3_4
XFILLER_52_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4918_ _4918_/A _4918_/B VGND VGND VPWR VPWR _4919_/D sky130_fd_sc_hd__nand2_1
X_5898_ _6563_/Q _5631_/X _5637_/X _6698_/Q _5897_/X VGND VGND VPWR VPWR _5906_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4849_ _4483_/Y _4846_/B _4535_/A VGND VGND VPWR VPWR _5073_/A sky130_fd_sc_hd__o21a_1
XFILLER_193_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6519_ _6668_/CLK _6519_/D _6400_/A VGND VGND VPWR VPWR _6519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3180_ _7101_/Q VGND VGND VPWR VPWR _5600_/A sky130_fd_sc_hd__inv_2
XFILLER_140_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6870_ _7051_/CLK _6870_/D fanout476/X VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5821_ _5821_/A1 _6279_/S _5819_/X _5820_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__o22a_1
XFILLER_62_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5752_ _7014_/Q _5630_/X _5645_/X _7030_/Q _5751_/X VGND VGND VPWR VPWR _5754_/B
+ sky130_fd_sc_hd__a221o_1
X_4703_ _4782_/A _4703_/B VGND VGND VPWR VPWR _4703_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5683_ _6923_/Q _5664_/X _5667_/X _6811_/Q _5682_/X VGND VGND VPWR VPWR _5690_/A
+ sky130_fd_sc_hd__a221o_1
X_4634_ _4716_/A _4635_/B _4661_/B VGND VGND VPWR VPWR _4753_/C sky130_fd_sc_hd__and3_1
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold601 _5516_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _4563_/D _4653_/B _4595_/A VGND VGND VPWR VPWR _4565_/X sky130_fd_sc_hd__a21o_1
Xhold612 _6672_/Q VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold623 _4111_/X VGND VGND VPWR VPWR _6525_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _6304_/A0 _6303_/X _6304_/S VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__mux2_1
Xhold634 _6971_/Q VGND VGND VPWR VPWR hold634/X sky130_fd_sc_hd__dlygate4sd3_1
X_3516_ _3573_/A _3814_/B VGND VGND VPWR VPWR _4032_/A sky130_fd_sc_hd__nor2_4
Xhold645 _5543_/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 _7015_/Q VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4496_ _4607_/A _4496_/B VGND VGND VPWR VPWR _4496_/Y sky130_fd_sc_hd__nand2_8
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold667 hold667/A VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__buf_8
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap386 _5646_/X VGND VGND VPWR VPWR _5814_/B1 sky130_fd_sc_hd__buf_8
Xhold678 _5417_/X VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 _6423_/Q VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlygate4sd3_1
X_6235_ _6687_/Q _5961_/X _6232_/X _6234_/X VGND VGND VPWR VPWR _6240_/A sky130_fd_sc_hd__a211o_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3447_ _3447_/A _3447_/B _3447_/C VGND VGND VPWR VPWR _3447_/Y sky130_fd_sc_hd__nand3_4
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6905_/Q _5976_/C _5971_/D _6833_/Q VGND VGND VPWR VPWR _6166_/X sky130_fd_sc_hd__a22o_1
X_3378_ _3586_/A hold75/X VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__nor2_8
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 _6434_/Q VGND VGND VPWR VPWR _3991_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 _3966_/X VGND VGND VPWR VPWR _6418_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1323 hold1416/X VGND VGND VPWR VPWR hold1323/X sky130_fd_sc_hd__dlygate4sd3_1
X_5117_ _4482_/B _4695_/Y _4858_/X _4823_/A VGND VGND VPWR VPWR _5118_/C sky130_fd_sc_hd__o211a_1
Xhold1334 hold1334/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6097_ hold79/A _5601_/X _5959_/X _6966_/Q VGND VGND VPWR VPWR _6097_/X sky130_fd_sc_hd__a22o_1
Xhold1345 hold1428/X VGND VGND VPWR VPWR hold1345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1356 hold1356/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xhold1367 _4190_/A1 VGND VGND VPWR VPWR hold1367/X sky130_fd_sc_hd__dlygate4sd3_1
X_5048_ _4672_/B _4496_/Y _4413_/Y VGND VGND VPWR VPWR _5057_/C sky130_fd_sc_hd__a21o_1
Xhold1378 hold1378/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
Xhold1389 _6788_/Q VGND VGND VPWR VPWR _5214_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6999_ _6999_/CLK _6999_/D fanout465/X VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4350_ _4661_/A _4357_/B _4631_/D VGND VGND VPWR VPWR _4351_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3301_ _3586_/A _3562_/A VGND VGND VPWR VPWR _5283_/A sky130_fd_sc_hd__nor2_8
X_4281_ _4281_/A0 _6353_/A1 _4285_/S VGND VGND VPWR VPWR _4281_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3232_ _3867_/A _3829_/A VGND VGND VPWR VPWR _3233_/S sky130_fd_sc_hd__nor2_1
X_6020_ _7019_/Q _5937_/X _5975_/D _6883_/Q VGND VGND VPWR VPWR _6020_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6922_ _6926_/CLK _6922_/D fanout458/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_82_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6853_ _6951_/CLK _6853_/D fanout474/X VGND VGND VPWR VPWR _6853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5804_ _6849_/Q _5616_/X _5655_/X _6801_/Q _5803_/X VGND VGND VPWR VPWR _5804_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6784_ _7076_/CLK _6784_/D fanout481/X VGND VGND VPWR VPWR _6784_/Q sky130_fd_sc_hd__dfrtp_1
X_3996_ hold574/X _5469_/A1 _3998_/S VGND VGND VPWR VPWR _3996_/X sky130_fd_sc_hd__mux2_1
X_5735_ _6507_/Q _5735_/A2 _6103_/B1 VGND VGND VPWR VPWR _5735_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5666_ _5664_/A _5666_/B _5666_/C VGND VGND VPWR VPWR _5666_/X sky130_fd_sc_hd__and3b_4
XFILLER_136_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4617_ _4627_/A _4846_/B VGND VGND VPWR VPWR _4646_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5597_ _5600_/A _5597_/B VGND VGND VPWR VPWR _5602_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold420 _5535_/X VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _6712_/Q VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlygate4sd3_1
X_4548_ _4500_/A _4947_/C _4464_/Y _4902_/A _5114_/A VGND VGND VPWR VPWR _4548_/X
+ sky130_fd_sc_hd__o221a_1
Xhold442 _5187_/X VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _6557_/Q VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold464 _4155_/X VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _6870_/Q VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _5351_/X VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4479_ _4653_/C VGND VGND VPWR VPWR _4479_/Y sky130_fd_sc_hd__inv_2
Xhold497 _7001_/Q VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__dlygate4sd3_1
X_6218_ _6218_/A _6218_/B _6218_/C VGND VGND VPWR VPWR _6226_/C sky130_fd_sc_hd__nor3_1
X_7198_ _7198_/A VGND VGND VPWR VPWR _7198_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1120 _5493_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6149_ _6816_/Q _5971_/B _5949_/X _6936_/Q _6148_/X VGND VGND VPWR VPWR _6150_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1131 _6580_/Q VGND VGND VPWR VPWR _4175_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1142 _5189_/X VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1153 _6826_/Q VGND VGND VPWR VPWR _5257_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1164 _4027_/X VGND VGND VPWR VPWR _6465_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 hold1590/X VGND VGND VPWR VPWR _4053_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1186 _5320_/X VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1197 _6888_/Q VGND VGND VPWR VPWR _5326_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3850_ _6488_/Q _3854_/S VGND VGND VPWR VPWR _3850_/Y sky130_fd_sc_hd__nor2_1
X_3781_ _6946_/Q _3781_/A2 _5523_/A _7063_/Q _3780_/X VGND VGND VPWR VPWR _3782_/D
+ sky130_fd_sc_hd__a221o_1
X_5520_ _5520_/A0 hold42/X hold87/A VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__mux2_1
XFILLER_9_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5451_ hold726/X _5469_/A1 _5453_/S VGND VGND VPWR VPWR _5451_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4402_ _4661_/A _4653_/B VGND VGND VPWR VPWR _4627_/B sky130_fd_sc_hd__nand2_4
X_5382_ _5382_/A hold17/X VGND VGND VPWR VPWR _5390_/S sky130_fd_sc_hd__and2_4
X_7121_ _7126_/CLK _7121_/D fanout456/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_1
X_4333_ hold902/X _6357_/A1 _4333_/S VGND VGND VPWR VPWR _4333_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7052_ _7086_/CLK _7052_/D fanout482/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_1
X_4264_ hold267/X _5534_/A1 _4267_/S VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6003_ _6001_/X _6002_/Y _6003_/B1 _6103_/B1 VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__a2bb2o_1
X_3215_ _6853_/Q VGND VGND VPWR VPWR _3215_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4195_ _3410_/Y _4195_/A1 _4195_/S VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6905_ _7076_/CLK _6905_/D fanout481/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6836_ _7065_/CLK _6836_/D fanout463/X VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6767_ _6890_/CLK _6767_/D fanout470/X VGND VGND VPWR VPWR _6767_/Q sky130_fd_sc_hd__dfrtp_1
X_3979_ hold20/X hold172/X _6624_/Q VGND VGND VPWR VPWR _3979_/X sky130_fd_sc_hd__mux2_1
X_5718_ _6821_/Q _5818_/A2 _5642_/X _6965_/Q VGND VGND VPWR VPWR _5718_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6698_ _6735_/CLK _6698_/D fanout445/X VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5649_ _5658_/B _5667_/C VGND VGND VPWR VPWR _5652_/B sky130_fd_sc_hd__and2_4
XFILLER_151_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold250 _5402_/X VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold261 _7072_/Q VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _5168_/X VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _6859_/Q VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _5285_/X VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _7157_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _7199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 _6428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _5513_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 hold99/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _3700_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_178 _6301_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_189 _6423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_174_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_2
XFILLER_49_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4951_ _5114_/A _4951_/B VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__and2_1
XFILLER_17_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3902_ _4337_/A _4337_/B VGND VGND VPWR VPWR _3907_/B sky130_fd_sc_hd__nor2_1
X_4882_ _5023_/D _4882_/B _4882_/C VGND VGND VPWR VPWR _4882_/X sky130_fd_sc_hd__and3_1
X_6621_ _6629_/CLK _6621_/D _6390_/A VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_189_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3833_ _6416_/Q _3838_/A VGND VGND VPWR VPWR _3836_/A sky130_fd_sc_hd__and2_1
X_6552_ _6632_/CLK _6552_/D fanout454/X VGND VGND VPWR VPWR _6552_/Q sky130_fd_sc_hd__dfstp_1
X_3764_ _3763_/X _3764_/A1 _3829_/B VGND VGND VPWR VPWR _3764_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5503_ hold910/X _5548_/A1 hold77/X VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6483_ _6704_/CLK _6483_/D fanout450/X VGND VGND VPWR VPWR _6483_/Q sky130_fd_sc_hd__dfrtp_1
X_3695_ _3251_/A _4083_/S _3358_/Y input13/X _3694_/X VGND VGND VPWR VPWR _3698_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5434_ hold521/X hold99/X _5435_/S VGND VGND VPWR VPWR _5434_/X sky130_fd_sc_hd__mux2_1
Xoutput300 _6754_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
Xoutput311 _7199_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
Xoutput322 hold1347/X VGND VGND VPWR VPWR hold1348/A sky130_fd_sc_hd__buf_12
XFILLER_133_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput333 hold1349/X VGND VGND VPWR VPWR hold1350/A sky130_fd_sc_hd__buf_12
Xoutput344 hold1329/X VGND VGND VPWR VPWR hold1330/A sky130_fd_sc_hd__buf_12
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5365_ _5365_/A0 _5524_/A1 _5372_/S VGND VGND VPWR VPWR _5365_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7104_ _7131_/CLK _7104_/D fanout460/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_3_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR _7001_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4316_ _4316_/A _6352_/B VGND VGND VPWR VPWR _4321_/S sky130_fd_sc_hd__and2_2
X_5296_ hold916/X _5509_/A1 _5300_/S VGND VGND VPWR VPWR _5296_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7035_ _7037_/CLK _7035_/D fanout455/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4247_ hold638/X _5544_/A1 _4249_/S VGND VGND VPWR VPWR _4247_/X sky130_fd_sc_hd__mux2_1
X_4178_ _6637_/Q _6307_/B VGND VGND VPWR VPWR _4186_/S sky130_fd_sc_hd__nand2_4
XFILLER_28_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6819_ _6884_/CLK _6819_/D fanout475/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3480_ _7060_/Q hold86/A _5505_/A _7052_/Q VGND VGND VPWR VPWR _3480_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ hold890/X _6354_/A1 _5153_/S VGND VGND VPWR VPWR _5150_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4101_ hold720/X _4100_/X _4101_/S VGND VGND VPWR VPWR _4101_/X sky130_fd_sc_hd__mux2_1
X_5081_ _4902_/A _4902_/B _4689_/A _4464_/Y VGND VGND VPWR VPWR _5082_/C sky130_fd_sc_hd__a31o_1
X_4032_ _4032_/A _5490_/B VGND VGND VPWR VPWR _4037_/S sky130_fd_sc_hd__and2_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5983_ _6842_/Q _5975_/A _5959_/X _6962_/Q VGND VGND VPWR VPWR _5983_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4934_ _4542_/D _4562_/Y _4620_/Y _4652_/Y _4770_/B VGND VGND VPWR VPWR _5003_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4865_ _4652_/Y _4700_/Y _4518_/C VGND VGND VPWR VPWR _5034_/A sky130_fd_sc_hd__o21a_1
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_12 _5265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _4220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6604_ _6746_/CLK _6604_/D fanout447/X VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_34 _3742_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3816_ _6826_/Q _5256_/A _4244_/A _6645_/Q _3815_/X VGND VGND VPWR VPWR _3817_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 _5627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_56 _5965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _4796_/A _5064_/A _4796_/C _4796_/D VGND VGND VPWR VPWR _4804_/A sky130_fd_sc_hd__and4_1
XANTENNA_67 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _6542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6925_/CLK _6535_/D fanout460/X VGND VGND VPWR VPWR _6535_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_89 _6664_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3747_ _7072_/Q _5532_/A _5490_/A _7035_/Q VGND VGND VPWR VPWR _3747_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6466_ _6653_/CLK _6466_/D _6401_/A VGND VGND VPWR VPWR _6466_/Q sky130_fd_sc_hd__dfrtp_4
X_3678_ _6980_/Q _5427_/A _4238_/A _6632_/Q _3677_/X VGND VGND VPWR VPWR _3679_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5417_ hold677/X _5540_/A1 _5417_/S VGND VGND VPWR VPWR _5417_/X sky130_fd_sc_hd__mux2_1
X_6397_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6397_/X sky130_fd_sc_hd__and2_1
Xoutput174 _3960_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
XFILLER_102_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5348_ hold572/X _5543_/A1 _5354_/S VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__mux2_1
Xoutput185 _3204_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3194_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5279_ hold467/X _5528_/A1 _5282_/S VGND VGND VPWR VPWR _5279_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7018_ _7051_/CLK _7018_/D fanout476/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout390 _4372_/X VGND VGND VPWR VPWR _4716_/A sky130_fd_sc_hd__buf_12
XFILLER_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4650_ _4650_/A _5043_/A VGND VGND VPWR VPWR _4650_/Y sky130_fd_sc_hd__nand2_1
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
X_3601_ _7050_/Q _5505_/A _5541_/A _7082_/Q VGND VGND VPWR VPWR _3601_/X sky130_fd_sc_hd__a22o_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4581_ _4810_/A _4581_/B VGND VGND VPWR VPWR _4581_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_1
X_6320_ _6320_/A _6320_/B VGND VGND VPWR VPWR _6320_/Y sky130_fd_sc_hd__nand2_1
Xhold805 _3992_/X VGND VGND VPWR VPWR _6435_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3532_ hold85/X _3714_/B VGND VGND VPWR VPWR _5148_/A sky130_fd_sc_hd__nor2_8
XFILLER_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7199_/A sky130_fd_sc_hd__clkbuf_4
Xinput76 qspi_enabled VGND VGND VPWR VPWR _3921_/S sky130_fd_sc_hd__clkbuf_8
Xhold816 _7083_/Q VGND VGND VPWR VPWR hold816/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7198_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold827 _4327_/X VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__clkbuf_2
Xhold838 _6694_/Q VGND VGND VPWR VPWR hold838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 _4046_/X VGND VGND VPWR VPWR _6481_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _6243_/X _6251_/B _6301_/C VGND VGND VPWR VPWR _6251_/X sky130_fd_sc_hd__and3b_1
XFILLER_143_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3463_ _6431_/Q _3981_/A _3381_/Y input31/X _3462_/X VGND VGND VPWR VPWR _3467_/B
+ sky130_fd_sc_hd__a221o_2
X_5202_ _6396_/B _5202_/B _5505_/B VGND VGND VPWR VPWR _5210_/S sky130_fd_sc_hd__and3b_4
X_6182_ _7151_/Q _5958_/X _5978_/X _6480_/Q VGND VGND VPWR VPWR _6182_/X sky130_fd_sc_hd__a22o_1
X_3394_ input42/X _5202_/B _3999_/A _6449_/Q VGND VGND VPWR VPWR _3394_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5133_ _4628_/Y _4970_/Y _5010_/Y _4631_/Y _4796_/D VGND VGND VPWR VPWR _5134_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1505 _6588_/Q VGND VGND VPWR VPWR _4184_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 _7105_/Q VGND VGND VPWR VPWR _5609_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 _7141_/Q VGND VGND VPWR VPWR _6325_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 hold97/A VGND VGND VPWR VPWR _3255_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5064_ _5064_/A _5064_/B _5064_/C VGND VGND VPWR VPWR _5106_/C sky130_fd_sc_hd__and3_1
Xhold1549 _7099_/Q VGND VGND VPWR VPWR _5592_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4015_ _4015_/A0 _6353_/A1 _4019_/S VGND VGND VPWR VPWR _4015_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5966_ _5966_/A _5981_/B _5981_/C VGND VGND VPWR VPWR _5971_/C sky130_fd_sc_hd__and3_4
XFILLER_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4917_ _4359_/Y _4887_/A _4384_/A _4887_/B _4872_/B VGND VGND VPWR VPWR _5033_/A
+ sky130_fd_sc_hd__o41a_1
X_5897_ _6648_/Q _5621_/X _5913_/B1 _6553_/Q VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4848_ _4469_/A _4689_/A _4490_/B VGND VGND VPWR VPWR _5029_/A sky130_fd_sc_hd__a21o_1
XFILLER_148_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4779_ _4902_/B _4611_/Y _4500_/A VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__a21o_1
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6518_ _6755_/CLK _6518_/D _6360_/A VGND VGND VPWR VPWR _6518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6449_ _7070_/CLK _6449_/D fanout473/X VGND VGND VPWR VPWR _6449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_csclk _6888_/CLK VGND VGND VPWR VPWR _6951_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5820_ _6507_/Q _5820_/A2 _5611_/Y VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5751_ _6950_/Q _5637_/X _5660_/X _6806_/Q VGND VGND VPWR VPWR _5751_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4702_ _4702_/A _4702_/B _4702_/C _4965_/B VGND VGND VPWR VPWR _4702_/Y sky130_fd_sc_hd__nand4_2
X_5682_ _6867_/Q _5628_/X _5666_/X _6891_/Q VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4633_ _4631_/D _4633_/B VGND VGND VPWR VPWR _4661_/B sky130_fd_sc_hd__and2b_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4564_ _4564_/A _4773_/A VGND VGND VPWR VPWR _4566_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold602 _7040_/Q VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 _4277_/X VGND VGND VPWR VPWR _6672_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6303_ _7130_/Q _6302_/X _6303_/S VGND VGND VPWR VPWR _6303_/X sky130_fd_sc_hd__mux2_2
Xhold624 _6849_/Q VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _3555_/A _3562_/B VGND VGND VPWR VPWR _4214_/A sky130_fd_sc_hd__nor2_4
Xhold635 _5420_/X VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ _4495_/A _4632_/B VGND VGND VPWR VPWR _5042_/B sky130_fd_sc_hd__nor2_4
Xhold646 _6445_/Q VGND VGND VPWR VPWR hold646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _5469_/X VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap376 _5611_/Y VGND VGND VPWR VPWR _6103_/B1 sky130_fd_sc_hd__buf_4
XFILLER_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold668 _5174_/X VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap387 _5631_/X VGND VGND VPWR VPWR _5818_/A2 sky130_fd_sc_hd__buf_8
X_6234_ _6477_/Q _5940_/X _5967_/X _6606_/Q _6231_/X VGND VGND VPWR VPWR _6234_/X
+ sky130_fd_sc_hd__a221o_1
Xhold679 _6833_/Q VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlygate4sd3_1
X_3446_ _3446_/A _3446_/B _3446_/C _3446_/D VGND VGND VPWR VPWR _3446_/Y sky130_fd_sc_hd__nor4_1
XFILLER_170_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6165_/A _6165_/B _6165_/C VGND VGND VPWR VPWR _6176_/C sky130_fd_sc_hd__nor3_2
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3377_ _3455_/A hold28/X VGND VGND VPWR VPWR _5541_/A sky130_fd_sc_hd__nor2_8
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _3991_/X VGND VGND VPWR VPWR _6434_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1313 _7034_/Q VGND VGND VPWR VPWR _5491_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5116_ _5116_/A VGND VGND VPWR VPWR _5116_/Y sky130_fd_sc_hd__inv_2
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 hold1324/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
X_6096_ _7030_/Q _5944_/X _5975_/A _6846_/Q _6095_/X VGND VGND VPWR VPWR _6099_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1335 hold1418/X VGND VGND VPWR VPWR hold1335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 hold1346/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1357 _6310_/A1 VGND VGND VPWR VPWR hold1357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 hold1368/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
X_5047_ _5047_/A _5096_/B VGND VGND VPWR VPWR _5122_/B sky130_fd_sc_hd__and2_1
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1379 hold1557/X VGND VGND VPWR VPWR hold1379/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6998_ _7065_/CLK _6998_/D fanout465/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfrtp_2
X_5949_ _5978_/A _5981_/A _5981_/B VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__and3_4
XFILLER_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3300_ _3355_/B _3311_/C VGND VGND VPWR VPWR _3300_/Y sky130_fd_sc_hd__nand2_8
XFILLER_140_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4280_ _4280_/A _5490_/B VGND VGND VPWR VPWR _4285_/S sky130_fd_sc_hd__and2_2
XFILLER_140_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3231_ _3837_/A _3234_/C VGND VGND VPWR VPWR _3829_/A sky130_fd_sc_hd__nand2_4
XFILLER_101_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6921_ _7001_/CLK _6921_/D fanout464/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6852_ _7049_/CLK _6852_/D fanout456/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5803_ _6993_/Q _5627_/X _5635_/X _6833_/Q VGND VGND VPWR VPWR _5803_/X sky130_fd_sc_hd__a22o_1
X_6783_ _6890_/CLK _6783_/D fanout476/X VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfrtp_1
X_3995_ hold586/X _6357_/A1 _3998_/S VGND VGND VPWR VPWR _3995_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5734_ _6789_/Q _5652_/Y _5728_/X _5733_/X _3178_/Y VGND VGND VPWR VPWR _5734_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_10_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5665_ _6858_/Q _5663_/X _5664_/X _6922_/Q VGND VGND VPWR VPWR _5665_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4616_ _4716_/A _4698_/C VGND VGND VPWR VPWR _4616_/Y sky130_fd_sc_hd__nand2_8
XFILLER_163_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5596_ _5596_/A1 _5574_/Y _5597_/B _5595_/X VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__a31o_1
XFILLER_135_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold410 _5517_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold421 _6671_/Q VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _4881_/B _4576_/B VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__nand2_4
Xhold432 _4325_/X VGND VGND VPWR VPWR _6712_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold443 _7193_/A VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _4148_/X VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold465 _6878_/Q VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold476 _5306_/X VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4642_/A _4739_/A VGND VGND VPWR VPWR _4653_/C sky130_fd_sc_hd__and2b_4
Xhold487 _6621_/Q VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 _5453_/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6217_ _6461_/Q _5945_/X _5975_/C _6579_/Q _6216_/X VGND VGND VPWR VPWR _6218_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3429_ input59/X _5193_/A _3358_/Y input18/X _3418_/X VGND VGND VPWR VPWR _3429_/X
+ sky130_fd_sc_hd__a221o_1
X_7197_ _7197_/A VGND VGND VPWR VPWR _7197_/X sky130_fd_sc_hd__clkbuf_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6448_/Q _5601_/X _5959_/X _6968_/Q VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__a22o_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1110 _5413_/X VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _6717_/Q VGND VGND VPWR VPWR _4331_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 _4175_/X VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 _6565_/Q VGND VGND VPWR VPWR _4158_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6079_ _7014_/Q _5940_/X _5967_/X _6854_/Q VGND VGND VPWR VPWR _6079_/X sky130_fd_sc_hd__a22o_1
Xhold1154 _5257_/X VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1165 hold1576/X VGND VGND VPWR VPWR _4110_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1176 _4053_/X VGND VGND VPWR VPWR _6490_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 _6442_/Q VGND VGND VPWR VPWR _4000_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _5326_/X VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3780_ input93/X _5190_/A _3355_/X _5283_/A _6850_/Q VGND VGND VPWR VPWR _3780_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5450_ hold152/X hold60/X _5453_/S VGND VGND VPWR VPWR _5450_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4401_ _4633_/B _4631_/D VGND VGND VPWR VPWR _4653_/B sky130_fd_sc_hd__and2b_4
X_5381_ hold307/X _5540_/A1 _5381_/S VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7131_/CLK sky130_fd_sc_hd__clkbuf_8
X_7120_ _7126_/CLK _7120_/D fanout466/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4332_ hold373/X _5494_/A1 _4333_/S VGND VGND VPWR VPWR _4332_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7051_ _7051_/CLK _7051_/D fanout485/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4263_ _4263_/A0 hold667/X _4267_/S VGND VGND VPWR VPWR _4263_/X sky130_fd_sc_hd__mux2_1
X_6002_ _6786_/Q _6226_/B _5610_/Y VGND VGND VPWR VPWR _6002_/Y sky130_fd_sc_hd__o21ai_1
X_3214_ _6861_/Q VGND VGND VPWR VPWR _3214_/Y sky130_fd_sc_hd__inv_2
X_4194_ _3447_/Y _4194_/A1 _4195_/S VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6904_ _7069_/CLK _6904_/D fanout482/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6835_ _7063_/CLK _6835_/D fanout463/X VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6766_ _6890_/CLK _6766_/D fanout470/X VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_4
X_3978_ _3978_/A0 hold99/X _3980_/S VGND VGND VPWR VPWR _3978_/X sky130_fd_sc_hd__mux2_1
X_5717_ _3207_/Y _5899_/B _5651_/B VGND VGND VPWR VPWR _5717_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6697_ _6755_/CLK _6697_/D fanout445/X VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3945_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5648_ _5664_/A _5658_/B _5663_/C VGND VGND VPWR VPWR _5648_/X sky130_fd_sc_hd__and3b_4
XFILLER_163_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5579_ _6508_/Q _5658_/B _5667_/C VGND VGND VPWR VPWR _5583_/S sky130_fd_sc_hd__and3_1
XFILLER_151_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold240 _4082_/X VGND VGND VPWR VPWR _6504_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _6787_/Q VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _5534_/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold273 _6620_/Q VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _5294_/X VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _6931_/Q VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_102 _7157_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_124 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _6431_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _5513_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 hold99/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _3700_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _4574_/A _4723_/B _4581_/Y _4810_/Y VGND VGND VPWR VPWR _4950_/X sky130_fd_sc_hd__a211o_1
X_3901_ _4374_/A _4702_/C _3901_/C _3901_/D VGND VGND VPWR VPWR _3907_/A sky130_fd_sc_hd__and4b_1
X_4881_ _4881_/A _4881_/B VGND VGND VPWR VPWR _4882_/C sky130_fd_sc_hd__nand2_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6620_ _6712_/CLK _6620_/D fanout470/X VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_4
X_3832_ _3837_/A _3832_/B VGND VGND VPWR VPWR _3838_/A sky130_fd_sc_hd__nor2_1
X_6551_ _6632_/CLK _6551_/D fanout454/X VGND VGND VPWR VPWR _6551_/Q sky130_fd_sc_hd__dfrtp_1
X_3763_ _3762_/Y _6727_/Q _3829_/A VGND VGND VPWR VPWR _3763_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5502_ _5502_/A0 hold42/X hold77/X VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__mux2_1
X_6482_ _6707_/CLK _6482_/D fanout450/X VGND VGND VPWR VPWR _6482_/Q sky130_fd_sc_hd__dfstp_2
X_3694_ _7057_/Q hold86/A _4232_/A _6627_/Q VGND VGND VPWR VPWR _3694_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5433_ hold698/X _5469_/A1 _5435_/S VGND VGND VPWR VPWR _5433_/X sky130_fd_sc_hd__mux2_1
Xoutput301 _3788_/Y VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
XFILLER_161_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput312 _7200_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
Xoutput323 hold1319/X VGND VGND VPWR VPWR hold1320/A sky130_fd_sc_hd__buf_12
X_5364_ _5364_/A hold17/X VGND VGND VPWR VPWR _5372_/S sky130_fd_sc_hd__and2_4
Xoutput334 hold1377/X VGND VGND VPWR VPWR hold1378/A sky130_fd_sc_hd__buf_12
Xoutput345 hold1341/X VGND VGND VPWR VPWR hold1342/A sky130_fd_sc_hd__buf_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7103_ _7131_/CLK _7103_/D fanout460/X VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4315_ hold614/X _6357_/A1 _4315_/S VGND VGND VPWR VPWR _4315_/X sky130_fd_sc_hd__mux2_1
X_5295_ hold407/X _5544_/A1 _5300_/S VGND VGND VPWR VPWR _5295_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7034_ _7037_/CLK _7034_/D fanout450/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_2
X_4246_ hold415/X _5534_/A1 _4249_/S VGND VGND VPWR VPWR _4246_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4177_ hold562/X _6357_/A1 _4177_/S VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6818_ _7067_/CLK _6818_/D fanout476/X VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_11_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6749_ _6749_/CLK _6749_/D fanout449/X VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4100_ hold341/X _5540_/A1 _5202_/B VGND VGND VPWR VPWR _4100_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5080_ _5080_/A _5080_/B _5080_/C VGND VGND VPWR VPWR _5087_/A sky130_fd_sc_hd__and3_1
XFILLER_96_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4031_ _4031_/A0 hold60/X hold68/X VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__mux2_1
XFILLER_96_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5982_ _6810_/Q _5971_/B _5946_/X _6890_/Q VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4933_ _5068_/C _5002_/C _4933_/C _5138_/A VGND VGND VPWR VPWR _4944_/A sky130_fd_sc_hd__and4_1
XFILLER_80_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4864_ _4618_/Y _4694_/Y _5084_/A VGND VGND VPWR VPWR _4864_/X sky130_fd_sc_hd__o21a_1
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 _5265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3815_ _7002_/Q _3370_/Y _5184_/A _6764_/Q VGND VGND VPWR VPWR _3815_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_24 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _6674_/CLK _6603_/D _6383_/A VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_35 _3828_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _5627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _4546_/Y _4631_/Y _4697_/Y VGND VGND VPWR VPWR _4796_/D sky130_fd_sc_hd__o21a_1
XANTENNA_57 _5971_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6534_ _6539_/CLK _6534_/D fanout461/X VGND VGND VPWR VPWR _6534_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_68 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ _6762_/Q _5182_/S _4304_/A _6696_/Q _3745_/X VGND VGND VPWR VPWR _3751_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA_79 _6787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6465_ _6654_/CLK _6465_/D _6401_/A VGND VGND VPWR VPWR _6465_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3677_ _7028_/Q hold49/A _5505_/A _7049_/Q VGND VGND VPWR VPWR _3677_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5416_ hold924/X _5548_/A1 _5417_/S VGND VGND VPWR VPWR _5416_/X sky130_fd_sc_hd__mux2_1
X_6396_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6396_/X sky130_fd_sc_hd__and2_1
X_5347_ _5347_/A0 _5473_/A1 _5354_/S VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__mux2_1
Xoutput175 _3935_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
XFILLER_142_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput186 _3934_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3220_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_102_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5278_ hold914/X _5509_/A1 _5282_/S VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__mux2_1
X_7017_ _7017_/CLK _7017_/D fanout461/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_1
X_4229_ _6640_/Q _4230_/B VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__and2b_4
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3600_ _6893_/Q _5328_/A _5166_/A _6754_/Q _3591_/X VGND VGND VPWR VPWR _3604_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4580_ _4561_/B _4611_/B _4948_/D _4578_/X _4575_/Y VGND VGND VPWR VPWR _4580_/X
+ sky130_fd_sc_hd__o32a_1
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_2
X_3531_ _6564_/Q _4151_/A _4262_/A _6664_/Q VGND VGND VPWR VPWR _3531_/X sky130_fd_sc_hd__a22o_2
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_2
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7200_/A sky130_fd_sc_hd__buf_4
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
Xhold806 _7075_/Q VGND VGND VPWR VPWR hold806/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 _5546_/X VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _6427_/Q VGND VGND VPWR VPWR hold828/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _3949_/B sky130_fd_sc_hd__buf_4
X_6250_ _6250_/A _6250_/B _6250_/C _6250_/D VGND VGND VPWR VPWR _6251_/B sky130_fd_sc_hd__nor4_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold839 _4303_/X VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR _4563_/A sky130_fd_sc_hd__clkbuf_16
X_3462_ _6975_/Q _5418_/A _5373_/A _6935_/Q VGND VGND VPWR VPWR _3462_/X sky130_fd_sc_hd__a22o_2
XFILLER_115_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5201_ hold395/X _5540_/A1 _5201_/S VGND VGND VPWR VPWR _5201_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6181_ _6609_/Q _5943_/X _5981_/X _6655_/Q VGND VGND VPWR VPWR _6181_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3393_ _6953_/Q _3781_/A2 _3358_/Y input19/X _3383_/X VGND VGND VPWR VPWR _3393_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5132_ _5087_/A _5120_/X _5131_/X _5116_/Y VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__a31o_1
XFILLER_123_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1506 _7131_/Q VGND VGND VPWR VPWR _6304_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1517 _7128_/Q VGND VGND VPWR VPWR _6229_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5063_ _4619_/Y _5010_/Y _4974_/B VGND VGND VPWR VPWR _5064_/C sky130_fd_sc_hd__o21a_1
Xhold1528 _7161_/Q VGND VGND VPWR VPWR _3259_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _7150_/Q VGND VGND VPWR VPWR _6351_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4014_ _4014_/A _6352_/B VGND VGND VPWR VPWR _4019_/S sky130_fd_sc_hd__and2_2
XFILLER_38_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5965_ _5979_/A _5981_/B _5969_/C VGND VGND VPWR VPWR _5965_/X sky130_fd_sc_hd__and3_4
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4916_ _5118_/A _4916_/B _4916_/C VGND VGND VPWR VPWR _4918_/B sky130_fd_sc_hd__and3_1
X_5896_ _5896_/A _5896_/B _5896_/C VGND VGND VPWR VPWR _5896_/Y sky130_fd_sc_hd__nor3_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4847_ _4847_/A VGND VGND VPWR VPWR _4847_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4778_ _5023_/B _5039_/B _4777_/X _4593_/Y VGND VGND VPWR VPWR _4884_/B sky130_fd_sc_hd__a31o_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3729_ _3729_/A _3729_/B _3729_/C _3729_/D VGND VGND VPWR VPWR _3730_/C sky130_fd_sc_hd__nor4_4
X_6517_ _7076_/CLK _6517_/D fanout481/X VGND VGND VPWR VPWR _6517_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6448_ _7086_/CLK _6448_/D fanout483/X VGND VGND VPWR VPWR _6448_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6379_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6379_/X sky130_fd_sc_hd__and2_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5750_ _6838_/Q _5928_/A2 _5740_/X _5749_/X VGND VGND VPWR VPWR _5754_/A sky130_fd_sc_hd__a211o_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4702_/A _4702_/B _4702_/C VGND VGND VPWR VPWR _4701_/Y sky130_fd_sc_hd__nand3_2
X_5681_ _5681_/A _5681_/B _5681_/C VGND VGND VPWR VPWR _5681_/Y sky130_fd_sc_hd__nor3_1
X_4632_ _4753_/B _4632_/B VGND VGND VPWR VPWR _4632_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4563_ _4563_/A _4631_/D _4633_/B _4563_/D VGND VGND VPWR VPWR _4773_/A sky130_fd_sc_hd__and4_1
Xhold603 _5498_/X VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6302_ _6289_/Y _6301_/X _6544_/Q _6226_/B VGND VGND VPWR VPWR _6302_/X sky130_fd_sc_hd__o2bb2a_1
Xhold614 _6704_/Q VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _6649_/Q _4244_/A _3511_/Y _3513_/X _3414_/Y VGND VGND VPWR VPWR _3523_/B
+ sky130_fd_sc_hd__a2111o_1
Xhold625 _5282_/X VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold636 _6952_/Q VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _5010_/A _4881_/B VGND VGND VPWR VPWR _4494_/Y sky130_fd_sc_hd__nand2_1
Xhold647 _4003_/X VGND VGND VPWR VPWR _6445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _6945_/Q VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ _6692_/Q _5954_/X _5976_/D _6621_/Q _6230_/X VGND VGND VPWR VPWR _6250_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold669 _6864_/Q VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlygate4sd3_1
X_3445_ _6968_/Q _5409_/A _3365_/Y input9/X _3444_/X VGND VGND VPWR VPWR _3446_/D
+ sky130_fd_sc_hd__a221o_1
Xmax_cap377 hold74/X VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__buf_12
XFILLER_171_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap388 _5616_/X VGND VGND VPWR VPWR _5902_/A2 sky130_fd_sc_hd__buf_8
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6985_/Q _5945_/X _5975_/C _6841_/Q _6157_/X VGND VGND VPWR VPWR _6165_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3717_/B _3376_/B VGND VGND VPWR VPWR _3964_/A sky130_fd_sc_hd__nor2_8
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5115_ _5115_/A _5115_/B _5115_/C _5115_/D VGND VGND VPWR VPWR _5116_/A sky130_fd_sc_hd__and4_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 _6540_/Q VGND VGND VPWR VPWR _4128_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 _5491_/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6095_ _7022_/Q _5937_/X _5975_/D _6886_/Q VGND VGND VPWR VPWR _6095_/X sky130_fd_sc_hd__a22o_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 hold1422/X VGND VGND VPWR VPWR hold1325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1336 hold1336/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
Xhold1347 hold1429/X VGND VGND VPWR VPWR hold1347/X sky130_fd_sc_hd__dlygate4sd3_1
X_5046_ _5046_/A _5046_/B _5046_/C VGND VGND VPWR VPWR _5096_/B sky130_fd_sc_hd__and3_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1358 hold1358/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
Xhold1369 _4191_/A1 VGND VGND VPWR VPWR hold1369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6997_ _6997_/CLK _6997_/D fanout465/X VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5948_ _5969_/A _5981_/A _5981_/C VGND VGND VPWR VPWR _5948_/X sky130_fd_sc_hd__and3_4
XFILLER_185_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5879_ _6452_/Q _5634_/X _5876_/X _5878_/X VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__a211o_1
XFILLER_178_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3230_ _6417_/Q _6416_/Q VGND VGND VPWR VPWR _3234_/C sky130_fd_sc_hd__nor2_1
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6920_ _6920_/CLK _6920_/D fanout473/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6851_ _6963_/CLK _6851_/D fanout456/X VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5802_ _3228_/Y _5899_/B _5651_/B VGND VGND VPWR VPWR _5802_/Y sky130_fd_sc_hd__a21oi_1
X_3994_ hold772/X _6356_/A1 _3998_/S VGND VGND VPWR VPWR _3994_/X sky130_fd_sc_hd__mux2_1
X_6782_ _6969_/CLK _6782_/D fanout481/X VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5733_ _6805_/Q _5660_/X _5729_/X _5731_/X _5732_/X VGND VGND VPWR VPWR _5733_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5664_ _5664_/A _5667_/C _5666_/C VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__and3_4
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4615_ _4661_/A _4615_/B VGND VGND VPWR VPWR _4615_/Y sky130_fd_sc_hd__nand2_1
X_5595_ _6508_/Q _5969_/A _5968_/A VGND VGND VPWR VPWR _5595_/X sky130_fd_sc_hd__and3_1
Xhold400 _5385_/X VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _7076_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _4562_/A _4753_/B VGND VGND VPWR VPWR _4546_/Y sky130_fd_sc_hd__nand2_1
Xhold422 _4276_/X VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold433 _6522_/Q VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold444 _5198_/X VGND VGND VPWR VPWR _6774_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _7022_/Q VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 _5315_/X VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _5010_/A _4650_/A VGND VGND VPWR VPWR _5088_/A sky130_fd_sc_hd__nand2_4
Xhold477 _6934_/Q VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold488 _4223_/X VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3428_ _6928_/Q _5364_/A _3981_/A _6432_/Q _3427_/X VGND VGND VPWR VPWR _3428_/X
+ sky130_fd_sc_hd__a221o_1
X_6216_ _6666_/Q _5938_/X _5952_/X _6706_/Q VGND VGND VPWR VPWR _6216_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_69_csclk _7001_/CLK VGND VGND VPWR VPWR _7026_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold499 _6658_/Q VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__dlygate4sd3_1
X_7196_ _7196_/A VGND VGND VPWR VPWR _7196_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _7032_/Q _5944_/X _5975_/A _6848_/Q _6146_/X VGND VGND VPWR VPWR _6150_/C
+ sky130_fd_sc_hd__a221o_1
X_3359_ _3562_/A hold28/X VGND VGND VPWR VPWR _5256_/A sky130_fd_sc_hd__nor2_8
Xhold1100 _5230_/X VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _6677_/Q VGND VGND VPWR VPWR _4283_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1122 _4331_/X VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 _6818_/Q VGND VGND VPWR VPWR _5248_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 _4158_/X VGND VGND VPWR VPWR _6565_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6078_ _6078_/A0 _6077_/X _6279_/S VGND VGND VPWR VPWR _6078_/X sky130_fd_sc_hd__mux2_1
Xhold1155 _6670_/Q VGND VGND VPWR VPWR _4275_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 _4110_/X VGND VGND VPWR VPWR _6524_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1177 _6665_/Q VGND VGND VPWR VPWR _4269_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5029_ _5029_/A _5029_/B VGND VGND VPWR VPWR _5083_/C sky130_fd_sc_hd__and2_1
Xhold1188 _4000_/X VGND VGND VPWR VPWR _6442_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 _6962_/Q VGND VGND VPWR VPWR _5410_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4400_ _4631_/D _4400_/B VGND VGND VPWR VPWR _4408_/B sky130_fd_sc_hd__xnor2_2
XFILLER_145_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5380_ hold930/X _5548_/A1 _5381_/S VGND VGND VPWR VPWR _5380_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4331_ _4331_/A0 _5493_/A1 _4333_/S VGND VGND VPWR VPWR _4331_/X sky130_fd_sc_hd__mux2_1
X_7050_ _7086_/CLK _7050_/D fanout483/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4262_ _4262_/A _4322_/B VGND VGND VPWR VPWR _4267_/S sky130_fd_sc_hd__and2_2
XFILLER_140_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6001_ _5992_/X _6226_/B _6001_/C _6001_/D VGND VGND VPWR VPWR _6001_/X sky130_fd_sc_hd__and4b_1
XFILLER_101_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3213_ _6869_/Q VGND VGND VPWR VPWR _3213_/Y sky130_fd_sc_hd__inv_2
X_4193_ _3486_/Y _4193_/A1 _4195_/S VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6903_ _7076_/CLK _6903_/D fanout481/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6834_ _7026_/CLK _6834_/D fanout463/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6765_ _6890_/CLK _6765_/D fanout470/X VGND VGND VPWR VPWR _6765_/Q sky130_fd_sc_hd__dfrtp_4
X_3977_ hold97/X hold106/X _6624_/Q VGND VGND VPWR VPWR _3977_/X sky130_fd_sc_hd__mux2_2
XFILLER_149_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5716_ _6445_/Q _5614_/X _5666_/X _6893_/Q VGND VGND VPWR VPWR _5716_/X sky130_fd_sc_hd__a22o_1
X_6696_ _6755_/CLK _6696_/D _6360_/A VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _7026_/Q _5645_/X _5646_/X _6906_/Q _5644_/X VGND VGND VPWR VPWR _5669_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5578_ _7095_/Q _7094_/Q VGND VGND VPWR VPWR _5667_/C sky130_fd_sc_hd__nor2_4
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold230 _4285_/X VGND VGND VPWR VPWR _6679_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold241 _6925_/Q VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _5213_/X VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4413_/Y _4724_/A VGND VGND VPWR VPWR _4529_/Y sky130_fd_sc_hd__nand2b_1
Xhold263 _6443_/Q VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold274 _4222_/X VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold285 _6827_/Q VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _5375_/X VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7179_ _7179_/A VGND VGND VPWR VPWR _7179_/X sky130_fd_sc_hd__clkbuf_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _7173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 _3957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_136 _6432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _6357_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 hold99/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _3803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_2
XFILLER_162_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3900_ input118/X input119/X _3900_/C _3900_/D VGND VGND VPWR VPWR _3901_/D sky130_fd_sc_hd__and4bb_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4880_ _4951_/B _5086_/B _5073_/A _4880_/D VGND VGND VPWR VPWR _4882_/B sky130_fd_sc_hd__and4_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3831_ _3837_/B _3837_/C VGND VGND VPWR VPWR _3832_/B sky130_fd_sc_hd__and2_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3762_ _3762_/A _3762_/B VGND VGND VPWR VPWR _3762_/Y sky130_fd_sc_hd__nand2_4
X_6550_ _6654_/CLK _6550_/D fanout454/X VGND VGND VPWR VPWR _6550_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5501_ hold182/X _5519_/A1 hold77/A VGND VGND VPWR VPWR _5501_/X sky130_fd_sc_hd__mux2_1
X_6481_ _6704_/CLK _6481_/D fanout450/X VGND VGND VPWR VPWR _6481_/Q sky130_fd_sc_hd__dfrtp_2
X_3693_ _6542_/Q _4127_/A _3692_/Y _6765_/Q _3691_/X VGND VGND VPWR VPWR _3698_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5432_ hold147/X hold60/X _5435_/S VGND VGND VPWR VPWR _5432_/X sky130_fd_sc_hd__mux2_1
Xoutput302 _3956_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
XFILLER_133_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput313 hold1379/X VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
X_5363_ hold489/X hold22/X _5363_/S VGND VGND VPWR VPWR _5363_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput324 hold1321/X VGND VGND VPWR VPWR hold1322/A sky130_fd_sc_hd__buf_12
Xoutput335 hold1361/X VGND VGND VPWR VPWR hold1362/A sky130_fd_sc_hd__buf_12
X_7102_ _7113_/CLK _7102_/D fanout464/X VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfrtp_4
X_4314_ hold782/X _6356_/A1 _4315_/S VGND VGND VPWR VPWR _4314_/X sky130_fd_sc_hd__mux2_1
X_5294_ hold283/X _5465_/A1 _5300_/S VGND VGND VPWR VPWR _5294_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7033_ _7033_/CLK _7033_/D fanout464/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_2
X_4245_ _4245_/A0 hold667/X _4249_/S VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4176_ hold734/X _6356_/A1 _4177_/S VGND VGND VPWR VPWR _4176_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ _7070_/CLK _6817_/D fanout473/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6748_ _6926_/CLK _6748_/D fanout449/X VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_137_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6679_ _7036_/CLK _6679_/D fanout455/X VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmgmt_gpio_14_buff_inst _3937_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_8
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4030_ _4030_/A0 _5494_/A1 hold68/X VGND VGND VPWR VPWR _4030_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5981_ _5981_/A _5981_/B _5981_/C VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__and3_4
XFILLER_80_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4932_ _4542_/A _4562_/Y _4673_/A _4628_/Y _4755_/X VGND VGND VPWR VPWR _5138_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4863_ _4542_/B _4496_/Y _4618_/Y _4700_/Y VGND VGND VPWR VPWR _4877_/C sky130_fd_sc_hd__o22a_1
XANTENNA_14 _5505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ _6769_/CLK _6602_/D fanout469/X VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_1
X_3814_ _3814_/A _3814_/B VGND VGND VPWR VPWR _5184_/A sky130_fd_sc_hd__nor2_1
XANTENNA_25 _4202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_36 _4084_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4846_/B _4616_/Y _4619_/Y _4689_/A VGND VGND VPWR VPWR _4796_/C sky130_fd_sc_hd__o22a_1
XANTENNA_47 _5631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _6301_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6533_ _6755_/CLK _6533_/D _6360_/A VGND VGND VPWR VPWR _6533_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_69 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ _6859_/Q _5292_/A _3370_/Y _7003_/Q VGND VGND VPWR VPWR _3745_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6464_ _6668_/CLK _6464_/D _6360_/A VGND VGND VPWR VPWR _6464_/Q sky130_fd_sc_hd__dfrtp_4
X_3676_ _6900_/Q _5337_/A _5301_/A _6868_/Q _3675_/X VGND VGND VPWR VPWR _3679_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5415_ hold469/X _5469_/A1 _5417_/S VGND VGND VPWR VPWR _5415_/X sky130_fd_sc_hd__mux2_1
X_6395_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6395_/X sky130_fd_sc_hd__and2_1
XFILLER_114_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5346_ _5346_/A _5541_/B VGND VGND VPWR VPWR _5354_/S sky130_fd_sc_hd__and2_4
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput176 _3213_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3203_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3193_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_102_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5277_ _5277_/A0 _5484_/A1 _5282_/S VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7016_ _7016_/CLK _7016_/D fanout474/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4228_ _6638_/Q _4228_/B VGND VGND VPWR VPWR _4228_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4159_ hold810/X _6354_/A1 _4162_/S VGND VGND VPWR VPWR _4159_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout392 hold22/X VGND VGND VPWR VPWR _5513_/A1 sky130_fd_sc_hd__buf_8
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_2
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_2
X_3530_ hold36/X hold66/X VGND VGND VPWR VPWR _4262_/A sky130_fd_sc_hd__nor2_8
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_2
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _3268_/C sky130_fd_sc_hd__buf_6
XFILLER_143_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold807 _5537_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold818 _6696_/Q VGND VGND VPWR VPWR hold818/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_2
Xhold829 _3983_/X VGND VGND VPWR VPWR _6427_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3461_ _6967_/Q _5409_/A _3964_/A _6423_/Q _3456_/X VGND VGND VPWR VPWR _3467_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5200_ hold365/X _5521_/A1 _5201_/S VGND VGND VPWR VPWR _5200_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3392_ _3392_/A _3392_/B _3392_/C _3392_/D VGND VGND VPWR VPWR _3392_/Y sky130_fd_sc_hd__nor4_1
X_6180_ _6660_/Q _5976_/B _5971_/C _6710_/Q VGND VGND VPWR VPWR _6180_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5131_ _5131_/A _5131_/B _5131_/C VGND VGND VPWR VPWR _5131_/X sky130_fd_sc_hd__and3_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1507 _7108_/Q VGND VGND VPWR VPWR _5735_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5062_ _5062_/A _5062_/B _5062_/C _5062_/D VGND VGND VPWR VPWR _5134_/B sky130_fd_sc_hd__and4_1
Xhold1518 _7111_/Q VGND VGND VPWR VPWR _5778_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _3258_/X VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4013_ hold978/X _5546_/A1 _4013_/S VGND VGND VPWR VPWR _4013_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5964_ _5964_/A _5969_/C _5981_/C VGND VGND VPWR VPWR _5975_/D sky130_fd_sc_hd__and3_4
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4915_ _4906_/Y _4915_/B _4915_/C _4915_/D VGND VGND VPWR VPWR _4916_/C sky130_fd_sc_hd__and4b_1
XFILLER_80_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5895_ _6688_/Q _5632_/X _5892_/X _5894_/X VGND VGND VPWR VPWR _5896_/C sky130_fd_sc_hd__a211o_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4846_ _4846_/A _4846_/B VGND VGND VPWR VPWR _4847_/A sky130_fd_sc_hd__nor2_1
XFILLER_166_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4777_ _4753_/A _4602_/Y _5114_/B _4776_/X VGND VGND VPWR VPWR _4777_/X sky130_fd_sc_hd__o211a_1
X_6516_ _7076_/CLK _6516_/D fanout481/X VGND VGND VPWR VPWR _6516_/Q sky130_fd_sc_hd__dfrtp_1
X_3728_ _6939_/Q _5382_/A _4196_/A _6600_/Q _3727_/X VGND VGND VPWR VPWR _3729_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_107_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6447_ _6447_/CLK _6447_/D fanout461/X VGND VGND VPWR VPWR _6447_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3659_ _6908_/Q _5346_/A _5355_/A _6916_/Q VGND VGND VPWR VPWR _3659_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6378_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6378_/X sky130_fd_sc_hd__and2_1
XFILLER_0_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5329_ _5329_/A0 _5473_/A1 _5336_/S VGND VGND VPWR VPWR _5329_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4716_/A _4911_/B VGND VGND VPWR VPWR _4700_/Y sky130_fd_sc_hd__nand2_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _7019_/Q _5619_/X _5677_/X _5679_/X VGND VGND VPWR VPWR _5681_/C sky130_fd_sc_hd__a211o_2
XFILLER_148_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4631_ _4633_/B _4716_/A _4653_/C _4631_/D VGND VGND VPWR VPWR _4631_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4562_ _4562_/A _4600_/B VGND VGND VPWR VPWR _4562_/Y sky130_fd_sc_hd__nand2_8
XFILLER_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6301_ _6292_/X _6301_/B _6301_/C VGND VGND VPWR VPWR _6301_/X sky130_fd_sc_hd__and3b_1
Xhold604 _6811_/Q VGND VGND VPWR VPWR hold604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 _4315_/X VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _7067_/Q _5523_/A _4020_/A _6464_/Q VGND VGND VPWR VPWR _3513_/X sky130_fd_sc_hd__a22o_1
Xhold626 _7017_/Q VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4493_ _5010_/A _4493_/B VGND VGND VPWR VPWR _5083_/A sky130_fd_sc_hd__nand2_1
Xhold637 _5398_/X VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _7007_/Q VGND VGND VPWR VPWR hold648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 _5390_/X VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _7153_/Q _5958_/X _5978_/X _6482_/Q VGND VGND VPWR VPWR _6232_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3444_ _6952_/Q _5391_/A hold29/A _7024_/Q VGND VGND VPWR VPWR _3444_/X sky130_fd_sc_hd__a22o_1
Xmax_cap378 _3543_/A VGND VGND VPWR VPWR _3573_/A sky130_fd_sc_hd__buf_12
XFILLER_103_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6977_/Q _5947_/X _5965_/X _6801_/Q _6162_/X VGND VGND VPWR VPWR _6165_/B
+ sky130_fd_sc_hd__a221o_1
X_3375_ _3375_/A _3415_/B VGND VGND VPWR VPWR _3814_/B sky130_fd_sc_hd__nand2_8
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A _5114_/B _5114_/C _5114_/D VGND VGND VPWR VPWR _5115_/D sky130_fd_sc_hd__and4_1
Xhold1304 _4128_/X VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _7067_/Q _5934_/X _5975_/B _6870_/Q _6093_/X VGND VGND VPWR VPWR _6094_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1315 hold1412/X VGND VGND VPWR VPWR hold1315/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1326 hold1326/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
Xhold1337 hold1421/X VGND VGND VPWR VPWR hold1337/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1348 hold1348/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
X_5045_ _4947_/B _4453_/B _4570_/Y VGND VGND VPWR VPWR _5046_/C sky130_fd_sc_hd__a21o_1
Xhold1359 _4168_/A1 VGND VGND VPWR VPWR hold1359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6996_ _7063_/CLK _6996_/D fanout463/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5947_ _5969_/A _5968_/A _5981_/A VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__and3_4
XFILLER_178_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5878_ _6647_/Q _5621_/X _5648_/X _6606_/Q _5877_/X VGND VGND VPWR VPWR _5878_/X
+ sky130_fd_sc_hd__a221o_1
X_4829_ _4456_/Y _4810_/B _4818_/X _4820_/X VGND VGND VPWR VPWR _4829_/X sky130_fd_sc_hd__o211a_1
XFILLER_138_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6850_ _6926_/CLK _6850_/D fanout457/X VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5801_ _6905_/Q _5621_/X _5648_/X _6857_/Q VGND VGND VPWR VPWR _5801_/X sky130_fd_sc_hd__a22o_1
X_6781_ _6969_/CLK _6781_/D fanout473/X VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtp_1
X_3993_ hold984/X _6355_/A1 _3998_/S VGND VGND VPWR VPWR _3993_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5732_ _6925_/Q _5664_/X _5716_/X _5718_/X VGND VGND VPWR VPWR _5732_/X sky130_fd_sc_hd__a211o_1
XFILLER_188_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5663_ _5664_/A _5666_/C _5663_/C VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__and3b_4
XFILLER_129_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4614_ _4661_/A _4615_/B VGND VGND VPWR VPWR _4698_/C sky130_fd_sc_hd__and2_2
X_5594_ _5594_/A _5964_/A VGND VGND VPWR VPWR _5597_/B sky130_fd_sc_hd__nand2_1
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold401 _6534_/Q VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4545_ _4562_/A _4753_/B VGND VGND VPWR VPWR _4576_/B sky130_fd_sc_hd__and2_2
Xhold412 _5538_/X VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _6769_/Q VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _4107_/X VGND VGND VPWR VPWR _6522_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold445 _6950_/Q VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold456 _5477_/X VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _4984_/A _4710_/A VGND VGND VPWR VPWR _4476_/Y sky130_fd_sc_hd__nand2_1
Xhold467 _6846_/Q VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _5378_/X VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6451_/Q _5947_/X _5965_/X _6546_/Q _6214_/X VGND VGND VPWR VPWR _6218_/B
+ sky130_fd_sc_hd__a221o_1
Xhold489 _6921_/Q VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__dlygate4sd3_1
X_3427_ input69/X _4083_/S _5532_/A _7077_/Q VGND VGND VPWR VPWR _3427_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7195_ _7195_/A VGND VGND VPWR VPWR _7195_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _7024_/Q _5937_/X _5975_/D _6888_/Q VGND VGND VPWR VPWR _6146_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _3511_/A _3573_/B VGND VGND VPWR VPWR _3358_/Y sky130_fd_sc_hd__nor2_8
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _6869_/Q VGND VGND VPWR VPWR _5305_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 _4283_/X VGND VGND VPWR VPWR _6677_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1123 _6632_/Q VGND VGND VPWR VPWR _4241_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _7121_/Q _6076_/X _6303_/S VGND VGND VPWR VPWR _6077_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1134 _5248_/X VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3289_ hold32/X _6488_/Q _3288_/Y VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__a21bo_1
Xhold1145 _6512_/Q VGND VGND VPWR VPWR _4091_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 _4275_/X VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1167 _6550_/Q VGND VGND VPWR VPWR _4140_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 _4269_/X VGND VGND VPWR VPWR _6665_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5028_ _4623_/Y _4695_/Y _4875_/A _4522_/D VGND VGND VPWR VPWR _5085_/B sky130_fd_sc_hd__o211a_1
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _7151_/Q VGND VGND VPWR VPWR _6353_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6979_ _7063_/CLK _6979_/D fanout463/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold990 _6763_/Q VGND VGND VPWR VPWR hold990/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4330_ _4330_/A0 _5492_/A1 _4333_/S VGND VGND VPWR VPWR _4330_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4261_ hold970/X _5546_/A1 _4261_/S VGND VGND VPWR VPWR _4261_/X sky130_fd_sc_hd__mux2_1
X_6000_ _6000_/A _6000_/B _6000_/C _6000_/D VGND VGND VPWR VPWR _6001_/D sky130_fd_sc_hd__nor4_1
XFILLER_86_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3212_ _6877_/Q VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4192_ _4192_/A0 _4192_/A1 _4195_/S VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6902_ _7079_/CLK _6902_/D fanout478/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfrtp_2
X_6833_ _6969_/CLK _6833_/D fanout473/X VGND VGND VPWR VPWR _6833_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6764_ _6926_/CLK _6764_/D fanout457/X VGND VGND VPWR VPWR _6764_/Q sky130_fd_sc_hd__dfrtp_1
X_3976_ hold689/X _5469_/A1 _3980_/S VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5715_ _6845_/Q _5902_/A2 _5928_/A2 _6837_/Q VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__a22o_1
X_6695_ _6735_/CLK _6695_/D fanout445/X VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5646_ _5664_/A _5667_/B _5666_/B VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__and3b_4
XFILLER_164_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5577_ _7094_/Q _5576_/B _5574_/Y _5576_/Y VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__a31o_1
XFILLER_117_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold220 _5449_/X VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 _6981_/Q VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4528_ _4542_/B _4947_/B _4902_/A _4413_/Y _4527_/X VGND VGND VPWR VPWR _4528_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_191_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold242 _5368_/X VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _7003_/Q VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _4001_/X VGND VGND VPWR VPWR _6443_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold275 _7011_/Q VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _5258_/X VGND VGND VPWR VPWR _6827_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _4459_/A _4459_/B VGND VGND VPWR VPWR _4542_/D sky130_fd_sc_hd__nand2_4
Xhold297 _6835_/Q VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7178_ _7178_/A VGND VGND VPWR VPWR _7178_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6129_ _6129_/A0 _6128_/X _6304_/S VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__mux2_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_115 _3251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _6433_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_148 _5528_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 hold666/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _3830_/A1 _3829_/B _3828_/Y _3829_/Y VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_68_csclk _7001_/CLK VGND VGND VPWR VPWR _7063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3761_ _3733_/X _3761_/B _3761_/C _3761_/D VGND VGND VPWR VPWR _3762_/B sky130_fd_sc_hd__and4b_1
XFILLER_13_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5500_ hold590/X _5509_/A1 hold77/X VGND VGND VPWR VPWR _5500_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6480_ _6707_/CLK _6480_/D fanout450/X VGND VGND VPWR VPWR _6480_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3692_ _3692_/A _3714_/B VGND VGND VPWR VPWR _3692_/Y sky130_fd_sc_hd__nor2_2
XFILLER_145_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5431_ hold231/X _5494_/A1 _5435_/S VGND VGND VPWR VPWR _5431_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput303 _5606_/A VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput314 hold1371/X VGND VGND VPWR VPWR hold1372/A sky130_fd_sc_hd__buf_12
X_5362_ hold718/X _5521_/A1 _5363_/S VGND VGND VPWR VPWR _5362_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput325 hold1365/X VGND VGND VPWR VPWR hold1366/A sky130_fd_sc_hd__buf_12
XFILLER_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput336 hold1367/X VGND VGND VPWR VPWR hold1368/A sky130_fd_sc_hd__buf_12
XFILLER_160_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7101_ _7113_/CLK _7101_/D fanout464/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfstp_2
X_4313_ hold972/X _6355_/A1 _4315_/S VGND VGND VPWR VPWR _4313_/X sky130_fd_sc_hd__mux2_1
X_5293_ _5293_/A0 _6353_/A1 _5300_/S VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7032_ _7086_/CLK _7032_/D fanout483/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_4
X_4244_ _4244_/A _4322_/B VGND VGND VPWR VPWR _4249_/S sky130_fd_sc_hd__and2_2
XFILLER_141_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4175_ _4175_/A0 _6355_/A1 _4177_/S VGND VGND VPWR VPWR _4175_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6816_ _7069_/CLK _6816_/D fanout482/X VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6747_ _6747_/CLK _6747_/D fanout447/X VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_4
X_3959_ _6768_/Q _3959_/B VGND VGND VPWR VPWR _3959_/X sky130_fd_sc_hd__and2_2
XFILLER_149_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6678_ _7037_/CLK _6678_/D fanout455/X VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5629_ _6986_/Q _5627_/X _5628_/X _6866_/Q _5626_/X VGND VGND VPWR VPWR _5641_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5980_ _6850_/Q _5967_/X _5979_/X _6986_/Q VGND VGND VPWR VPWR _5980_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4931_ _4741_/A _4741_/B _4921_/Y _4612_/Y _4663_/Y VGND VGND VPWR VPWR _4933_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_33_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4862_ _4456_/Y _4496_/Y _4689_/Y VGND VGND VPWR VPWR _4872_/B sky130_fd_sc_hd__o21ba_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6601_ _6601_/CLK _6601_/D fanout469/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfstp_2
X_3813_ _6858_/Q _5292_/A _5328_/A _6890_/Q _3812_/X VGND VGND VPWR VPWR _3817_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_15 _5505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _4127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4846_/B _4619_/Y _4645_/Y _4689_/A VGND VGND VPWR VPWR _5064_/A sky130_fd_sc_hd__o22a_1
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_37 _4108_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _5637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6532_ _6735_/CLK _6532_/D _3946_/B VGND VGND VPWR VPWR _6532_/Q sky130_fd_sc_hd__dfrtp_1
X_3744_ _6743_/Q _5154_/A _4214_/A _6615_/Q _3743_/X VGND VGND VPWR VPWR _3751_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA_59 _6301_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6463_ _6668_/CLK _6463_/D _6400_/A VGND VGND VPWR VPWR _6463_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3675_ _6924_/Q _5364_/A _4316_/A _6707_/Q VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5414_ hold802/X _5546_/A1 _5417_/S VGND VGND VPWR VPWR _5414_/X sky130_fd_sc_hd__mux2_1
X_6394_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6394_/X sky130_fd_sc_hd__and2_1
X_5345_ hold331/X _5540_/A1 _5345_/S VGND VGND VPWR VPWR _5345_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput177 _3212_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3202_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
X_5276_ hold560/X _5543_/A1 _5282_/S VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__mux2_1
Xoutput199 _3192_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7015_ _7017_/CLK _7015_/D fanout461/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4227_ _6636_/Q _6637_/Q _6639_/Q VGND VGND VPWR VPWR _4228_/B sky130_fd_sc_hd__nor3_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ _4158_/A0 _5491_/A1 _4162_/S VGND VGND VPWR VPWR _4158_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4089_ hold610/X _4088_/X _4101_/S VGND VGND VPWR VPWR _4089_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout393 hold22/X VGND VGND VPWR VPWR _5540_/A1 sky130_fd_sc_hd__buf_6
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_2
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_2
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__buf_2
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _3956_/A sky130_fd_sc_hd__clkbuf_4
Xhold808 _6541_/Q VGND VGND VPWR VPWR hold808/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold819 _4306_/X VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput79 spi_enabled VGND VGND VPWR VPWR _3957_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3460_ input49/X _4058_/S _5523_/A _7068_/Q VGND VGND VPWR VPWR _3460_/X sky130_fd_sc_hd__a22o_1
X_3391_ _6921_/Q _5355_/A _5274_/A _6849_/Q _3390_/X VGND VGND VPWR VPWR _3392_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5130_ _4691_/A _4631_/Y _4855_/Y _4895_/B _4518_/B VGND VGND VPWR VPWR _5131_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_123_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1508 _6586_/Q VGND VGND VPWR VPWR _4182_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5061_ _5061_/A1 _4229_/X _5022_/Y _5060_/X VGND VGND VPWR VPWR _6723_/D sky130_fd_sc_hd__a211o_1
XFILLER_96_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1519 _5778_/X VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4012_ hold507/X _5518_/A1 _4013_/S VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5963_ _5978_/A _5969_/A _5969_/C VGND VGND VPWR VPWR _5975_/C sky130_fd_sc_hd__and3_4
Xclkbuf_opt_4_0_csclk _6888_/CLK VGND VGND VPWR VPWR clkbuf_opt_4_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_52_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4914_ _5114_/B _5083_/B _5114_/C VGND VGND VPWR VPWR _4915_/D sky130_fd_sc_hd__and3_1
X_5894_ _6568_/Q _5635_/X _5654_/X _6678_/Q _5893_/X VGND VGND VPWR VPWR _5894_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4845_ _4907_/B _5042_/B _4644_/B _4911_/B VGND VGND VPWR VPWR _4845_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4776_ _5088_/A _5114_/A _4776_/C VGND VGND VPWR VPWR _4776_/X sky130_fd_sc_hd__and3_1
XFILLER_165_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6515_ _6890_/CLK _6515_/D fanout476/X VGND VGND VPWR VPWR _6515_/Q sky130_fd_sc_hd__dfrtp_1
X_3727_ _7040_/Q hold76/A _6352_/A _7152_/Q VGND VGND VPWR VPWR _3727_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6446_ _7081_/CLK hold80/X fanout478/X VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__dfrtp_2
X_3658_ _6796_/Q _3326_/Y _5154_/A _6744_/Q _3657_/X VGND VGND VPWR VPWR _3661_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_161_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6377_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6377_/X sky130_fd_sc_hd__and2_1
X_3589_ _7058_/Q hold86/A _4274_/A _6673_/Q VGND VGND VPWR VPWR _3589_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5328_ _5328_/A _5541_/B VGND VGND VPWR VPWR _5336_/S sky130_fd_sc_hd__and2_4
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5259_ hold844/X _5484_/A1 _5264_/S VGND VGND VPWR VPWR _5259_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4630_ _4633_/B _4716_/A _4653_/C _4631_/D VGND VGND VPWR VPWR _4630_/X sky130_fd_sc_hd__and4b_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4561_ _4690_/A _4561_/B VGND VGND VPWR VPWR _5043_/A sky130_fd_sc_hd__nor2_4
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6300_ _6300_/A _6300_/B _6300_/C _6300_/D VGND VGND VPWR VPWR _6301_/B sky130_fd_sc_hd__nor4_1
X_3512_ _3546_/A _3573_/A VGND VGND VPWR VPWR _4020_/A sky130_fd_sc_hd__nor2_4
Xhold605 _5240_/X VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _6459_/Q VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4492_ _4739_/A _4911_/A _4896_/A _4492_/D VGND VGND VPWR VPWR _4881_/B sky130_fd_sc_hd__and4b_4
Xhold627 _5471_/X VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _6647_/Q VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 _5460_/X VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _6611_/Q _5943_/X _5981_/X _6657_/Q VGND VGND VPWR VPWR _6231_/X sky130_fd_sc_hd__a22o_1
X_3443_ input41/X _5202_/B _5274_/A _6848_/Q _3442_/X VGND VGND VPWR VPWR _3446_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap368 _5391_/A VGND VGND VPWR VPWR _3781_/A2 sky130_fd_sc_hd__buf_8
XFILLER_143_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6897_/Q _5946_/X _5955_/X _6809_/Q VGND VGND VPWR VPWR _6162_/X sky130_fd_sc_hd__a22o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3374_ _3374_/A hold85/X VGND VGND VPWR VPWR _5301_/A sky130_fd_sc_hd__nor2_8
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A1 _4229_/X _5109_/Y _5112_/X VGND VGND VPWR VPWR _5113_/X sky130_fd_sc_hd__a22o_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6093_ _7051_/Q _5971_/A _5979_/X _6990_/Q VGND VGND VPWR VPWR _6093_/X sky130_fd_sc_hd__a22o_1
Xhold1305 _6518_/Q VGND VGND VPWR VPWR _4103_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 hold1316/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1327 hold1424/X VGND VGND VPWR VPWR hold1327/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _4948_/C _5042_/Y _5043_/Y _4948_/B VGND VGND VPWR VPWR _5058_/A sky130_fd_sc_hd__o22a_1
XFILLER_38_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1338 hold1338/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1349 _6311_/A1 VGND VGND VPWR VPWR hold1349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6995_ _7017_/CLK _6995_/D fanout458/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5946_ _5979_/A _5964_/A _5969_/C VGND VGND VPWR VPWR _5946_/X sky130_fd_sc_hd__and3_4
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5877_ _6616_/Q _5628_/X _5910_/B1 _6627_/Q VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4828_ _4948_/B _4562_/Y _4827_/X _5027_/A VGND VGND VPWR VPWR _4828_/X sky130_fd_sc_hd__o211a_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4759_ _4542_/A _4672_/B _4626_/Y _4689_/B VGND VGND VPWR VPWR _4999_/A sky130_fd_sc_hd__o22a_1
XFILLER_153_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6429_ _7155_/CLK _6429_/D fanout449/X VGND VGND VPWR VPWR _6429_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 hold5/X VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__buf_8
XFILLER_181_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5800_ _5799_/Y _5798_/X _6279_/S _5820_/A2 VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6780_ _6969_/CLK _6780_/D fanout473/X VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfrtp_1
X_3992_ hold804/X _6354_/A1 _3998_/S VGND VGND VPWR VPWR _3992_/X sky130_fd_sc_hd__mux2_1
X_5731_ _6797_/Q _5905_/A2 _5715_/X _5730_/X VGND VGND VPWR VPWR _5731_/X sky130_fd_sc_hd__a211o_1
XFILLER_31_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5662_ _6802_/Q _5913_/B1 _5661_/X _6874_/Q _5659_/X VGND VGND VPWR VPWR _5669_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4613_ _4716_/A _4636_/A VGND VGND VPWR VPWR _4613_/Y sky130_fd_sc_hd__nand2_4
X_5593_ _7100_/Q _7099_/Q VGND VGND VPWR VPWR _5964_/A sky130_fd_sc_hd__and2_2
XFILLER_175_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4544_ _4948_/A _4413_/Y _4561_/B _4562_/A VGND VGND VPWR VPWR _4589_/B sky130_fd_sc_hd__a211o_1
Xhold402 _4121_/X VGND VGND VPWR VPWR _6534_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold413 _6626_/Q VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 _5192_/X VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _7067_/Q VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _5396_/X VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4984_/A _4710_/A VGND VGND VPWR VPWR _4650_/A sky130_fd_sc_hd__and2_1
XFILLER_144_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold457 _6692_/Q VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _5279_/X VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6214_ _6631_/Q _5946_/X _5955_/X _6551_/Q VGND VGND VPWR VPWR _6214_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3426_ _6832_/Q _5256_/A _3423_/X _3425_/X VGND VGND VPWR VPWR _3426_/X sky130_fd_sc_hd__a211o_1
Xhold479 _6894_/Q VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlygate4sd3_1
X_7194_ hold91/A VGND VGND VPWR VPWR _7194_/X sky130_fd_sc_hd__clkbuf_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _7069_/Q _5934_/X _5975_/B _6872_/Q _6144_/X VGND VGND VPWR VPWR _6145_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3357_ hold65/X _3454_/A VGND VGND VPWR VPWR _3573_/B sky130_fd_sc_hd__nand2_8
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _5305_/X VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1113 _7187_/A VGND VGND VPWR VPWR _4065_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6789_/Q _6226_/B _6075_/X VGND VGND VPWR VPWR _6076_/X sky130_fd_sc_hd__o21ba_1
Xhold1124 _4241_/X VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 _6799_/Q VGND VGND VPWR VPWR _5226_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3288_ _6488_/Q _6414_/Q VGND VGND VPWR VPWR _3288_/Y sky130_fd_sc_hd__nand2b_1
Xhold1146 _4091_/X VGND VGND VPWR VPWR _6512_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5027_ _5027_/A _5027_/B _5027_/C VGND VGND VPWR VPWR _5080_/B sky130_fd_sc_hd__and3_1
Xhold1157 _6874_/Q VGND VGND VPWR VPWR _5311_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _4140_/X VGND VGND VPWR VPWR _6550_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 _6858_/Q VGND VGND VPWR VPWR _5293_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6978_ _7012_/CLK _6978_/D fanout458/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfstp_1
X_5929_ _6544_/Q _5652_/Y _5920_/X _5928_/X _6303_/S VGND VGND VPWR VPWR _5929_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold980 _7153_/Q VGND VGND VPWR VPWR hold980/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 _5182_/X VGND VGND VPWR VPWR _5183_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4260_ hold499/X _5518_/A1 _4261_/S VGND VGND VPWR VPWR _4260_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3211_ _6885_/Q VGND VGND VPWR VPWR _3211_/Y sky130_fd_sc_hd__inv_2
X_4191_ _3640_/Y _4191_/A1 _4195_/S VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6901_ _7076_/CLK _6901_/D fanout481/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6832_ _6951_/CLK _6832_/D fanout474/X VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6763_ _6953_/CLK _6763_/D fanout460/X VGND VGND VPWR VPWR _6763_/Q sky130_fd_sc_hd__dfrtp_1
X_3975_ hold40/X hold52/X _3975_/S VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__mux2_1
X_5714_ _5735_/A2 _5713_/X _6279_/S VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__mux2_1
X_6694_ _6714_/CLK _6694_/D fanout470/X VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5645_ _5664_/A _5666_/B _5660_/C VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__and3_4
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5576_ _7094_/Q _5576_/B VGND VGND VPWR VPWR _5576_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold210 _5177_/X VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _6957_/Q VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4527_ _4542_/B _4453_/B _4525_/X _5084_/B VGND VGND VPWR VPWR _4527_/X sky130_fd_sc_hd__o211a_1
Xhold232 _5431_/X VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold254 _5456_/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _6711_/Q VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _5465_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4458_ _4551_/A _4813_/A _4459_/B VGND VGND VPWR VPWR _4953_/A sky130_fd_sc_hd__and3_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold287 _6819_/Q VGND VGND VPWR VPWR hold287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold298 _5267_/X VGND VGND VPWR VPWR _6835_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _3409_/A _3409_/B wire357/X VGND VGND VPWR VPWR _3410_/B sky130_fd_sc_hd__nor3b_1
XFILLER_132_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7177_ _7177_/A VGND VGND VPWR VPWR _7177_/X sky130_fd_sc_hd__clkbuf_1
X_4389_ _4631_/D _4661_/A _4441_/B VGND VGND VPWR VPWR _4389_/Y sky130_fd_sc_hd__nand3_1
X_6128_ _6128_/A0 _6127_/X _6303_/S VGND VGND VPWR VPWR _6128_/X sky130_fd_sc_hd__mux2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6059_ _7058_/Q _5954_/X _5976_/D _6877_/Q _6058_/X VGND VGND VPWR VPWR _6074_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 _3251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _6440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_149 _5494_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3760_ _3760_/A _3760_/B _3760_/C _3760_/D VGND VGND VPWR VPWR _3761_/D sky130_fd_sc_hd__nor4_1
XFILLER_9_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3691_ _7004_/Q _3370_/Y _4038_/A _6477_/Q VGND VGND VPWR VPWR _3691_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5430_ hold357/X _5526_/A1 _5435_/S VGND VGND VPWR VPWR _5430_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput304 _3450_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
X_5361_ hold708/X _5469_/A1 _5363_/S VGND VGND VPWR VPWR _5361_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput315 hold1325/X VGND VGND VPWR VPWR hold1326/A sky130_fd_sc_hd__buf_12
XFILLER_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput326 hold1359/X VGND VGND VPWR VPWR hold1360/A sky130_fd_sc_hd__buf_12
Xoutput337 hold1327/X VGND VGND VPWR VPWR hold1328/A sky130_fd_sc_hd__buf_12
XFILLER_160_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4312_ hold834/X _6354_/A1 _4315_/S VGND VGND VPWR VPWR _4312_/X sky130_fd_sc_hd__mux2_1
X_7100_ _7113_/CLK _7100_/D fanout464/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5292_ _5292_/A _5505_/B VGND VGND VPWR VPWR _5300_/S sky130_fd_sc_hd__and2_4
XFILLER_114_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7031_ _7086_/CLK hold51/X fanout484/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4243_ hold974/X _5546_/A1 _4243_/S VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4174_ _4174_/A0 _5492_/A1 _4177_/S VGND VGND VPWR VPWR _4174_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6815_ _6969_/CLK _6815_/D fanout473/X VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6746_ _6746_/CLK _6746_/D fanout447/X VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfstp_4
X_3958_ _3958_/A input1/X VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__and2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3889_ _7097_/Q _7098_/Q VGND VGND VPWR VPWR _5978_/A sky130_fd_sc_hd__and2b_4
X_6677_ _6677_/CLK _6677_/D fanout450/X VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_109_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5628_ _5638_/A _5660_/C _5663_/C VGND VGND VPWR VPWR _5628_/X sky130_fd_sc_hd__and3b_4
XFILLER_191_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5559_ _7088_/Q _7089_/Q VGND VGND VPWR VPWR _5604_/B sky130_fd_sc_hd__nand2_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_27_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ _4482_/B _4562_/Y _4741_/A _5099_/B _4758_/X VGND VGND VPWR VPWR _4930_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_18_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4861_ _4465_/B _4845_/X _4847_/A VGND VGND VPWR VPWR _4869_/C sky130_fd_sc_hd__a21oi_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6600_ _7036_/CLK _6600_/D fanout455/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfrtp_4
X_3812_ _7173_/A _3320_/X _3355_/X _4268_/A _6665_/Q VGND VGND VPWR VPWR _3812_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_16 _3571_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4792_ _4576_/B _4703_/B _4689_/Y VGND VGND VPWR VPWR _4796_/A sky130_fd_sc_hd__a21oi_2
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 _4304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_38 _4108_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3743_ _6819_/Q _5247_/A _4032_/A _6471_/Q VGND VGND VPWR VPWR _3743_/X sky130_fd_sc_hd__a22o_1
XANTENNA_49 _5643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ _6990_/CLK hold39/X fanout479/X VGND VGND VPWR VPWR _6531_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3674_ input22/X _3367_/Y _4310_/A _6702_/Q _3673_/X VGND VGND VPWR VPWR _3679_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6462_ _6668_/CLK _6462_/D _6400_/A VGND VGND VPWR VPWR _6462_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5413_ _5413_/A0 _5545_/A1 _5417_/S VGND VGND VPWR VPWR _5413_/X sky130_fd_sc_hd__mux2_1
X_6393_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6393_/X sky130_fd_sc_hd__and2_1
X_5344_ hold932/X _5548_/A1 _5345_/S VGND VGND VPWR VPWR _5344_/X sky130_fd_sc_hd__mux2_1
Xoutput178 _3211_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
X_5275_ _5275_/A0 hold666/X _5282_/S VGND VGND VPWR VPWR _5275_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput189 _3201_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7014_ _7049_/CLK _7014_/D fanout457/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfrtp_4
X_4226_ _6643_/Q _6642_/Q _6644_/Q VGND VGND VPWR VPWR _4230_/B sky130_fd_sc_hd__nor3_4
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4157_ _4157_/A _6352_/B VGND VGND VPWR VPWR _4162_/S sky130_fd_sc_hd__and2_2
XFILLER_95_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4088_ hold257/X _5534_/A1 _5202_/B VGND VGND VPWR VPWR _4088_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6729_ _3945_/A1 _6729_/D _6381_/X VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_csclk _7001_/CLK VGND VGND VPWR VPWR _6537_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout394 hold174/X VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__buf_6
XFILLER_47_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _3958_/A sky130_fd_sc_hd__buf_6
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_2
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _3251_/A sky130_fd_sc_hd__buf_12
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold809 _4129_/X VGND VGND VPWR VPWR _6541_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3390_ _6873_/Q _5301_/A _5541_/A _7086_/Q VGND VGND VPWR VPWR _3390_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5060_ _5069_/A _5004_/Y _5038_/X _5059_/X VGND VGND VPWR VPWR _5060_/X sky130_fd_sc_hd__a211o_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 _7106_/Q VGND VGND VPWR VPWR _5672_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4011_ _4011_/A0 _6355_/A1 _4013_/S VGND VGND VPWR VPWR _4011_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5962_ _5978_/A _5969_/C _5979_/C VGND VGND VPWR VPWR _5975_/B sky130_fd_sc_hd__and3_4
X_4913_ _5051_/A _4782_/A _4881_/B VGND VGND VPWR VPWR _5114_/C sky130_fd_sc_hd__o21ai_1
X_5893_ _7037_/Q _5614_/X _5630_/X _6478_/Q VGND VGND VPWR VPWR _5893_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4844_ _4686_/Y _5041_/C _4887_/A VGND VGND VPWR VPWR _4869_/B sky130_fd_sc_hd__a21o_1
XFILLER_178_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4775_ _4912_/A _4775_/B _5074_/A _4775_/D VGND VGND VPWR VPWR _4776_/C sky130_fd_sc_hd__and4_1
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6514_ _6969_/CLK _6514_/D fanout473/X VGND VGND VPWR VPWR _7180_/A sky130_fd_sc_hd__dfrtp_1
X_3726_ _6971_/Q _5418_/A _3585_/Y input96/X _3725_/X VGND VGND VPWR VPWR _3729_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6445_ _7082_/CLK _6445_/D fanout483/X VGND VGND VPWR VPWR _6445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3657_ _7153_/Q _6352_/A _4014_/A _6457_/Q VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6376_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6376_/X sky130_fd_sc_hd__and2_1
X_3588_ _6813_/Q _5238_/A _4157_/A _6568_/Q VGND VGND VPWR VPWR _3588_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5327_ hold681/X _5540_/A1 _5327_/S VGND VGND VPWR VPWR _5327_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5258_ hold285/X _5534_/A1 _5264_/S VGND VGND VPWR VPWR _5258_/X sky130_fd_sc_hd__mux2_1
X_4209_ _4209_/A0 _6353_/A1 _4213_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5189_ _5189_/A0 hold667/X _5189_/S VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4560_ _4563_/A _4631_/D _4563_/D VGND VGND VPWR VPWR _4595_/A sky130_fd_sc_hd__nand3_1
XFILLER_175_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3511_ _3511_/A _3571_/B VGND VGND VPWR VPWR _3511_/Y sky130_fd_sc_hd__nor2_1
Xhold606 _6865_/Q VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ _4739_/A _4492_/D VGND VGND VPWR VPWR _4491_/Y sky130_fd_sc_hd__nand2b_1
Xhold617 _4019_/X VGND VGND VPWR VPWR _6459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _6877_/Q VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 _4247_/X VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3442_ _6888_/Q _5319_/A _5301_/A _6872_/Q VGND VGND VPWR VPWR _3442_/X sky130_fd_sc_hd__a22o_1
X_6230_ _6662_/Q _5976_/B _5971_/C _6712_/Q VGND VGND VPWR VPWR _6230_/X sky130_fd_sc_hd__a22o_1
Xmax_cap369 _3814_/A VGND VGND VPWR VPWR _3455_/A sky130_fd_sc_hd__buf_12
XFILLER_170_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6161_ _6945_/Q _5961_/X _6159_/X _6160_/X VGND VGND VPWR VPWR _6165_/A sky130_fd_sc_hd__a211o_1
XFILLER_97_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3373_ _3374_/A _3373_/B VGND VGND VPWR VPWR _5319_/A sky130_fd_sc_hd__nor2_8
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5112_ _5112_/A _5112_/B _5112_/C _5112_/D VGND VGND VPWR VPWR _5112_/X sky130_fd_sc_hd__and4_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6822_/Q _5953_/X _5960_/X _7075_/Q _6091_/X VGND VGND VPWR VPWR _6092_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 _4103_/X VGND VGND VPWR VPWR _6518_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A _5043_/B VGND VGND VPWR VPWR _5043_/Y sky130_fd_sc_hd__nor2_1
Xhold1317 hold1413/X VGND VGND VPWR VPWR hold1317/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 hold1328/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
Xhold1339 hold1423/X VGND VGND VPWR VPWR hold1339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wbbd_sck _7149_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6994_ _7012_/CLK _6994_/D fanout458/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5945_ _5981_/A _5981_/C _5979_/C VGND VGND VPWR VPWR _5945_/X sky130_fd_sc_hd__and3_4
XFILLER_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5876_ _6462_/Q _5624_/X _5654_/X _6677_/Q _5866_/Y VGND VGND VPWR VPWR _5876_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4827_ _4948_/C _4810_/B _4825_/Y _4826_/X _4574_/Y VGND VGND VPWR VPWR _4827_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_138_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4758_ _4607_/A _4413_/Y _4947_/A _4611_/Y _4616_/Y VGND VGND VPWR VPWR _4758_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3709_ _3709_/A _3709_/B _3709_/C VGND VGND VPWR VPWR _3730_/A sky130_fd_sc_hd__nor3_1
X_4689_ _4689_/A _4689_/B VGND VGND VPWR VPWR _4689_/Y sky130_fd_sc_hd__nor2_4
XFILLER_161_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6428_ _7155_/CLK _6428_/D fanout449/X VGND VGND VPWR VPWR _6428_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_161_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6359_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6359_/X sky130_fd_sc_hd__and2_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3991_ _3991_/A0 _5491_/A1 _3998_/S VGND VGND VPWR VPWR _3991_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5730_ _6989_/Q _5627_/X _5635_/X _6829_/Q VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5661_ _5638_/A _5667_/B _5663_/C VGND VGND VPWR VPWR _5661_/X sky130_fd_sc_hd__and3b_4
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4612_ _4975_/A _5010_/B VGND VGND VPWR VPWR _4612_/Y sky130_fd_sc_hd__nor2_1
X_5592_ _5592_/A1 _5594_/A _5591_/Y VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__a21oi_1
XFILLER_191_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4543_ _4948_/C _4456_/Y _4542_/X _4561_/B VGND VGND VPWR VPWR _4589_/A sky130_fd_sc_hd__a31o_1
XFILLER_128_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold403 _7052_/Q VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold414 _4234_/X VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold425 _6631_/Q VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold436 _5528_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4474_ _4615_/B _4638_/A VGND VGND VPWR VPWR _4710_/A sky130_fd_sc_hd__and2_1
Xhold447 _6613_/Q VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold458 _4301_/X VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _6686_/Q _5961_/X _6207_/X _6212_/X VGND VGND VPWR VPWR _6218_/A sky130_fd_sc_hd__a211o_1
Xhold469 _6967_/Q VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3425_ input50/X _4058_/S _5211_/A _6792_/Q _3424_/X VGND VGND VPWR VPWR _3425_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7193_ _7193_/A VGND VGND VPWR VPWR _7193_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3356_/A _3356_/B VGND VGND VPWR VPWR _3511_/A sky130_fd_sc_hd__nand2_8
X_6144_ _7053_/Q _5971_/A _5979_/X _6992_/Q VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__a22o_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1103 _7066_/Q VGND VGND VPWR VPWR _5527_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _4065_/X VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3975_/S hold101/X _3285_/X VGND VGND VPWR VPWR _3287_/Y sky130_fd_sc_hd__a21oi_4
X_6075_ _6069_/X _6301_/C _6075_/C _6075_/D VGND VGND VPWR VPWR _6075_/X sky130_fd_sc_hd__and4b_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _6452_/Q VGND VGND VPWR VPWR _4011_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1136 _5226_/X VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 _6914_/Q VGND VGND VPWR VPWR _5356_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5026_ _4638_/Y _4695_/Y _4915_/B VGND VGND VPWR VPWR _5027_/C sky130_fd_sc_hd__o21a_1
Xhold1158 _5311_/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 hold1593/X VGND VGND VPWR VPWR _4070_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7033_/CLK _6977_/D fanout464/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5928_ _6582_/Q _5928_/A2 _5923_/X _5927_/X VGND VGND VPWR VPWR _5928_/X sky130_fd_sc_hd__a211o_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5859_ _6686_/Q _5632_/X _5642_/X _6716_/Q _5858_/X VGND VGND VPWR VPWR _5862_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold970 _6659_/Q VGND VGND VPWR VPWR hold970/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 _6355_/X VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold992 _5183_/X VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3210_ _6893_/Q VGND VGND VPWR VPWR _3210_/Y sky130_fd_sc_hd__inv_2
X_4190_ _3700_/Y _4190_/A1 _4195_/S VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6900_ _6990_/CLK _6900_/D fanout479/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6831_ _6951_/CLK _6831_/D fanout474/X VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6762_ _6953_/CLK _6762_/D fanout460/X VGND VGND VPWR VPWR _6762_/Q sky130_fd_sc_hd__dfrtp_4
X_3974_ hold640/X _6357_/A1 _3980_/S VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__mux2_1
X_5713_ _5713_/A0 _5712_/X _6303_/S VGND VGND VPWR VPWR _5713_/X sky130_fd_sc_hd__mux2_1
X_6693_ _6714_/CLK _6693_/D fanout470/X VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5644_ _6962_/Q _5642_/X _5643_/X _6994_/Q VGND VGND VPWR VPWR _5644_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5575_ _5610_/B _5658_/B _5667_/B _5575_/B1 _5568_/Y VGND VGND VPWR VPWR _7093_/D
+ sky130_fd_sc_hd__o32a_1
Xhold200 _6797_/Q VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold211 _6754_/Q VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4526_ _4542_/B _4531_/B VGND VGND VPWR VPWR _5084_/B sky130_fd_sc_hd__nand2b_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold222 _5404_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _6569_/Q VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _4122_/X VGND VGND VPWR VPWR _6535_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold255 _6762_/Q VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _4459_/A _4724_/A _4579_/B VGND VGND VPWR VPWR _4508_/C sky130_fd_sc_hd__nand3_1
Xhold266 _4324_/X VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold277 _6691_/Q VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold288 _5249_/X VGND VGND VPWR VPWR _6819_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _6979_/Q VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3408_ _3408_/A _3408_/B _3408_/C _3408_/D VGND VGND VPWR VPWR _3408_/Y sky130_fd_sc_hd__nor4_1
X_7176_ _7176_/A VGND VGND VPWR VPWR _7176_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4388_ _4642_/A _4441_/B VGND VGND VPWR VPWR _4396_/A sky130_fd_sc_hd__and2_1
XFILLER_98_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6127_ _6791_/Q _6226_/B _6126_/X VGND VGND VPWR VPWR _6127_/X sky130_fd_sc_hd__o21ba_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ hold36/X _3692_/A VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__nor2_8
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6058_ _7082_/Q _5976_/B _5971_/C _7042_/Q VGND VGND VPWR VPWR _6058_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _4625_/B _4702_/Y _4981_/A VGND VGND VPWR VPWR _5112_/C sky130_fd_sc_hd__o21a_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 input45/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _3581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3690_ _7065_/Q _5523_/A _3365_/Y input5/X _3689_/X VGND VGND VPWR VPWR _3698_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput305 _3417_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
X_5360_ hold473/X _5528_/A1 _5363_/S VGND VGND VPWR VPWR _5360_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput316 hold1333/X VGND VGND VPWR VPWR hold1334/A sky130_fd_sc_hd__buf_12
Xoutput327 hold1323/X VGND VGND VPWR VPWR hold1324/A sky130_fd_sc_hd__buf_12
X_4311_ _4311_/A0 _6353_/A1 _4315_/S VGND VGND VPWR VPWR _4311_/X sky130_fd_sc_hd__mux2_1
Xoutput338 hold1355/X VGND VGND VPWR VPWR hold1356/A sky130_fd_sc_hd__buf_12
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5291_ hold327/X _5540_/A1 _5291_/S VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7030_ _7080_/CLK _7030_/D fanout478/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0__f__1177_ clkbuf_0__1177_/X VGND VGND VPWR VPWR _4192_/A0 sky130_fd_sc_hd__clkbuf_16
X_4242_ hold509/X _5518_/A1 _4243_/S VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4173_ hold999/X hold666/X _4177_/S VGND VGND VPWR VPWR _4173_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6814_ _7058_/CLK _6814_/D fanout480/X VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6745_ _6746_/CLK _6745_/D fanout447/X VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfrtp_4
X_3957_ _3957_/A _3957_/B VGND VGND VPWR VPWR _3957_/X sky130_fd_sc_hd__and2_1
X_6676_ _7036_/CLK _6676_/D fanout455/X VGND VGND VPWR VPWR _6676_/Q sky130_fd_sc_hd__dfrtp_1
X_3888_ _6303_/S _3887_/Y _5610_/B VGND VGND VPWR VPWR _6507_/D sky130_fd_sc_hd__o21ai_1
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5627_ _5638_/A _5666_/C _5663_/C VGND VGND VPWR VPWR _5627_/X sky130_fd_sc_hd__and3_4
X_5558_ _5555_/Y _5564_/A _5558_/C VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__and3b_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4509_ _4947_/B _4948_/C _4456_/Y _4496_/Y VGND VGND VPWR VPWR _4509_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5489_ hold690/X _5513_/A1 hold50/X VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7159_ _3927_/A1 _7159_/D _6389_/X VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4860_ _4685_/A _5042_/B _4504_/X VGND VGND VPWR VPWR _5023_/D sky130_fd_sc_hd__a21oi_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ _3958_/A _4118_/B _4250_/A _6650_/Q _3810_/X VGND VGND VPWR VPWR _3817_/B
+ sky130_fd_sc_hd__a221o_1
X_4791_ _4791_/A _4791_/B _5106_/A _4791_/D VGND VGND VPWR VPWR _4791_/X sky130_fd_sc_hd__and4_1
XANTENNA_17 _5154_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _3585_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_39 _5291_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _6990_/CLK _6530_/D fanout479/X VGND VGND VPWR VPWR _6530_/Q sky130_fd_sc_hd__dfrtp_1
X_3742_ _3742_/A _3742_/B _3742_/C _3742_/D VGND VGND VPWR VPWR _3761_/B sky130_fd_sc_hd__nor4_1
XFILLER_146_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6461_ _6668_/CLK _6461_/D _6400_/A VGND VGND VPWR VPWR _6461_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3673_ _6452_/Q _4008_/A _4304_/A _6697_/Q VGND VGND VPWR VPWR _3673_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5412_ hold321/X _5526_/A1 _5417_/S VGND VGND VPWR VPWR _5412_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6392_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6392_/X sky130_fd_sc_hd__and2_1
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5343_ hold429/X _5538_/A1 _5345_/S VGND VGND VPWR VPWR _5343_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput179 _3210_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
X_5274_ _5274_/A _5541_/B VGND VGND VPWR VPWR _5282_/S sky130_fd_sc_hd__and2_4
X_7013_ _7082_/CLK _7013_/D fanout480/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfrtp_4
X_4225_ hold820/X _5546_/A1 _4225_/S VGND VGND VPWR VPWR _4225_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4156_ hold946/X _5546_/A1 _4156_/S VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4087_ _4087_/A0 _4086_/X _4101_/S VGND VGND VPWR VPWR _4087_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4989_ _4542_/A _4428_/Y _4846_/B _4628_/Y VGND VGND VPWR VPWR _4999_/C sky130_fd_sc_hd__o22a_1
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6728_ _3945_/A1 _6728_/D _6380_/X VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6659_ _6659_/CLK _6659_/D fanout468/X VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout395 _5521_/A1 VGND VGND VPWR VPWR _5548_/A1 sky130_fd_sc_hd__buf_6
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4010_ _4010_/A0 _5492_/A1 _4013_/S VGND VGND VPWR VPWR _4010_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5961_ _5968_/A _5981_/A _5981_/B VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__and3_4
XFILLER_80_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4912_ _4912_/A _5073_/A _4912_/C VGND VGND VPWR VPWR _5083_/B sky130_fd_sc_hd__and3_1
XFILLER_33_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5892_ _6483_/Q _5643_/X _5910_/B1 _6628_/Q VGND VGND VPWR VPWR _5892_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4843_ _4959_/A _4843_/B VGND VGND VPWR VPWR _5041_/C sky130_fd_sc_hd__nand2_1
XFILLER_33_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4774_ _5002_/A _4774_/B _4774_/C _5002_/B VGND VGND VPWR VPWR _4775_/D sky130_fd_sc_hd__and4_1
XFILLER_165_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6513_ _6969_/CLK _6513_/D fanout473/X VGND VGND VPWR VPWR _7179_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3725_ _6716_/Q _4328_/A _4322_/A _6711_/Q VGND VGND VPWR VPWR _3725_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6444_ _7081_/CLK _6444_/D fanout479/X VGND VGND VPWR VPWR _6444_/Q sky130_fd_sc_hd__dfrtp_2
X_3656_ _6828_/Q _5256_/A _3654_/Y _3655_/X VGND VGND VPWR VPWR _3661_/B sky130_fd_sc_hd__a211o_1
XFILLER_174_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6375_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__and2_1
X_3587_ _6997_/Q _5445_/A hold67/A _6468_/Q VGND VGND VPWR VPWR _3587_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5326_ _5326_/A0 _5548_/A1 _5327_/S VGND VGND VPWR VPWR _5326_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5257_ _5257_/A0 _5473_/A1 _5264_/S VGND VGND VPWR VPWR _5257_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4208_ _4208_/A _4322_/B VGND VGND VPWR VPWR _4213_/S sky130_fd_sc_hd__and2_2
XFILLER_180_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5188_ hold279/X _5534_/A1 _5189_/S VGND VGND VPWR VPWR _5188_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4139_ _4139_/A _4322_/B VGND VGND VPWR VPWR _4144_/S sky130_fd_sc_hd__and2_2
XFILLER_56_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3510_ _3555_/A _3577_/B VGND VGND VPWR VPWR _4244_/A sky130_fd_sc_hd__nor2_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4490_ _4689_/A _4490_/B VGND VGND VPWR VPWR _4490_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold607 _5300_/X VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _6899_/Q VGND VGND VPWR VPWR hold618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 _5314_/X VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _6976_/Q _5418_/A _3326_/Y _6800_/Q _3440_/X VGND VGND VPWR VPWR _3446_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6160_ _7017_/Q _5940_/X _5967_/X _6857_/Q _6158_/X VGND VGND VPWR VPWR _6160_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3546_/A _3717_/B VGND VGND VPWR VPWR _3372_/Y sky130_fd_sc_hd__nor2_8
XFILLER_170_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5111_ _4482_/A _4625_/B _4615_/Y _4650_/Y _5110_/X VGND VGND VPWR VPWR _5112_/D
+ sky130_fd_sc_hd__o311a_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6910_/Q _5973_/A _5948_/X _6950_/Q _6090_/X VGND VGND VPWR VPWR _6091_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _6545_/Q VGND VGND VPWR VPWR _4134_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1318 hold1318/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
X_5042_ _5051_/A _5042_/B VGND VGND VPWR VPWR _5042_/Y sky130_fd_sc_hd__nor2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1329 hold1425/X VGND VGND VPWR VPWR hold1329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6993_ _7053_/CLK _6993_/D fanout459/X VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_csclk _7001_/CLK VGND VGND VPWR VPWR _6865_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5944_ _5978_/A _5964_/A _5981_/A VGND VGND VPWR VPWR _5944_/X sky130_fd_sc_hd__and3_4
X_5875_ _6557_/Q _5667_/X _5870_/X _5872_/X _5874_/X VGND VGND VPWR VPWR _5875_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4826_ _4902_/A _4810_/B _4948_/B VGND VGND VPWR VPWR _4826_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_66_csclk _6447_/CLK VGND VGND VPWR VPWR _7012_/CLK sky130_fd_sc_hd__clkbuf_16
X_4757_ _4581_/B _4542_/D _4611_/Y _4653_/Y VGND VGND VPWR VPWR _4770_/B sky130_fd_sc_hd__o22a_1
X_3708_ _6947_/Q _3781_/A2 _3964_/A _6419_/Q _3707_/X VGND VGND VPWR VPWR _3709_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4688_ _4689_/A _4619_/Y _4631_/Y _4902_/B _5108_/A VGND VGND VPWR VPWR _4722_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6427_ _6747_/CLK _6427_/D fanout449/X VGND VGND VPWR VPWR _6427_/Q sky130_fd_sc_hd__dfstp_2
X_3639_ _3639_/A _3639_/B _3639_/C VGND VGND VPWR VPWR _3640_/D sky130_fd_sc_hd__and3_2
XFILLER_162_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6358_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6358_/X sky130_fd_sc_hd__and2_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5309_ hold738/X _5540_/A1 _5309_/S VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__mux2_1
X_6289_ _6289_/A _6289_/B _6289_/C VGND VGND VPWR VPWR _6289_/Y sky130_fd_sc_hd__nor3_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6890_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xnet399_2 net399_2/A VGND VGND VPWR VPWR _3941_/B sky130_fd_sc_hd__inv_2
X_3990_ _3990_/A _6352_/B VGND VGND VPWR VPWR _3998_/S sky130_fd_sc_hd__and2_2
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5660_ _5664_/A _5667_/C _5660_/C VGND VGND VPWR VPWR _5660_/X sky130_fd_sc_hd__and3b_4
XFILLER_176_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4611_ _4753_/B _4611_/B VGND VGND VPWR VPWR _4611_/Y sky130_fd_sc_hd__nand2_8
X_5591_ _7099_/Q _5574_/Y _5594_/A VGND VGND VPWR VPWR _5591_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4542_ _4542_/A _4542_/B _4948_/B _4542_/D VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__and4_1
XFILLER_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold404 _5511_/X VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold415 _6646_/Q VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 _4240_/X VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4739_/A _4642_/A VGND VGND VPWR VPWR _4638_/A sky130_fd_sc_hd__and2b_1
XFILLER_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold437 _6974_/Q VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _4213_/X VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6476_/Q _5940_/X _5967_/X _6605_/Q _6206_/X VGND VGND VPWR VPWR _6212_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold459 _6854_/Q VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_3424_ _6856_/Q _5283_/A _3370_/Y _7008_/Q VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7192_ _7192_/A VGND VGND VPWR VPWR _7192_/X sky130_fd_sc_hd__clkbuf_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6824_/Q _5953_/X _5960_/X _7077_/Q _6142_/X VGND VGND VPWR VPWR _6143_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3355_ _3356_/A _3355_/B hold72/X VGND VGND VPWR VPWR _3355_/X sky130_fd_sc_hd__and3_4
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6074_ _6074_/A _6074_/B _6074_/C _6074_/D VGND VGND VPWR VPWR _6075_/D sky130_fd_sc_hd__nor4_1
Xhold1104 _5527_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3975_/S hold101/X hold204/X VGND VGND VPWR VPWR _3286_/X sky130_fd_sc_hd__a21o_4
Xhold1115 _7179_/A VGND VGND VPWR VPWR _4093_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _4011_/X VGND VGND VPWR VPWR _6452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 _7192_/A VGND VGND VPWR VPWR _5197_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5025_ _4413_/Y _4902_/A _4616_/Y _4691_/A _4877_/B VGND VGND VPWR VPWR _5118_/B
+ sky130_fd_sc_hd__o221a_1
Xhold1148 _5356_/X VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _7189_/A VGND VGND VPWR VPWR _5194_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6976_ _7082_/CLK _6976_/D fanout483/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5927_ _6689_/Q _5632_/X _5924_/X _5926_/X VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__a211o_1
XFILLER_179_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5858_ _6561_/Q _5631_/X _5667_/X _6556_/Q VGND VGND VPWR VPWR _5858_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4809_ _4992_/A _4886_/B VGND VGND VPWR VPWR _4810_/B sky130_fd_sc_hd__nor2_4
X_5789_ _7016_/Q _5630_/X _5658_/X _6888_/Q _5788_/X VGND VGND VPWR VPWR _5797_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold960 _6457_/Q VGND VGND VPWR VPWR hold960/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 _4261_/X VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold982 _6618_/Q VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _6428_/Q VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6830_ _6884_/CLK _6830_/D fanout475/X VGND VGND VPWR VPWR _6830_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6761_ _6953_/CLK _6761_/D fanout459/X VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3973_ hold58/X _3973_/A1 _3975_/S VGND VGND VPWR VPWR _3973_/X sky130_fd_sc_hd__mux2_4
XFILLER_50_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5712_ _5706_/Y _5711_/Y _6788_/Q _5652_/Y VGND VGND VPWR VPWR _5712_/X sky130_fd_sc_hd__o2bb2a_1
X_6692_ _6714_/CLK _6692_/D fanout470/X VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5643_ _5664_/A _5660_/C _5663_/C VGND VGND VPWR VPWR _5643_/X sky130_fd_sc_hd__and3_4
XFILLER_31_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5574_ _6506_/Q _5610_/B VGND VGND VPWR VPWR _5574_/Y sky130_fd_sc_hd__nand2_1
Xhold201 _5224_/X VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4525_ _4948_/A _4453_/B _4522_/X _5084_/A VGND VGND VPWR VPWR _4525_/X sky130_fd_sc_hd__o211a_1
Xhold212 _5170_/X VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _6837_/Q VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold234 _4162_/X VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _6923_/Q VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _5181_/X VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4456_ _4456_/A _4579_/B VGND VGND VPWR VPWR _4456_/Y sky130_fd_sc_hd__nand2_8
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold267 _6661_/Q VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _4300_/X VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _6795_/Q VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ _6913_/Q _5346_/A _5238_/A _6817_/Q _3406_/X VGND VGND VPWR VPWR _3408_/D
+ sky130_fd_sc_hd__a221o_1
X_7175_ _7175_/A VGND VGND VPWR VPWR _7175_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4387_ _4661_/A _4441_/B VGND VGND VPWR VPWR _4400_/B sky130_fd_sc_hd__nand2_2
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _6118_/X _6226_/B _6126_/C _6126_/D VGND VGND VPWR VPWR _6126_/X sky130_fd_sc_hd__and4b_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3338_ _3454_/B _3415_/B VGND VGND VPWR VPWR _3692_/A sky130_fd_sc_hd__nand2_8
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6057_ _6813_/Q _5971_/B _5949_/X _6933_/Q _6056_/X VGND VGND VPWR VPWR _6074_/A
+ sky130_fd_sc_hd__a221o_1
X_3269_ _6390_/A _6396_/B VGND VGND VPWR VPWR _3269_/X sky130_fd_sc_hd__and2_1
XFILLER_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5008_ _5008_/A _5008_/B _5008_/C _5008_/D VGND VGND VPWR VPWR _5112_/B sky130_fd_sc_hd__and4_1
XFILLER_39_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6959_ _6999_/CLK _6959_/D fanout465/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold790 _6831_/Q VGND VGND VPWR VPWR hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1490 _6078_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3927_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput306 _3940_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
Xoutput317 hold1353/X VGND VGND VPWR VPWR hold1354/A sky130_fd_sc_hd__buf_12
X_4310_ _4310_/A _6352_/B VGND VGND VPWR VPWR _4315_/S sky130_fd_sc_hd__and2_2
Xoutput328 hold1315/X VGND VGND VPWR VPWR hold1316/A sky130_fd_sc_hd__buf_12
X_5290_ hold141/X hold99/X _5291_/S VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__mux2_1
Xoutput339 hold1369/X VGND VGND VPWR VPWR hold1370/A sky130_fd_sc_hd__buf_12
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4241_ _4241_/A0 _5493_/A1 _4243_/S VGND VGND VPWR VPWR _4241_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ _4172_/A _5490_/B VGND VGND VPWR VPWR _4177_/S sky130_fd_sc_hd__and2_2
XFILLER_68_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6813_ _7076_/CLK _6813_/D fanout481/X VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3956_ _3956_/A _3956_/B VGND VGND VPWR VPWR _3956_/X sky130_fd_sc_hd__and2_1
X_6744_ _6746_/CLK _6744_/D _3946_/B VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6675_ _7036_/CLK _6675_/D fanout455/X VGND VGND VPWR VPWR _6675_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3887_ _5606_/A _3887_/B VGND VGND VPWR VPWR _3887_/Y sky130_fd_sc_hd__nor2_1
X_5626_ _6978_/Q _5624_/X _5625_/X _7002_/Q VGND VGND VPWR VPWR _5626_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5557_ _7088_/Q _5562_/D VGND VGND VPWR VPWR _5558_/C sky130_fd_sc_hd__nand2_1
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4508_ _4507_/X _5027_/A _4508_/C _4508_/D VGND VGND VPWR VPWR _4508_/X sky130_fd_sc_hd__and4b_1
XFILLER_117_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5488_ hold894/X _5548_/A1 hold50/X VGND VGND VPWR VPWR _5488_/X sky130_fd_sc_hd__mux2_1
X_4439_ _4615_/B _4635_/B VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__nand2_8
XFILLER_160_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7158_ _3927_/A1 _7158_/D _6388_/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6109_ _7015_/Q _5940_/X _5967_/X _6855_/Q _6107_/X VGND VGND VPWR VPWR _6109_/X
+ sky130_fd_sc_hd__a221o_1
X_7089_ _7113_/CLK _7089_/D fanout460/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3810_ input71/X _3331_/Y _4196_/A _6599_/Q VGND VGND VPWR VPWR _3810_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4790_ _4556_/A _4632_/B _4482_/A _4672_/A _4789_/X VGND VGND VPWR VPWR _4791_/D
+ sky130_fd_sc_hd__o41a_1
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _5164_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ input47/X _4118_/B _4310_/A _6701_/Q _3740_/X VGND VGND VPWR VPWR _3742_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_29 _5166_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6460_ _6668_/CLK _6460_/D _6400_/A VGND VGND VPWR VPWR _6460_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ _6547_/Q _4133_/A _5490_/A _7036_/Q _3671_/X VGND VGND VPWR VPWR _3679_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5411_ _5411_/A0 hold13/X _5417_/S VGND VGND VPWR VPWR _5411_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6391_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6391_/X sky130_fd_sc_hd__and2_1
X_5342_ hold184/X _5519_/A1 _5345_/S VGND VGND VPWR VPWR _5342_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5273_ hold632/X _5513_/A1 _5273_/S VGND VGND VPWR VPWR _5273_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7012_ _7012_/CLK _7012_/D fanout466/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4224_ hold309/X _5518_/A1 _4225_/S VGND VGND VPWR VPWR _4224_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4155_ hold463/X _5518_/A1 _4156_/S VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4086_ _5203_/A0 _5473_/A1 _5202_/B VGND VGND VPWR VPWR _4086_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4988_ _4919_/X _4945_/Y _4987_/X _5006_/A _4988_/B2 VGND VGND VPWR VPWR _6722_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_168_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6727_ _3568_/A1 _6727_/D _6379_/X VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfrtn_1
X_3939_ _7103_/Q _6759_/Q _6762_/Q VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6658_ _6659_/CLK _6658_/D fanout469/X VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_2
X_5609_ _5609_/A1 _5606_/B _5608_/X _3886_/B VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6589_ _7137_/CLK _6589_/D VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout396 hold99/X VGND VGND VPWR VPWR _5521_/A1 sky130_fd_sc_hd__buf_6
XFILLER_143_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5960_ _5969_/A _5966_/A _5981_/C VGND VGND VPWR VPWR _5960_/X sky130_fd_sc_hd__and3_4
XFILLER_80_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4911_ _4911_/A _4911_/B _4911_/C VGND VGND VPWR VPWR _4912_/C sky130_fd_sc_hd__nand3_1
X_5891_ _6473_/Q _5627_/X _5667_/X _6558_/Q _5890_/X VGND VGND VPWR VPWR _5896_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4842_ _4947_/B _4542_/D _4623_/Y _4694_/Y VGND VGND VPWR VPWR _4875_/A sky130_fd_sc_hd__o22a_1
XFILLER_193_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4773_ _4773_/A _4928_/A VGND VGND VPWR VPWR _5002_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6512_ _6969_/CLK _6512_/D fanout473/X VGND VGND VPWR VPWR _6512_/Q sky130_fd_sc_hd__dfrtp_1
X_3724_ input53/X _5193_/A _4145_/A _6556_/Q _3723_/X VGND VGND VPWR VPWR _3729_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6443_ _7017_/CLK _6443_/D fanout458/X VGND VGND VPWR VPWR _6443_/Q sky130_fd_sc_hd__dfstp_1
X_3655_ _6844_/Q _5274_/A _5166_/A _6753_/Q VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6374_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6374_/X sky130_fd_sc_hd__and2_1
X_3586_ _3586_/A _3814_/A VGND VGND VPWR VPWR _5166_/A sky130_fd_sc_hd__nor2_8
X_5325_ hold788/X _5538_/A1 _5327_/S VGND VGND VPWR VPWR _5325_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5256_ _5256_/A _5505_/B VGND VGND VPWR VPWR _5264_/S sky130_fd_sc_hd__and2_4
XFILLER_130_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4207_ hold529/X _6357_/A1 _4207_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5187_ hold441/X _5544_/A1 _5189_/S VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4138_ hold962/X _5546_/A1 _4138_/S VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4069_ _4119_/A0 _5491_/A1 _4118_/B VGND VGND VPWR VPWR _4069_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold608 _6544_/Q VGND VGND VPWR VPWR hold608/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3440_ _6992_/Q _5436_/A _5373_/A _6936_/Q VGND VGND VPWR VPWR _3440_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold619 _5339_/X VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3371_ _3586_/A _3717_/B VGND VGND VPWR VPWR _3981_/A sky130_fd_sc_hd__nor2_8
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _4483_/Y _4625_/B _4716_/Y _4484_/Y _5006_/A VGND VGND VPWR VPWR _5110_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ _6902_/Q _5976_/C _5971_/D _6830_/Q VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__a22o_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A _5041_/B _5041_/C VGND VGND VPWR VPWR _5041_/Y sky130_fd_sc_hd__nand3_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 _4134_/X VGND VGND VPWR VPWR _6545_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1319 hold1414/X VGND VGND VPWR VPWR hold1319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6992_ _7069_/CLK _6992_/D fanout482/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5943_ _5979_/A _5969_/C _5979_/C VGND VGND VPWR VPWR _5943_/X sky130_fd_sc_hd__and3_4
XFILLER_34_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5874_ _6482_/Q _5643_/X _5664_/X _6667_/Q _5873_/X VGND VGND VPWR VPWR _5874_/X
+ sky130_fd_sc_hd__a221o_1
X_4825_ _4551_/A _4815_/Y _4812_/Y VGND VGND VPWR VPWR _4825_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4756_ _4542_/B _4672_/B _4626_/Y _4645_/Y VGND VGND VPWR VPWR _4771_/C sky130_fd_sc_hd__o22a_1
X_3707_ _6851_/Q _5283_/A _5409_/A _6963_/Q VGND VGND VPWR VPWR _3707_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4687_ _4469_/A _4644_/Y _4663_/Y _4689_/A VGND VGND VPWR VPWR _5108_/A sky130_fd_sc_hd__o22a_1
XFILLER_162_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3638_ _3638_/A _3638_/B _3638_/C _3638_/D VGND VGND VPWR VPWR _3639_/C sky130_fd_sc_hd__nor4_1
X_6426_ _6747_/CLK _6426_/D fanout449/X VGND VGND VPWR VPWR _6426_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6357_ hold566/X _6357_/A1 _6357_/S VGND VGND VPWR VPWR _6357_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3569_ _3573_/A _3692_/A VGND VGND VPWR VPWR _4008_/A sky130_fd_sc_hd__nor2_8
XFILLER_161_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5308_ hold716/X _5521_/A1 _5309_/S VGND VGND VPWR VPWR _5308_/X sky130_fd_sc_hd__mux2_1
X_6288_ _6464_/Q _5945_/X _5975_/C _6582_/Q _6287_/X VGND VGND VPWR VPWR _6289_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5239_ _5239_/A0 hold667/X _5246_/S VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4610_ _4753_/B _4611_/B VGND VGND VPWR VPWR _5010_/B sky130_fd_sc_hd__and2_2
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5590_ _5610_/B _5978_/A _5979_/A _5568_/Y _5590_/B2 VGND VGND VPWR VPWR _7098_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_30_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4541_ _4661_/A _4724_/A _4959_/B _3962_/A VGND VGND VPWR VPWR _4541_/X sky130_fd_sc_hd__a31o_1
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold405 hold405/A VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire380 _4674_/Y VGND VGND VPWR VPWR wire380/X sky130_fd_sc_hd__clkbuf_1
Xhold416 _4246_/X VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4472_ _4472_/A _4489_/B VGND VGND VPWR VPWR _4472_/X sky130_fd_sc_hd__and2_1
Xhold427 _6656_/Q VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold438 _5423_/X VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _6864_/Q _5292_/A _5337_/A _6904_/Q VGND VGND VPWR VPWR _3423_/X sky130_fd_sc_hd__a22o_1
Xhold449 _6911_/Q VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_6211_ _6691_/Q _5954_/X _5976_/D _6620_/Q _6210_/X VGND VGND VPWR VPWR _6225_/B
+ sky130_fd_sc_hd__a221o_2
X_7191_ _7191_/A VGND VGND VPWR VPWR _7191_/X sky130_fd_sc_hd__clkbuf_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _6912_/Q _5973_/A _5948_/X _6952_/Q _6141_/X VGND VGND VPWR VPWR _6142_/X
+ sky130_fd_sc_hd__a221o_1
X_3354_ _3571_/A _3373_/B VGND VGND VPWR VPWR _5247_/A sky130_fd_sc_hd__nor2_8
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _7029_/Q _5944_/X _5975_/A _6845_/Q _6072_/X VGND VGND VPWR VPWR _6074_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3285_ _3975_/S _3285_/B VGND VGND VPWR VPWR _3285_/X sky130_fd_sc_hd__and2b_1
Xhold1105 _6917_/Q VGND VGND VPWR VPWR _5359_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1116 _4093_/X VGND VGND VPWR VPWR _6513_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _6552_/Q VGND VGND VPWR VPWR _4142_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5024_ _5051_/B _5024_/B VGND VGND VPWR VPWR _5086_/C sky130_fd_sc_hd__nand2_1
Xhold1138 _5197_/X VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 _6906_/Q VGND VGND VPWR VPWR _5347_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6975_ _7016_/CLK _6975_/D fanout474/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5926_ _6479_/Q _5630_/X _5638_/X _6709_/Q _5925_/X VGND VGND VPWR VPWR _5926_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5857_ _6651_/Q _5646_/X _5928_/A2 _6579_/Q _5856_/X VGND VGND VPWR VPWR _5862_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4808_ _5068_/B _4805_/X _4964_/A VGND VGND VPWR VPWR _4884_/C sky130_fd_sc_hd__a21bo_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5788_ _6448_/Q _5614_/X _5814_/B1 _6912_/Q VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4739_ _4739_/A _4739_/B VGND VGND VPWR VPWR _4740_/B sky130_fd_sc_hd__and2_1
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6409_ _3568_/A1 _6409_/D _6365_/X VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__dfrtp_1
Xhold950 _6744_/Q VGND VGND VPWR VPWR hold950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 _4017_/X VGND VGND VPWR VPWR _6457_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold972 _6702_/Q VGND VGND VPWR VPWR hold972/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold983 _4219_/X VGND VGND VPWR VPWR _6618_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 _3984_/X VGND VGND VPWR VPWR _6428_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_csclk _7001_/CLK VGND VGND VPWR VPWR _6999_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_csclk _6447_/CLK VGND VGND VPWR VPWR _7006_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6760_ _6953_/CLK _6760_/D fanout459/X VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfrtp_1
X_3972_ hold784/X _6356_/A1 _3980_/S VGND VGND VPWR VPWR _3972_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5711_ _5711_/A _5711_/B _5711_/C VGND VGND VPWR VPWR _5711_/Y sky130_fd_sc_hd__nor3_1
XFILLER_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6691_ _6712_/CLK _6691_/D fanout470/X VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5642_ _5664_/A _5657_/B _5660_/C VGND VGND VPWR VPWR _5642_/X sky130_fd_sc_hd__and3_4
XFILLER_31_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5573_ _6506_/Q _5610_/B VGND VGND VPWR VPWR _5602_/A sky130_fd_sc_hd__and2_1
XFILLER_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold202 _6488_/Q VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _4584_/A _4724_/A VGND VGND VPWR VPWR _5084_/A sky130_fd_sc_hd__nand2_1
Xhold213 _6464_/Q VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _5269_/X VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7083_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold235 _7038_/Q VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold246 _5366_/X VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4455_ _4498_/A _4579_/B VGND VGND VPWR VPWR _4948_/C sky130_fd_sc_hd__nand2_8
Xhold257 _6779_/Q VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold268 _4264_/X VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _6766_/Q VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _6881_/Q _5310_/A _5229_/A _6809_/Q VGND VGND VPWR VPWR _3406_/X sky130_fd_sc_hd__a22o_1
X_7174_ _7174_/A VGND VGND VPWR VPWR _7174_/X sky130_fd_sc_hd__clkbuf_1
X_4386_ _4661_/A _4441_/B VGND VGND VPWR VPWR _4563_/D sky130_fd_sc_hd__and2_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6125_ _6125_/A _6125_/B _6125_/C _6125_/D VGND VGND VPWR VPWR _6126_/D sky130_fd_sc_hd__nor4_1
X_3337_ _3453_/A hold64/X _3415_/B VGND VGND VPWR VPWR _5186_/A sky130_fd_sc_hd__and3_4
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3268_ _6764_/Q _6813_/Q _3268_/C VGND VGND VPWR VPWR _3268_/Y sky130_fd_sc_hd__nor3_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6056_ _6445_/Q _5601_/X _5959_/X _6965_/Q VGND VGND VPWR VPWR _6056_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5007_ _4576_/Y _4710_/Y _4482_/A VGND VGND VPWR VPWR _5008_/D sky130_fd_sc_hd__a21o_1
XFILLER_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3199_ _6981_/Q VGND VGND VPWR VPWR _3199_/Y sky130_fd_sc_hd__inv_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_108 input92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 _3899_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _7065_/CLK _6958_/D fanout465/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5909_ _5908_/Y _5907_/X _6279_/S _5909_/B2 VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__o2bb2a_1
X_6889_ _6969_/CLK _6889_/D fanout475/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold780 _6847_/Q VGND VGND VPWR VPWR hold780/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold791 _5262_/X VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1480 _6638_/Q VGND VGND VPWR VPWR _3880_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1491 _7121_/Q VGND VGND VPWR VPWR _6053_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput307 _3939_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
XFILLER_160_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput318 hold1343/X VGND VGND VPWR VPWR hold1344/A sky130_fd_sc_hd__buf_12
XFILLER_153_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput329 hold1317/X VGND VGND VPWR VPWR hold1318/A sky130_fd_sc_hd__buf_12
XFILLER_114_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ hold425/X _5534_/A1 _4243_/S VGND VGND VPWR VPWR _4240_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4171_ _3410_/Y _4171_/A1 _4171_/S VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6812_ _6990_/CLK _6812_/D fanout478/X VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6743_ _6746_/CLK _6743_/D _3946_/B VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfstp_2
X_3955_ _6643_/Q _3961_/B VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__and2_1
X_6674_ _6674_/CLK _6674_/D fanout468/X VGND VGND VPWR VPWR _6674_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_176_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3886_ _7088_/Q _3886_/B _7090_/Q _7091_/Q VGND VGND VPWR VPWR _3887_/B sky130_fd_sc_hd__nand4b_1
X_5625_ _5638_/A _5667_/B _5663_/C VGND VGND VPWR VPWR _5625_/X sky130_fd_sc_hd__and3_4
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5556_ _5552_/B _3887_/B _5554_/Y _6509_/Q VGND VGND VPWR VPWR _5564_/A sky130_fd_sc_hd__a211o_1
XFILLER_129_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4507_ _4782_/A _4493_/B _4472_/X _4502_/X _4450_/Y VGND VGND VPWR VPWR _4507_/X
+ sky130_fd_sc_hd__a2111o_1
X_5487_ _5487_/A0 hold42/X hold50/X VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__mux2_1
XFILLER_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4438_ _4615_/B _4635_/B VGND VGND VPWR VPWR _4965_/B sky130_fd_sc_hd__and2_4
XFILLER_59_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7157_ _7157_/CLK _7157_/D _3269_/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfstp_2
X_4369_ _4556_/A _4441_/A VGND VGND VPWR VPWR _4454_/A sky130_fd_sc_hd__and2_4
XFILLER_98_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6108_ _7007_/Q _5958_/X _5978_/X _6999_/Q VGND VGND VPWR VPWR _6108_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7113_/CLK _7088_/D fanout460/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6039_ _6980_/Q _5945_/X _5975_/C _6836_/Q _6038_/X VGND VGND VPWR VPWR _6040_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_19 _5164_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _6795_/Q _3326_/Y _4292_/A _6686_/Q VGND VGND VPWR VPWR _3740_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3671_ _6932_/Q _5373_/A _4274_/A _6672_/Q VGND VGND VPWR VPWR _3671_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5410_ _5410_/A0 _5524_/A1 _5417_/S VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6390_ _6390_/A _6396_/B VGND VGND VPWR VPWR _6390_/X sky130_fd_sc_hd__and2_1
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ _5341_/A0 _5545_/A1 _5345_/S VGND VGND VPWR VPWR _5341_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ hold135/X hold99/X _5273_/S VGND VGND VPWR VPWR _5272_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7011_ _7011_/CLK _7011_/D fanout456/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfstp_2
X_4223_ hold487/X _5544_/A1 _4225_/S VGND VGND VPWR VPWR _4223_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4154_ hold596/X _5544_/A1 _4156_/S VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4085_ _6367_/B _3379_/A _5202_/B _4050_/X _4322_/B VGND VGND VPWR VPWR _4101_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4987_ _5039_/A _5039_/C _4963_/Y _4986_/X VGND VGND VPWR VPWR _4987_/X sky130_fd_sc_hd__a31o_1
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6726_ _7140_/CLK _6726_/D _6307_/B VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3938_ _6515_/Q input93/X _6767_/Q VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__mux2_2
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6657_ _6659_/CLK _6657_/D fanout468/X VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_177_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3869_ _3911_/B1 _3869_/A2 _3832_/B _6405_/Q VGND VGND VPWR VPWR _6405_/D sky130_fd_sc_hd__a31o_1
XFILLER_164_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5608_ _7088_/Q _6509_/Q _5608_/C VGND VGND VPWR VPWR _5608_/X sky130_fd_sc_hd__and3_1
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6588_ _7137_/CLK _6588_/D VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ hold898/X _5548_/A1 _5540_/S VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout375 _6304_/S VGND VGND VPWR VPWR _6279_/S sky130_fd_sc_hd__buf_6
XFILLER_101_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout397 hold108/X VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__buf_12
XFILLER_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _3960_/B sky130_fd_sc_hd__buf_2
XFILLER_155_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4910_ _4691_/A _4482_/A _4672_/A _4964_/B _4909_/Y VGND VGND VPWR VPWR _4915_/C
+ sky130_fd_sc_hd__o311a_1
X_5890_ _6708_/Q _5638_/X _5928_/A2 _6581_/Q VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4841_ _4493_/B _4911_/B _4472_/X VGND VGND VPWR VPWR _4841_/X sky130_fd_sc_hd__a21o_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4772_ _4772_/A _5099_/C _4772_/C _4772_/D VGND VGND VPWR VPWR _4774_/C sky130_fd_sc_hd__and4_1
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6511_ _6969_/CLK _6511_/D fanout473/X VGND VGND VPWR VPWR _6511_/Q sky130_fd_sc_hd__dfrtp_1
X_3723_ _6769_/Q _5190_/A _5190_/B _4274_/A _6671_/Q VGND VGND VPWR VPWR _3723_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_158_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6442_ _6926_/CLK _6442_/D fanout458/X VGND VGND VPWR VPWR _6442_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_146_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3654_ hold85/A _3562_/B _3511_/A VGND VGND VPWR VPWR _3654_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6373_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6373_/X sky130_fd_sc_hd__and2_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7126_/CLK sky130_fd_sc_hd__clkbuf_8
X_3585_ hold48/A _3714_/B VGND VGND VPWR VPWR _3585_/Y sky130_fd_sc_hd__nor2_4
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5324_ hold798/X _5528_/A1 _5327_/S VGND VGND VPWR VPWR _5324_/X sky130_fd_sc_hd__mux2_1
X_5255_ hold746/X _5540_/A1 _5255_/S VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4206_ hold730/X _6356_/A1 _4207_/S VGND VGND VPWR VPWR _4206_/X sky130_fd_sc_hd__mux2_1
X_5186_ _5186_/A _5190_/B hold16/X VGND VGND VPWR VPWR _5189_/S sky130_fd_sc_hd__and3_1
XFILLER_56_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4137_ hold760/X _6356_/A1 _4138_/S VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4068_ _6396_/B _3546_/A _4118_/B _4050_/X _4322_/B VGND VGND VPWR VPWR _4084_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_83_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6709_ _6709_/CLK _6709_/D fanout445/X VGND VGND VPWR VPWR _6709_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold609 _4132_/X VGND VGND VPWR VPWR _6544_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3370_ _3370_/A hold74/X VGND VGND VPWR VPWR _3370_/Y sky130_fd_sc_hd__nor2_8
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _4574_/A _4816_/Y _4950_/X VGND VGND VPWR VPWR _5089_/B sky130_fd_sc_hd__a21oi_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1309 _6470_/Q VGND VGND VPWR VPWR _4033_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6991_ _7086_/CLK _6991_/D fanout484/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5942_ _7099_/Q _7100_/Q VGND VGND VPWR VPWR _5979_/C sky130_fd_sc_hd__and2b_2
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5873_ _6562_/Q _5631_/X _5646_/X _6652_/Q VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__a22o_1
X_4824_ _4542_/D _4562_/Y _4522_/D VGND VGND VPWR VPWR _4824_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4755_ _4542_/A _4581_/B _4611_/Y _4628_/Y VGND VGND VPWR VPWR _4755_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3706_ input35/X _3365_/Y _5301_/A _6867_/Q _3705_/X VGND VGND VPWR VPWR _3709_/B
+ sky130_fd_sc_hd__a221o_1
X_4686_ _4911_/B _4686_/B VGND VGND VPWR VPWR _4686_/Y sky130_fd_sc_hd__nand2_1
XFILLER_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6425_ _6926_/CLK _6425_/D fanout457/X VGND VGND VPWR VPWR _6425_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_162_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3637_ _7029_/Q hold49/A _4328_/A _6718_/Q _3636_/X VGND VGND VPWR VPWR _3638_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_174_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6356_ hold768/X _6356_/A1 _6357_/S VGND VGND VPWR VPWR _6356_/X sky130_fd_sc_hd__mux2_1
X_3568_ _3568_/A1 _4118_/B hold37/A input48/X _3567_/X VGND VGND VPWR VPWR _3580_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5307_ hold513/X _5538_/A1 _5309_/S VGND VGND VPWR VPWR _5307_/X sky130_fd_sc_hd__mux2_1
X_6287_ _6669_/Q _5938_/X _5952_/X _6709_/Q VGND VGND VPWR VPWR _6287_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3499_ _3573_/A _3562_/B VGND VGND VPWR VPWR _4280_/A sky130_fd_sc_hd__nor2_4
XFILLER_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5238_ _5238_/A _5541_/B VGND VGND VPWR VPWR _5246_/S sky130_fd_sc_hd__and2_4
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5169_ hold367/X _5526_/A1 _5170_/S VGND VGND VPWR VPWR _5169_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__buf_8
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4540_ _4661_/A _4724_/A _4959_/B _3962_/A VGND VGND VPWR VPWR _5039_/A sky130_fd_sc_hd__a31oi_4
XFILLER_156_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire381 _5975_/Y VGND VGND VPWR VPWR _5977_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_171_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold406 _4080_/X VGND VGND VPWR VPWR _6503_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4471_ _4702_/C _4471_/B _4471_/C VGND VGND VPWR VPWR _4489_/B sky130_fd_sc_hd__and3_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold417 _6895_/Q VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 _4258_/X VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6661_/Q _5976_/B _5971_/C _6711_/Q VGND VGND VPWR VPWR _6210_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold439 _6990_/Q VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_3422_ _6840_/Q _5265_/A _3414_/Y _3419_/X _3421_/X VGND VGND VPWR VPWR _3431_/A
+ sky130_fd_sc_hd__a2111o_1
X_7190_ _7190_/A VGND VGND VPWR VPWR _7190_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _6904_/Q _5976_/C _5971_/D _6832_/Q VGND VGND VPWR VPWR _6141_/X sky130_fd_sc_hd__a22o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3814_/A _3373_/B VGND VGND VPWR VPWR _5532_/A sky130_fd_sc_hd__nor2_8
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6072_ _7021_/Q _5937_/X _5975_/D _6885_/Q VGND VGND VPWR VPWR _6072_/X sky130_fd_sc_hd__a22o_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ hold62/X hold202/X _3283_/Y VGND VGND VPWR VPWR _3284_/X sky130_fd_sc_hd__a21bo_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _5359_/X VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _6667_/Q VGND VGND VPWR VPWR _4271_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 _4142_/X VGND VGND VPWR VPWR _6552_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5023_ _5023_/A _5023_/B _5023_/C _5023_/D VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__and4_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1139 _6768_/Q VGND VGND VPWR VPWR _5191_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6974_ _6990_/CLK _6974_/D fanout480/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfrtp_4
X_5925_ _7155_/Q _5625_/X _5661_/X _6623_/Q VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5856_ _6551_/Q _5913_/B1 _5855_/Y _5652_/B VGND VGND VPWR VPWR _5856_/X sky130_fd_sc_hd__a22o_1
X_4807_ _4846_/B _4645_/Y _4653_/Y _4689_/A VGND VGND VPWR VPWR _4807_/X sky130_fd_sc_hd__o22a_1
X_5787_ _5787_/A _5787_/B _5787_/C VGND VGND VPWR VPWR _5787_/Y sky130_fd_sc_hd__nor3_2
XFILLER_119_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4738_ _4738_/A VGND VGND VPWR VPWR _4738_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4669_ _4739_/A _5043_/A _4747_/B _4739_/B VGND VGND VPWR VPWR _4676_/B sky130_fd_sc_hd__and4b_1
XFILLER_174_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6408_ _3568_/A1 _6408_/D _6364_/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfrtp_2
Xhold940 _6896_/Q VGND VGND VPWR VPWR hold940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold951 _5157_/X VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 _6549_/Q VGND VGND VPWR VPWR hold962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 _4313_/X VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold984 _6436_/Q VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ _6642_/Q _6339_/A2 _6339_/B1 _6350_/A2 _6338_/X VGND VGND VPWR VPWR _6339_/X
+ sky130_fd_sc_hd__a221o_1
Xhold995 _6739_/Q VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3971_ hold93/X hold154/X _3975_/S VGND VGND VPWR VPWR _3971_/X sky130_fd_sc_hd__mux2_8
XFILLER_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5710_ _7012_/Q _5630_/X _5645_/X _7028_/Q _5709_/X VGND VGND VPWR VPWR _5711_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6690_ _6714_/CLK _6690_/D fanout470/X VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5641_ _5641_/A _5641_/B _5641_/C VGND VGND VPWR VPWR _5670_/A sky130_fd_sc_hd__nor3_1
XFILLER_148_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5572_ _7093_/Q _7092_/Q VGND VGND VPWR VPWR _5667_/B sky130_fd_sc_hd__and2_2
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_116_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4523_ _4584_/A _5042_/B VGND VGND VPWR VPWR _4523_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold203 _3284_/X VGND VGND VPWR VPWR _3285_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _4025_/X VGND VGND VPWR VPWR _6464_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _6789_/Q VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _5495_/X VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _4454_/A _4626_/B VGND VGND VPWR VPWR _4947_/C sky130_fd_sc_hd__nand2_8
XFILLER_171_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold247 _6419_/Q VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold258 _5204_/X VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _6681_/Q VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ input51/X _4058_/S _5337_/A _6905_/Q _3404_/X VGND VGND VPWR VPWR _3408_/C
+ sky130_fd_sc_hd__a221o_1
X_7173_ _7173_/A VGND VGND VPWR VPWR _7173_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4385_ _4556_/A _4753_/A _4607_/A VGND VGND VPWR VPWR _4441_/B sky130_fd_sc_hd__and3_4
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _7060_/Q _5954_/X _5976_/D _6879_/Q _6106_/X VGND VGND VPWR VPWR _6125_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ hold26/X hold46/X VGND VGND VPWR VPWR _3415_/B sky130_fd_sc_hd__and2_4
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _7005_/Q _5958_/X _5978_/X _6997_/Q VGND VGND VPWR VPWR _6055_/X sky130_fd_sc_hd__a22o_1
X_3267_ _3868_/A1 _3265_/X _3870_/S _3251_/A VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__a22o_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5006_ _5006_/A _5112_/A VGND VGND VPWR VPWR _5006_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3198_ _6989_/Q VGND VGND VPWR VPWR _3198_/Y sky130_fd_sc_hd__inv_2
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _6997_/CLK _6957_/D fanout463/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ _5552_/B _7116_/Q _6103_/B1 VGND VGND VPWR VPWR _5908_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6888_ _6888_/CLK _6888_/D fanout473/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5839_ _6685_/Q _5632_/X _5835_/X _5838_/X VGND VGND VPWR VPWR _5839_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold770 _6429_/Q VGND VGND VPWR VPWR hold770/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _5280_/X VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _7186_/A VGND VGND VPWR VPWR hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1470 _7107_/Q VGND VGND VPWR VPWR _5713_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 _6575_/Q VGND VGND VPWR VPWR _4169_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 _6053_/X VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput308 _3957_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
XFILLER_5_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput319 hold1345/X VGND VGND VPWR VPWR hold1346/A sky130_fd_sc_hd__buf_12
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4170_ _3447_/Y _4170_/A1 _4171_/S VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6811_ _7080_/CLK _6811_/D fanout479/X VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6742_ _6746_/CLK _6742_/D _3946_/B VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfrtp_4
X_3954_ _3954_/A _3961_/B VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__and2_1
XFILLER_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6673_ _6674_/CLK _6673_/D fanout468/X VGND VGND VPWR VPWR _6673_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_176_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3885_ _5552_/B _5606_/A VGND VGND VPWR VPWR _3885_/Y sky130_fd_sc_hd__nand2_1
X_5624_ _5638_/A _5658_/B _5663_/C VGND VGND VPWR VPWR _5624_/X sky130_fd_sc_hd__and3_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5555_ _7088_/Q _5562_/D VGND VGND VPWR VPWR _5555_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4506_ _4469_/A _4887_/A _4672_/A _4846_/A _4672_/B VGND VGND VPWR VPWR _4508_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5486_ hold503/X _5528_/A1 hold50/X VGND VGND VPWR VPWR _5486_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4437_ _4739_/A _4642_/A VGND VGND VPWR VPWR _4635_/B sky130_fd_sc_hd__nor2_8
X_7156_ _3945_/A1 _7156_/D _6387_/X VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfrtn_1
XFILLER_86_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4368_ _4500_/A _4469_/A _6644_/Q VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__o21a_1
XFILLER_59_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6107_ _6863_/Q _5943_/X _5981_/X _6919_/Q VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3319_ _3453_/A hold64/X VGND VGND VPWR VPWR _3454_/B sky130_fd_sc_hd__and2_4
X_7087_ _7131_/CLK _7087_/D fanout460/X VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4299_ _4299_/A0 hold667/X _4303_/S VGND VGND VPWR VPWR _4299_/X sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _6924_/Q _5938_/X _5952_/X _6956_/Q VGND VGND VPWR VPWR _6038_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_csclk _6447_/CLK VGND VGND VPWR VPWR _7049_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_79_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6735_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ _3670_/A _3670_/B _3670_/C _3670_/D VGND VGND VPWR VPWR _3670_/Y sky130_fd_sc_hd__nor4_1
XFILLER_185_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5340_ hold862/X _5484_/A1 _5345_/S VGND VGND VPWR VPWR _5340_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5271_ hold704/X _5469_/A1 _5273_/S VGND VGND VPWR VPWR _5271_/X sky130_fd_sc_hd__mux2_1
X_7010_ _7049_/CLK _7010_/D fanout457/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_141_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4222_ hold273/X _5534_/A1 _4225_/S VGND VGND VPWR VPWR _4222_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4153_ _4153_/A0 _5492_/A1 _4156_/S VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4084_ hold986/X _4083_/X _4084_/S VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4986_ _5005_/B _4985_/Y _4229_/X VGND VGND VPWR VPWR _4986_/X sky130_fd_sc_hd__a21o_1
X_6725_ _7140_/CLK _6725_/D _6307_/B VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfrtp_1
X_3937_ _6516_/Q _3937_/A1 _6765_/Q VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6656_ _6659_/CLK _6656_/D fanout469/X VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfrtp_4
X_3868_ _6406_/Q _3868_/A1 _3868_/S VGND VGND VPWR VPWR _6406_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5607_ _5607_/A1 _5606_/B _5606_/Y _5552_/B VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__a22o_1
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6587_ _7137_/CLK _6587_/D VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3799_ _6737_/Q _5148_/A hold67/A _6465_/Q VGND VGND VPWR VPWR _3799_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5538_ hold411/X _5538_/A1 _5540_/S VGND VGND VPWR VPWR _5538_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5469_ hold656/X _5469_/A1 _5471_/S VGND VGND VPWR VPWR _5469_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7139_ _7140_/CLK _7139_/D VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout398 hold42/X VGND VGND VPWR VPWR _5469_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_86_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4840_ _5051_/B _4911_/B VGND VGND VPWR VPWR _5086_/B sky130_fd_sc_hd__nand2_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _4771_/A _4995_/A _4771_/C _4771_/D VGND VGND VPWR VPWR _4772_/D sky130_fd_sc_hd__and4_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6510_ _6951_/CLK _6510_/D fanout473/X VGND VGND VPWR VPWR _6510_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3722_ _6907_/Q _5346_/A _4058_/S input44/X _3721_/X VGND VGND VPWR VPWR _3729_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6441_ _6747_/CLK _6441_/D fanout449/X VGND VGND VPWR VPWR _6441_/Q sky130_fd_sc_hd__dfstp_2
X_3653_ _6860_/Q _5292_/A _4151_/A _6562_/Q _3652_/X VGND VGND VPWR VPWR _3661_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6372_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6372_/X sky130_fd_sc_hd__and2_1
X_3584_ _3583_/X _6731_/Q _3829_/B VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__mux2_1
X_5323_ hold896/X _5509_/A1 _5327_/S VGND VGND VPWR VPWR _5323_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5254_ hold714/X _5521_/A1 _5255_/S VGND VGND VPWR VPWR _5254_/X sky130_fd_sc_hd__mux2_1
X_4205_ hold936/X _6355_/A1 _4207_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5185_ _6353_/A1 _5185_/A1 _5185_/S VGND VGND VPWR VPWR _5185_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR _6888_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4136_ hold866/X _5493_/A1 _4138_/S VGND VGND VPWR VPWR _4136_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4067_ hold732/X _4066_/X _4067_/S VGND VGND VPWR VPWR _4067_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4969_ _4969_/A _4969_/B VGND VGND VPWR VPWR _4969_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6708_ _6709_/CLK _6708_/D fanout445/X VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6639_ _3937_/A1 _6639_/D fanout487/X VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6990_ _6990_/CLK _6990_/D fanout480/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5941_ _5968_/A _5964_/A _5969_/C VGND VGND VPWR VPWR _5973_/A sky130_fd_sc_hd__and3_4
X_5872_ _7036_/Q _5614_/X _5871_/X VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4823_ _4823_/A _5099_/A VGND VGND VPWR VPWR _4823_/X sky130_fd_sc_hd__and2_1
XFILLER_179_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4754_ _4581_/B _4456_/Y _4611_/Y _4689_/B VGND VGND VPWR VPWR _4768_/C sky130_fd_sc_hd__o22a_1
XFILLER_119_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3705_ _7056_/Q hold86/A _5436_/A _6987_/Q VGND VGND VPWR VPWR _3705_/X sky130_fd_sc_hd__a22o_1
X_4685_ _4685_/A _5042_/B VGND VGND VPWR VPWR _4964_/B sky130_fd_sc_hd__nand2_2
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6424_ _6926_/CLK _6424_/D fanout457/X VGND VGND VPWR VPWR _6424_/Q sky130_fd_sc_hd__dfstp_2
X_3636_ _3268_/C _4118_/B _4262_/A _6663_/Q _3635_/X VGND VGND VPWR VPWR _3636_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6355_ hold980/X _6355_/A1 _6357_/S VGND VGND VPWR VPWR _6355_/X sky130_fd_sc_hd__mux2_1
X_3567_ _3960_/B _3331_/Y _4316_/A _6709_/Q VGND VGND VPWR VPWR _3567_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5306_ hold475/X _5528_/A1 _5309_/S VGND VGND VPWR VPWR _5306_/X sky130_fd_sc_hd__mux2_1
X_6286_ _6454_/Q _5947_/X _5965_/X _6549_/Q _6285_/X VGND VGND VPWR VPWR _6289_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_115_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3498_ _6894_/Q _5328_/A _4220_/A _6623_/Q VGND VGND VPWR VPWR _3498_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5237_ hold391/X _5540_/A1 _5237_/S VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5168_ hold271/X _5465_/A1 _5170_/S VGND VGND VPWR VPWR _5168_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4119_ _4119_/A0 _5491_/A1 _4126_/S VGND VGND VPWR VPWR _4119_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5099_ _5099_/A _5099_/B _5099_/C _5099_/D VGND VGND VPWR VPWR _5099_/X sky130_fd_sc_hd__and4_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire360 _5906_/Y VGND VGND VPWR VPWR wire360/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4470_ _4702_/C _4471_/C VGND VGND VPWR VPWR _4664_/A sky130_fd_sc_hd__nand2_1
Xhold407 _6860_/Q VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold418 _5334_/X VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3421_ _6944_/Q _5382_/A _3372_/Y _6440_/Q _3420_/X VGND VGND VPWR VPWR _3421_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold429 _6903_/Q VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6140_ _6140_/A _6140_/B _6140_/C VGND VGND VPWR VPWR _6140_/Y sky130_fd_sc_hd__nor3_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _3374_/A hold28/X VGND VGND VPWR VPWR _5328_/A sky130_fd_sc_hd__nor2_8
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _7066_/Q _5934_/X _5975_/B _6869_/Q _6070_/X VGND VGND VPWR VPWR _6074_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ hold202/X hold70/X VGND VGND VPWR VPWR _3283_/Y sky130_fd_sc_hd__nand2b_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _6462_/Q VGND VGND VPWR VPWR _4023_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5022_ _5112_/B _5021_/X _5006_/Y VGND VGND VPWR VPWR _5022_/Y sky130_fd_sc_hd__a21oi_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _4271_/X VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 _6567_/Q VGND VGND VPWR VPWR _4160_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6973_ _6990_/CLK _6973_/D fanout480/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5924_ _6699_/Q _5637_/X _5645_/X _6459_/Q VGND VGND VPWR VPWR _5924_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5855_ _6656_/Q _5899_/B VGND VGND VPWR VPWR _5855_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4806_ _4504_/X _5039_/B VGND VGND VPWR VPWR _4964_/C sky130_fd_sc_hd__and2b_1
X_5786_ _7008_/Q _5625_/X _5783_/X _5785_/X VGND VGND VPWR VPWR _5787_/C sky130_fd_sc_hd__a211o_1
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4737_ _4737_/A _4737_/B VGND VGND VPWR VPWR _4738_/A sky130_fd_sc_hd__and2_1
XFILLER_119_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4668_ _4921_/A _4928_/A _4668_/C VGND VGND VPWR VPWR _5002_/A sky130_fd_sc_hd__nand3_1
XFILLER_134_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3619_ _6740_/Q _5148_/A _4014_/A _6458_/Q _3618_/X VGND VGND VPWR VPWR _3620_/D
+ sky130_fd_sc_hd__a221o_1
X_6407_ _3568_/A1 _6407_/D _6363_/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfrtp_2
XFILLER_134_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold930 _6936_/Q VGND VGND VPWR VPWR hold930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _5335_/X VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _4563_/A _4396_/A _4598_/Y VGND VGND VPWR VPWR _4739_/B sky130_fd_sc_hd__a21oi_2
XFILLER_190_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold952 _6542_/Q VGND VGND VPWR VPWR hold952/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold963 _4138_/X VGND VGND VPWR VPWR _6549_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold974 _6634_/Q VGND VGND VPWR VPWR hold974/X sky130_fd_sc_hd__dlygate4sd3_1
X_6338_ _6644_/Q _6338_/A2 _6338_/B1 _6643_/Q VGND VGND VPWR VPWR _6338_/X sky130_fd_sc_hd__a22o_1
Xhold985 _3993_/X VGND VGND VPWR VPWR _6436_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold996 _5151_/X VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6269_ _6683_/Q _5934_/X _5975_/B _6617_/Q _6268_/X VGND VGND VPWR VPWR _6275_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3970_ hold988/X _6355_/A1 _3980_/S VGND VGND VPWR VPWR _3970_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5640_ _7010_/Q _5630_/X _5633_/X _5639_/X VGND VGND VPWR VPWR _5641_/C sky130_fd_sc_hd__a211o_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5571_ _6508_/Q _5658_/B VGND VGND VPWR VPWR _5576_/B sky130_fd_sc_hd__nand2_1
X_4522_ _4522_/A _4522_/B _4522_/C _4522_/D VGND VGND VPWR VPWR _4522_/X sky130_fd_sc_hd__and4_1
XFILLER_117_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold204 _3285_/X VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _7081_/Q VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _5215_/X VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _4607_/A _4453_/B VGND VGND VPWR VPWR _4886_/B sky130_fd_sc_hd__nor2_4
XFILLER_172_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold237 hold237/A VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _3968_/X VGND VGND VPWR VPWR _6419_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold259 _6995_/Q VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _6897_/Q _5328_/A _5247_/A _6825_/Q VGND VGND VPWR VPWR _3404_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4384_ _4384_/A _4892_/A VGND VGND VPWR VPWR _4907_/B sky130_fd_sc_hd__nor2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6815_/Q _5971_/B _5949_/X _6935_/Q _6122_/X VGND VGND VPWR VPWR _6125_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3335_ _3370_/A _3573_/A VGND VGND VPWR VPWR _5382_/A sky130_fd_sc_hd__nor2_8
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6861_/Q _5943_/X _5981_/X _6917_/Q VGND VGND VPWR VPWR _6054_/X sky130_fd_sc_hd__a22o_1
X_3266_ _6415_/Q _3266_/B VGND VGND VPWR VPWR _3870_/S sky130_fd_sc_hd__nor2_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5068_/B _5005_/B _5069_/B VGND VGND VPWR VPWR _5112_/A sky130_fd_sc_hd__and3_1
XFILLER_100_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3197_ _6997_/Q VGND VGND VPWR VPWR _3197_/Y sky130_fd_sc_hd__inv_2
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _6981_/CLK _6956_/D fanout463/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_1
X_5907_ _3223_/Y _5651_/Y _5896_/Y wire360/X _5552_/B VGND VGND VPWR VPWR _5907_/X
+ sky130_fd_sc_hd__a221o_1
X_6887_ _6951_/CLK _6887_/D fanout474/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5838_ _7034_/Q _5614_/X _5836_/X _5837_/X VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__a211o_1
XFILLER_182_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5769_ _6815_/Q _5667_/X _5764_/X _5765_/X _5768_/X VGND VGND VPWR VPWR _5769_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_108_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold760 _6548_/Q VGND VGND VPWR VPWR hold760/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold771 _3985_/X VGND VGND VPWR VPWR _6429_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 _6703_/Q VGND VGND VPWR VPWR hold782/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold793 _4063_/X VGND VGND VPWR VPWR _6495_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1460 _3488_/X VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1471 _5693_/X VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1482 _7127_/Q VGND VGND VPWR VPWR _6204_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 _7171_/Q VGND VGND VPWR VPWR _3233_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput309 _3952_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
XFILLER_5_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6810_ _7058_/CLK _6810_/D _6396_/A VGND VGND VPWR VPWR _6810_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6741_ _6746_/CLK _6741_/D _3946_/B VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3953_ _6403_/Q _3953_/B VGND VGND VPWR VPWR _3953_/X sky130_fd_sc_hd__and2b_4
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3884_ _3894_/B2 _3174_/Y _3883_/X VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__a21o_1
X_6672_ _6674_/CLK _6672_/D fanout468/X VGND VGND VPWR VPWR _6672_/Q sky130_fd_sc_hd__dfrtp_1
X_5623_ _7094_/Q _7095_/Q VGND VGND VPWR VPWR _5663_/C sky130_fd_sc_hd__and2b_2
XFILLER_164_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5554_ _5562_/D VGND VGND VPWR VPWR _5554_/Y sky130_fd_sc_hd__inv_2
X_4505_ _5010_/A _4972_/A VGND VGND VPWR VPWR _4912_/A sky130_fd_sc_hd__nand2_1
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5485_ _5485_/A0 _5545_/A1 hold50/X VGND VGND VPWR VPWR _5485_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4436_ _4631_/D _4633_/B VGND VGND VPWR VPWR _4615_/B sky130_fd_sc_hd__nor2_4
XFILLER_144_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7155_ _7155_/CLK _7155_/D fanout450/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_4
X_4367_ _4562_/A _4690_/B VGND VGND VPWR VPWR _4469_/A sky130_fd_sc_hd__nand2_4
X_3318_ _3555_/A _3714_/A VGND VGND VPWR VPWR _5292_/A sky130_fd_sc_hd__nor2_8
X_6106_ _7084_/Q _5976_/B _5971_/C _7044_/Q VGND VGND VPWR VPWR _6106_/X sky130_fd_sc_hd__a22o_1
X_7086_ _7086_/CLK hold23/X fanout483/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4298_ _4298_/A _4322_/B VGND VGND VPWR VPWR _4303_/S sky130_fd_sc_hd__and2_2
XFILLER_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3249_/A _3249_/B VGND VGND VPWR VPWR _3250_/B sky130_fd_sc_hd__nor2_1
X_6037_ _6972_/Q _5947_/X _5965_/X _6796_/Q _6036_/X VGND VGND VPWR VPWR _6040_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _6981_/CLK _6939_/D fanout463/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfstp_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_csclk _3942_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_135_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold590 _7042_/Q VGND VGND VPWR VPWR hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1290 _4281_/X VGND VGND VPWR VPWR _6675_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5270_ hold166/X hold60/X _5273_/S VGND VGND VPWR VPWR _5270_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4221_ _4221_/A0 hold667/X _4225_/S VGND VGND VPWR VPWR _4221_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4152_ _4152_/A0 _6353_/A1 _4156_/S VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__mux2_1
X_4083_ hold555/X _5513_/A1 _4083_/S VGND VGND VPWR VPWR _4083_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4985_ _5068_/B _5069_/B _5008_/B _4985_/D VGND VGND VPWR VPWR _4985_/Y sky130_fd_sc_hd__nand4_1
XFILLER_168_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6724_ _7150_/CLK _6724_/D _6307_/B VGND VGND VPWR VPWR _6724_/Q sky130_fd_sc_hd__dfrtp_2
X_3936_ _6517_/Q user_clock _6766_/Q VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR _6447_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6655_ _6655_/CLK _6655_/D fanout468/X VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfrtp_2
X_3867_ _3867_/A _3867_/B VGND VGND VPWR VPWR _3868_/S sky130_fd_sc_hd__nor2_1
XFILLER_137_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5606_ _5606_/A _5606_/B VGND VGND VPWR VPWR _5606_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6586_ _7137_/CLK _6586_/D VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfxtp_1
X_3798_ _6434_/Q _3372_/Y _3511_/Y _3796_/X _3797_/X VGND VGND VPWR VPWR _3798_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_118_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5537_ hold806/X _5546_/A1 _5540_/S VGND VGND VPWR VPWR _5537_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5468_ hold131/X hold60/X _5471_/S VGND VGND VPWR VPWR _5468_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4419_ _4556_/A _4563_/A VGND VGND VPWR VPWR _4561_/B sky130_fd_sc_hd__nand2_4
X_5399_ hold592/X _5513_/A1 _5399_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7138_ _7140_/CLK _7138_/D VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7069_ _7069_/CLK _7069_/D fanout482/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout399 hold42/X VGND VGND VPWR VPWR _5538_/A1 sky130_fd_sc_hd__buf_6
XFILLER_86_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _4942_/C _4770_/B _5003_/A _4770_/D VGND VGND VPWR VPWR _4771_/D sky130_fd_sc_hd__and4_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3721_ _6899_/Q _5337_/A _5166_/A _6752_/Q VGND VGND VPWR VPWR _3721_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6440_ _6747_/CLK _6440_/D fanout447/X VGND VGND VPWR VPWR _6440_/Q sky130_fd_sc_hd__dfstp_4
X_3652_ _6657_/Q _4256_/A _4214_/A _6616_/Q VGND VGND VPWR VPWR _3652_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6371_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6371_/X sky130_fd_sc_hd__and2_1
X_3583_ _4192_/A0 _3642_/A1 _3829_/A VGND VGND VPWR VPWR _3583_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5322_ _5322_/A0 _5484_/A1 _5327_/S VGND VGND VPWR VPWR _5322_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ hold800/X _5538_/A1 _5255_/S VGND VGND VPWR VPWR _5253_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4204_ hold822/X _6354_/A1 _4207_/S VGND VGND VPWR VPWR _4204_/X sky130_fd_sc_hd__mux2_1
X_5184_ _5184_/A _6352_/B VGND VGND VPWR VPWR _5185_/S sky130_fd_sc_hd__nand2_1
X_4135_ _4135_/A0 _5492_/A1 _4138_/S VGND VGND VPWR VPWR _4135_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_csclk _6447_/CLK VGND VGND VPWR VPWR _7011_/CLK sky130_fd_sc_hd__clkbuf_16
X_4066_ _4117_/A0 _5540_/A1 hold37/X VGND VGND VPWR VPWR _4066_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_78_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6739_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4968_ _4627_/A _5041_/A _4789_/X VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__o21a_1
X_6707_ _6707_/CLK _6707_/D fanout445/X VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_20_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3919_ _6522_/Q input89/X _3921_/S VGND VGND VPWR VPWR _3919_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4899_ _4899_/A _4899_/B _4877_/A VGND VGND VPWR VPWR _5118_/A sky130_fd_sc_hd__nor3b_1
XFILLER_177_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6638_ _7150_/CLK _6638_/D fanout487/X VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6569_ _6653_/CLK _6569_/D fanout454/X VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7058_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5940_ _5964_/A _5981_/A _5981_/C VGND VGND VPWR VPWR _5940_/X sky130_fd_sc_hd__and3_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5871_ _6717_/Q _5642_/X _5666_/X _6632_/Q VGND VGND VPWR VPWR _5871_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4822_ _5084_/B _4942_/A VGND VGND VPWR VPWR _5092_/A sky130_fd_sc_hd__and2_1
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4753_ _4753_/A _4753_/B _4753_/C VGND VGND VPWR VPWR _5062_/C sky130_fd_sc_hd__nand3_1
X_3704_ _6666_/Q _4268_/A _4316_/A _6706_/Q _3703_/X VGND VGND VPWR VPWR _3709_/A
+ sky130_fd_sc_hd__a221o_1
X_4684_ _4482_/A _4672_/A _4626_/Y _4230_/B VGND VGND VPWR VPWR _4964_/A sky130_fd_sc_hd__o31a_1
X_6423_ _7049_/CLK _6423_/D fanout457/X VGND VGND VPWR VPWR _6423_/Q sky130_fd_sc_hd__dfstp_4
X_3635_ _7074_/Q _5532_/A _4202_/A _6607_/Q VGND VGND VPWR VPWR _3635_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6354_ hold836/X _6354_/A1 _6357_/S VGND VGND VPWR VPWR _6354_/X sky130_fd_sc_hd__mux2_1
X_3566_ _3573_/A hold66/X VGND VGND VPWR VPWR _4316_/A sky130_fd_sc_hd__nor2_8
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5305_ _5305_/A0 _5545_/A1 _5309_/S VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6285_ _6634_/Q _5946_/X _5955_/X _6554_/Q VGND VGND VPWR VPWR _6285_/X sky130_fd_sc_hd__a22o_1
X_3497_ _3554_/A _3571_/B VGND VGND VPWR VPWR _4220_/A sky130_fd_sc_hd__nor2_4
XFILLER_115_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5236_ hold908/X _5548_/A1 _5237_/S VGND VGND VPWR VPWR _5236_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5167_ _5167_/A0 _5524_/A1 _5170_/S VGND VGND VPWR VPWR _5167_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4118_ _6400_/B _4118_/B _6352_/B VGND VGND VPWR VPWR _4126_/S sky130_fd_sc_hd__and3b_4
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5098_ _4810_/A _4582_/Y _4616_/Y _4626_/Y _4658_/C VGND VGND VPWR VPWR _5099_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_44_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4049_ hold539/X _6357_/A1 _4049_/S VGND VGND VPWR VPWR _4049_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire350 _3661_/Y VGND VGND VPWR VPWR _3700_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_190_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire372 _3554_/A VGND VGND VPWR VPWR _3374_/A sky130_fd_sc_hd__buf_12
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold408 _5295_/X VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 _7073_/Q VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ _7085_/Q _5541_/A hold76/A _7045_/Q VGND VGND VPWR VPWR _3420_/X sky130_fd_sc_hd__a22o_2
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3351_ _3586_/A _3573_/A VGND VGND VPWR VPWR _5427_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3282_ hold47/X _3313_/A VGND VGND VPWR VPWR _3586_/A sky130_fd_sc_hd__nand2_8
X_6070_ _7050_/Q _5971_/A _5979_/X _6989_/Q VGND VGND VPWR VPWR _6070_/X sky130_fd_sc_hd__a22o_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _4023_/X VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5021_ _5021_/A _5021_/B _5021_/C _5021_/D VGND VGND VPWR VPWR _5021_/X sky130_fd_sc_hd__and4_1
Xhold1119 _7036_/Q VGND VGND VPWR VPWR _5493_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6972_ _7080_/CLK _6972_/D fanout479/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5923_ _6608_/Q _5648_/X _5910_/X _5922_/X VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5854_ _6706_/Q _5638_/X _5654_/X _6676_/Q _5853_/X VGND VGND VPWR VPWR _5862_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4805_ _4690_/A _4741_/A _4601_/B _4791_/X _4804_/X VGND VGND VPWR VPWR _4805_/X
+ sky130_fd_sc_hd__o311a_1
X_5785_ _6904_/Q _5621_/X _5645_/X _7032_/Q _5784_/X VGND VGND VPWR VPWR _5785_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4736_ _5010_/B _4644_/B _4735_/X _4921_/A VGND VGND VPWR VPWR _4737_/B sky130_fd_sc_hd__a22o_1
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4667_ _4739_/B _4733_/B _4747_/B VGND VGND VPWR VPWR _4668_/C sky130_fd_sc_hd__and3b_1
XFILLER_107_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6406_ _3945_/A1 _6406_/D _6362_/X VGND VGND VPWR VPWR _6406_/Q sky130_fd_sc_hd__dfrtp_4
X_3618_ _6989_/Q _5436_/A _5463_/A _7013_/Q VGND VGND VPWR VPWR _3618_/X sky130_fd_sc_hd__a22o_2
XFILLER_134_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold920 _6816_/Q VGND VGND VPWR VPWR hold920/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold931 _5380_/X VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4598_ _4642_/A _5043_/A VGND VGND VPWR VPWR _4598_/Y sky130_fd_sc_hd__nor2_1
Xhold942 _6603_/Q VGND VGND VPWR VPWR hold942/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold953 _4130_/X VGND VGND VPWR VPWR _6542_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold964 _6674_/Q VGND VGND VPWR VPWR hold964/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6337_ _6336_/X _6337_/A1 _6346_/S VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__mux2_1
Xhold975 _4243_/X VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3549_ _6822_/Q _5247_/A hold49/A _7030_/Q VGND VGND VPWR VPWR _3549_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold986 _7178_/A VGND VGND VPWR VPWR hold986/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold997 _7184_/A VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6268_ _6703_/Q _5971_/A _5979_/X _6473_/Q VGND VGND VPWR VPWR _6268_/X sky130_fd_sc_hd__a22o_2
XFILLER_88_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5219_ hold660/X _5513_/A1 hold18/X VGND VGND VPWR VPWR _5219_/X sky130_fd_sc_hd__mux2_1
X_6199_ _6690_/Q _5954_/X _5976_/D _6619_/Q _6180_/X VGND VGND VPWR VPWR _6200_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_29_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5570_ _7093_/Q _7092_/Q VGND VGND VPWR VPWR _5658_/B sky130_fd_sc_hd__nor2_8
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4521_ _4584_/A _4531_/B VGND VGND VPWR VPWR _4522_/D sky130_fd_sc_hd__nand2_1
XFILLER_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold205 _3286_/X VGND VGND VPWR VPWR _3347_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ _4753_/A _4454_/A VGND VGND VPWR VPWR _4453_/B sky130_fd_sc_hd__nand2b_4
Xhold216 _5544_/X VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _6669_/Q VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _4105_/X VGND VGND VPWR VPWR _6520_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _6955_/Q VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3403_ _6977_/Q _5418_/A _3381_/Y input33/X _3402_/X VGND VGND VPWR VPWR _3408_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7171_ _3945_/A1 _7171_/D _6401_/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4383_ _4892_/A VGND VGND VPWR VPWR _4462_/B sky130_fd_sc_hd__inv_2
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6447_/Q _5601_/X _5959_/X _6967_/Q VGND VGND VPWR VPWR _6122_/X sky130_fd_sc_hd__a22o_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3571_/A _3370_/A VGND VGND VPWR VPWR _5238_/A sky130_fd_sc_hd__nor2_8
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A0 _6052_/X _6279_/S VGND VGND VPWR VPWR _6053_/X sky130_fd_sc_hd__mux2_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _7159_/Q _6415_/Q _3266_/B VGND VGND VPWR VPWR _3265_/X sky130_fd_sc_hd__a21o_1
XFILLER_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5004_/A _5004_/B _5074_/B _5071_/B VGND VGND VPWR VPWR _5004_/Y sky130_fd_sc_hd__nand4_1
X_3196_ _7005_/Q VGND VGND VPWR VPWR _3196_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _7012_/CLK _6955_/D fanout458/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5906_ _5906_/A _5906_/B _5906_/C _5906_/D VGND VGND VPWR VPWR _5906_/Y sky130_fd_sc_hd__nor4_1
XFILLER_62_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6886_ _6890_/CLK _6886_/D fanout476/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5837_ _6650_/Q _5646_/X _5667_/X _6555_/Q VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5768_ _6447_/Q _5614_/X _5766_/X _5767_/X VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__a211o_1
XFILLER_108_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4719_ _4469_/A _4639_/Y _4673_/B _4694_/Y VGND VGND VPWR VPWR _4719_/X sky130_fd_sc_hd__o22a_1
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5699_ _6868_/Q _5628_/X _5634_/X _6972_/Q _5698_/X VGND VGND VPWR VPWR _5706_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold750 _7016_/Q VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 _4137_/X VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold772 _6437_/Q VGND VGND VPWR VPWR hold772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 _4314_/X VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _6686_/Q VGND VGND VPWR VPWR hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1450 _3313_/A VGND VGND VPWR VPWR _3375_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _6733_/Q VGND VGND VPWR VPWR _3449_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1472 _6576_/Q VGND VGND VPWR VPWR _4170_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1483 _7125_/Q VGND VGND VPWR VPWR _6178_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1494 _6571_/Q VGND VGND VPWR VPWR _4165_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6740_ _6746_/CLK _6740_/D _3946_/B VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3952_ _6404_/Q _3952_/B VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__and2b_4
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6671_ _6671_/CLK _6671_/D fanout468/X VGND VGND VPWR VPWR _6671_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_189_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3883_ _7088_/Q _7089_/Q _6509_/Q _5608_/C VGND VGND VPWR VPWR _3883_/X sky130_fd_sc_hd__and4b_1
X_5622_ _7018_/Q _5619_/X _5621_/X _6898_/Q _5617_/X VGND VGND VPWR VPWR _5641_/A
+ sky130_fd_sc_hd__a221o_1
X_5553_ _6509_/Q _5552_/B _6508_/Q _3885_/Y VGND VGND VPWR VPWR _5562_/D sky130_fd_sc_hd__o31a_1
XFILLER_129_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4504_ _4969_/A _4984_/A _4965_/B VGND VGND VPWR VPWR _4504_/X sky130_fd_sc_hd__and3_1
X_5484_ hold878/X _5484_/A1 hold50/X VGND VGND VPWR VPWR _5484_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4435_ _4566_/A _4591_/A VGND VGND VPWR VPWR _4482_/A sky130_fd_sc_hd__nand2_4
XFILLER_132_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7154_ _7155_/CLK _7154_/D fanout449/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfrtp_2
X_4366_ _4690_/A _4460_/A VGND VGND VPWR VPWR _5010_/A sky130_fd_sc_hd__nor2_4
XFILLER_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6105_ _7068_/Q _5934_/X _5975_/B _6871_/Q VGND VGND VPWR VPWR _6105_/X sky130_fd_sc_hd__a22o_1
X_3317_ hold27/X hold84/X VGND VGND VPWR VPWR _3714_/A sky130_fd_sc_hd__nand2_8
X_7085_ _7085_/CLK _7085_/D fanout483/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfrtp_1
X_4297_ hold531/X _6357_/A1 _4297_/S VGND VGND VPWR VPWR _4297_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6892_/Q _5946_/X _5955_/X _6804_/Q VGND VGND VPWR VPWR _6036_/X sky130_fd_sc_hd__a22o_1
X_3248_ _3248_/A1 _3249_/B _3247_/Y _7168_/Q VGND VGND VPWR VPWR _3248_/X sky130_fd_sc_hd__o22a_1
XFILLER_73_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3179_ _6508_/Q VGND VGND VPWR VPWR _5610_/B sky130_fd_sc_hd__clkinv_2
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7026_/CLK _6938_/D fanout463/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfstp_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ _7085_/CLK _6869_/D fanout477/X VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold580 _6709_/Q VGND VGND VPWR VPWR hold580/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 _5500_/X VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1280 _4021_/X VGND VGND VPWR VPWR _6460_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 _6560_/Q VGND VGND VPWR VPWR _4152_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4220_ _4220_/A _4322_/B VGND VGND VPWR VPWR _4225_/S sky130_fd_sc_hd__and2_2
XFILLER_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4151_ _4151_/A _4322_/B VGND VGND VPWR VPWR _4156_/S sky130_fd_sc_hd__and2_2
XFILLER_95_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4082_ hold239/X _4081_/X _4084_/S VGND VGND VPWR VPWR _4082_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4984_ _4984_/A _4984_/B VGND VGND VPWR VPWR _4997_/C sky130_fd_sc_hd__nand2_1
X_6723_ _7150_/CLK _6723_/D _6307_/B VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3935_ _3222_/Y input2/X input1/X VGND VGND VPWR VPWR _3935_/X sky130_fd_sc_hd__mux2_4
X_6654_ _6654_/CLK hold61/X fanout454/X VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfrtp_1
X_3866_ _3865_/X _3866_/A1 _3866_/S VGND VGND VPWR VPWR _6407_/D sky130_fd_sc_hd__mux2_1
X_5605_ _5552_/Y _5567_/Y _5604_/Y _6509_/Q VGND VGND VPWR VPWR _5606_/B sky130_fd_sc_hd__a22o_1
XFILLER_137_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6585_ _7137_/CLK _6585_/D VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfxtp_1
X_3797_ _6882_/Q _5319_/A _4238_/A _6630_/Q VGND VGND VPWR VPWR _3797_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5536_ _5536_/A0 _5545_/A1 _5540_/S VGND VGND VPWR VPWR _5536_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5467_ _5467_/A0 _5545_/A1 _5471_/S VGND VGND VPWR VPWR _5467_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4418_ _4556_/A _4563_/A VGND VGND VPWR VPWR _4600_/B sky130_fd_sc_hd__and2_4
X_5398_ hold636/X _5521_/A1 _5399_/S VGND VGND VPWR VPWR _5398_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7137_ _7137_/CLK _7137_/D VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4349_ _4471_/B _4591_/A VGND VGND VPWR VPWR _4911_/A sky130_fd_sc_hd__and2b_2
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7068_ _7078_/CLK _7068_/D fanout482/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout389 _4546_/Y VGND VGND VPWR VPWR _4846_/B sky130_fd_sc_hd__buf_6
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6019_ _7064_/Q _5934_/X _5975_/B _6867_/Q _6018_/X VGND VGND VPWR VPWR _6024_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3720_ _3720_/A _3720_/B _3720_/C _3720_/D VGND VGND VPWR VPWR _3730_/B sky130_fd_sc_hd__nor4_1
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3651_ _3651_/A _3651_/B _3651_/C _3651_/D VGND VGND VPWR VPWR _3651_/Y sky130_fd_sc_hd__nor4_1
XFILLER_158_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6370_ _6383_/A _6396_/B VGND VGND VPWR VPWR _6370_/X sky130_fd_sc_hd__and2_1
X_3582_ _3582_/A _3582_/B _3582_/C VGND VGND VPWR VPWR _3582_/Y sky130_fd_sc_hd__nand3_2
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5321_ hold535/X _5543_/A1 _5327_/S VGND VGND VPWR VPWR _5321_/X sky130_fd_sc_hd__mux2_1
X_5252_ hold188/X _5519_/A1 _5255_/S VGND VGND VPWR VPWR _5252_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4203_ _4203_/A0 _5491_/A1 _4207_/S VGND VGND VPWR VPWR _4203_/X sky130_fd_sc_hd__mux2_1
X_5183_ hold17/X _5183_/B VGND VGND VPWR VPWR _5183_/X sky130_fd_sc_hd__and2_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4134_ _4134_/A0 _5491_/A1 _4138_/S VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4065_ _4065_/A0 _4064_/X _4067_/S VGND VGND VPWR VPWR _4065_/X sky130_fd_sc_hd__mux2_1
X_4967_ _4967_/A _4967_/B VGND VGND VPWR VPWR _5066_/A sky130_fd_sc_hd__and2_1
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6706_ _6709_/CLK _6706_/D fanout445/X VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfrtp_2
X_3918_ _6523_/Q input91/X _3921_/S VGND VGND VPWR VPWR _3918_/X sky130_fd_sc_hd__mux2_2
X_4898_ _4359_/Y _4892_/B _4877_/C VGND VGND VPWR VPWR _4899_/B sky130_fd_sc_hd__o21ai_1
XFILLER_149_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6637_ _7150_/CLK _6637_/D fanout487/X VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_4
X_3849_ _3849_/A1 _3851_/C _3848_/X _3292_/X VGND VGND VPWR VPWR _6413_/D sky130_fd_sc_hd__o22a_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6568_ _6755_/CLK _6568_/D fanout445/X VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5519_ hold178/X _5519_/A1 hold87/A VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__mux2_1
X_6499_ _6755_/CLK _6499_/D _6360_/A VGND VGND VPWR VPWR _6499_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5870_ _6477_/Q _5630_/X _5867_/X _5868_/X _5869_/X VGND VGND VPWR VPWR _5870_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4821_ _4542_/A _4562_/Y _4518_/B VGND VGND VPWR VPWR _4821_/X sky130_fd_sc_hd__o21a_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4752_ _4413_/Y _4672_/B _4619_/Y _4626_/Y VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__o22a_1
XFILLER_147_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3703_ _6461_/Q _4020_/A _4014_/A _6456_/Q VGND VGND VPWR VPWR _3703_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4683_ _4424_/Y _4430_/Y _4504_/X _4682_/Y _4920_/B VGND VGND VPWR VPWR _4683_/X
+ sky130_fd_sc_hd__o41a_1
X_6422_ _6749_/CLK _6422_/D fanout449/X VGND VGND VPWR VPWR _6422_/Q sky130_fd_sc_hd__dfstp_1
X_3634_ _6973_/Q _5418_/A _5364_/A _6925_/Q _3633_/X VGND VGND VPWR VPWR _3638_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_147_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6353_ _6353_/A0 _6353_/A1 _6357_/S VGND VGND VPWR VPWR _6353_/X sky130_fd_sc_hd__mux2_1
X_3565_ _3565_/A _3565_/B _3565_/C VGND VGND VPWR VPWR _3581_/C sky130_fd_sc_hd__nor3_1
X_5304_ hold966/X _5484_/A1 _5309_/S VGND VGND VPWR VPWR _5304_/X sky130_fd_sc_hd__mux2_1
X_6284_ _6689_/Q _5961_/X _6282_/X _6283_/X VGND VGND VPWR VPWR _6289_/A sky130_fd_sc_hd__a211o_1
X_3496_ _6757_/Q _5182_/S _4310_/A _6704_/Q _3494_/X VGND VGND VPWR VPWR _3504_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5235_ hold511/X _5538_/A1 _5237_/S VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5166_ _5166_/A hold17/X VGND VGND VPWR VPWR _5170_/S sky130_fd_sc_hd__and2_1
XFILLER_68_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4117_ _4117_/A0 hold22/X hold38/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__mux2_1
XFILLER_29_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5097_ _5115_/A _5087_/Y _5096_/X _5078_/X VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__a211o_1
X_4048_ hold774/X _6356_/A1 _4049_/S VGND VGND VPWR VPWR _4048_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5999_ _6802_/Q _5955_/X _5975_/B _6866_/Q _5983_/X VGND VGND VPWR VPWR _6000_/D
+ sky130_fd_sc_hd__a221o_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput290 _6437_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_58_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__buf_6
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire351 _3651_/Y VGND VGND VPWR VPWR _3700_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_62_csclk _6447_/CLK VGND VGND VPWR VPWR _6963_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold409 _7057_/Q VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3350_ hold48/X _3543_/A VGND VGND VPWR VPWR _5409_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6746_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ hold83/X hold64/X VGND VGND VPWR VPWR _3313_/A sky130_fd_sc_hd__and2_4
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5021_/A _5021_/B _5021_/D VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__and3_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1109 _6965_/Q VGND VGND VPWR VPWR _5413_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6971_ _7080_/CLK _6971_/D fanout480/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5922_ _6649_/Q _5621_/X _5654_/X _6679_/Q _5921_/X VGND VGND VPWR VPWR _5922_/X
+ sky130_fd_sc_hd__a221o_1
X_5853_ _7152_/Q _5625_/X _5666_/X _6631_/Q VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6712_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4804_ _4804_/A _4804_/B _4804_/C VGND VGND VPWR VPWR _4804_/X sky130_fd_sc_hd__and3_1
X_5784_ _6944_/Q _5632_/X _5664_/X _6928_/Q VGND VGND VPWR VPWR _5784_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4735_ _4735_/A _4735_/B _4747_/C VGND VGND VPWR VPWR _4735_/X sky130_fd_sc_hd__and3_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4666_ _4441_/A _4400_/B _4665_/X VGND VGND VPWR VPWR _4733_/B sky130_fd_sc_hd__o21ai_1
X_6405_ _3945_/A1 _6405_/D _6361_/X VGND VGND VPWR VPWR _6405_/Q sky130_fd_sc_hd__dfrtp_4
X_3617_ _6949_/Q _3781_/A2 _4280_/A _6678_/Q _3616_/X VGND VGND VPWR VPWR _3620_/C
+ sky130_fd_sc_hd__a221o_1
Xhold910 _7045_/Q VGND VGND VPWR VPWR hold910/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 _5245_/X VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4597_ _4735_/B _4735_/A VGND VGND VPWR VPWR _4747_/B sky130_fd_sc_hd__and2b_1
Xhold932 _6904_/Q VGND VGND VPWR VPWR hold932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _4201_/X VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 _6707_/Q VGND VGND VPWR VPWR hold954/X sky130_fd_sc_hd__dlygate4sd3_1
X_6336_ _6642_/Q _6336_/A2 _6336_/B1 _6350_/A2 _6335_/X VGND VGND VPWR VPWR _6336_/X
+ sky130_fd_sc_hd__a221o_1
X_3548_ input24/X _3367_/Y _5463_/A _7014_/Q _3547_/X VGND VGND VPWR VPWR _3552_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold965 _4279_/X VGND VGND VPWR VPWR _6674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _6599_/Q VGND VGND VPWR VPWR hold976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 _4084_/X VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _4059_/X VGND VGND VPWR VPWR _6493_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6267_ _6563_/Q _5953_/X _5960_/X _6673_/Q _6266_/X VGND VGND VPWR VPWR _6267_/X
+ sky130_fd_sc_hd__a221o_1
X_3479_ _6807_/Q _5229_/A _5301_/A _6871_/Q _3478_/X VGND VGND VPWR VPWR _3484_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5218_ hold139/X hold99/X hold18/X VGND VGND VPWR VPWR _5218_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6198_ _6555_/Q _5971_/B _5949_/X _6675_/Q _6197_/X VGND VGND VPWR VPWR _6200_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5149_ _5149_/A0 _5491_/A1 _5153_/S VGND VGND VPWR VPWR _5149_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4520_ _4724_/A _4953_/A VGND VGND VPWR VPWR _4522_/C sky130_fd_sc_hd__nand2_1
XFILLER_117_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold206 _3370_/Y VGND VGND VPWR VPWR _5454_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _4753_/A _4495_/A VGND VGND VPWR VPWR _4496_/B sky130_fd_sc_hd__nor2_2
XFILLER_172_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold217 _6941_/Q VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _4273_/X VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold239 _6504_/Q VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _6961_/Q _5400_/A _5256_/A _6833_/Q VGND VGND VPWR VPWR _3402_/X sky130_fd_sc_hd__a22o_1
X_7170_ _3927_/A1 _7170_/D _6400_/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_1
X_4382_ _4359_/B _4382_/B VGND VGND VPWR VPWR _4892_/A sky130_fd_sc_hd__nand2b_2
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6121_ _7031_/Q _5944_/X _5975_/A _6847_/Q _6120_/X VGND VGND VPWR VPWR _6125_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ hold85/X hold75/X VGND VGND VPWR VPWR _5445_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _7120_/Q _6051_/X _6303_/S VGND VGND VPWR VPWR _6052_/X sky130_fd_sc_hd__mux2_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _6485_/Q _3264_/B VGND VGND VPWR VPWR _3266_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5003_ _5003_/A _5003_/B _5003_/C VGND VGND VPWR VPWR _5071_/B sky130_fd_sc_hd__and3_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3195_ _7013_/Q VGND VGND VPWR VPWR _3195_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6954_ _7012_/CLK _6954_/D fanout458/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfstp_1
X_5905_ _6548_/Q _5905_/A2 _5666_/X _6633_/Q _5904_/X VGND VGND VPWR VPWR _5906_/D
+ sky130_fd_sc_hd__a221o_1
X_6885_ _6969_/CLK _6885_/D fanout475/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5836_ _6715_/Q _5642_/X _5666_/X _6630_/Q VGND VGND VPWR VPWR _5836_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5767_ _6999_/Q _5643_/X _5664_/X _6927_/Q VGND VGND VPWR VPWR _5767_/X sky130_fd_sc_hd__a22o_1
X_4718_ _4645_/Y _4690_/Y _4716_/Y _4717_/X VGND VGND VPWR VPWR _4721_/B sky130_fd_sc_hd__o211a_1
X_5698_ _6980_/Q _5624_/X _5654_/X _6932_/Q VGND VGND VPWR VPWR _5698_/X sky130_fd_sc_hd__a22o_1
X_4649_ _4612_/Y _4613_/Y _4616_/Y _4609_/Y _4621_/X VGND VGND VPWR VPWR _4660_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold740 _6708_/Q VGND VGND VPWR VPWR hold740/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold751 _5470_/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _6817_/Q VGND VGND VPWR VPWR hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _3994_/X VGND VGND VPWR VPWR _6437_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold784 _6421_/Q VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__dlygate4sd3_1
X_6319_ _6320_/B _6319_/B VGND VGND VPWR VPWR _6319_/Y sky130_fd_sc_hd__nand2_1
Xhold795 _4294_/X VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1440 _6591_/Q VGND VGND VPWR VPWR _4188_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 _3814_/B VGND VGND VPWR VPWR _3376_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1462 _6721_/Q VGND VGND VPWR VPWR _4885_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1473 _6572_/Q VGND VGND VPWR VPWR _4166_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 _6154_/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1495 _6589_/Q VGND VGND VPWR VPWR _4185_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3951_ input85/X _3251_/A _6404_/Q VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__mux2_2
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6670_ _6671_/CLK _6670_/D fanout468/X VGND VGND VPWR VPWR _6670_/Q sky130_fd_sc_hd__dfrtp_2
X_3882_ _7090_/Q _7091_/Q VGND VGND VPWR VPWR _5608_/C sky130_fd_sc_hd__nor2_1
XFILLER_149_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5621_ _5664_/A _5666_/B _5660_/C VGND VGND VPWR VPWR _5621_/X sky130_fd_sc_hd__and3b_4
X_5552_ _6509_/Q _5552_/B VGND VGND VPWR VPWR _5552_/Y sky130_fd_sc_hd__nor2_1
X_4503_ _4582_/B _4881_/B VGND VGND VPWR VPWR _4925_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5483_ hold588/X _5543_/A1 hold50/X VGND VGND VPWR VPWR _5483_/X sky130_fd_sc_hd__mux2_1
X_4434_ _4566_/A _4434_/B VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__and2_2
XFILLER_104_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7153_ _7155_/CLK _7153_/D fanout449/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_132_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4365_ _4556_/A _4563_/A VGND VGND VPWR VPWR _4460_/A sky130_fd_sc_hd__nand2b_4
XFILLER_113_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6104_ _6103_/Y _6102_/X _6279_/S _6104_/B2 VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__o2bb2a_1
X_3316_ hold27/X hold84/X VGND VGND VPWR VPWR _5161_/A sky130_fd_sc_hd__and2_1
XFILLER_113_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7084_ _7086_/CLK hold43/X fanout482/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_1
X_4296_ hold724/X _6356_/A1 _4297_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6035_ _6940_/Q _5961_/X _6031_/X _6034_/X VGND VGND VPWR VPWR _6040_/A sky130_fd_sc_hd__a211o_1
X_3247_ _3249_/B _3250_/A VGND VGND VPWR VPWR _3247_/Y sky130_fd_sc_hd__nor2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3178_ _5552_/B VGND VGND VPWR VPWR _3178_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6937_ _7086_/CLK _6937_/D fanout483/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6868_ _6882_/CLK _6868_/D fanout475/X VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5819_ _6793_/Q _5652_/Y _5811_/X _5818_/X _6303_/S VGND VGND VPWR VPWR _5819_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6799_ _6888_/CLK _6799_/D fanout474/X VGND VGND VPWR VPWR _6799_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold570 _6987_/Q VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 _4321_/X VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold592 _6953_/Q VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1270 _4239_/X VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1281 _6650_/Q VGND VGND VPWR VPWR _4251_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1292 _4152_/X VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4150_ hold192/X _5519_/A1 _4150_/S VGND VGND VPWR VPWR _4150_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4081_ _4125_/A0 hold99/X _4118_/B VGND VGND VPWR VPWR _4081_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4983_ _5066_/A _4983_/B _4983_/C VGND VGND VPWR VPWR _4985_/D sky130_fd_sc_hd__and3_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6722_ _7150_/CLK _6722_/D fanout487/X VGND VGND VPWR VPWR _6722_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3934_ _3221_/Y _7157_/Q _6400_/B VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_2
X_6653_ _6653_/CLK _6653_/D _6401_/A VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfrtp_4
X_3865_ _3167_/Y _3251_/A _6488_/Q VGND VGND VPWR VPWR _3865_/X sky130_fd_sc_hd__mux2_1
X_5604_ _5608_/C _5604_/B VGND VGND VPWR VPWR _5604_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3796_ _6914_/Q _5355_/A _5541_/A _7079_/Q _3795_/X VGND VGND VPWR VPWR _3796_/X
+ sky130_fd_sc_hd__a221o_1
X_6584_ _7137_/CLK _6584_/D VGND VGND VPWR VPWR _6584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5535_ hold419/X _5544_/A1 _5540_/S VGND VGND VPWR VPWR _5535_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5466_ hold353/X _5526_/A1 _5471_/S VGND VGND VPWR VPWR _5466_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4417_ _4459_/B _4456_/A VGND VGND VPWR VPWR _4542_/B sky130_fd_sc_hd__nand2_4
X_5397_ hold786/X _5538_/A1 _5399_/S VGND VGND VPWR VPWR _5397_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7136_ _7140_/CLK _7136_/D VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4348_ _4376_/A _4376_/B VGND VGND VPWR VPWR _4471_/B sky130_fd_sc_hd__and2_1
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7067_ _7067_/CLK _7067_/D fanout477/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_2
X_4279_ hold964/X _5546_/A1 _4279_/S VGND VGND VPWR VPWR _4279_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6018_ _7048_/Q _5971_/A _5979_/X _6987_/Q VGND VGND VPWR VPWR _6018_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3650_ _6892_/Q _5328_/A _3981_/A _6428_/Q _3649_/X VGND VGND VPWR VPWR _3651_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3581_ _3581_/A _3581_/B _3581_/C _3581_/D VGND VGND VPWR VPWR _3582_/C sky130_fd_sc_hd__and4_2
XFILLER_115_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5320_ _5320_/A0 _5473_/A1 _5327_/S VGND VGND VPWR VPWR _5320_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5251_ _5251_/A0 _5545_/A1 _5255_/S VGND VGND VPWR VPWR _5251_/X sky130_fd_sc_hd__mux2_1
X_4202_ _4202_/A _6352_/B VGND VGND VPWR VPWR _4207_/S sky130_fd_sc_hd__and2_2
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5182_ hold990/X _5524_/A1 _5182_/S VGND VGND VPWR VPWR _5182_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4133_ _4133_/A _6352_/B VGND VGND VPWR VPWR _4138_/S sky130_fd_sc_hd__and2_2
XFILLER_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4064_ hold900/X _5548_/A1 hold37/X VGND VGND VPWR VPWR _4064_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4966_ _5088_/A _5114_/A _5088_/C VGND VGND VPWR VPWR _5008_/B sky130_fd_sc_hd__and3_1
X_6705_ _6707_/CLK _6705_/D fanout445/X VGND VGND VPWR VPWR _6705_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3917_ _6487_/Q _3916_/Y _3829_/B VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__o21a_2
X_4897_ _4900_/B _4911_/C VGND VGND VPWR VPWR _4899_/A sky130_fd_sc_hd__and2_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6636_ _7150_/CLK _6636_/D fanout487/X VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfrtp_4
X_3848_ _3866_/S _3845_/S _3847_/X _3860_/B VGND VGND VPWR VPWR _3848_/X sky130_fd_sc_hd__o211a_1
XFILLER_164_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3779_ _6426_/Q _3981_/A _6352_/A _7151_/Q _3778_/X VGND VGND VPWR VPWR _3782_/C
+ sky130_fd_sc_hd__a221o_1
X_6567_ _6653_/CLK _6567_/D _6401_/A VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5518_ hold323/X _5518_/A1 hold87/A VGND VGND VPWR VPWR _5518_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6498_ _6735_/CLK _6498_/D _3946_/B VGND VGND VPWR VPWR _6498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5449_ hold219/X _5494_/A1 _5453_/S VGND VGND VPWR VPWR _5449_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7119_ _7126_/CLK _7119_/D fanout466/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6347_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4820_ _4542_/A _4902_/A _4456_/Y _4562_/Y VGND VGND VPWR VPWR _4820_/X sky130_fd_sc_hd__o22a_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4581_/B _4948_/C _4611_/Y _4639_/Y VGND VGND VPWR VPWR _4768_/B sky130_fd_sc_hd__o22a_1
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3702_ _3701_/X _3702_/A1 _3829_/B VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__mux2_1
X_4682_ _4682_/A _4682_/B _4682_/C VGND VGND VPWR VPWR _4682_/Y sky130_fd_sc_hd__nand3_1
XFILLER_147_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6421_ _6749_/CLK _6421_/D fanout449/X VGND VGND VPWR VPWR _6421_/Q sky130_fd_sc_hd__dfstp_1
X_3633_ _6957_/Q _5400_/A _4008_/A _6453_/Q VGND VGND VPWR VPWR _3633_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6352_ _6352_/A _6352_/B VGND VGND VPWR VPWR _6357_/S sky130_fd_sc_hd__and2_2
X_3564_ _6998_/Q _5445_/A _5238_/A _6814_/Q _3563_/X VGND VGND VPWR VPWR _3565_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5303_ hold551/X _5543_/A1 _5309_/S VGND VGND VPWR VPWR _5303_/X sky130_fd_sc_hd__mux2_1
X_6283_ _6479_/Q _5940_/X _5967_/X _6608_/Q _6281_/X VGND VGND VPWR VPWR _6283_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3495_ hold74/X _3814_/B VGND VGND VPWR VPWR _4310_/A sky130_fd_sc_hd__nor2_2
X_5234_ hold451/X _5528_/A1 _5237_/S VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__mux2_1
X_5165_ _5165_/A0 _5524_/A1 _5165_/S VGND VGND VPWR VPWR _5165_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4116_ hold900/X _5548_/A1 hold38/X VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5096_ _5122_/A _5096_/B _5096_/C VGND VGND VPWR VPWR _5096_/X sky130_fd_sc_hd__and3_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4047_ hold934/X _6355_/A1 _4049_/S VGND VGND VPWR VPWR _4047_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5998_ _6858_/Q _5943_/X _5952_/X _6954_/Q _5997_/X VGND VGND VPWR VPWR _6000_/C
+ sky130_fd_sc_hd__a221o_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4949_ _4542_/A _4456_/Y _4948_/X _4946_/X VGND VGND VPWR VPWR _4963_/A sky130_fd_sc_hd__a31o_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6619_ _6712_/CLK _6619_/D fanout470/X VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput280 _6420_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
Xoutput291 _6438_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire352 _3611_/Y VGND VGND VPWR VPWR _3640_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3280_ hold63/X _6723_/Q _3975_/S VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__mux2_8
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6970_ _7063_/CLK _6970_/D fanout463/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5921_ _6464_/Q _5624_/X _5634_/X _6454_/Q _5911_/Y VGND VGND VPWR VPWR _5921_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5852_ _5852_/A _5852_/B _5852_/C VGND VGND VPWR VPWR _5852_/Y sky130_fd_sc_hd__nor3_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ _5088_/A _5088_/C _4803_/C VGND VGND VPWR VPWR _4804_/C sky130_fd_sc_hd__and3_1
XFILLER_179_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5783_ _6808_/Q _5660_/X _5667_/X _6816_/Q VGND VGND VPWR VPWR _5783_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4734_ _4735_/A _4735_/B VGND VGND VPWR VPWR _4740_/A sky130_fd_sc_hd__and2_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _4563_/A _4642_/A _4441_/B _4739_/A VGND VGND VPWR VPWR _4665_/X sky130_fd_sc_hd__a31o_1
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6404_ _3927_/A1 _6404_/D _6360_/X VGND VGND VPWR VPWR _6404_/Q sky130_fd_sc_hd__dfrtp_4
X_3616_ _6478_/Q _4038_/A _6352_/A _7154_/Q VGND VGND VPWR VPWR _3616_/X sky130_fd_sc_hd__a22o_1
Xhold900 _6530_/Q VGND VGND VPWR VPWR hold900/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold911 _5503_/X VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 _6848_/Q VGND VGND VPWR VPWR hold922/X sky130_fd_sc_hd__dlygate4sd3_1
X_4596_ _4627_/B _4562_/Y _4595_/A _4633_/B VGND VGND VPWR VPWR _4735_/B sky130_fd_sc_hd__a2bb2o_1
Xhold933 _5344_/X VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 _6554_/Q VGND VGND VPWR VPWR hold944/X sky130_fd_sc_hd__dlygate4sd3_1
X_6335_ _6644_/Q _6335_/A2 _6335_/B1 _6643_/Q VGND VGND VPWR VPWR _6335_/X sky130_fd_sc_hd__a22o_1
Xhold955 _4319_/X VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3547_ _7051_/Q _5505_/A _4322_/A _6714_/Q VGND VGND VPWR VPWR _3547_/X sky130_fd_sc_hd__a22o_1
Xhold966 _6868_/Q VGND VGND VPWR VPWR hold966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _4197_/X VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold988 _6420_/Q VGND VGND VPWR VPWR hold988/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 _6578_/Q VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__dlygate4sd3_1
X_3478_ _6959_/Q _5400_/A hold29/A hold56/A VGND VGND VPWR VPWR _3478_/X sky130_fd_sc_hd__a22o_1
X_6266_ _6653_/Q _5973_/A _5948_/X _6698_/Q _6265_/X VGND VGND VPWR VPWR _6266_/X
+ sky130_fd_sc_hd__a221o_1
X_5217_ hold683/X _5469_/A1 hold18/X VGND VGND VPWR VPWR _5217_/X sky130_fd_sc_hd__mux2_1
Xhold1600 _6535_/Q VGND VGND VPWR VPWR hold243/A sky130_fd_sc_hd__dlygate4sd3_1
X_6197_ _7034_/Q _5601_/X _5959_/X _6715_/Q VGND VGND VPWR VPWR _6197_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5148_ _5148_/A _6352_/B VGND VGND VPWR VPWR _5153_/S sky130_fd_sc_hd__and2_2
XFILLER_57_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5079_ _4902_/A _4456_/Y _4689_/B _4691_/A _4872_/A VGND VGND VPWR VPWR _5080_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4450_ _4902_/A _4948_/B _4442_/Y VGND VGND VPWR VPWR _4450_/Y sky130_fd_sc_hd__o21ai_1
Xhold207 _5461_/S VGND VGND VPWR VPWR _5462_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold218 _5386_/X VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold229 _6679_/Q VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _7062_/Q hold86/A _3981_/A _6433_/Q _3400_/X VGND VGND VPWR VPWR _3408_/A
+ sky130_fd_sc_hd__a221o_1
X_4381_ _4739_/A _4492_/D VGND VGND VPWR VPWR _4381_/Y sky130_fd_sc_hd__nand2_1
X_6120_ hold56/A _5937_/X _5975_/D _6887_/Q VGND VGND VPWR VPWR _6120_/X sky130_fd_sc_hd__a22o_1
X_3332_ _3347_/A hold73/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__nand2_8
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3263_ _3834_/B2 _3262_/Y _3261_/X VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__a21bo_1
X_6051_ _6040_/Y _6050_/X _6788_/Q _6226_/B VGND VGND VPWR VPWR _6051_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A _5002_/B _5002_/C VGND VGND VPWR VPWR _5074_/B sky130_fd_sc_hd__and3_1
X_3194_ _7021_/Q VGND VGND VPWR VPWR _3194_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6953_ _6953_/CLK _6953_/D fanout460/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5904_ _6463_/Q _5624_/X _5664_/X _6668_/Q VGND VGND VPWR VPWR _5904_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6884_ _6884_/CLK _6884_/D fanout477/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_1
X_5835_ _6705_/Q _5638_/X _5834_/X VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5766_ _6823_/Q _5818_/A2 _5814_/B1 _6911_/Q VGND VGND VPWR VPWR _5766_/X sky130_fd_sc_hd__a22o_1
X_4717_ _4482_/A _4672_/A _4902_/A _4476_/Y _4609_/Y VGND VGND VPWR VPWR _4717_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5697_ _6988_/Q _5627_/X _5635_/X _6828_/Q VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4648_ _4556_/A _4563_/A _4689_/B _5062_/A _4647_/X VGND VGND VPWR VPWR _4648_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold730 _6607_/Q VGND VGND VPWR VPWR hold730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _4320_/X VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4579_ _4579_/A _4579_/B VGND VGND VPWR VPWR _4948_/D sky130_fd_sc_hd__nand2_1
XFILLER_190_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold752 _6521_/Q VGND VGND VPWR VPWR hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _5246_/X VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 _6483_/Q VGND VGND VPWR VPWR hold774/X sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ _6320_/B _6318_/B VGND VGND VPWR VPWR _6318_/Y sky130_fd_sc_hd__nand2_1
Xhold785 _3972_/X VGND VGND VPWR VPWR _6421_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 _6476_/Q VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6249_ _7036_/Q _5601_/X _5959_/X _6717_/Q _6248_/X VGND VGND VPWR VPWR _6250_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1430 _7136_/Q VGND VGND VPWR VPWR _6311_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _7134_/Q VGND VGND VPWR VPWR _6309_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 _3976_/X VGND VGND VPWR VPWR _6423_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1463 _3303_/Y VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1474 _7139_/Q VGND VGND VPWR VPWR _6314_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk _6447_/CLK VGND VGND VPWR VPWR _7017_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1485 _7129_/Q VGND VGND VPWR VPWR _6278_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _6639_/Q VGND VGND VPWR VPWR _3881_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6707_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6629_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7080_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3950_ _3950_/A VGND VGND VPWR VPWR _3950_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3881_ _6644_/Q _3962_/B _3881_/B1 VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__a21o_1
XFILLER_149_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5620_ _7092_/Q _7093_/Q VGND VGND VPWR VPWR _5660_/C sky130_fd_sc_hd__and2b_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ _6506_/Q _6763_/Q _3177_/Y _5551_/B1 _5550_/Y VGND VGND VPWR VPWR _7087_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4502_ _4896_/B _4462_/B _4496_/B _4900_/A _4465_/B VGND VGND VPWR VPWR _4502_/X
+ sky130_fd_sc_hd__o2111a_1
X_5482_ _5482_/A0 hold666/X hold50/X VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4433_ _4607_/A _4881_/A VGND VGND VPWR VPWR _4691_/A sky130_fd_sc_hd__nand2_4
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7152_ _7155_/CLK _7152_/D fanout449/X VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4364_ _4556_/A _4441_/A VGND VGND VPWR VPWR _4690_/B sky130_fd_sc_hd__nor2_8
XFILLER_113_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6103_ _6507_/Q _7122_/Q _6103_/B1 VGND VGND VPWR VPWR _6103_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3315_ hold83/X hold64/X VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__nor2_8
X_4295_ hold958/X _6355_/A1 _4297_/S VGND VGND VPWR VPWR _4295_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7083_ _7083_/CLK _7083_/D fanout485/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3246_ _7167_/Q _3253_/S VGND VGND VPWR VPWR _3250_/A sky130_fd_sc_hd__nor2_1
X_6034_ _7012_/Q _5940_/X _5967_/X _6852_/Q _6030_/X VGND VGND VPWR VPWR _6034_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3177_ _6509_/Q VGND VGND VPWR VPWR _3177_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _7069_/CLK _6936_/D fanout482/X VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6867_ _7067_/CLK _6867_/D fanout477/X VGND VGND VPWR VPWR _6867_/Q sky130_fd_sc_hd__dfstp_1
X_5818_ _6825_/Q _5818_/A2 _5812_/X _5815_/X _5817_/X VGND VGND VPWR VPWR _5818_/X
+ sky130_fd_sc_hd__a2111o_4
X_6798_ _7049_/CLK _6798_/D fanout457/X VGND VGND VPWR VPWR _6798_/Q sky130_fd_sc_hd__dfrtp_4
X_5749_ _6846_/Q _5902_/A2 _5905_/A2 _6798_/Q _5739_/X VGND VGND VPWR VPWR _5749_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold560 _6843_/Q VGND VGND VPWR VPWR hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold571 _5438_/X VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _6474_/Q VGND VGND VPWR VPWR hold582/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold593 _5399_/X VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1260 _4087_/X VGND VGND VPWR VPWR _6510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 _6685_/Q VGND VGND VPWR VPWR _4293_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _4251_/X VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1293 _6715_/Q VGND VGND VPWR VPWR _4329_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4080_ hold405/X _4079_/X _4084_/S VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4982_ _4902_/B _4673_/A _4969_/Y _4689_/B VGND VGND VPWR VPWR _4982_/X sky130_fd_sc_hd__a31o_1
X_6721_ _3937_/A1 _6721_/D fanout487/X VGND VGND VPWR VPWR _6721_/Q sky130_fd_sc_hd__dfrtp_1
X_3933_ _6498_/Q input3/X input1/X VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__mux2_4
XFILLER_51_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6652_ _6654_/CLK _6652_/D fanout454/X VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfstp_1
X_3864_ _3866_/A1 _3863_/Y _3862_/X VGND VGND VPWR VPWR _6408_/D sky130_fd_sc_hd__a21o_1
X_5603_ _6508_/Q _5601_/X _5602_/Y _7102_/Q VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6583_ _7137_/CLK _6583_/D VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3795_ _6460_/Q _4020_/A _4008_/A _6450_/Q VGND VGND VPWR VPWR _3795_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5534_ hold261/X _5534_/A1 _5540_/S VGND VGND VPWR VPWR _5534_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5465_ hold275/X _5465_/A1 _5471_/S VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4416_ _4551_/A _4549_/B VGND VGND VPWR VPWR _4456_/A sky130_fd_sc_hd__and2_2
X_5396_ hold445/X _5528_/A1 _5399_/S VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7135_ _7140_/CLK _7135_/D VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4347_ _4702_/B _4564_/A _4347_/C VGND VGND VPWR VPWR _4376_/B sky130_fd_sc_hd__nand3_1
XFILLER_99_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7066_ _7069_/CLK _7066_/D fanout477/X VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_4
X_4278_ hold481/X _5518_/A1 _4279_/S VGND VGND VPWR VPWR _4278_/X sky130_fd_sc_hd__mux2_1
X_6017_ _6819_/Q _5953_/X _5960_/X _7072_/Q _6016_/X VGND VGND VPWR VPWR _6017_/X
+ sky130_fd_sc_hd__a221o_1
X_3229_ _4563_/A VGND VGND VPWR VPWR _4441_/A sky130_fd_sc_hd__inv_6
XFILLER_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3942_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6919_ _6999_/CLK _6919_/D fanout465/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold390 _4254_/X VGND VGND VPWR VPWR _6653_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1090 _5233_/X VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3580_ _3580_/A _3580_/B _3580_/C _3580_/D VGND VGND VPWR VPWR _3581_/D sky130_fd_sc_hd__nor4_2
XFILLER_127_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5250_ _5250_/A0 _5484_/A1 _5255_/S VGND VGND VPWR VPWR _5250_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4201_ hold942/X _5546_/A1 _4201_/S VGND VGND VPWR VPWR _4201_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5181_ hold255/X _5465_/A1 _5181_/S VGND VGND VPWR VPWR _5181_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4132_ hold608/X _6357_/A1 _4132_/S VGND VGND VPWR VPWR _4132_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4063_ hold792/X _4062_/X _4067_/S VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4965_ _4984_/A _4965_/B _5051_/A VGND VGND VPWR VPWR _5069_/B sky130_fd_sc_hd__nand3_1
X_6704_ _6704_/CLK _6704_/D fanout450/X VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_1
X_3916_ _6486_/Q _6489_/Q VGND VGND VPWR VPWR _3916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_189_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4896_ _4896_/A _4896_/B VGND VGND VPWR VPWR _4911_/C sky130_fd_sc_hd__and2_1
XFILLER_177_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6635_ _7150_/CLK _6635_/D fanout487/X VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ _6412_/Q hold70/A _3854_/S hold32/A VGND VGND VPWR VPWR _3847_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6566_ _6755_/CLK _6566_/D fanout445/X VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfrtp_4
X_3778_ _6906_/Q _5346_/A _4310_/A _6700_/Q VGND VGND VPWR VPWR _3778_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5517_ hold409/X _5544_/A1 hold87/A VGND VGND VPWR VPWR _5517_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6497_ _6990_/CLK _6497_/D fanout479/X VGND VGND VPWR VPWR _7188_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5448_ hold385/X _5526_/A1 _5453_/S VGND VGND VPWR VPWR _5448_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5379_ hold694/X _5469_/A1 _5381_/S VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7118_ _7130_/CLK _7118_/D fanout447/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7049_ _7049_/CLK _7049_/D fanout456/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4542_/D _4672_/B _4626_/Y _4628_/Y VGND VGND VPWR VPWR _4769_/A sky130_fd_sc_hd__o22a_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3701_ _3700_/Y _3764_/A1 _3829_/A VGND VGND VPWR VPWR _3701_/X sky130_fd_sc_hd__mux2_1
X_4681_ _5010_/B _4686_/B VGND VGND VPWR VPWR _4681_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6420_ _6749_/CLK _6420_/D fanout457/X VGND VGND VPWR VPWR _6420_/Q sky130_fd_sc_hd__dfstp_4
X_3632_ _6941_/Q _5382_/A _3358_/Y input14/X _3631_/X VGND VGND VPWR VPWR _3638_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6351_ _6641_/Q _6351_/A2 _5006_/A _6350_/X VGND VGND VPWR VPWR _6351_/X sky130_fd_sc_hd__o31a_1
X_3563_ _6966_/Q _5409_/A _4139_/A _6554_/Q VGND VGND VPWR VPWR _3563_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5302_ _5302_/A0 _5473_/A1 _5309_/S VGND VGND VPWR VPWR _5302_/X sky130_fd_sc_hd__mux2_1
X_6282_ _7155_/Q _5958_/X _5978_/X _6484_/Q VGND VGND VPWR VPWR _6282_/X sky130_fd_sc_hd__a22o_1
X_3494_ _6613_/Q _4208_/A _4157_/A _6569_/Q VGND VGND VPWR VPWR _3494_/X sky130_fd_sc_hd__a22o_2
XFILLER_103_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5233_ _5233_/A0 _5545_/A1 _5237_/S VGND VGND VPWR VPWR _5233_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_opt_3_0_csclk _6888_/CLK VGND VGND VPWR VPWR clkbuf_opt_3_0_csclk/X sky130_fd_sc_hd__clkbuf_16
X_5164_ _5171_/B _5164_/B hold17/X VGND VGND VPWR VPWR _5164_/X sky130_fd_sc_hd__and3_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4115_ _4115_/A0 hold42/X hold38/X VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__mux2_1
X_5095_ _5122_/C _5126_/B _5142_/B VGND VGND VPWR VPWR _5096_/C sky130_fd_sc_hd__nand3_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4046_ hold848/X _6354_/A1 _4049_/S VGND VGND VPWR VPWR _4046_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _7002_/Q _5958_/X _5975_/D _6882_/Q VGND VGND VPWR VPWR _5997_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4948_ _4948_/A _4948_/B _4948_/C _4948_/D VGND VGND VPWR VPWR _4948_/X sky130_fd_sc_hd__and4_1
X_4879_ _4902_/B _4613_/Y _4877_/X _4878_/X _4529_/Y VGND VGND VPWR VPWR _4880_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6618_ _6655_/CLK _6618_/D fanout469/X VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6549_ _6674_/CLK _6549_/D _6383_/A VGND VGND VPWR VPWR _6549_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput270 _6744_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
XFILLER_121_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput281 _6421_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
Xoutput292 _6439_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_160_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire353 _3604_/Y VGND VGND VPWR VPWR _3640_/B sky130_fd_sc_hd__clkbuf_1
Xwire364 _6225_/Y VGND VGND VPWR VPWR _6226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5920_ _6559_/Q _5667_/X _5915_/X _5916_/X _5919_/X VGND VGND VPWR VPWR _5920_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5851_ _6696_/Q _5637_/X _5848_/X _5850_/X VGND VGND VPWR VPWR _5852_/C sky130_fd_sc_hd__a211o_1
XFILLER_179_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4802_ _4689_/A _4631_/Y _4645_/Y _4846_/B VGND VGND VPWR VPWR _4803_/C sky130_fd_sc_hd__o22a_1
X_5782_ _6992_/Q _5627_/X _5637_/X _6952_/Q _5781_/X VGND VGND VPWR VPWR _5787_/B
+ sky130_fd_sc_hd__a221o_1
X_4733_ _4739_/B _4733_/B VGND VGND VPWR VPWR _4747_/C sky130_fd_sc_hd__nor2_1
XFILLER_174_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4664_ _4664_/A _4664_/B VGND VGND VPWR VPWR _4928_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6403_ _3927_/A1 _6403_/D _6359_/X VGND VGND VPWR VPWR _6403_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3615_ _7042_/Q hold76/A _5182_/S _6758_/Q _3614_/X VGND VGND VPWR VPWR _3620_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4595_ _4595_/A _4595_/B VGND VGND VPWR VPWR _4735_/A sky130_fd_sc_hd__nand2_1
Xhold901 _4116_/X VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 _6853_/Q VGND VGND VPWR VPWR hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _5281_/X VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold934 _6482_/Q VGND VGND VPWR VPWR hold934/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6334_ _6333_/X _6334_/A1 _6346_/S VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__mux2_1
Xhold945 _4144_/X VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3546_ _3546_/A hold75/X VGND VGND VPWR VPWR _4322_/A sky130_fd_sc_hd__nor2_4
XFILLER_89_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold956 _6697_/Q VGND VGND VPWR VPWR hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _5304_/X VGND VGND VPWR VPWR _6868_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold978 _6454_/Q VGND VGND VPWR VPWR hold978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 _3970_/X VGND VGND VPWR VPWR _6420_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ _6648_/Q _5976_/C _5971_/D _6568_/Q VGND VGND VPWR VPWR _6265_/X sky130_fd_sc_hd__a22o_1
X_3477_ _6999_/Q _5445_/A _5211_/A _6791_/Q _3459_/X VGND VGND VPWR VPWR _3484_/A
+ sky130_fd_sc_hd__a221o_1
X_5216_ hold118/X hold60/X hold18/X VGND VGND VPWR VPWR _5216_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6196_ _6455_/Q _5944_/X _5975_/A _6599_/Q _6195_/X VGND VGND VPWR VPWR _6200_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1601 _7132_/Q VGND VGND VPWR VPWR _6306_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5147_ hold884/X _6354_/A1 _5147_/S VGND VGND VPWR VPWR _5147_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5078_ _6724_/Q _4229_/X _5103_/B _5077_/Y _5067_/Y VGND VGND VPWR VPWR _5078_/X
+ sky130_fd_sc_hd__a221o_1
X_4029_ hold870/X _5493_/A1 hold68/X VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold208 _5458_/X VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold219 _6997_/Q VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3400_ _7070_/Q _5523_/A _5319_/A _6889_/Q VGND VGND VPWR VPWR _3400_/X sky130_fd_sc_hd__a22o_1
X_4380_ _4739_/A _4492_/D VGND VGND VPWR VPWR _4896_/B sky130_fd_sc_hd__and2_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3331_ _3379_/A hold36/X VGND VGND VPWR VPWR _3331_/Y sky130_fd_sc_hd__nor2_4
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6043_/X _6045_/X _6050_/C _6301_/C VGND VGND VPWR VPWR _6050_/X sky130_fd_sc_hd__and4bb_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _6416_/Q _3837_/A _3262_/C VGND VGND VPWR VPWR _3262_/Y sky130_fd_sc_hd__nor3_1
XFILLER_112_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5001_ _5001_/A _5001_/B _5076_/B VGND VGND VPWR VPWR _5004_/B sky130_fd_sc_hd__and3_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3193_ _7029_/Q VGND VGND VPWR VPWR _3193_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6952_ _6969_/CLK _6952_/D fanout475/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_1
X_5903_ _6617_/Q _5628_/X _5661_/X _6622_/Q _5902_/X VGND VGND VPWR VPWR _5906_/C
+ sky130_fd_sc_hd__a221o_1
X_6883_ _7067_/CLK _6883_/D fanout477/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_179_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ _7151_/Q _5625_/X _5661_/X _6619_/Q VGND VGND VPWR VPWR _5834_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5765_ _6967_/Q _5642_/X _5666_/X _6895_/Q VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4716_ _4716_/A _4965_/B _4969_/B VGND VGND VPWR VPWR _4716_/Y sky130_fd_sc_hd__nand3_2
X_5696_ _6940_/Q _5632_/X _5638_/X _6956_/Q _5694_/X VGND VGND VPWR VPWR _5711_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4647_ _4846_/B _4673_/A _4611_/Y _4628_/Y VGND VGND VPWR VPWR _4647_/X sky130_fd_sc_hd__a31o_1
XFILLER_107_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold720 _6517_/Q VGND VGND VPWR VPWR hold720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 _4206_/X VGND VGND VPWR VPWR _6607_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4578_ _4947_/B _4902_/A _4846_/B _4672_/A VGND VGND VPWR VPWR _4578_/X sky130_fd_sc_hd__a31o_1
Xhold742 _6537_/Q VGND VGND VPWR VPWR hold742/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold753 _4106_/X VGND VGND VPWR VPWR _6521_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 _6815_/Q VGND VGND VPWR VPWR hold764/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6317_ _6317_/A VGND VGND VPWR VPWR _6317_/Y sky130_fd_sc_hd__inv_2
X_3529_ _3562_/A _3573_/B VGND VGND VPWR VPWR _4151_/A sky130_fd_sc_hd__nor2_4
Xhold775 _4048_/X VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 _6951_/Q VGND VGND VPWR VPWR hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _4040_/X VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6248_ _6557_/Q _5971_/B _5949_/X _6677_/Q VGND VGND VPWR VPWR _6248_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6179_ _6179_/A0 _6178_/X _6304_/S VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1420 _6596_/Q VGND VGND VPWR VPWR hold1420/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1431 _6587_/Q VGND VGND VPWR VPWR _4183_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 _6432_/Q VGND VGND VPWR VPWR hold151/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _6947_/Q VGND VGND VPWR VPWR _5393_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 _6727_/Q VGND VGND VPWR VPWR _3830_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1475 _6590_/Q VGND VGND VPWR VPWR _4186_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 _6254_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1497 _6583_/Q VGND VGND VPWR VPWR _4179_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3880_ _6643_/Q _3962_/B _3880_/B1 VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__a21o_1
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5550_ _6506_/Q _3177_/Y _3883_/X VGND VGND VPWR VPWR _5550_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4501_ _4782_/A _5051_/B VGND VGND VPWR VPWR _4535_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5481_ hold49/X _5505_/B VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__and2_4
XFILLER_172_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4432_ _4460_/A _4632_/B VGND VGND VPWR VPWR _4969_/A sky130_fd_sc_hd__nor2_4
X_7151_ _7155_/CLK _7151_/D fanout450/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4363_ _4556_/A _4690_/A VGND VGND VPWR VPWR _4817_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6102_ _6089_/Y _6100_/X _6101_/Y _5552_/B VGND VGND VPWR VPWR _6102_/X sky130_fd_sc_hd__a211o_1
X_3314_ hold36/X _3546_/A VGND VGND VPWR VPWR _4118_/B sky130_fd_sc_hd__nor2_8
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7082_ _7082_/CLK _7082_/D fanout479/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfrtp_2
X_4294_ hold794/X _6354_/A1 _4297_/S VGND VGND VPWR VPWR _4294_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6033_ _7081_/Q _5976_/B _5971_/C _7041_/Q VGND VGND VPWR VPWR _6049_/B sky130_fd_sc_hd__a22o_1
X_3245_ _3875_/B _3244_/Y _3249_/B VGND VGND VPWR VPWR _3253_/S sky130_fd_sc_hd__a21oi_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _3176_/A VGND VGND VPWR VPWR _3176_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _6997_/CLK _6935_/D fanout465/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6866_ _6908_/CLK _6866_/D fanout475/X VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_167_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5817_ _6841_/Q _5657_/X _5660_/X _6809_/Q _5816_/X VGND VGND VPWR VPWR _5817_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6797_ _7012_/CLK _6797_/D fanout458/X VGND VGND VPWR VPWR _6797_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5748_ _5748_/A _5748_/B _5748_/C _5748_/D VGND VGND VPWR VPWR _5748_/Y sky130_fd_sc_hd__nor4_1
X_5679_ _6843_/Q _5902_/A2 _5814_/B1 _6907_/Q _5678_/X VGND VGND VPWR VPWR _5679_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold550 _5330_/X VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _5276_/X VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold572 _6907_/Q VGND VGND VPWR VPWR hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _4037_/X VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _7019_/Q VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1250 _5524_/X VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 _6680_/Q VGND VGND VPWR VPWR _4287_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1272 _4293_/X VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _6735_/Q VGND VGND VPWR VPWR _5146_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1294 _4329_/X VGND VGND VPWR VPWR _6715_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput170 wb_we_i VGND VGND VPWR VPWR _6320_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4981_ _4981_/A _4981_/B _4981_/C _4981_/D VGND VGND VPWR VPWR _4983_/C sky130_fd_sc_hd__and4_1
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3932_ _3931_/X _3953_/B _6403_/Q VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_4
XFILLER_17_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6720_ _3937_/A1 _6720_/D fanout487/X VGND VGND VPWR VPWR _6720_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6651_ _6668_/CLK _6651_/D fanout452/X VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfrtp_1
X_3863_ hold24/A _3860_/B _3866_/S VGND VGND VPWR VPWR _3863_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_176_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5602_ _5602_/A _5602_/B VGND VGND VPWR VPWR _5602_/Y sky130_fd_sc_hd__nor2_1
X_6582_ _6709_/CLK _6582_/D _6360_/A VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3794_ _3794_/A _3794_/B _3794_/C VGND VGND VPWR VPWR _3828_/A sky130_fd_sc_hd__and3_1
XFILLER_192_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5533_ _5533_/A0 hold667/X _5540_/S VGND VGND VPWR VPWR _5533_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_csclk _6447_/CLK VGND VGND VPWR VPWR _7054_/CLK sky130_fd_sc_hd__clkbuf_16
X_5464_ _5464_/A0 _5524_/A1 _5471_/S VGND VGND VPWR VPWR _5464_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4415_ _4415_/A _4415_/B VGND VGND VPWR VPWR _4549_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5395_ _5395_/A0 _5545_/A1 _5399_/S VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__mux2_1
X_7134_ _7137_/CLK _7134_/D VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfxtp_1
X_4346_ _4564_/A _4347_/C _4702_/B VGND VGND VPWR VPWR _4376_/A sky130_fd_sc_hd__a21o_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_75_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6704_/CLK sky130_fd_sc_hd__clkbuf_16
X_7065_ _7065_/CLK _7065_/D fanout465/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout359 _6301_/C VGND VGND VPWR VPWR _6226_/B sky130_fd_sc_hd__buf_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4277_ hold612/X _5544_/A1 _4279_/S VGND VGND VPWR VPWR _4277_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6016_ _6907_/Q _5973_/A _5948_/X _6947_/Q _6015_/X VGND VGND VPWR VPWR _6016_/X
+ sky130_fd_sc_hd__a221o_1
X_3228_ _6921_/Q VGND VGND VPWR VPWR _3228_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _7081_/CLK _6918_/D fanout478/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6849_ _6865_/CLK _6849_/D fanout464/X VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6990_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold380 _5442_/X VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold391 _6809_/Q VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1080 _5242_/X VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1091 _7074_/Q VGND VGND VPWR VPWR _5536_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4200_ hold501/X _5518_/A1 _4201_/S VGND VGND VPWR VPWR _4200_/X sky130_fd_sc_hd__mux2_1
X_5180_ hold129/X hold99/X _5181_/S VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4131_ hold758/X _6356_/A1 _4132_/S VGND VGND VPWR VPWR _4131_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4062_ _4115_/A0 _5538_/A1 hold37/X VGND VGND VPWR VPWR _4062_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4964_ _4964_/A _4964_/B _4964_/C VGND VGND VPWR VPWR _5005_/B sky130_fd_sc_hd__and3_1
X_6703_ _6704_/CLK _6703_/D fanout450/X VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3915_ _3954_/A _3962_/B _3908_/Y _6635_/Q VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__a22o_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4895_ _5084_/D _4895_/B _5029_/B _5085_/A VGND VGND VPWR VPWR _4918_/A sky130_fd_sc_hd__and4_1
XFILLER_149_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3846_ _3845_/X _3846_/A1 _3866_/S VGND VGND VPWR VPWR _6414_/D sky130_fd_sc_hd__mux2_1
X_6634_ _6659_/CLK _6634_/D _6383_/A VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3777_ _6970_/Q _5418_/A _3358_/Y input11/X _3776_/X VGND VGND VPWR VPWR _3782_/B
+ sky130_fd_sc_hd__a221o_1
X_6565_ _6755_/CLK _6565_/D _6360_/A VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5516_ hold600/X _5543_/A1 hold87/X VGND VGND VPWR VPWR _5516_/X sky130_fd_sc_hd__mux2_1
X_6496_ _6990_/CLK _6496_/D fanout479/X VGND VGND VPWR VPWR _7187_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5447_ hold259/X _5465_/A1 _5453_/S VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5378_ hold477/X _5528_/A1 _5381_/S VGND VGND VPWR VPWR _5378_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7117_ _7130_/CLK _7117_/D fanout447/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfrtp_1
X_4329_ _4329_/A0 _6353_/A1 _4333_/S VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7048_ _7067_/CLK _7048_/D fanout485/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3700_/A _3700_/B _3700_/C VGND VGND VPWR VPWR _3700_/Y sky130_fd_sc_hd__nand3_4
X_4680_ _4773_/A _4737_/A VGND VGND VPWR VPWR _4774_/B sky130_fd_sc_hd__nand2_1
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3631_ _6703_/Q _4310_/A _4133_/A _6548_/Q VGND VGND VPWR VPWR _3631_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6350_ _3910_/A _6350_/A2 _6317_/A _6349_/X _6320_/B VGND VGND VPWR VPWR _6350_/X
+ sky130_fd_sc_hd__a32o_1
X_3562_ _3562_/A _3562_/B VGND VGND VPWR VPWR _4139_/A sky130_fd_sc_hd__nor2_4
XFILLER_127_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5301_ _5301_/A _5505_/B VGND VGND VPWR VPWR _5309_/S sky130_fd_sc_hd__and2_4
X_6281_ _6613_/Q _5943_/X _5981_/X _6659_/Q VGND VGND VPWR VPWR _6281_/X sky130_fd_sc_hd__a22o_1
X_3493_ _3571_/A hold66/X VGND VGND VPWR VPWR _4157_/A sky130_fd_sc_hd__nor2_8
X_5232_ hold850/X _5484_/A1 _5237_/S VGND VGND VPWR VPWR _5232_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5163_ hold852/X _6354_/A1 _5163_/S VGND VGND VPWR VPWR _5163_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4114_ hold812/X _5546_/A1 hold38/X VGND VGND VPWR VPWR _4114_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5094_ _4948_/C _4946_/X _5058_/A _5093_/X _4818_/X VGND VGND VPWR VPWR _5142_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4045_ _4045_/A0 _5491_/A1 _4049_/S VGND VGND VPWR VPWR _4045_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5996_ _7079_/Q _5976_/B _5975_/C _6834_/Q _5995_/X VGND VGND VPWR VPWR _6000_/B
+ sky130_fd_sc_hd__a221o_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4947_ _4947_/A _4947_/B _4947_/C VGND VGND VPWR VPWR _5043_/B sky130_fd_sc_hd__nand3_2
X_4878_ _5083_/A _5029_/A _4878_/C VGND VGND VPWR VPWR _4878_/X sky130_fd_sc_hd__and3_1
X_6617_ _6769_/CLK _6617_/D fanout469/X VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3829_ _3829_/A _3829_/B VGND VGND VPWR VPWR _3829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6548_ _6735_/CLK _6548_/D fanout445/X VGND VGND VPWR VPWR _6548_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_192_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6479_ _6707_/CLK _6479_/D _3946_/B VGND VGND VPWR VPWR _6479_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_161_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput260 _6750_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
Xoutput271 _6434_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
Xoutput282 _6435_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
XFILLER_121_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput293 _6440_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XFILLER_181_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire354 _3504_/Y VGND VGND VPWR VPWR _3582_/A sky130_fd_sc_hd__clkbuf_1
Xwire365 _6200_/Y VGND VGND VPWR VPWR _6201_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_183_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5850_ _6566_/Q _5635_/X _5661_/X _6620_/Q _5849_/X VGND VGND VPWR VPWR _5850_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _4673_/B _4700_/Y _4707_/Y _4799_/X _4800_/X VGND VGND VPWR VPWR _4804_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5781_ _6848_/Q _5902_/A2 _5654_/X _6936_/Q VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4732_ _4428_/Y _4611_/Y _4500_/A VGND VGND VPWR VPWR _5114_/B sky130_fd_sc_hd__a21o_1
XFILLER_159_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4663_ _4716_/A _4686_/B VGND VGND VPWR VPWR _4663_/Y sky130_fd_sc_hd__nand2_2
X_3614_ _6745_/Q _5154_/A _3585_/Y input95/X VGND VGND VPWR VPWR _3614_/X sky130_fd_sc_hd__a22o_1
X_6402_ _3927_/A1 _6402_/D _6358_/X VGND VGND VPWR VPWR _6402_/Q sky130_fd_sc_hd__dfrtp_4
X_4594_ _4563_/A _4661_/A _4441_/B _4631_/D VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__a31o_1
XFILLER_190_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold902 _6719_/Q VGND VGND VPWR VPWR hold902/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 _5287_/X VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3545_ _6958_/Q _5400_/A _4127_/A _6544_/Q _3544_/X VGND VGND VPWR VPWR _3552_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold924 _6968_/Q VGND VGND VPWR VPWR hold924/X sky130_fd_sc_hd__dlygate4sd3_1
X_6333_ _6642_/Q _6333_/A2 _6333_/B1 _6350_/A2 _6332_/X VGND VGND VPWR VPWR _6333_/X
+ sky130_fd_sc_hd__a221o_1
Xhold935 _4047_/X VGND VGND VPWR VPWR _6482_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _6564_/Q VGND VGND VPWR VPWR hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _4307_/X VGND VGND VPWR VPWR _6697_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _6477_/Q VGND VGND VPWR VPWR hold968/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6264_ _6264_/A _6264_/B _6264_/C VGND VGND VPWR VPWR _6276_/C sky130_fd_sc_hd__nor3_1
XFILLER_142_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3476_ _6879_/Q _5310_/A hold49/A _7031_/Q _3475_/X VGND VGND VPWR VPWR _3485_/B
+ sky130_fd_sc_hd__a221oi_1
Xhold979 _4013_/X VGND VGND VPWR VPWR _6454_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5215_ hold225/X _5494_/A1 hold18/X VGND VGND VPWR VPWR _5215_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6195_ _6465_/Q _5937_/X _5975_/D _6625_/Q VGND VGND VPWR VPWR _6195_/X sky130_fd_sc_hd__a22o_1
X_5146_ _5146_/A0 _5491_/A1 _5147_/S VGND VGND VPWR VPWR _5146_/X sky130_fd_sc_hd__mux2_1
Xhold1602 _7123_/Q VGND VGND VPWR VPWR _6128_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5077_ _5077_/A _5103_/C _5077_/C VGND VGND VPWR VPWR _5077_/Y sky130_fd_sc_hd__nand3_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4028_ _4028_/A0 _5492_/A1 hold68/X VGND VGND VPWR VPWR _4028_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5979_ _5979_/A _5981_/A _5979_/C VGND VGND VPWR VPWR _5979_/X sky130_fd_sc_hd__and3_4
XFILLER_40_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 _6758_/Q VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_166_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3330_ _3543_/A _3373_/B VGND VGND VPWR VPWR _5391_/A sky130_fd_sc_hd__nor2_8
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _6417_/Q _6415_/Q _6485_/Q _3164_/Y VGND VGND VPWR VPWR _3261_/X sky130_fd_sc_hd__a31o_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _4948_/C _4582_/Y _4941_/D _4991_/X VGND VGND VPWR VPWR _5076_/B sky130_fd_sc_hd__o211a_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3192_ _6445_/Q VGND VGND VPWR VPWR _3192_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6951_ _6951_/CLK _6951_/D fanout474/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5902_ _6602_/Q _5902_/A2 _5634_/X _6453_/Q VGND VGND VPWR VPWR _5902_/X sky130_fd_sc_hd__a22o_1
X_6882_ _6882_/CLK _6882_/D fanout475/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfstp_1
X_5833_ _6560_/Q _5631_/X _5830_/X _5832_/X VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__a211o_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5764_ _7015_/Q _5630_/X _5761_/X _5762_/X _5763_/X VGND VGND VPWR VPWR _5764_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_147_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4715_ _4469_/A _4714_/X _4713_/X _5084_/C _5062_/B VGND VGND VPWR VPWR _4722_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_30_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5695_ _7020_/Q _5619_/X _5663_/X _6860_/Q VGND VGND VPWR VPWR _5695_/X sky130_fd_sc_hd__a22o_1
X_4646_ _4646_/A _4707_/C VGND VGND VPWR VPWR _4646_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold710 _6959_/Q VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4577_ _4672_/A _4902_/A VGND VGND VPWR VPWR _4723_/B sky130_fd_sc_hd__nor2_1
Xhold721 _4101_/X VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 _7188_/A VGND VGND VPWR VPWR hold732/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold743 _4124_/X VGND VGND VPWR VPWR _6537_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 _6745_/Q VGND VGND VPWR VPWR hold754/X sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ _6320_/B _6316_/A2 _6640_/Q VGND VGND VPWR VPWR _6317_/A sky130_fd_sc_hd__a21bo_1
X_3528_ _6438_/Q _3372_/Y hold76/A _7043_/Q _3527_/X VGND VGND VPWR VPWR _3538_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold765 _5244_/X VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 _6478_/Q VGND VGND VPWR VPWR hold776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _5397_/X VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold798 _6886_/Q VGND VGND VPWR VPWR hold798/X sky130_fd_sc_hd__dlygate4sd3_1
X_6247_ _6457_/Q _5944_/X _5975_/A _6601_/Q _6246_/X VGND VGND VPWR VPWR _6250_/C
+ sky130_fd_sc_hd__a221o_1
X_3459_ _6799_/Q _3326_/Y _4102_/A _7200_/A VGND VGND VPWR VPWR _3459_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6178_ _6178_/A0 _6177_/X _6303_/S VGND VGND VPWR VPWR _6178_/X sky130_fd_sc_hd__mux2_1
Xhold1410 _6424_/Q VGND VGND VPWR VPWR _3978_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1421 _6598_/Q VGND VGND VPWR VPWR hold1421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 _6574_/Q VGND VGND VPWR VPWR _4168_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1443 _3988_/X VGND VGND VPWR VPWR _6432_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5129_ _5113_/X _5129_/B _5129_/C _5129_/D VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__nand4b_1
Xhold1454 _6730_/Q VGND VGND VPWR VPWR _3642_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 _6433_/Q VGND VGND VPWR VPWR hold557/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1476 _6597_/Q VGND VGND VPWR VPWR _4194_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _6414_/Q VGND VGND VPWR VPWR _3846_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 _6486_/Q VGND VGND VPWR VPWR _3911_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4500_ _4500_/A _4689_/A VGND VGND VPWR VPWR _4500_/Y sky130_fd_sc_hd__nor2_1
XFILLER_191_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5480_ _5480_/A0 hold22/X hold30/X VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__mux2_1
XFILLER_184_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 _7157_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4431_ _4753_/A _4460_/A VGND VGND VPWR VPWR _4881_/A sky130_fd_sc_hd__nor2_2
XFILLER_172_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4362_ _4911_/A _4489_/A VGND VGND VPWR VPWR _4500_/A sky130_fd_sc_hd__nand2_8
X_7150_ _7150_/CLK _7150_/D _6307_/B VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfrtp_1
X_6101_ _6790_/Q _6226_/B VGND VGND VPWR VPWR _6101_/Y sky130_fd_sc_hd__nor2_1
X_3313_ _3313_/A _3454_/A VGND VGND VPWR VPWR _3546_/A sky130_fd_sc_hd__nand2_8
X_7081_ _7081_/CLK _7081_/D fanout485/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_1
X_4293_ _4293_/A0 _5491_/A1 _4297_/S VGND VGND VPWR VPWR _4293_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3244_ _3875_/C _3260_/S VGND VGND VPWR VPWR _3244_/Y sky130_fd_sc_hd__nor2_1
X_6032_ _7057_/Q _5954_/X _5976_/D _6876_/Q VGND VGND VPWR VPWR _6049_/A sky130_fd_sc_hd__a22o_1
XFILLER_140_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3175_ _7089_/Q VGND VGND VPWR VPWR _3886_/B sky130_fd_sc_hd__inv_2
XFILLER_67_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6934_ _7081_/CLK _6934_/D fanout478/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6865_ _6865_/CLK _6865_/D fanout465/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5816_ _7025_/Q _5619_/X _5663_/X _6865_/Q VGND VGND VPWR VPWR _5816_/X sky130_fd_sc_hd__a22o_1
X_6796_ _7011_/CLK _6796_/D fanout456/X VGND VGND VPWR VPWR _6796_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5747_ _6822_/Q _5818_/A2 _5814_/B1 _6910_/Q _5746_/X VGND VGND VPWR VPWR _5748_/D
+ sky130_fd_sc_hd__a221o_1
X_5678_ _6899_/Q _5621_/X _5818_/A2 _6819_/Q VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4629_ _4716_/A _4975_/A _4698_/C VGND VGND VPWR VPWR _5099_/B sky130_fd_sc_hd__nand3_2
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold540 _4049_/X VGND VGND VPWR VPWR _6484_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold551 _6867_/Q VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _6582_/Q VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold573 _5348_/X VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _7009_/Q VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold595 _5474_/X VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1240 _5515_/X VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1251 _6625_/Q VGND VGND VPWR VPWR _4233_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1262 _4287_/X VGND VGND VPWR VPWR _6680_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 _6705_/Q VGND VGND VPWR VPWR _4317_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1284 _5146_/X VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1295 _6604_/Q VGND VGND VPWR VPWR _4203_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6342_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4980_ _4619_/Y _4970_/Y _4975_/Y _4644_/Y _5062_/A VGND VGND VPWR VPWR _4981_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3931_ _3930_/X input38/X _6405_/Q VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_1
X_6650_ _6668_/CLK _6650_/D fanout452/X VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfrtp_2
X_3862_ _3167_/Y _3866_/S _3860_/B hold24/A VGND VGND VPWR VPWR _3862_/X sky130_fd_sc_hd__o211a_1
X_5601_ _5968_/A _5964_/A _5981_/A VGND VGND VPWR VPWR _5601_/X sky130_fd_sc_hd__and3_4
XFILLER_176_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6581_ _6709_/CLK _6581_/D fanout445/X VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfrtp_4
X_3793_ _3793_/A _3793_/B _3793_/C _3793_/D VGND VGND VPWR VPWR _3794_/C sky130_fd_sc_hd__nor4_1
XFILLER_118_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5532_ _5532_/A _5541_/B VGND VGND VPWR VPWR _5540_/S sky130_fd_sc_hd__and2_4
XFILLER_192_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_csclk _6601_/CLK VGND VGND VPWR VPWR _6659_/CLK sky130_fd_sc_hd__clkbuf_16
X_5463_ _5463_/A hold17/X VGND VGND VPWR VPWR _5471_/S sky130_fd_sc_hd__and2_4
XFILLER_132_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4414_ _4459_/B _4579_/A VGND VGND VPWR VPWR _4542_/A sky130_fd_sc_hd__nand2_8
X_5394_ hold363/X _5526_/A1 _5399_/S VGND VGND VPWR VPWR _5394_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7133_ _7137_/CLK _7133_/D VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4345_ _4631_/D _4633_/B _4661_/A _4357_/B VGND VGND VPWR VPWR _4347_/C sky130_fd_sc_hd__and4_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4276_ hold421/X _5534_/A1 _4279_/S VGND VGND VPWR VPWR _4276_/X sky130_fd_sc_hd__mux2_1
X_7064_ _7067_/CLK _7064_/D fanout477/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_100_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3227_ _6792_/Q VGND VGND VPWR VPWR _3227_/Y sky130_fd_sc_hd__inv_2
X_6015_ _6899_/Q _5976_/C _5971_/D _6827_/Q VGND VGND VPWR VPWR _6015_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6917_ _7085_/CLK _6917_/D fanout477/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6848_ _7069_/CLK _6848_/D fanout482/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6779_ _6969_/CLK _6779_/D fanout473/X VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold370 _5268_/X VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _6796_/Q VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold392 _5237_/X VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1070 _5377_/X VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 _7082_/Q VGND VGND VPWR VPWR _5545_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 _5536_/X VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4130_ hold952/X _6355_/A1 _4132_/S VGND VGND VPWR VPWR _4130_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4061_ _4061_/A0 _4060_/X _4067_/S VGND VGND VPWR VPWR _4061_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4963_ _4963_/A _4963_/B VGND VGND VPWR VPWR _4963_/Y sky130_fd_sc_hd__nand2_1
X_6702_ _7155_/CLK _6702_/D fanout450/X VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfstp_1
X_3914_ _3837_/B _3875_/X _3875_/B _6488_/Q VGND VGND VPWR VPWR _6487_/D sky130_fd_sc_hd__a2bb2o_1
X_4894_ _4689_/A _4631_/Y _5034_/B _4518_/C VGND VGND VPWR VPWR _5085_/A sky130_fd_sc_hd__o211a_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6633_ _6659_/CLK _6633_/D fanout469/X VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3845_ _3288_/Y hold33/A _3845_/S VGND VGND VPWR VPWR _3845_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6564_ _6674_/CLK _6564_/D _6383_/A VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfrtp_1
X_3776_ _6994_/Q _5445_/A _3367_/Y input20/X VGND VGND VPWR VPWR _3776_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5515_ _5515_/A0 hold667/X hold87/A VGND VGND VPWR VPWR _5515_/X sky130_fd_sc_hd__mux2_1
X_6495_ _6990_/CLK _6495_/D fanout478/X VGND VGND VPWR VPWR _7186_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5446_ _5446_/A0 _5524_/A1 _5453_/S VGND VGND VPWR VPWR _5446_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5377_ _5377_/A0 _5545_/A1 _5381_/S VGND VGND VPWR VPWR _5377_/X sky130_fd_sc_hd__mux2_1
X_7116_ _7130_/CLK _7116_/D fanout447/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4328_ _4328_/A _5490_/B VGND VGND VPWR VPWR _4333_/S sky130_fd_sc_hd__and2_2
XFILLER_87_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7047_ _7049_/CLK _7047_/D fanout457/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfstp_1
X_4259_ hold642/X _5544_/A1 _4261_/S VGND VGND VPWR VPWR _4259_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6747_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3630_ _6789_/Q _5211_/A _4044_/A _6483_/Q _3629_/X VGND VGND VPWR VPWR _3638_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3561_ _6934_/Q _5373_/A _5154_/A _6746_/Q _3560_/X VGND VGND VPWR VPWR _3565_/B
+ sky130_fd_sc_hd__a221o_1
X_5300_ hold606/X _5513_/A1 _5300_/S VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3492_ _3562_/A _3814_/B VGND VGND VPWR VPWR _4208_/A sky130_fd_sc_hd__nor2_8
X_6280_ _6664_/Q _5976_/B _5971_/C _6714_/Q VGND VGND VPWR VPWR _6280_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5231_ hold537/X _5543_/A1 _5237_/S VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5162_ _5162_/A0 _6353_/A1 _5163_/S VGND VGND VPWR VPWR _5162_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_csclk _6601_/CLK VGND VGND VPWR VPWR _6671_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4113_ hold692/X _5509_/A1 hold38/X VGND VGND VPWR VPWR _4113_/X sky130_fd_sc_hd__mux2_1
X_5093_ _4672_/B _4496_/Y _4456_/Y VGND VGND VPWR VPWR _5093_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4044_ _4044_/A _6352_/B VGND VGND VPWR VPWR _4049_/S sky130_fd_sc_hd__and2_2
XFILLER_83_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7081_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5995_ _7055_/Q _5954_/X _5976_/C _6898_/Q VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4946_ _4947_/A _4947_/B _4947_/C VGND VGND VPWR VPWR _4946_/X sky130_fd_sc_hd__and3_2
XFILLER_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _4877_/A _4877_/B _4877_/C _4877_/D VGND VGND VPWR VPWR _4877_/X sky130_fd_sc_hd__and4_1
X_6616_ _6655_/CLK _6616_/D fanout469/X VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfstp_1
X_3828_ _3828_/A _3828_/B VGND VGND VPWR VPWR _3828_/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6547_ _6654_/CLK _6547_/D fanout454/X VGND VGND VPWR VPWR _6547_/Q sky130_fd_sc_hd__dfrtp_2
X_3759_ input72/X _3331_/Y _4238_/A _6631_/Q _3758_/X VGND VGND VPWR VPWR _3760_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6478_ _6704_/CLK _6478_/D fanout448/X VGND VGND VPWR VPWR _6478_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5429_ hold299/X _5465_/A1 _5435_/S VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput250 _3944_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
Xoutput261 _6736_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
Xoutput272 _6428_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
Xoutput283 _6422_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
Xoutput294 _6441_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XFILLER_58_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire355 _3467_/Y VGND VGND VPWR VPWR _3486_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire366 _6049_/Y VGND VGND VPWR VPWR _6050_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_183_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_124_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4902_/B _4673_/A _4616_/Y VGND VGND VPWR VPWR _4800_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5780_ _6832_/Q _5635_/X _5928_/A2 _6840_/Q _5779_/X VGND VGND VPWR VPWR _5787_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4538_/X _4683_/X _4730_/X _5006_/A _4731_/B2 VGND VGND VPWR VPWR _6720_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4662_ _4686_/B VGND VGND VPWR VPWR _4662_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6401_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__and2_1
X_3613_ _6965_/Q _5409_/A _3367_/Y input23/X _3612_/X VGND VGND VPWR VPWR _3620_/A
+ sky130_fd_sc_hd__a221o_1
X_4593_ _4920_/B VGND VGND VPWR VPWR _4593_/Y sky130_fd_sc_hd__inv_2
Xhold903 _4333_/X VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold914 _6845_/Q VGND VGND VPWR VPWR hold914/X sky130_fd_sc_hd__dlygate4sd3_1
X_6332_ _6644_/Q _6332_/A2 _6332_/B1 _6643_/Q VGND VGND VPWR VPWR _6332_/X sky130_fd_sc_hd__a22o_1
X_3544_ _6878_/Q _5310_/A _4328_/A _6719_/Q VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__a22o_1
Xhold925 _5416_/X VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _6606_/Q VGND VGND VPWR VPWR hold936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 _4156_/X VGND VGND VPWR VPWR _6564_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold958 _6687_/Q VGND VGND VPWR VPWR hold958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 _4041_/X VGND VGND VPWR VPWR _6477_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6263_ _6463_/Q _5945_/X _5975_/C _6581_/Q _6262_/X VGND VGND VPWR VPWR _6264_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3475_ _6919_/Q _5355_/A _5238_/A _6815_/Q _3474_/X VGND VGND VPWR VPWR _3475_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5214_ _5214_/A0 hold6/X hold18/X VGND VGND VPWR VPWR _5214_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6194_ _6680_/Q _5934_/X _5975_/B _6614_/Q _6193_/X VGND VGND VPWR VPWR _6200_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1603 _7126_/Q VGND VGND VPWR VPWR _6203_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5145_ _5145_/A _6352_/B VGND VGND VPWR VPWR _5147_/S sky130_fd_sc_hd__and2_1
XFILLER_57_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5076_ _5076_/A _5076_/B _5076_/C VGND VGND VPWR VPWR _5077_/C sky130_fd_sc_hd__and3_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4027_ _4027_/A0 _6353_/A1 hold68/X VGND VGND VPWR VPWR _4027_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5978_ _5978_/A _5981_/A _5979_/C VGND VGND VPWR VPWR _5978_/X sky130_fd_sc_hd__and3_4
XFILLER_52_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4929_ _4673_/A _4613_/Y _4772_/A _4928_/Y VGND VGND VPWR VPWR _5002_/C sky130_fd_sc_hd__o211a_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmgmt_gpio_9_buff_inst _3927_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_8
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3260_ _3251_/A _3260_/A1 _3260_/S VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__mux2_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _7042_/Q VGND VGND VPWR VPWR _3191_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6950_ _7067_/CLK _6950_/D fanout476/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5901_ _6607_/Q _5648_/X _5663_/X _6612_/Q _5900_/X VGND VGND VPWR VPWR _5906_/B
+ sky130_fd_sc_hd__a221o_1
X_6881_ _7070_/CLK _6881_/D fanout473/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_4
X_5832_ _6645_/Q _5621_/X _5648_/X _6604_/Q _5831_/X VGND VGND VPWR VPWR _5832_/X
+ sky130_fd_sc_hd__a221o_1
X_5763_ _6951_/Q _5637_/X _5645_/X _7031_/Q VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4714_ _4633_/B _4627_/A _4479_/Y _4619_/Y _4645_/Y VGND VGND VPWR VPWR _4714_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5694_ _7004_/Q _5625_/X _5661_/X _6876_/Q VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4645_ _4716_/A _4645_/B VGND VGND VPWR VPWR _4645_/Y sky130_fd_sc_hd__nand2_8
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold700 _6977_/Q VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 _5406_/X VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4576_ _4965_/B _4576_/B VGND VGND VPWR VPWR _4576_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold722 _6800_/Q VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold733 _4067_/X VGND VGND VPWR VPWR _6497_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6315_ _3410_/Y _6315_/A1 _6315_/S VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__mux2_1
Xhold744 _6449_/Q VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__dlygate4sd3_1
X_3527_ _6942_/Q _5382_/A _5211_/A _6790_/Q VGND VGND VPWR VPWR _3527_/X sky130_fd_sc_hd__a22o_1
Xhold755 _5158_/X VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold766 _6782_/Q VGND VGND VPWR VPWR hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _4042_/X VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold788 _6887_/Q VGND VGND VPWR VPWR hold788/X sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _6467_/Q _5937_/X _5975_/D _6627_/Q VGND VGND VPWR VPWR _6246_/X sky130_fd_sc_hd__a22o_1
Xhold799 _5324_/X VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3458_ input17/X _3358_/Y _3372_/Y _6439_/Q VGND VGND VPWR VPWR _3458_/X sky130_fd_sc_hd__a22o_2
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6177_ _6793_/Q _6226_/B _6176_/X VGND VGND VPWR VPWR _6177_/X sky130_fd_sc_hd__o21ba_1
XFILLER_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3389_ _6929_/Q _5364_/A _3365_/Y input10/X _3386_/X VGND VGND VPWR VPWR _3392_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1400 _7031_/Q VGND VGND VPWR VPWR _5487_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 _7173_/A VGND VGND VPWR VPWR _5173_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 _6585_/Q VGND VGND VPWR VPWR hold1422/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5128_ _5142_/A _5126_/X _5142_/C _5123_/Y VGND VGND VPWR VPWR _5129_/C sky130_fd_sc_hd__a31o_1
Xhold1433 _7140_/Q VGND VGND VPWR VPWR _6315_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1444 _6624_/Q VGND VGND VPWR VPWR _3963_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 _3642_/X VGND VGND VPWR VPWR _6730_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 _3989_/X VGND VGND VPWR VPWR _6433_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1477 _6734_/Q VGND VGND VPWR VPWR _3413_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5059_ _5058_/X _5122_/A VGND VGND VPWR VPWR _5059_/X sky130_fd_sc_hd__and2b_1
Xhold1488 _6636_/Q VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _3911_/X VGND VGND VPWR VPWR _6486_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__buf_12
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4430_ _5068_/A VGND VGND VPWR VPWR _4430_/Y sky130_fd_sc_hd__inv_2
XANTENNA_2 _5190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4361_ _4911_/A _4489_/A VGND VGND VPWR VPWR _4685_/A sky130_fd_sc_hd__and2_1
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6100_ _6092_/X _6094_/X _6100_/C _6301_/C VGND VGND VPWR VPWR _6100_/X sky130_fd_sc_hd__and4bb_2
XFILLER_125_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3312_ hold26/X hold46/X VGND VGND VPWR VPWR _3454_/A sky130_fd_sc_hd__and2b_4
XFILLER_112_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7080_ _7080_/CLK _7080_/D fanout479/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfstp_1
X_4292_ _4292_/A _5490_/B VGND VGND VPWR VPWR _4297_/S sky130_fd_sc_hd__and2_2
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6031_ _7004_/Q _5958_/X _5978_/X _6996_/Q VGND VGND VPWR VPWR _6031_/X sky130_fd_sc_hd__a22o_1
X_3243_ _6487_/Q _3837_/C VGND VGND VPWR VPWR _3260_/S sky130_fd_sc_hd__nand2_8
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3174_ _6763_/Q VGND VGND VPWR VPWR _3174_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6933_ _7082_/CLK _6933_/D fanout483/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6864_ _6951_/CLK _6864_/D fanout474/X VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5815_ _6817_/Q _5667_/X _5813_/X _5814_/X VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__a211o_1
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6795_ _6963_/CLK _6795_/D fanout456/X VGND VGND VPWR VPWR _6795_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5746_ _6998_/Q _5643_/X _5652_/B _6918_/Q _5651_/Y VGND VGND VPWR VPWR _5746_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5677_ _6795_/Q _5905_/A2 _5660_/X _6803_/Q VGND VGND VPWR VPWR _5677_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4628_ _4661_/A _4716_/A _4653_/B VGND VGND VPWR VPWR _4628_/Y sky130_fd_sc_hd__nand3_4
XFILLER_190_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold530 _4207_/X VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4559_ _5088_/B _4559_/B _4721_/A VGND VGND VPWR VPWR _4559_/X sky130_fd_sc_hd__and3_1
Xhold541 _6875_/Q VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold552 _5303_/X VGND VGND VPWR VPWR _6867_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _4177_/X VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_9_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold574 _6439_/Q VGND VGND VPWR VPWR hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold585 _5462_/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold596 _6562_/Q VGND VGND VPWR VPWR hold596/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6229_ _6229_/A0 _6228_/X _6279_/S VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1230 _5497_/X VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1241 _6710_/Q VGND VGND VPWR VPWR _4323_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _4233_/X VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1263 _6480_/Q VGND VGND VPWR VPWR _4045_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1274 _4317_/X VGND VGND VPWR VPWR _6705_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 _6609_/Q VGND VGND VPWR VPWR _4209_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 _4203_/X VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6330_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6345_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3930_ _6499_/Q _6734_/Q _6400_/B VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3861_ _3861_/A _3861_/B VGND VGND VPWR VPWR _6409_/D sky130_fd_sc_hd__xnor2_1
XFILLER_189_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5600_ _5600_/A _7102_/Q VGND VGND VPWR VPWR _5981_/A sky130_fd_sc_hd__nor2_8
XFILLER_176_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6580_ _6677_/CLK _6580_/D fanout452/X VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3792_ _6442_/Q _3999_/A _5182_/S _7087_/Q _3791_/X VGND VGND VPWR VPWR _3793_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5531_ hold176/X hold22/X _5531_/S VGND VGND VPWR VPWR _5531_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5462_ hold584/X _5513_/A1 _5462_/S VGND VGND VPWR VPWR _5462_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4413_ _4549_/A _4579_/A VGND VGND VPWR VPWR _4413_/Y sky130_fd_sc_hd__nand2_8
X_5393_ _5393_/A0 hold13/X _5399_/S VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__mux2_1
X_7132_ _7150_/CLK _7132_/D fanout487/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_141_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4344_ _4631_/D _4661_/A _4357_/B VGND VGND VPWR VPWR _4352_/B sky130_fd_sc_hd__nand3_1
XFILLER_125_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7063_ _7063_/CLK _7063_/D fanout463/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_98_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4275_ _4275_/A0 hold667/X _4279_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6014_ _6014_/A _6014_/B _6014_/C VGND VGND VPWR VPWR _6014_/Y sky130_fd_sc_hd__nor3_1
X_3226_ _6919_/Q VGND VGND VPWR VPWR _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6916_ _7081_/CLK _6916_/D fanout478/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6847_ _6951_/CLK _6847_/D fanout474/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6778_ _6969_/CLK _6778_/D fanout473/X VGND VGND VPWR VPWR _6778_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5729_ _7021_/Q _5619_/X _5663_/X _6861_/Q VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold360 _5178_/X VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold371 _7065_/Q VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _5223_/X VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _7180_/A VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1060 _5341_/X VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 _6821_/Q VGND VGND VPWR VPWR _5251_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 _5545_/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 _6748_/Q VGND VGND VPWR VPWR _5162_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_200 _4102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4060_ hold812/X _5546_/A1 hold37/X VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4962_ _4950_/X _4962_/B _4962_/C VGND VGND VPWR VPWR _4963_/B sky130_fd_sc_hd__and3b_1
XFILLER_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6701_ _7155_/CLK _6701_/D fanout449/X VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_1
X_3913_ _3164_/Y _3165_/Y _3868_/S _3867_/B _6488_/Q VGND VGND VPWR VPWR _6488_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4893_ _4893_/A VGND VGND VPWR VPWR _5034_/B sky130_fd_sc_hd__inv_2
X_6632_ _6632_/CLK _6632_/D fanout454/X VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfstp_2
X_3844_ hold32/A _6412_/Q hold70/A _3854_/S VGND VGND VPWR VPWR _3845_/S sky130_fd_sc_hd__nand4_1
XFILLER_149_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6563_ _6674_/CLK _6563_/D _6383_/A VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfrtp_1
X_3775_ _6922_/Q _5364_/A _5274_/A _6842_/Q _3774_/X VGND VGND VPWR VPWR _3782_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5514_ hold86/X _5541_/B VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__and2_4
XFILLER_118_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6494_ _7079_/CLK _6494_/D fanout478/X VGND VGND VPWR VPWR _7185_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5445_ _5445_/A hold17/X VGND VGND VPWR VPWR _5453_/S sky130_fd_sc_hd__and2_4
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5376_ hold864/X _5484_/A1 _5381_/S VGND VGND VPWR VPWR _5376_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7115_ _7130_/CLK _7115_/D fanout447/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4327_ hold826/X _5546_/A1 _4327_/S VGND VGND VPWR VPWR _4327_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7046_ _7086_/CLK _7046_/D fanout483/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfrtp_4
X_4258_ hold427/X _5534_/A1 _4261_/S VGND VGND VPWR VPWR _4258_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3209_ _6901_/Q VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__inv_2
X_4189_ _3762_/Y _4189_/A1 _4195_/S VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold190 _6830_/Q VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_csclk _6601_/CLK VGND VGND VPWR VPWR _6769_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3560_ _6674_/Q _4274_/A _4133_/A _6549_/Q VGND VGND VPWR VPWR _3560_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3491_ input56/X _5193_/A _5274_/A _6846_/Q _3490_/X VGND VGND VPWR VPWR _3504_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5230_ _5230_/A0 _5473_/A1 _5237_/S VGND VGND VPWR VPWR _5230_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5161_ _5161_/A _5190_/B hold16/X VGND VGND VPWR VPWR _5163_/S sky130_fd_sc_hd__and3_4
XFILLER_170_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4112_ _4112_/A0 hold6/X hold38/A VGND VGND VPWR VPWR _4112_/X sky130_fd_sc_hd__mux2_1
X_5092_ _5092_/A _5092_/B _5092_/C VGND VGND VPWR VPWR _5126_/B sky130_fd_sc_hd__and3_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4043_ hold533/X _6357_/A1 _4043_/S VGND VGND VPWR VPWR _4043_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5994_ _7063_/Q _5934_/X _5973_/A _6906_/Q _5993_/X VGND VGND VPWR VPWR _6000_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4945_ _4930_/X _4944_/X _5069_/A VGND VGND VPWR VPWR _4945_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4876_ _4623_/Y _4700_/Y _4864_/X _4875_/X _4523_/Y VGND VGND VPWR VPWR _4877_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_149_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3827_ _3798_/X _3827_/B _3827_/C _3827_/D VGND VGND VPWR VPWR _3828_/B sky130_fd_sc_hd__and4b_1
X_6615_ _7036_/CLK _6615_/D fanout455/X VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6546_ _6677_/CLK _6546_/D fanout452/X VGND VGND VPWR VPWR _6546_/Q sky130_fd_sc_hd__dfrtp_1
X_3758_ _6891_/Q _5328_/A _5541_/A _7080_/Q VGND VGND VPWR VPWR _3758_/X sky130_fd_sc_hd__a22o_2
XFILLER_180_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6477_ _6707_/CLK _6477_/D fanout450/X VGND VGND VPWR VPWR _6477_/Q sky130_fd_sc_hd__dfstp_1
X_3689_ _6948_/Q _5391_/A _5400_/A _6956_/Q VGND VGND VPWR VPWR _3689_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5428_ _5428_/A0 _5524_/A1 _5435_/S VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput240 _3919_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
Xoutput251 _3951_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
Xoutput262 _6737_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
Xoutput273 _6429_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
Xoutput284 _6423_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
X_5359_ _5359_/A0 _5545_/A1 _5363_/S VGND VGND VPWR VPWR _5359_/X sky130_fd_sc_hd__mux2_1
Xoutput295 _6426_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7029_ _7082_/CLK _7029_/D fanout483/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire356 _3446_/Y VGND VGND VPWR VPWR _3447_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_137_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire367 _5748_/Y VGND VGND VPWR VPWR wire367/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4730_ _5039_/A _4589_/Y _4729_/X VGND VGND VPWR VPWR _4730_/X sky130_fd_sc_hd__a21o_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4661_ _4661_/A _4661_/B VGND VGND VPWR VPWR _4686_/B sky130_fd_sc_hd__and2_2
XFILLER_187_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6400_ _6400_/A _6400_/B VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__and2_1
X_3612_ _6445_/Q _3999_/A _4322_/A _6713_/Q VGND VGND VPWR VPWR _3612_/X sky130_fd_sc_hd__a22o_2
X_4592_ _4565_/X _4601_/A _6643_/Q VGND VGND VPWR VPWR _4920_/B sky130_fd_sc_hd__o21a_1
XFILLER_190_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold904 _6781_/Q VGND VGND VPWR VPWR hold904/X sky130_fd_sc_hd__dlygate4sd3_1
X_6331_ _6330_/X _6331_/A1 _6346_/S VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__mux2_1
X_3543_ _3543_/A _3577_/B VGND VGND VPWR VPWR _4328_/A sky130_fd_sc_hd__nor2_4
Xhold915 _5278_/X VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _7085_/Q VGND VGND VPWR VPWR hold926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _4205_/X VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 _6472_/Q VGND VGND VPWR VPWR hold948/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 _4295_/X VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _6668_/Q _5938_/X _5952_/X _6708_/Q VGND VGND VPWR VPWR _6262_/X sky130_fd_sc_hd__a22o_1
X_3474_ _6927_/Q _5364_/A _3999_/A _6447_/Q _3473_/X VGND VGND VPWR VPWR _3474_/X
+ sky130_fd_sc_hd__a221o_2
X_5213_ hold251/X _5465_/A1 hold18/X VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6193_ _6700_/Q _5971_/A _5979_/X _6470_/Q VGND VGND VPWR VPWR _6193_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5144_ _5123_/A _5142_/Y _5143_/Y _5136_/X VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__a211o_1
XFILLER_130_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5075_ _4428_/Y _4456_/Y _4846_/B _4689_/B _4768_/A VGND VGND VPWR VPWR _5076_/C
+ sky130_fd_sc_hd__o221a_1
X_4026_ hold67/X _5490_/B VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__and2_2
XFILLER_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ _5977_/A _5977_/B _5977_/C VGND VGND VPWR VPWR _6301_/C sky130_fd_sc_hd__nand3_4
X_4928_ _4928_/A _4984_/B VGND VGND VPWR VPWR _4928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4859_ _4947_/C _4689_/A _4500_/A VGND VGND VPWR VPWR _5023_/C sky130_fd_sc_hd__a21o_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6529_ _6990_/CLK hold55/X fanout478/X VGND VGND VPWR VPWR _6529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_73_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7155_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_csclk _6601_/CLK VGND VGND VPWR VPWR _6674_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7051_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _7050_/Q VGND VGND VPWR VPWR _3190_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5900_ _6468_/Q _5619_/X _5652_/B _5899_/Y VGND VGND VPWR VPWR _5900_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6880_ _7069_/CLK _6880_/D fanout482/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5831_ _6614_/Q _5628_/X _5910_/B1 _6625_/Q VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5762_ _6943_/Q _5632_/X _5638_/X _6959_/Q _5759_/X VGND VGND VPWR VPWR _5762_/X
+ sky130_fd_sc_hd__a221o_1
X_4713_ _5041_/B _4576_/Y _4712_/X _4711_/X VGND VGND VPWR VPWR _4713_/X sky130_fd_sc_hd__a31o_1
X_5693_ _5713_/A0 _5692_/X _6279_/S VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4644_ _4716_/A _4644_/B VGND VGND VPWR VPWR _4644_/Y sky130_fd_sc_hd__nand2_4
XFILLER_147_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold701 _5426_/X VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ _4574_/A _4574_/B _4551_/A VGND VGND VPWR VPWR _4575_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_162_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold712 _6943_/Q VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 _5227_/X VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 _6581_/Q VGND VGND VPWR VPWR hold734/X sky130_fd_sc_hd__dlygate4sd3_1
X_3526_ _6798_/Q _3326_/Y _3981_/A _6430_/Q _3525_/X VGND VGND VPWR VPWR _3538_/A
+ sky130_fd_sc_hd__a221o_1
X_6314_ _3447_/Y _6314_/A1 _6315_/S VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold745 _4007_/X VGND VGND VPWR VPWR _6449_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 _6458_/Q VGND VGND VPWR VPWR hold756/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 _5207_/X VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _6473_/Q VGND VGND VPWR VPWR hold778/X sky130_fd_sc_hd__dlygate4sd3_1
X_6245_ _6682_/Q _5934_/X _5975_/B _6616_/Q _6244_/X VGND VGND VPWR VPWR _6250_/B
+ sky130_fd_sc_hd__a221o_1
X_3457_ input8/X _3365_/Y _3367_/Y input25/X VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__a22o_1
Xhold789 _5325_/X VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6176_ _6168_/X _6226_/B _6176_/C _6176_/D VGND VGND VPWR VPWR _6176_/X sky130_fd_sc_hd__and4b_2
XFILLER_162_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3388_ input60/X _5193_/A _3326_/Y _6801_/Q _3385_/X VGND VGND VPWR VPWR _3392_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1401 _6881_/Q VGND VGND VPWR VPWR _5318_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 _6576_/Q VGND VGND VPWR VPWR hold1412/X sky130_fd_sc_hd__dlygate4sd3_1
X_5127_ _4948_/B _5042_/Y _5043_/Y _4948_/D VGND VGND VPWR VPWR _5142_/C sky130_fd_sc_hd__o22a_1
Xhold1423 _6590_/Q VGND VGND VPWR VPWR hold1423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _7135_/Q VGND VGND VPWR VPWR _6310_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1445 _3965_/X VGND VGND VPWR VPWR hold665/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1456 _6728_/Q VGND VGND VPWR VPWR _3764_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1467 _6440_/Q VGND VGND VPWR VPWR _3997_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5058_ _5058_/A _5122_/B _5058_/C _5058_/D VGND VGND VPWR VPWR _5058_/X sky130_fd_sc_hd__and4_1
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1478 _6596_/Q VGND VGND VPWR VPWR _4193_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1489 _7122_/Q VGND VGND VPWR VPWR _6078_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _4009_/A0 _6353_/A1 _4013_/S VGND VGND VPWR VPWR _4009_/X sky130_fd_sc_hd__mux2_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__buf_6
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__buf_6
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 _5346_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4360_ _4359_/Y _4360_/B _4379_/B VGND VGND VPWR VPWR _4489_/A sky130_fd_sc_hd__and3b_2
X_3311_ hold34/X _3323_/B _3311_/C VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__nand3_2
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4291_ hold186/X _5519_/A1 _4291_/S VGND VGND VPWR VPWR _4291_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6030_ _6860_/Q _5943_/X _5981_/X _6916_/Q VGND VGND VPWR VPWR _6030_/X sky130_fd_sc_hd__a22o_1
X_3242_ _6488_/Q _6485_/Q VGND VGND VPWR VPWR _3837_/C sky130_fd_sc_hd__nor2_4
XFILLER_79_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3173_ _6813_/Q VGND VGND VPWR VPWR _3173_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6932_ _7067_/CLK _6932_/D fanout476/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6863_ _6865_/CLK _6863_/D fanout465/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5814_ _6449_/Q _5614_/X _5814_/B1 _6913_/Q VGND VGND VPWR VPWR _5814_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6794_ _7006_/CLK _6794_/D fanout458/X VGND VGND VPWR VPWR _6794_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_10_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5745_ hold79/A _5614_/X _5664_/X _6926_/Q _5738_/X VGND VGND VPWR VPWR _5748_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5676_ _6443_/Q _5614_/X _5625_/X _7003_/Q _5675_/X VGND VGND VPWR VPWR _5681_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4627_ _4627_/A _4627_/B VGND VGND VPWR VPWR _4703_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold520 _4289_/X VGND VGND VPWR VPWR _6682_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _6689_/Q VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _4563_/A _4484_/Y _5088_/C VGND VGND VPWR VPWR _4721_/A sky130_fd_sc_hd__o21a_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold542 _5312_/X VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _6746_/Q VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _6741_/Q VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold575 _3996_/X VGND VGND VPWR VPWR _6439_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _6484_/Q _4044_/A _4250_/A _6654_/Q _3508_/X VGND VGND VPWR VPWR _3523_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold586 _6438_/Q VGND VGND VPWR VPWR hold586/X sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _4489_/A _4489_/B VGND VGND VPWR VPWR _4490_/B sky130_fd_sc_hd__nand2_1
Xhold597 _4154_/X VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6228_ _7127_/Q _6227_/X _6303_/S VGND VGND VPWR VPWR _6228_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _7009_/Q _5958_/X _5978_/X _7001_/Q VGND VGND VPWR VPWR _6159_/X sky130_fd_sc_hd__a22o_1
Xhold1220 _5506_/X VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1231 _7071_/Q VGND VGND VPWR VPWR _5533_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 _4323_/X VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1253 _6778_/Q VGND VGND VPWR VPWR _5203_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 _4045_/X VGND VGND VPWR VPWR _6480_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 _6695_/Q VGND VGND VPWR VPWR _4305_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1286 _4209_/X VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1297 hold1589/X VGND VGND VPWR VPWR _4119_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6326_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6332_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6324_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3860_ hold81/A _3860_/B VGND VGND VPWR VPWR _3861_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3791_ _6750_/Q _3355_/X _5164_/B _3365_/Y input34/X VGND VGND VPWR VPWR _3791_/X
+ sky130_fd_sc_hd__a32o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5530_ hold938/X _5548_/A1 _5531_/S VGND VGND VPWR VPWR _5530_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5461_ hold164/X hold99/X _5461_/S VGND VGND VPWR VPWR _5461_/X sky130_fd_sc_hd__mux2_1
X_4412_ _4551_/A _4959_/A VGND VGND VPWR VPWR _4579_/A sky130_fd_sc_hd__and2_4
X_7200_ _7200_/A VGND VGND VPWR VPWR _7200_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5392_ _5392_/A0 _5524_/A1 _5399_/S VGND VGND VPWR VPWR _5392_/X sky130_fd_sc_hd__mux2_1
X_7131_ _7131_/CLK _7131_/D fanout459/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_1
X_4343_ _4556_/A _4563_/A _4753_/A _4607_/A VGND VGND VPWR VPWR _4357_/B sky130_fd_sc_hd__o211a_2
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7062_ _7086_/CLK _7062_/D fanout483/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfrtp_1
X_4274_ _4274_/A _4322_/B VGND VGND VPWR VPWR _4279_/S sky130_fd_sc_hd__and2_2
XFILLER_98_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6013_ _6979_/Q _5945_/X _5975_/C _6835_/Q _6012_/X VGND VGND VPWR VPWR _6014_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3225_ _6659_/Q VGND VGND VPWR VPWR _3225_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6915_ _6981_/CLK _6915_/D fanout463/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6846_ _7051_/CLK _6846_/D fanout476/X VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6777_ _6777_/CLK _6777_/D fanout483/X VGND VGND VPWR VPWR _7196_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3989_ hold557/X _5513_/A1 _3989_/S VGND VGND VPWR VPWR _3989_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5728_ _6973_/Q _5634_/X _5722_/X _5723_/X _5727_/X VGND VGND VPWR VPWR _5728_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5659_ _6834_/Q _5928_/A2 _5910_/B1 _6882_/Q VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold350 _4078_/X VGND VGND VPWR VPWR _6502_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold361 _6628_/Q VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold372 _5526_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _6523_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _4095_/X VGND VGND VPWR VPWR _6514_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1050 _5277_/X VGND VGND VPWR VPWR _6844_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 _6938_/Q VGND VGND VPWR VPWR _5383_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _5251_/X VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 _7029_/Q VGND VGND VPWR VPWR _5485_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 _5162_/X VGND VGND VPWR VPWR _6748_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _5614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4961_ _4957_/Y _5046_/B _5088_/D _5039_/D VGND VGND VPWR VPWR _4962_/C sky130_fd_sc_hd__and4b_1
XFILLER_17_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6700_ _6704_/CLK _6700_/D fanout449/X VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3912_ _3912_/A1 _6485_/Q _3875_/B _3912_/B1 VGND VGND VPWR VPWR _6489_/D sky130_fd_sc_hd__a31o_1
X_4892_ _4892_/A _4892_/B VGND VGND VPWR VPWR _4893_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6631_ _6632_/CLK _6631_/D fanout454/X VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfrtp_4
X_3843_ hold62/A hold81/A hold24/A hold44/A VGND VGND VPWR VPWR _3854_/S sky130_fd_sc_hd__and4_1
XFILLER_177_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6562_ _6674_/CLK _6562_/D _6383_/A VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfstp_2
X_3774_ _6818_/Q _5247_/A _4298_/A _6690_/Q VGND VGND VPWR VPWR _3774_/X sky130_fd_sc_hd__a22o_2
XFILLER_164_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5513_ hold650/X _5513_/A1 _5513_/S VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__mux2_1
X_6493_ _6527_/CLK _6493_/D fanout484/X VGND VGND VPWR VPWR _7184_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_118_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5444_ hold685/X _5513_/A1 _5444_/S VGND VGND VPWR VPWR _5444_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5375_ hold295/X _5465_/A1 _5381_/S VGND VGND VPWR VPWR _5375_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7114_ _7130_/CLK _7114_/D fanout448/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4326_ hold303/X _5518_/A1 _4327_/S VGND VGND VPWR VPWR _4326_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4257_ _4257_/A0 hold667/X _4261_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
X_7045_ _7085_/CLK _7045_/D fanout485/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfrtp_1
X_3208_ _6909_/Q VGND VGND VPWR VPWR _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4188_ _3828_/Y _4188_/A1 _4195_/S VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6829_ _6967_/CLK _6829_/D fanout474/X VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold180 _6862_/Q VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _5261_/X VGND VGND VPWR VPWR _6830_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3490_ _6902_/Q _5337_/A _4232_/A _6629_/Q VGND VGND VPWR VPWR _3490_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5160_ hold545/X _5469_/A1 _5160_/S VGND VGND VPWR VPWR _5160_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4111_ hold622/X _5543_/A1 hold38/X VGND VGND VPWR VPWR _4111_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5091_ _4584_/A _5043_/B _5090_/Y VGND VGND VPWR VPWR _5092_/C sky130_fd_sc_hd__a21oi_1
XFILLER_96_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4042_ hold776/X _6356_/A1 _4043_/S VGND VGND VPWR VPWR _4042_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5993_ _6978_/Q _5945_/X _5978_/X _6994_/Q VGND VGND VPWR VPWR _5993_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4944_ _4944_/A _4944_/B _4944_/C VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__and3_1
X_4875_ _4875_/A _5034_/A _4875_/C VGND VGND VPWR VPWR _4875_/X sky130_fd_sc_hd__and3_1
XFILLER_177_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6614_ _7036_/CLK _6614_/D fanout455/X VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfrtp_1
X_3826_ _3826_/A _3826_/B _3826_/C _3826_/D VGND VGND VPWR VPWR _3826_/Y sky130_fd_sc_hd__nor4_1
XFILLER_165_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6545_ _6709_/CLK _6545_/D fanout445/X VGND VGND VPWR VPWR _6545_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3757_ input21/X _3367_/Y _4038_/A _6476_/Q _3756_/X VGND VGND VPWR VPWR _3760_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6476_ _6746_/CLK _6476_/D _3946_/B VGND VGND VPWR VPWR _6476_/Q sky130_fd_sc_hd__dfrtp_4
X_3688_ _3688_/A _3688_/B _3688_/C VGND VGND VPWR VPWR _3699_/C sky130_fd_sc_hd__nor3_1
X_5427_ _5427_/A hold17/X VGND VGND VPWR VPWR _5435_/S sky130_fd_sc_hd__and2_4
Xoutput230 _7192_/X VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
Xoutput241 _3918_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
Xoutput252 _3948_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput263 _6738_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
Xoutput274 _6430_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput285 _6424_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5358_ hold874/X _5484_/A1 _5363_/S VGND VGND VPWR VPWR _5358_/X sky130_fd_sc_hd__mux2_1
Xoutput296 _6427_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4309_ hold578/X _6357_/A1 _4309_/S VGND VGND VPWR VPWR _4309_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5289_ hold702/X _5469_/A1 _5291_/S VGND VGND VPWR VPWR _5289_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7028_ _7080_/CLK _7028_/D fanout479/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire346 _3538_/Y VGND VGND VPWR VPWR _3581_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire357 _3408_/Y VGND VGND VPWR VPWR wire357/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire379 _5976_/Y VGND VGND VPWR VPWR _5977_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_152_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4660_ _4660_/A _4660_/B _4660_/C _4660_/D VGND VGND VPWR VPWR _4660_/X sky130_fd_sc_hd__and4_1
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3611_ _3611_/A _3611_/B _3611_/C _3611_/D VGND VGND VPWR VPWR _3611_/Y sky130_fd_sc_hd__nor4_1
XFILLER_175_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4591_ _4591_/A _4664_/B VGND VGND VPWR VPWR _4601_/A sky130_fd_sc_hd__nand2_1
XFILLER_190_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6330_ _6644_/Q _6330_/A2 _6330_/B1 _6643_/Q _6329_/X VGND VGND VPWR VPWR _6330_/X
+ sky130_fd_sc_hd__a221o_1
X_3542_ _3546_/A _3714_/B VGND VGND VPWR VPWR _4127_/A sky130_fd_sc_hd__nor2_4
Xhold905 _5206_/X VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold916 _6861_/Q VGND VGND VPWR VPWR hold916/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold927 _5548_/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold938 _7069_/Q VGND VGND VPWR VPWR hold938/X sky130_fd_sc_hd__dlygate4sd3_1
X_3473_ _7007_/Q _3370_/Y _5182_/S _3450_/X VGND VGND VPWR VPWR _3473_/X sky130_fd_sc_hd__a22o_1
Xhold949 _4035_/X VGND VGND VPWR VPWR _6472_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6261_ _6453_/Q _5947_/X _5965_/X _6548_/Q _6260_/X VGND VGND VPWR VPWR _6264_/B
+ sky130_fd_sc_hd__a221o_1
X_5212_ _5212_/A0 _5524_/A1 hold18/X VGND VGND VPWR VPWR _5212_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6192_ _6560_/Q _5953_/X _5960_/X _6670_/Q _6191_/X VGND VGND VPWR VPWR _6192_/X
+ sky130_fd_sc_hd__a221o_1
X_5143_ _5143_/A _5143_/B VGND VGND VPWR VPWR _5143_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5074_ _5074_/A _5074_/B _5074_/C VGND VGND VPWR VPWR _5103_/C sky130_fd_sc_hd__and3_1
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4025_ hold213/X hold60/X _4025_/S VGND VGND VPWR VPWR _4025_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5976_ _5981_/A _5976_/B _5976_/C _5976_/D VGND VGND VPWR VPWR _5976_/Y sky130_fd_sc_hd__nor4_1
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4927_ _4542_/B _4562_/Y _4771_/A VGND VGND VPWR VPWR _4995_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4858_ _4482_/B _4694_/Y _4529_/Y VGND VGND VPWR VPWR _4858_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3809_ _6930_/Q _5373_/A _4151_/A _6560_/Q _3808_/X VGND VGND VPWR VPWR _3817_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4789_ _4672_/A _4620_/Y _4701_/Y _4710_/Y VGND VGND VPWR VPWR _4789_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6528_ _7079_/CLK _6528_/D fanout478/X VGND VGND VPWR VPWR _6528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7038_/CLK sky130_fd_sc_hd__clkbuf_16
X_6459_ _6704_/CLK _6459_/D fanout448/X VGND VGND VPWR VPWR _6459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5830_ _6480_/Q _5643_/X _5664_/X _6665_/Q VGND VGND VPWR VPWR _5830_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5761_ _6847_/Q _5902_/A2 _5905_/A2 _6799_/Q _5760_/X VGND VGND VPWR VPWR _5761_/X
+ sky130_fd_sc_hd__a221o_1
X_4712_ _4691_/A _4673_/B _4710_/Y VGND VGND VPWR VPWR _4712_/X sky130_fd_sc_hd__o21a_1
X_5692_ _7106_/Q _5691_/X _6303_/S VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4643_ _4653_/C _4661_/B VGND VGND VPWR VPWR _4643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4574_ _4574_/A _4574_/B VGND VGND VPWR VPWR _4574_/Y sky130_fd_sc_hd__nand2_1
Xhold702 _6855_/Q VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _5388_/X VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold724 _6688_/Q VGND VGND VPWR VPWR hold724/X sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ _3486_/Y _6313_/A1 _6315_/S VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold735 _4176_/X VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3525_ input16/X _3358_/Y _4202_/A _6608_/Q VGND VGND VPWR VPWR _3525_/X sky130_fd_sc_hd__a22o_1
Xhold746 _6825_/Q VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 _4018_/X VGND VGND VPWR VPWR _6458_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold768 _7154_/Q VGND VGND VPWR VPWR hold768/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6244_ _6702_/Q _5971_/A _5979_/X _6472_/Q VGND VGND VPWR VPWR _6244_/X sky130_fd_sc_hd__a22o_2
Xhold779 _4036_/X VGND VGND VPWR VPWR _6473_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3456_ _6991_/Q _5436_/A hold76/A _7044_/Q VGND VGND VPWR VPWR _3456_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3387_ _7001_/Q _5445_/A _5373_/A _6937_/Q _3382_/X VGND VGND VPWR VPWR _3392_/A
+ sky130_fd_sc_hd__a221o_1
X_6175_ _6175_/A _6175_/B _6175_/C _6175_/D VGND VGND VPWR VPWR _6176_/D sky130_fd_sc_hd__nor4_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1402 _6468_/Q VGND VGND VPWR VPWR _4030_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5126_ _5126_/A _5126_/B _5126_/C VGND VGND VPWR VPWR _5126_/X sky130_fd_sc_hd__and3_1
Xhold1413 _6577_/Q VGND VGND VPWR VPWR hold1413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 _7139_/Q VGND VGND VPWR VPWR hold1424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 _6570_/Q VGND VGND VPWR VPWR _4164_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1446 _7133_/Q VGND VGND VPWR VPWR _6308_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1457 _3764_/X VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5057_ _5057_/A _5057_/B _5057_/C VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__and3_1
Xhold1468 _6577_/Q VGND VGND VPWR VPWR _4171_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1479 _6585_/Q VGND VGND VPWR VPWR _4181_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4008_ _4008_/A _4322_/B VGND VGND VPWR VPWR _4013_/S sky130_fd_sc_hd__and2_2
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5959_ _5959_/A _5981_/A VGND VGND VPWR VPWR _5959_/X sky130_fd_sc_hd__and2_4
XFILLER_185_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__buf_6
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_4 _5310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3310_ _3374_/A _3370_/A VGND VGND VPWR VPWR _5310_/A sky130_fd_sc_hd__nor2_8
X_4290_ hold377/X _5518_/A1 _4291_/S VGND VGND VPWR VPWR _4290_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3241_ _7169_/Q _7168_/Q VGND VGND VPWR VPWR _3875_/C sky130_fd_sc_hd__nor2_1
XFILLER_112_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3172_ _6485_/Q VGND VGND VPWR VPWR _3867_/A sky130_fd_sc_hd__inv_2
XFILLER_79_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6931_ _6963_/CLK _6931_/D fanout458/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6862_ _7079_/CLK _6862_/D fanout480/X VGND VGND VPWR VPWR _6862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5813_ _6969_/Q _5642_/X _5666_/X _6897_/Q VGND VGND VPWR VPWR _5813_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6793_ _7053_/CLK _6793_/D fanout459/X VGND VGND VPWR VPWR _6793_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5744_ _6854_/Q _5648_/X _5666_/X _6894_/Q _5743_/X VGND VGND VPWR VPWR _5748_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5675_ _6995_/Q _5643_/X _5645_/X _7027_/Q VGND VGND VPWR VPWR _5675_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_72_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6749_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4626_ _4753_/B _4626_/B VGND VGND VPWR VPWR _4626_/Y sky130_fd_sc_hd__nand2_8
Xhold510 _4242_/X VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold521 _6984_/Q VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _4557_/A VGND VGND VPWR VPWR _4967_/A sky130_fd_sc_hd__inv_2
Xhold532 _4297_/X VGND VGND VPWR VPWR _6689_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _7064_/Q VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold554 _5159_/X VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _7006_/Q _3370_/Y _4292_/A _6689_/Q VGND VGND VPWR VPWR _3508_/X sky130_fd_sc_hd__a22o_2
Xhold565 _5153_/X VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 _6961_/Q VGND VGND VPWR VPWR hold576/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4488_ _4600_/B _4611_/B VGND VGND VPWR VPWR _4672_/B sky130_fd_sc_hd__nand2_8
Xhold587 _3995_/X VGND VGND VPWR VPWR _6438_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold598 _7050_/Q VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ _6541_/Q _6226_/B _6226_/X VGND VGND VPWR VPWR _6227_/X sky130_fd_sc_hd__o21ba_1
X_3439_ _6920_/Q _5355_/A _5247_/A _6824_/Q _3438_/X VGND VGND VPWR VPWR _3446_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6865_/Q _5943_/X _5981_/X _6921_/Q VGND VGND VPWR VPWR _6158_/X sky130_fd_sc_hd__a22o_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _5221_/X VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _6986_/Q VGND VGND VPWR VPWR _5437_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_csclk _6601_/CLK VGND VGND VPWR VPWR _6655_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1232 _5533_/X VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 _6655_/Q VGND VGND VPWR VPWR _4257_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5109_ _5135_/A _5109_/B _5135_/B VGND VGND VPWR VPWR _5109_/Y sky130_fd_sc_hd__nand3_2
X_6089_ _6089_/A _6089_/B _6089_/C VGND VGND VPWR VPWR _6089_/Y sky130_fd_sc_hd__nor3_2
Xhold1254 _5203_/X VGND VGND VPWR VPWR _6778_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1265 _6614_/Q VGND VGND VPWR VPWR _4215_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 _4305_/X VGND VGND VPWR VPWR _6695_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 _6450_/Q VGND VGND VPWR VPWR _4009_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _4119_/X VGND VGND VPWR VPWR _6532_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7067_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4337_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6329_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6335_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6326_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3790_ _6986_/Q _5436_/A _5145_/A _6735_/Q _3789_/X VGND VGND VPWR VPWR _3793_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5460_ hold648/X _5469_/A1 _5462_/S VGND VGND VPWR VPWR _5460_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4411_ _4739_/A _4415_/A VGND VGND VPWR VPWR _4959_/A sky130_fd_sc_hd__and2_1
X_5391_ _5391_/A _5505_/B VGND VGND VPWR VPWR _5399_/S sky130_fd_sc_hd__and2_4
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7130_ _7130_/CLK _7130_/D fanout486/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4342_ _4556_/A _4563_/A VGND VGND VPWR VPWR _4753_/B sky130_fd_sc_hd__nor2_8
XFILLER_99_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7061_ _7082_/CLK _7061_/D fanout483/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfrtp_1
X_4273_ hold227/X hold60/X _4273_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6012_ _6923_/Q _5938_/X _5952_/X _6955_/Q VGND VGND VPWR VPWR _6012_/X sky130_fd_sc_hd__a22o_1
.ends

