magic
tech sky130A
magscale 1 2
timestamp 1675162573
<< viali >>
rect 3249 8585 3283 8619
rect 5825 8585 5859 8619
rect 3893 8517 3927 8551
rect 6469 8517 6503 8551
rect 1777 8449 1811 8483
rect 2605 8381 2639 8415
rect 4721 8381 4755 8415
rect 7297 8381 7331 8415
rect 1777 8041 1811 8075
rect 2237 7837 2271 7871
rect 3893 7837 3927 7871
rect 5733 7837 5767 7871
rect 3065 7769 3099 7803
rect 4721 7769 4755 7803
rect 6561 7769 6595 7803
rect 7113 7701 7147 7735
rect 1593 7497 1627 7531
rect 4077 7497 4111 7531
rect 5549 7497 5583 7531
rect 3525 7429 3559 7463
rect 2697 7361 2731 7395
rect 6469 7361 6503 7395
rect 4629 7293 4663 7327
rect 7297 7293 7331 7327
rect 2145 7225 2179 7259
rect 4905 6817 4939 6851
rect 6561 6817 6595 6851
rect 1869 6749 1903 6783
rect 2697 6749 2731 6783
rect 4077 6681 4111 6715
rect 6009 6681 6043 6715
rect 7389 6681 7423 6715
rect 3249 6613 3283 6647
rect 1685 6409 1719 6443
rect 3617 6341 3651 6375
rect 4261 6341 4295 6375
rect 7297 6341 7331 6375
rect 2789 6273 2823 6307
rect 5917 6273 5951 6307
rect 6469 6273 6503 6307
rect 5365 6137 5399 6171
rect 2329 6069 2363 6103
rect 4813 6069 4847 6103
rect 5917 5865 5951 5899
rect 3985 5729 4019 5763
rect 6469 5661 6503 5695
rect 4813 5593 4847 5627
rect 5273 5593 5307 5627
rect 7297 5593 7331 5627
rect 1501 5525 1535 5559
rect 2237 5525 2271 5559
rect 2789 5525 2823 5559
rect 3249 5525 3283 5559
rect 4445 5253 4479 5287
rect 5181 5253 5215 5287
rect 6561 5253 6595 5287
rect 3617 5185 3651 5219
rect 5917 5185 5951 5219
rect 7389 5185 7423 5219
rect 2053 5049 2087 5083
rect 2605 4981 2639 5015
rect 3065 4981 3099 5015
rect 5365 4777 5399 4811
rect 3249 4641 3283 4675
rect 2421 4573 2455 4607
rect 6469 4573 6503 4607
rect 3893 4505 3927 4539
rect 4721 4505 4755 4539
rect 7205 4505 7239 4539
rect 1869 4437 1903 4471
rect 6009 4437 6043 4471
rect 4445 4165 4479 4199
rect 6469 4165 6503 4199
rect 3617 4097 3651 4131
rect 5089 4097 5123 4131
rect 5825 4097 5859 4131
rect 3065 4029 3099 4063
rect 7297 4029 7331 4063
rect 1961 3893 1995 3927
rect 2513 3893 2547 3927
rect 5457 3689 5491 3723
rect 4721 3553 4755 3587
rect 7297 3553 7331 3587
rect 3341 3485 3375 3519
rect 6469 3485 6503 3519
rect 2605 3417 2639 3451
rect 3893 3417 3927 3451
rect 1961 3349 1995 3383
rect 6009 3349 6043 3383
rect 2329 3077 2363 3111
rect 3341 3077 3375 3111
rect 4169 3077 4203 3111
rect 6469 3077 6503 3111
rect 1501 3009 1535 3043
rect 4629 3009 4663 3043
rect 7297 3009 7331 3043
rect 5457 2941 5491 2975
rect 5457 2601 5491 2635
rect 6009 2533 6043 2567
rect 2605 2465 2639 2499
rect 4721 2465 4755 2499
rect 7297 2465 7331 2499
rect 3341 2397 3375 2431
rect 6469 2397 6503 2431
rect 3893 2329 3927 2363
rect 1961 2261 1995 2295
rect 1777 2057 1811 2091
rect 3617 1989 3651 2023
rect 4353 1989 4387 2023
rect 5181 1989 5215 2023
rect 5917 1989 5951 2023
rect 6469 1989 6503 2023
rect 7297 1989 7331 2023
rect 2237 1921 2271 1955
rect 3065 1921 3099 1955
rect 2605 1377 2639 1411
rect 4169 1377 4203 1411
rect 1961 1309 1995 1343
rect 4905 1309 4939 1343
rect 7297 1309 7331 1343
rect 3341 1241 3375 1275
rect 6469 1241 6503 1275
rect 5365 1173 5399 1207
<< metal1 >>
rect 3418 8848 3424 8900
rect 3476 8888 3482 8900
rect 7374 8888 7380 8900
rect 3476 8860 7380 8888
rect 3476 8848 3482 8860
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 1012 8730 8071 8752
rect 1012 8678 2582 8730
rect 2634 8678 2646 8730
rect 2698 8678 2710 8730
rect 2762 8678 2774 8730
rect 2826 8678 2838 8730
rect 2890 8678 4307 8730
rect 4359 8678 4371 8730
rect 4423 8678 4435 8730
rect 4487 8678 4499 8730
rect 4551 8678 4563 8730
rect 4615 8678 6032 8730
rect 6084 8678 6096 8730
rect 6148 8678 6160 8730
rect 6212 8678 6224 8730
rect 6276 8678 6288 8730
rect 6340 8678 7757 8730
rect 7809 8678 7821 8730
rect 7873 8678 7885 8730
rect 7937 8678 7949 8730
rect 8001 8678 8013 8730
rect 8065 8678 8071 8730
rect 1012 8656 8071 8678
rect 934 8576 940 8628
rect 992 8616 998 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 992 8588 3249 8616
rect 992 8576 998 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 3252 8548 3280 8579
rect 3694 8576 3700 8628
rect 3752 8616 3758 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 3752 8588 5825 8616
rect 3752 8576 3758 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 5813 8579 5871 8585
rect 3881 8551 3939 8557
rect 3881 8548 3893 8551
rect 3252 8520 3893 8548
rect 3881 8517 3893 8520
rect 3927 8517 3939 8551
rect 5828 8548 5856 8579
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 5828 8520 6469 8548
rect 3881 8511 3939 8517
rect 6457 8517 6469 8520
rect 6503 8517 6515 8551
rect 6457 8511 6515 8517
rect 1762 8480 1768 8492
rect 1723 8452 1768 8480
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 4614 8412 4620 8424
rect 2639 8384 4620 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 5442 8412 5448 8424
rect 4755 8384 5448 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7466 8412 7472 8424
rect 7331 8384 7472 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 5258 8276 5264 8288
rect 5040 8248 5264 8276
rect 5040 8236 5046 8248
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 1012 8186 7912 8208
rect 1012 8134 1720 8186
rect 1772 8134 1784 8186
rect 1836 8134 1848 8186
rect 1900 8134 1912 8186
rect 1964 8134 1976 8186
rect 2028 8134 3445 8186
rect 3497 8134 3509 8186
rect 3561 8134 3573 8186
rect 3625 8134 3637 8186
rect 3689 8134 3701 8186
rect 3753 8134 5170 8186
rect 5222 8134 5234 8186
rect 5286 8134 5298 8186
rect 5350 8134 5362 8186
rect 5414 8134 5426 8186
rect 5478 8134 6895 8186
rect 6947 8134 6959 8186
rect 7011 8134 7023 8186
rect 7075 8134 7087 8186
rect 7139 8134 7151 8186
rect 7203 8134 7912 8186
rect 1012 8112 7912 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 2038 8072 2044 8084
rect 1811 8044 2044 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 5626 8072 5632 8084
rect 5224 8044 5632 8072
rect 5224 8032 5230 8044
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 3142 7896 3148 7948
rect 3200 7936 3206 7948
rect 3200 7908 4752 7936
rect 3200 7896 3206 7908
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 2096 7840 2237 7868
rect 2096 7828 2102 7840
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 2464 7840 3893 7868
rect 2464 7828 2470 7840
rect 3881 7837 3893 7840
rect 3927 7868 3939 7871
rect 4062 7868 4068 7880
rect 3927 7840 4068 7868
rect 3927 7837 3939 7840
rect 3881 7831 3939 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 4724 7868 4752 7908
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5626 7936 5632 7948
rect 4856 7908 5632 7936
rect 4856 7896 4862 7908
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5350 7868 5356 7880
rect 4724 7840 5356 7868
rect 5350 7828 5356 7840
rect 5408 7868 5414 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 5408 7840 5733 7868
rect 5408 7828 5414 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 3053 7803 3111 7809
rect 3053 7769 3065 7803
rect 3099 7769 3111 7803
rect 3053 7763 3111 7769
rect 4709 7803 4767 7809
rect 4709 7769 4721 7803
rect 4755 7800 4767 7803
rect 4798 7800 4804 7812
rect 4755 7772 4804 7800
rect 4755 7769 4767 7772
rect 4709 7763 4767 7769
rect 3068 7732 3096 7763
rect 4798 7760 4804 7772
rect 4856 7760 4862 7812
rect 6546 7800 6552 7812
rect 6507 7772 6552 7800
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 5534 7732 5540 7744
rect 3068 7704 5540 7732
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 7098 7732 7104 7744
rect 7059 7704 7104 7732
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 1012 7642 8071 7664
rect 1012 7590 2582 7642
rect 2634 7590 2646 7642
rect 2698 7590 2710 7642
rect 2762 7590 2774 7642
rect 2826 7590 2838 7642
rect 2890 7590 4307 7642
rect 4359 7590 4371 7642
rect 4423 7590 4435 7642
rect 4487 7590 4499 7642
rect 4551 7590 4563 7642
rect 4615 7590 6032 7642
rect 6084 7590 6096 7642
rect 6148 7590 6160 7642
rect 6212 7590 6224 7642
rect 6276 7590 6288 7642
rect 6340 7590 7757 7642
rect 7809 7590 7821 7642
rect 7873 7590 7885 7642
rect 7937 7590 7949 7642
rect 8001 7590 8013 7642
rect 8065 7590 8071 7642
rect 1012 7568 8071 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 4062 7528 4068 7540
rect 4023 7500 4068 7528
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 5074 7528 5080 7540
rect 4672 7500 5080 7528
rect 4672 7488 4678 7500
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 5408 7500 5549 7528
rect 5408 7488 5414 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 5537 7491 5595 7497
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7742 7528 7748 7540
rect 7616 7500 7748 7528
rect 7616 7488 7622 7500
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 3513 7463 3571 7469
rect 3513 7429 3525 7463
rect 3559 7460 3571 7463
rect 4706 7460 4712 7472
rect 3559 7432 4712 7460
rect 3559 7429 3571 7432
rect 3513 7423 3571 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 7374 7420 7380 7472
rect 7432 7460 7438 7472
rect 7432 7432 7604 7460
rect 7432 7420 7438 7432
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 2148 7364 2697 7392
rect 1486 7216 1492 7268
rect 1544 7256 1550 7268
rect 2148 7265 2176 7364
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 6457 7395 6515 7401
rect 6457 7392 6469 7395
rect 4028 7364 6469 7392
rect 4028 7352 4034 7364
rect 6457 7361 6469 7364
rect 6503 7392 6515 7395
rect 7098 7392 7104 7404
rect 6503 7364 7104 7392
rect 6503 7361 6515 7364
rect 6457 7355 6515 7361
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7576 7336 7604 7432
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 4120 7296 4629 7324
rect 4120 7284 4126 7296
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 7374 7324 7380 7336
rect 7331 7296 7380 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7558 7284 7564 7336
rect 7616 7284 7622 7336
rect 2133 7259 2191 7265
rect 2133 7256 2145 7259
rect 1544 7228 2145 7256
rect 1544 7216 1550 7228
rect 2133 7225 2145 7228
rect 2179 7225 2191 7259
rect 2133 7219 2191 7225
rect 1012 7098 7912 7120
rect 1012 7046 1720 7098
rect 1772 7046 1784 7098
rect 1836 7046 1848 7098
rect 1900 7046 1912 7098
rect 1964 7046 1976 7098
rect 2028 7046 3445 7098
rect 3497 7046 3509 7098
rect 3561 7046 3573 7098
rect 3625 7046 3637 7098
rect 3689 7046 3701 7098
rect 3753 7046 5170 7098
rect 5222 7046 5234 7098
rect 5286 7046 5298 7098
rect 5350 7046 5362 7098
rect 5414 7046 5426 7098
rect 5478 7046 6895 7098
rect 6947 7046 6959 7098
rect 7011 7046 7023 7098
rect 7075 7046 7087 7098
rect 7139 7046 7151 7098
rect 7203 7046 7912 7098
rect 1012 7024 7912 7046
rect 3326 6876 3332 6928
rect 3384 6916 3390 6928
rect 3384 6888 6592 6916
rect 3384 6876 3390 6888
rect 4893 6851 4951 6857
rect 4893 6817 4905 6851
rect 4939 6848 4951 6851
rect 5074 6848 5080 6860
rect 4939 6820 5080 6848
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 6564 6857 6592 6888
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 1857 6783 1915 6789
rect 1857 6780 1869 6783
rect 1360 6752 1869 6780
rect 1360 6740 1366 6752
rect 1857 6749 1869 6752
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 4522 6780 4528 6792
rect 2731 6752 4528 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4065 6715 4123 6721
rect 4065 6681 4077 6715
rect 4111 6681 4123 6715
rect 4065 6675 4123 6681
rect 5997 6715 6055 6721
rect 5997 6681 6009 6715
rect 6043 6712 6055 6715
rect 7377 6715 7435 6721
rect 7377 6712 7389 6715
rect 6043 6684 7389 6712
rect 6043 6681 6055 6684
rect 5997 6675 6055 6681
rect 7377 6681 7389 6684
rect 7423 6712 7435 6715
rect 8202 6712 8208 6724
rect 7423 6684 8208 6712
rect 7423 6681 7435 6684
rect 7377 6675 7435 6681
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 3108 6616 3249 6644
rect 3108 6604 3114 6616
rect 3237 6613 3249 6616
rect 3283 6644 3295 6647
rect 4080 6644 4108 6675
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 3283 6616 4108 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 5902 6644 5908 6656
rect 5132 6616 5908 6644
rect 5132 6604 5138 6616
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6362 6604 6368 6656
rect 6420 6644 6426 6656
rect 7742 6644 7748 6656
rect 6420 6616 7748 6644
rect 6420 6604 6426 6616
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 1012 6554 8071 6576
rect 1012 6502 2582 6554
rect 2634 6502 2646 6554
rect 2698 6502 2710 6554
rect 2762 6502 2774 6554
rect 2826 6502 2838 6554
rect 2890 6502 4307 6554
rect 4359 6502 4371 6554
rect 4423 6502 4435 6554
rect 4487 6502 4499 6554
rect 4551 6502 4563 6554
rect 4615 6502 6032 6554
rect 6084 6502 6096 6554
rect 6148 6502 6160 6554
rect 6212 6502 6224 6554
rect 6276 6502 6288 6554
rect 6340 6502 7757 6554
rect 7809 6502 7821 6554
rect 7873 6502 7885 6554
rect 7937 6502 7949 6554
rect 8001 6502 8013 6554
rect 8065 6502 8071 6554
rect 1012 6480 8071 6502
rect 1302 6400 1308 6452
rect 1360 6440 1366 6452
rect 1673 6443 1731 6449
rect 1673 6440 1685 6443
rect 1360 6412 1685 6440
rect 1360 6400 1366 6412
rect 1673 6409 1685 6412
rect 1719 6409 1731 6443
rect 1673 6403 1731 6409
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6730 6440 6736 6452
rect 5960 6412 6736 6440
rect 5960 6400 5966 6412
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 3605 6375 3663 6381
rect 3605 6341 3617 6375
rect 3651 6372 3663 6375
rect 3878 6372 3884 6384
rect 3651 6344 3884 6372
rect 3651 6341 3663 6344
rect 3605 6335 3663 6341
rect 3878 6332 3884 6344
rect 3936 6332 3942 6384
rect 4249 6375 4307 6381
rect 4249 6341 4261 6375
rect 4295 6372 4307 6375
rect 6362 6372 6368 6384
rect 4295 6344 6368 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 7285 6375 7343 6381
rect 7285 6341 7297 6375
rect 7331 6372 7343 6375
rect 7558 6372 7564 6384
rect 7331 6344 7564 6372
rect 7331 6341 7343 6344
rect 7285 6335 7343 6341
rect 7558 6332 7564 6344
rect 7616 6332 7622 6384
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6457 6307 6515 6313
rect 6457 6304 6469 6307
rect 5951 6276 6469 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6457 6273 6469 6276
rect 6503 6304 6515 6307
rect 6730 6304 6736 6316
rect 6503 6276 6736 6304
rect 6503 6273 6515 6276
rect 6457 6267 6515 6273
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2792 6100 2820 6267
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 5534 6236 5540 6248
rect 3016 6208 5540 6236
rect 3016 6196 3022 6208
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 5353 6171 5411 6177
rect 5353 6137 5365 6171
rect 5399 6168 5411 6171
rect 7558 6168 7564 6180
rect 5399 6140 7564 6168
rect 5399 6137 5411 6140
rect 5353 6131 5411 6137
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 2958 6100 2964 6112
rect 2363 6072 2964 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 5902 6100 5908 6112
rect 4847 6072 5908 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 1012 6010 7912 6032
rect 1012 5958 1720 6010
rect 1772 5958 1784 6010
rect 1836 5958 1848 6010
rect 1900 5958 1912 6010
rect 1964 5958 1976 6010
rect 2028 5958 3445 6010
rect 3497 5958 3509 6010
rect 3561 5958 3573 6010
rect 3625 5958 3637 6010
rect 3689 5958 3701 6010
rect 3753 5958 5170 6010
rect 5222 5958 5234 6010
rect 5286 5958 5298 6010
rect 5350 5958 5362 6010
rect 5414 5958 5426 6010
rect 5478 5958 6895 6010
rect 6947 5958 6959 6010
rect 7011 5958 7023 6010
rect 7075 5958 7087 6010
rect 7139 5958 7151 6010
rect 7203 5958 7912 6010
rect 1012 5936 7912 5958
rect 1026 5856 1032 5908
rect 1084 5896 1090 5908
rect 5166 5896 5172 5908
rect 1084 5868 5172 5896
rect 1084 5856 1090 5868
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 5905 5899 5963 5905
rect 5905 5896 5917 5899
rect 5684 5868 5917 5896
rect 5684 5856 5690 5868
rect 5905 5865 5917 5868
rect 5951 5865 5963 5899
rect 5905 5859 5963 5865
rect 2498 5720 2504 5772
rect 2556 5760 2562 5772
rect 3973 5763 4031 5769
rect 3973 5760 3985 5763
rect 2556 5732 3985 5760
rect 2556 5720 2562 5732
rect 3973 5729 3985 5732
rect 4019 5729 4031 5763
rect 3973 5723 4031 5729
rect 2130 5652 2136 5704
rect 2188 5692 2194 5704
rect 5442 5692 5448 5704
rect 2188 5664 5448 5692
rect 2188 5652 2194 5664
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5920 5692 5948 5859
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 7558 5896 7564 5908
rect 7248 5868 7564 5896
rect 7248 5856 7254 5868
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7558 5760 7564 5772
rect 7340 5732 7564 5760
rect 7340 5720 7346 5732
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 6457 5695 6515 5701
rect 6457 5692 6469 5695
rect 5920 5664 6469 5692
rect 6457 5661 6469 5664
rect 6503 5661 6515 5695
rect 6457 5655 6515 5661
rect 1394 5584 1400 5636
rect 1452 5624 1458 5636
rect 3326 5624 3332 5636
rect 1452 5596 3332 5624
rect 1452 5584 1458 5596
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 4798 5624 4804 5636
rect 4759 5596 4804 5624
rect 4798 5584 4804 5596
rect 4856 5624 4862 5636
rect 5261 5627 5319 5633
rect 5261 5624 5273 5627
rect 4856 5596 5273 5624
rect 4856 5584 4862 5596
rect 5261 5593 5273 5596
rect 5307 5593 5319 5627
rect 5261 5587 5319 5593
rect 5626 5584 5632 5636
rect 5684 5624 5690 5636
rect 5902 5624 5908 5636
rect 5684 5596 5908 5624
rect 5684 5584 5690 5596
rect 5902 5584 5908 5596
rect 5960 5584 5966 5636
rect 7282 5624 7288 5636
rect 7243 5596 7288 5624
rect 7282 5584 7288 5596
rect 7340 5584 7346 5636
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2222 5556 2228 5568
rect 2183 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 3142 5556 3148 5568
rect 2823 5528 3148 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3878 5556 3884 5568
rect 3283 5528 3884 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 1012 5466 8071 5488
rect 1012 5414 2582 5466
rect 2634 5414 2646 5466
rect 2698 5414 2710 5466
rect 2762 5414 2774 5466
rect 2826 5414 2838 5466
rect 2890 5414 4307 5466
rect 4359 5414 4371 5466
rect 4423 5414 4435 5466
rect 4487 5414 4499 5466
rect 4551 5414 4563 5466
rect 4615 5414 6032 5466
rect 6084 5414 6096 5466
rect 6148 5414 6160 5466
rect 6212 5414 6224 5466
rect 6276 5414 6288 5466
rect 6340 5414 7757 5466
rect 7809 5414 7821 5466
rect 7873 5414 7885 5466
rect 7937 5414 7949 5466
rect 8001 5414 8013 5466
rect 8065 5414 8071 5466
rect 1012 5392 8071 5414
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6454 5352 6460 5364
rect 6328 5324 6460 5352
rect 6328 5312 6334 5324
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 4433 5287 4491 5293
rect 4433 5253 4445 5287
rect 4479 5284 4491 5287
rect 4890 5284 4896 5296
rect 4479 5256 4896 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 5166 5284 5172 5296
rect 5127 5256 5172 5284
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 5592 5256 6561 5284
rect 5592 5244 5598 5256
rect 6549 5253 6561 5256
rect 6595 5253 6607 5287
rect 6549 5247 6607 5253
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 3108 5188 3617 5216
rect 3108 5176 3114 5188
rect 3605 5185 3617 5188
rect 3651 5185 3663 5219
rect 5902 5216 5908 5228
rect 5863 5188 5908 5216
rect 3605 5179 3663 5185
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 7190 5176 7196 5228
rect 7248 5216 7254 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 7248 5188 7389 5216
rect 7248 5176 7254 5188
rect 7377 5185 7389 5188
rect 7423 5216 7435 5219
rect 7423 5188 7512 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 2041 5083 2099 5089
rect 2041 5049 2053 5083
rect 2087 5080 2099 5083
rect 4890 5080 4896 5092
rect 2087 5052 4896 5080
rect 2087 5049 2099 5052
rect 2041 5043 2099 5049
rect 4890 5040 4896 5052
rect 4948 5040 4954 5092
rect 7484 5024 7512 5188
rect 2593 5015 2651 5021
rect 2593 4981 2605 5015
rect 2639 5012 2651 5015
rect 2774 5012 2780 5024
rect 2639 4984 2780 5012
rect 2639 4981 2651 4984
rect 2593 4975 2651 4981
rect 2774 4972 2780 4984
rect 2832 4972 2838 5024
rect 3050 5012 3056 5024
rect 3011 4984 3056 5012
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 7466 4972 7472 5024
rect 7524 4972 7530 5024
rect 1012 4922 7912 4944
rect 1012 4870 1720 4922
rect 1772 4870 1784 4922
rect 1836 4870 1848 4922
rect 1900 4870 1912 4922
rect 1964 4870 1976 4922
rect 2028 4870 3445 4922
rect 3497 4870 3509 4922
rect 3561 4870 3573 4922
rect 3625 4870 3637 4922
rect 3689 4870 3701 4922
rect 3753 4870 5170 4922
rect 5222 4870 5234 4922
rect 5286 4870 5298 4922
rect 5350 4870 5362 4922
rect 5414 4870 5426 4922
rect 5478 4870 6895 4922
rect 6947 4870 6959 4922
rect 7011 4870 7023 4922
rect 7075 4870 7087 4922
rect 7139 4870 7151 4922
rect 7203 4870 7912 4922
rect 1012 4848 7912 4870
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3878 4808 3884 4820
rect 3752 4780 3884 4808
rect 3752 4768 3758 4780
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4706 4768 4712 4820
rect 4764 4808 4770 4820
rect 5353 4811 5411 4817
rect 5353 4808 5365 4811
rect 4764 4780 5365 4808
rect 4764 4768 4770 4780
rect 5353 4777 5365 4780
rect 5399 4777 5411 4811
rect 5353 4771 5411 4777
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3786 4672 3792 4684
rect 3283 4644 3792 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2774 4604 2780 4616
rect 2455 4576 2780 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2774 4564 2780 4576
rect 2832 4604 2838 4616
rect 3970 4604 3976 4616
rect 2832 4576 3976 4604
rect 2832 4564 2838 4576
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 5368 4604 5396 4771
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 5368 4576 6469 4604
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 3881 4539 3939 4545
rect 3881 4505 3893 4539
rect 3927 4505 3939 4539
rect 3881 4499 3939 4505
rect 4709 4539 4767 4545
rect 4709 4505 4721 4539
rect 4755 4536 4767 4539
rect 6638 4536 6644 4548
rect 4755 4508 6644 4536
rect 4755 4505 4767 4508
rect 4709 4499 4767 4505
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1636 4440 1869 4468
rect 1636 4428 1642 4440
rect 1857 4437 1869 4440
rect 1903 4468 1915 4471
rect 3896 4468 3924 4499
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 6822 4496 6828 4548
rect 6880 4536 6886 4548
rect 7193 4539 7251 4545
rect 7193 4536 7205 4539
rect 6880 4508 7205 4536
rect 6880 4496 6886 4508
rect 7193 4505 7205 4508
rect 7239 4505 7251 4539
rect 7193 4499 7251 4505
rect 1903 4440 3924 4468
rect 1903 4437 1915 4440
rect 1857 4431 1915 4437
rect 5902 4428 5908 4480
rect 5960 4468 5966 4480
rect 5997 4471 6055 4477
rect 5997 4468 6009 4471
rect 5960 4440 6009 4468
rect 5960 4428 5966 4440
rect 5997 4437 6009 4440
rect 6043 4468 6055 4471
rect 6362 4468 6368 4480
rect 6043 4440 6368 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 1012 4378 8071 4400
rect 1012 4326 2582 4378
rect 2634 4326 2646 4378
rect 2698 4326 2710 4378
rect 2762 4326 2774 4378
rect 2826 4326 2838 4378
rect 2890 4326 4307 4378
rect 4359 4326 4371 4378
rect 4423 4326 4435 4378
rect 4487 4326 4499 4378
rect 4551 4326 4563 4378
rect 4615 4326 6032 4378
rect 6084 4326 6096 4378
rect 6148 4326 6160 4378
rect 6212 4326 6224 4378
rect 6276 4326 6288 4378
rect 6340 4326 7757 4378
rect 7809 4326 7821 4378
rect 7873 4326 7885 4378
rect 7937 4326 7949 4378
rect 8001 4326 8013 4378
rect 8065 4326 8071 4378
rect 1012 4304 8071 4326
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 4246 4264 4252 4276
rect 4120 4236 4252 4264
rect 4120 4224 4126 4236
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 4890 4224 4896 4276
rect 4948 4264 4954 4276
rect 6638 4264 6644 4276
rect 4948 4236 6644 4264
rect 4948 4224 4954 4236
rect 6638 4224 6644 4236
rect 6696 4264 6702 4276
rect 8110 4264 8116 4276
rect 6696 4236 8116 4264
rect 6696 4224 6702 4236
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4196 4491 4199
rect 4706 4196 4712 4208
rect 4479 4168 4712 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3605 4131 3663 4137
rect 3605 4128 3617 4131
rect 3292 4100 3617 4128
rect 3292 4088 3298 4100
rect 3605 4097 3617 4100
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4060 3111 4063
rect 4448 4060 4476 4159
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 5718 4156 5724 4208
rect 5776 4196 5782 4208
rect 6457 4199 6515 4205
rect 6457 4196 6469 4199
rect 5776 4168 6469 4196
rect 5776 4156 5782 4168
rect 6457 4165 6469 4168
rect 6503 4165 6515 4199
rect 6457 4159 6515 4165
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5442 4128 5448 4140
rect 5123 4100 5448 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5810 4128 5816 4140
rect 5771 4100 5816 4128
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 7282 4060 7288 4072
rect 3099 4032 4476 4060
rect 7243 4032 7288 4060
rect 3099 4029 3111 4032
rect 3053 4023 3111 4029
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 3694 3992 3700 4004
rect 3292 3964 3700 3992
rect 3292 3952 3298 3964
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2038 3924 2044 3936
rect 1995 3896 2044 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 3786 3924 3792 3936
rect 2547 3896 3792 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 1012 3834 7912 3856
rect 1012 3782 1720 3834
rect 1772 3782 1784 3834
rect 1836 3782 1848 3834
rect 1900 3782 1912 3834
rect 1964 3782 1976 3834
rect 2028 3782 3445 3834
rect 3497 3782 3509 3834
rect 3561 3782 3573 3834
rect 3625 3782 3637 3834
rect 3689 3782 3701 3834
rect 3753 3782 5170 3834
rect 5222 3782 5234 3834
rect 5286 3782 5298 3834
rect 5350 3782 5362 3834
rect 5414 3782 5426 3834
rect 5478 3782 6895 3834
rect 6947 3782 6959 3834
rect 7011 3782 7023 3834
rect 7075 3782 7087 3834
rect 7139 3782 7151 3834
rect 7203 3782 7912 3834
rect 1012 3760 7912 3782
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 4246 3720 4252 3732
rect 3752 3692 4252 3720
rect 3752 3680 3758 3692
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 5445 3723 5503 3729
rect 5445 3689 5457 3723
rect 5491 3720 5503 3723
rect 5718 3720 5724 3732
rect 5491 3692 5724 3720
rect 5491 3689 5503 3692
rect 5445 3683 5503 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 4709 3587 4767 3593
rect 4709 3553 4721 3587
rect 4755 3584 4767 3587
rect 4982 3584 4988 3596
rect 4755 3556 4988 3584
rect 4755 3553 4767 3556
rect 4709 3547 4767 3553
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 7650 3584 7656 3596
rect 7331 3556 7656 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 2096 3488 3341 3516
rect 2096 3476 2102 3488
rect 3329 3485 3341 3488
rect 3375 3516 3387 3519
rect 5442 3516 5448 3528
rect 3375 3488 5448 3516
rect 3375 3485 3387 3488
rect 3329 3479 3387 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 5776 3488 6469 3516
rect 5776 3476 5782 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 2593 3451 2651 3457
rect 2593 3417 2605 3451
rect 2639 3448 2651 3451
rect 2958 3448 2964 3460
rect 2639 3420 2964 3448
rect 2639 3417 2651 3420
rect 2593 3411 2651 3417
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 3881 3451 3939 3457
rect 3881 3417 3893 3451
rect 3927 3417 3939 3451
rect 3881 3411 3939 3417
rect 1949 3383 2007 3389
rect 1949 3349 1961 3383
rect 1995 3380 2007 3383
rect 2498 3380 2504 3392
rect 1995 3352 2504 3380
rect 1995 3349 2007 3352
rect 1949 3343 2007 3349
rect 2498 3340 2504 3352
rect 2556 3380 2562 3392
rect 3896 3380 3924 3411
rect 2556 3352 3924 3380
rect 2556 3340 2562 3352
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 5810 3380 5816 3392
rect 5132 3352 5816 3380
rect 5132 3340 5138 3352
rect 5810 3340 5816 3352
rect 5868 3380 5874 3392
rect 5997 3383 6055 3389
rect 5997 3380 6009 3383
rect 5868 3352 6009 3380
rect 5868 3340 5874 3352
rect 5997 3349 6009 3352
rect 6043 3349 6055 3383
rect 5997 3343 6055 3349
rect 1012 3290 8071 3312
rect 1012 3238 2582 3290
rect 2634 3238 2646 3290
rect 2698 3238 2710 3290
rect 2762 3238 2774 3290
rect 2826 3238 2838 3290
rect 2890 3238 4307 3290
rect 4359 3238 4371 3290
rect 4423 3238 4435 3290
rect 4487 3238 4499 3290
rect 4551 3238 4563 3290
rect 4615 3238 6032 3290
rect 6084 3238 6096 3290
rect 6148 3238 6160 3290
rect 6212 3238 6224 3290
rect 6276 3238 6288 3290
rect 6340 3238 7757 3290
rect 7809 3238 7821 3290
rect 7873 3238 7885 3290
rect 7937 3238 7949 3290
rect 8001 3238 8013 3290
rect 8065 3238 8071 3290
rect 1012 3216 8071 3238
rect 8386 3176 8392 3188
rect 2332 3148 8392 3176
rect 2332 3117 2360 3148
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 2317 3111 2375 3117
rect 2317 3077 2329 3111
rect 2363 3077 2375 3111
rect 3326 3108 3332 3120
rect 3287 3080 3332 3108
rect 2317 3071 2375 3077
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 3786 3068 3792 3120
rect 3844 3108 3850 3120
rect 4157 3111 4215 3117
rect 4157 3108 4169 3111
rect 3844 3080 4169 3108
rect 3844 3068 3850 3080
rect 4157 3077 4169 3080
rect 4203 3108 4215 3111
rect 5810 3108 5816 3120
rect 4203 3080 5816 3108
rect 4203 3077 4215 3080
rect 4157 3071 4215 3077
rect 5810 3068 5816 3080
rect 5868 3068 5874 3120
rect 6454 3108 6460 3120
rect 6415 3080 6460 3108
rect 6454 3068 6460 3080
rect 6512 3068 6518 3120
rect 290 3000 296 3052
rect 348 3040 354 3052
rect 1486 3040 1492 3052
rect 348 3012 1492 3040
rect 348 3000 354 3012
rect 1486 3000 1492 3012
rect 1544 3000 1550 3052
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3040 4675 3043
rect 4798 3040 4804 3052
rect 4663 3012 4804 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 7558 2972 7564 2984
rect 5491 2944 7564 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 3234 2864 3240 2916
rect 3292 2904 3298 2916
rect 8570 2904 8576 2916
rect 3292 2876 8576 2904
rect 3292 2864 3298 2876
rect 8570 2864 8576 2876
rect 8628 2864 8634 2916
rect 750 2796 756 2848
rect 808 2836 814 2848
rect 5718 2836 5724 2848
rect 808 2808 5724 2836
rect 808 2796 814 2808
rect 5718 2796 5724 2808
rect 5776 2836 5782 2848
rect 5994 2836 6000 2848
rect 5776 2808 6000 2836
rect 5776 2796 5782 2808
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 1012 2746 7912 2768
rect 1012 2694 1720 2746
rect 1772 2694 1784 2746
rect 1836 2694 1848 2746
rect 1900 2694 1912 2746
rect 1964 2694 1976 2746
rect 2028 2694 3445 2746
rect 3497 2694 3509 2746
rect 3561 2694 3573 2746
rect 3625 2694 3637 2746
rect 3689 2694 3701 2746
rect 3753 2694 5170 2746
rect 5222 2694 5234 2746
rect 5286 2694 5298 2746
rect 5350 2694 5362 2746
rect 5414 2694 5426 2746
rect 5478 2694 6895 2746
rect 6947 2694 6959 2746
rect 7011 2694 7023 2746
rect 7075 2694 7087 2746
rect 7139 2694 7151 2746
rect 7203 2694 7912 2746
rect 1012 2672 7912 2694
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 5166 2632 5172 2644
rect 3936 2604 5172 2632
rect 3936 2592 3942 2604
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 6454 2632 6460 2644
rect 5491 2604 6460 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 5994 2564 6000 2576
rect 5955 2536 6000 2564
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 2593 2499 2651 2505
rect 2593 2465 2605 2499
rect 2639 2496 2651 2499
rect 2774 2496 2780 2508
rect 2639 2468 2780 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 4709 2499 4767 2505
rect 4709 2465 4721 2499
rect 4755 2496 4767 2499
rect 5902 2496 5908 2508
rect 4755 2468 5908 2496
rect 4755 2465 4767 2468
rect 4709 2459 4767 2465
rect 5902 2456 5908 2468
rect 5960 2456 5966 2508
rect 7282 2496 7288 2508
rect 7243 2468 7288 2496
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3292 2400 3341 2428
rect 3292 2388 3298 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 6457 2431 6515 2437
rect 6457 2428 6469 2431
rect 5684 2400 6469 2428
rect 5684 2388 5690 2400
rect 6457 2397 6469 2400
rect 6503 2397 6515 2431
rect 6457 2391 6515 2397
rect 3881 2363 3939 2369
rect 3881 2329 3893 2363
rect 3927 2329 3939 2363
rect 3881 2323 3939 2329
rect 1949 2295 2007 2301
rect 1949 2261 1961 2295
rect 1995 2292 2007 2295
rect 2130 2292 2136 2304
rect 1995 2264 2136 2292
rect 1995 2261 2007 2264
rect 1949 2255 2007 2261
rect 2130 2252 2136 2264
rect 2188 2292 2194 2304
rect 3896 2292 3924 2323
rect 2188 2264 3924 2292
rect 2188 2252 2194 2264
rect 1012 2202 8071 2224
rect 1012 2150 2582 2202
rect 2634 2150 2646 2202
rect 2698 2150 2710 2202
rect 2762 2150 2774 2202
rect 2826 2150 2838 2202
rect 2890 2150 4307 2202
rect 4359 2150 4371 2202
rect 4423 2150 4435 2202
rect 4487 2150 4499 2202
rect 4551 2150 4563 2202
rect 4615 2150 6032 2202
rect 6084 2150 6096 2202
rect 6148 2150 6160 2202
rect 6212 2150 6224 2202
rect 6276 2150 6288 2202
rect 6340 2150 7757 2202
rect 7809 2150 7821 2202
rect 7873 2150 7885 2202
rect 7937 2150 7949 2202
rect 8001 2150 8013 2202
rect 8065 2150 8071 2202
rect 1012 2128 8071 2150
rect 1765 2091 1823 2097
rect 1765 2057 1777 2091
rect 1811 2088 1823 2091
rect 8110 2088 8116 2100
rect 1811 2060 8116 2088
rect 1811 2057 1823 2060
rect 1765 2051 1823 2057
rect 3142 1980 3148 2032
rect 3200 2020 3206 2032
rect 3605 2023 3663 2029
rect 3605 2020 3617 2023
rect 3200 1992 3617 2020
rect 3200 1980 3206 1992
rect 3605 1989 3617 1992
rect 3651 1989 3663 2023
rect 3605 1983 3663 1989
rect 4154 1980 4160 2032
rect 4212 2020 4218 2032
rect 4341 2023 4399 2029
rect 4341 2020 4353 2023
rect 4212 1992 4353 2020
rect 4212 1980 4218 1992
rect 4341 1989 4353 1992
rect 4387 1989 4399 2023
rect 5166 2020 5172 2032
rect 5127 1992 5172 2020
rect 4341 1983 4399 1989
rect 5166 1980 5172 1992
rect 5224 1980 5230 2032
rect 5920 2029 5948 2060
rect 8110 2048 8116 2060
rect 8168 2048 8174 2100
rect 5905 2023 5963 2029
rect 5905 1989 5917 2023
rect 5951 1989 5963 2023
rect 5905 1983 5963 1989
rect 6457 2023 6515 2029
rect 6457 1989 6469 2023
rect 6503 2020 6515 2023
rect 6546 2020 6552 2032
rect 6503 1992 6552 2020
rect 6503 1989 6515 1992
rect 6457 1983 6515 1989
rect 6546 1980 6552 1992
rect 6604 1980 6610 2032
rect 7282 2020 7288 2032
rect 7243 1992 7288 2020
rect 7282 1980 7288 1992
rect 7340 1980 7346 2032
rect 2225 1955 2283 1961
rect 2225 1921 2237 1955
rect 2271 1921 2283 1955
rect 2225 1915 2283 1921
rect 3053 1955 3111 1961
rect 3053 1921 3065 1955
rect 3099 1952 3111 1955
rect 4982 1952 4988 1964
rect 3099 1924 4988 1952
rect 3099 1921 3111 1924
rect 3053 1915 3111 1921
rect 1486 1844 1492 1896
rect 1544 1884 1550 1896
rect 2240 1884 2268 1915
rect 4982 1912 4988 1924
rect 5040 1912 5046 1964
rect 3786 1884 3792 1896
rect 1544 1856 3792 1884
rect 1544 1844 1550 1856
rect 3786 1844 3792 1856
rect 3844 1844 3850 1896
rect 1012 1658 7912 1680
rect 1012 1606 1720 1658
rect 1772 1606 1784 1658
rect 1836 1606 1848 1658
rect 1900 1606 1912 1658
rect 1964 1606 1976 1658
rect 2028 1606 3445 1658
rect 3497 1606 3509 1658
rect 3561 1606 3573 1658
rect 3625 1606 3637 1658
rect 3689 1606 3701 1658
rect 3753 1606 5170 1658
rect 5222 1606 5234 1658
rect 5286 1606 5298 1658
rect 5350 1606 5362 1658
rect 5414 1606 5426 1658
rect 5478 1606 6895 1658
rect 6947 1606 6959 1658
rect 7011 1606 7023 1658
rect 7075 1606 7087 1658
rect 7139 1606 7151 1658
rect 7203 1606 7912 1658
rect 1012 1584 7912 1606
rect 7190 1504 7196 1556
rect 7248 1544 7254 1556
rect 8202 1544 8208 1556
rect 7248 1516 8208 1544
rect 7248 1504 7254 1516
rect 8202 1504 8208 1516
rect 8260 1504 8266 1556
rect 2593 1411 2651 1417
rect 2593 1377 2605 1411
rect 2639 1408 2651 1411
rect 2774 1408 2780 1420
rect 2639 1380 2780 1408
rect 2639 1377 2651 1380
rect 2593 1371 2651 1377
rect 2774 1368 2780 1380
rect 2832 1368 2838 1420
rect 4154 1408 4160 1420
rect 4115 1380 4160 1408
rect 4154 1368 4160 1380
rect 4212 1368 4218 1420
rect 1949 1343 2007 1349
rect 1949 1309 1961 1343
rect 1995 1340 2007 1343
rect 4893 1343 4951 1349
rect 4893 1340 4905 1343
rect 1995 1312 4905 1340
rect 1995 1309 2007 1312
rect 1949 1303 2007 1309
rect 4893 1309 4905 1312
rect 4939 1340 4951 1343
rect 6822 1340 6828 1352
rect 4939 1312 6828 1340
rect 4939 1309 4951 1312
rect 4893 1303 4951 1309
rect 6822 1300 6828 1312
rect 6880 1300 6886 1352
rect 7282 1340 7288 1352
rect 7243 1312 7288 1340
rect 7282 1300 7288 1312
rect 7340 1300 7346 1352
rect 2222 1232 2228 1284
rect 2280 1272 2286 1284
rect 3329 1275 3387 1281
rect 3329 1272 3341 1275
rect 2280 1244 3341 1272
rect 2280 1232 2286 1244
rect 3329 1241 3341 1244
rect 3375 1272 3387 1275
rect 4982 1272 4988 1284
rect 3375 1244 4988 1272
rect 3375 1241 3387 1244
rect 3329 1235 3387 1241
rect 4982 1232 4988 1244
rect 5040 1232 5046 1284
rect 6457 1275 6515 1281
rect 6457 1241 6469 1275
rect 6503 1272 6515 1275
rect 6638 1272 6644 1284
rect 6503 1244 6644 1272
rect 6503 1241 6515 1244
rect 6457 1235 6515 1241
rect 6638 1232 6644 1244
rect 6696 1232 6702 1284
rect 1210 1164 1216 1216
rect 1268 1204 1274 1216
rect 4798 1204 4804 1216
rect 1268 1176 4804 1204
rect 1268 1164 1274 1176
rect 4798 1164 4804 1176
rect 4856 1204 4862 1216
rect 5353 1207 5411 1213
rect 5353 1204 5365 1207
rect 4856 1176 5365 1204
rect 4856 1164 4862 1176
rect 5353 1173 5365 1176
rect 5399 1173 5411 1207
rect 5353 1167 5411 1173
rect 1012 1114 8071 1136
rect 1012 1062 2582 1114
rect 2634 1062 2646 1114
rect 2698 1062 2710 1114
rect 2762 1062 2774 1114
rect 2826 1062 2838 1114
rect 2890 1062 4307 1114
rect 4359 1062 4371 1114
rect 4423 1062 4435 1114
rect 4487 1062 4499 1114
rect 4551 1062 4563 1114
rect 4615 1062 6032 1114
rect 6084 1062 6096 1114
rect 6148 1062 6160 1114
rect 6212 1062 6224 1114
rect 6276 1062 6288 1114
rect 6340 1062 7757 1114
rect 7809 1062 7821 1114
rect 7873 1062 7885 1114
rect 7937 1062 7949 1114
rect 8001 1062 8013 1114
rect 8065 1062 8071 1114
rect 1012 1040 8071 1062
<< via1 >>
rect 3424 8848 3476 8900
rect 7380 8848 7432 8900
rect 2582 8678 2634 8730
rect 2646 8678 2698 8730
rect 2710 8678 2762 8730
rect 2774 8678 2826 8730
rect 2838 8678 2890 8730
rect 4307 8678 4359 8730
rect 4371 8678 4423 8730
rect 4435 8678 4487 8730
rect 4499 8678 4551 8730
rect 4563 8678 4615 8730
rect 6032 8678 6084 8730
rect 6096 8678 6148 8730
rect 6160 8678 6212 8730
rect 6224 8678 6276 8730
rect 6288 8678 6340 8730
rect 7757 8678 7809 8730
rect 7821 8678 7873 8730
rect 7885 8678 7937 8730
rect 7949 8678 8001 8730
rect 8013 8678 8065 8730
rect 940 8576 992 8628
rect 3700 8576 3752 8628
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 4620 8372 4672 8424
rect 5448 8372 5500 8424
rect 7472 8372 7524 8424
rect 4988 8236 5040 8288
rect 5264 8236 5316 8288
rect 1720 8134 1772 8186
rect 1784 8134 1836 8186
rect 1848 8134 1900 8186
rect 1912 8134 1964 8186
rect 1976 8134 2028 8186
rect 3445 8134 3497 8186
rect 3509 8134 3561 8186
rect 3573 8134 3625 8186
rect 3637 8134 3689 8186
rect 3701 8134 3753 8186
rect 5170 8134 5222 8186
rect 5234 8134 5286 8186
rect 5298 8134 5350 8186
rect 5362 8134 5414 8186
rect 5426 8134 5478 8186
rect 6895 8134 6947 8186
rect 6959 8134 7011 8186
rect 7023 8134 7075 8186
rect 7087 8134 7139 8186
rect 7151 8134 7203 8186
rect 2044 8032 2096 8084
rect 5172 8032 5224 8084
rect 5632 8032 5684 8084
rect 3148 7896 3200 7948
rect 2044 7828 2096 7880
rect 2412 7828 2464 7880
rect 4068 7828 4120 7880
rect 4804 7896 4856 7948
rect 5632 7896 5684 7948
rect 5356 7828 5408 7880
rect 4804 7760 4856 7812
rect 6552 7803 6604 7812
rect 6552 7769 6561 7803
rect 6561 7769 6595 7803
rect 6595 7769 6604 7803
rect 6552 7760 6604 7769
rect 5540 7692 5592 7744
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 2582 7590 2634 7642
rect 2646 7590 2698 7642
rect 2710 7590 2762 7642
rect 2774 7590 2826 7642
rect 2838 7590 2890 7642
rect 4307 7590 4359 7642
rect 4371 7590 4423 7642
rect 4435 7590 4487 7642
rect 4499 7590 4551 7642
rect 4563 7590 4615 7642
rect 6032 7590 6084 7642
rect 6096 7590 6148 7642
rect 6160 7590 6212 7642
rect 6224 7590 6276 7642
rect 6288 7590 6340 7642
rect 7757 7590 7809 7642
rect 7821 7590 7873 7642
rect 7885 7590 7937 7642
rect 7949 7590 8001 7642
rect 8013 7590 8065 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 4068 7531 4120 7540
rect 4068 7497 4077 7531
rect 4077 7497 4111 7531
rect 4111 7497 4120 7531
rect 4068 7488 4120 7497
rect 4620 7488 4672 7540
rect 5080 7488 5132 7540
rect 5356 7488 5408 7540
rect 7564 7488 7616 7540
rect 7748 7488 7800 7540
rect 4712 7420 4764 7472
rect 7380 7420 7432 7472
rect 1492 7216 1544 7268
rect 3976 7352 4028 7404
rect 7104 7352 7156 7404
rect 4068 7284 4120 7336
rect 7380 7284 7432 7336
rect 7564 7284 7616 7336
rect 1720 7046 1772 7098
rect 1784 7046 1836 7098
rect 1848 7046 1900 7098
rect 1912 7046 1964 7098
rect 1976 7046 2028 7098
rect 3445 7046 3497 7098
rect 3509 7046 3561 7098
rect 3573 7046 3625 7098
rect 3637 7046 3689 7098
rect 3701 7046 3753 7098
rect 5170 7046 5222 7098
rect 5234 7046 5286 7098
rect 5298 7046 5350 7098
rect 5362 7046 5414 7098
rect 5426 7046 5478 7098
rect 6895 7046 6947 7098
rect 6959 7046 7011 7098
rect 7023 7046 7075 7098
rect 7087 7046 7139 7098
rect 7151 7046 7203 7098
rect 3332 6876 3384 6928
rect 5080 6808 5132 6860
rect 1308 6740 1360 6792
rect 4528 6740 4580 6792
rect 3056 6604 3108 6656
rect 8208 6672 8260 6724
rect 5080 6604 5132 6656
rect 5908 6604 5960 6656
rect 6368 6604 6420 6656
rect 7748 6604 7800 6656
rect 2582 6502 2634 6554
rect 2646 6502 2698 6554
rect 2710 6502 2762 6554
rect 2774 6502 2826 6554
rect 2838 6502 2890 6554
rect 4307 6502 4359 6554
rect 4371 6502 4423 6554
rect 4435 6502 4487 6554
rect 4499 6502 4551 6554
rect 4563 6502 4615 6554
rect 6032 6502 6084 6554
rect 6096 6502 6148 6554
rect 6160 6502 6212 6554
rect 6224 6502 6276 6554
rect 6288 6502 6340 6554
rect 7757 6502 7809 6554
rect 7821 6502 7873 6554
rect 7885 6502 7937 6554
rect 7949 6502 8001 6554
rect 8013 6502 8065 6554
rect 1308 6400 1360 6452
rect 5908 6400 5960 6452
rect 6736 6400 6788 6452
rect 3884 6332 3936 6384
rect 6368 6332 6420 6384
rect 7564 6332 7616 6384
rect 6736 6264 6788 6316
rect 2964 6196 3016 6248
rect 5540 6196 5592 6248
rect 7564 6128 7616 6180
rect 2964 6060 3016 6112
rect 5908 6060 5960 6112
rect 1720 5958 1772 6010
rect 1784 5958 1836 6010
rect 1848 5958 1900 6010
rect 1912 5958 1964 6010
rect 1976 5958 2028 6010
rect 3445 5958 3497 6010
rect 3509 5958 3561 6010
rect 3573 5958 3625 6010
rect 3637 5958 3689 6010
rect 3701 5958 3753 6010
rect 5170 5958 5222 6010
rect 5234 5958 5286 6010
rect 5298 5958 5350 6010
rect 5362 5958 5414 6010
rect 5426 5958 5478 6010
rect 6895 5958 6947 6010
rect 6959 5958 7011 6010
rect 7023 5958 7075 6010
rect 7087 5958 7139 6010
rect 7151 5958 7203 6010
rect 1032 5856 1084 5908
rect 5172 5856 5224 5908
rect 5632 5856 5684 5908
rect 2504 5720 2556 5772
rect 2136 5652 2188 5704
rect 5448 5652 5500 5704
rect 7196 5856 7248 5908
rect 7564 5856 7616 5908
rect 7288 5720 7340 5772
rect 7564 5720 7616 5772
rect 1400 5584 1452 5636
rect 3332 5584 3384 5636
rect 4804 5627 4856 5636
rect 4804 5593 4813 5627
rect 4813 5593 4847 5627
rect 4847 5593 4856 5627
rect 4804 5584 4856 5593
rect 5632 5584 5684 5636
rect 5908 5584 5960 5636
rect 7288 5627 7340 5636
rect 7288 5593 7297 5627
rect 7297 5593 7331 5627
rect 7331 5593 7340 5627
rect 7288 5584 7340 5593
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 3148 5516 3200 5568
rect 3884 5516 3936 5568
rect 2582 5414 2634 5466
rect 2646 5414 2698 5466
rect 2710 5414 2762 5466
rect 2774 5414 2826 5466
rect 2838 5414 2890 5466
rect 4307 5414 4359 5466
rect 4371 5414 4423 5466
rect 4435 5414 4487 5466
rect 4499 5414 4551 5466
rect 4563 5414 4615 5466
rect 6032 5414 6084 5466
rect 6096 5414 6148 5466
rect 6160 5414 6212 5466
rect 6224 5414 6276 5466
rect 6288 5414 6340 5466
rect 7757 5414 7809 5466
rect 7821 5414 7873 5466
rect 7885 5414 7937 5466
rect 7949 5414 8001 5466
rect 8013 5414 8065 5466
rect 6276 5312 6328 5364
rect 6460 5312 6512 5364
rect 4896 5244 4948 5296
rect 5172 5287 5224 5296
rect 5172 5253 5181 5287
rect 5181 5253 5215 5287
rect 5215 5253 5224 5287
rect 5172 5244 5224 5253
rect 5540 5244 5592 5296
rect 3056 5176 3108 5228
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 7196 5176 7248 5228
rect 4896 5040 4948 5092
rect 2780 4972 2832 5024
rect 3056 5015 3108 5024
rect 3056 4981 3065 5015
rect 3065 4981 3099 5015
rect 3099 4981 3108 5015
rect 3056 4972 3108 4981
rect 7472 4972 7524 5024
rect 1720 4870 1772 4922
rect 1784 4870 1836 4922
rect 1848 4870 1900 4922
rect 1912 4870 1964 4922
rect 1976 4870 2028 4922
rect 3445 4870 3497 4922
rect 3509 4870 3561 4922
rect 3573 4870 3625 4922
rect 3637 4870 3689 4922
rect 3701 4870 3753 4922
rect 5170 4870 5222 4922
rect 5234 4870 5286 4922
rect 5298 4870 5350 4922
rect 5362 4870 5414 4922
rect 5426 4870 5478 4922
rect 6895 4870 6947 4922
rect 6959 4870 7011 4922
rect 7023 4870 7075 4922
rect 7087 4870 7139 4922
rect 7151 4870 7203 4922
rect 3700 4768 3752 4820
rect 3884 4768 3936 4820
rect 4712 4768 4764 4820
rect 3792 4632 3844 4684
rect 2780 4564 2832 4616
rect 3976 4564 4028 4616
rect 1584 4428 1636 4480
rect 6644 4496 6696 4548
rect 6828 4496 6880 4548
rect 5908 4428 5960 4480
rect 6368 4428 6420 4480
rect 2582 4326 2634 4378
rect 2646 4326 2698 4378
rect 2710 4326 2762 4378
rect 2774 4326 2826 4378
rect 2838 4326 2890 4378
rect 4307 4326 4359 4378
rect 4371 4326 4423 4378
rect 4435 4326 4487 4378
rect 4499 4326 4551 4378
rect 4563 4326 4615 4378
rect 6032 4326 6084 4378
rect 6096 4326 6148 4378
rect 6160 4326 6212 4378
rect 6224 4326 6276 4378
rect 6288 4326 6340 4378
rect 7757 4326 7809 4378
rect 7821 4326 7873 4378
rect 7885 4326 7937 4378
rect 7949 4326 8001 4378
rect 8013 4326 8065 4378
rect 4068 4224 4120 4276
rect 4252 4224 4304 4276
rect 4896 4224 4948 4276
rect 6644 4224 6696 4276
rect 8116 4224 8168 4276
rect 3240 4088 3292 4140
rect 4712 4156 4764 4208
rect 5724 4156 5776 4208
rect 5448 4088 5500 4140
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 3240 3952 3292 4004
rect 3700 3952 3752 4004
rect 2044 3884 2096 3936
rect 3792 3884 3844 3936
rect 1720 3782 1772 3834
rect 1784 3782 1836 3834
rect 1848 3782 1900 3834
rect 1912 3782 1964 3834
rect 1976 3782 2028 3834
rect 3445 3782 3497 3834
rect 3509 3782 3561 3834
rect 3573 3782 3625 3834
rect 3637 3782 3689 3834
rect 3701 3782 3753 3834
rect 5170 3782 5222 3834
rect 5234 3782 5286 3834
rect 5298 3782 5350 3834
rect 5362 3782 5414 3834
rect 5426 3782 5478 3834
rect 6895 3782 6947 3834
rect 6959 3782 7011 3834
rect 7023 3782 7075 3834
rect 7087 3782 7139 3834
rect 7151 3782 7203 3834
rect 3700 3680 3752 3732
rect 4252 3680 4304 3732
rect 5724 3680 5776 3732
rect 4988 3544 5040 3596
rect 7656 3544 7708 3596
rect 2044 3476 2096 3528
rect 5448 3476 5500 3528
rect 5724 3476 5776 3528
rect 2964 3408 3016 3460
rect 2504 3340 2556 3392
rect 5080 3340 5132 3392
rect 5816 3340 5868 3392
rect 2582 3238 2634 3290
rect 2646 3238 2698 3290
rect 2710 3238 2762 3290
rect 2774 3238 2826 3290
rect 2838 3238 2890 3290
rect 4307 3238 4359 3290
rect 4371 3238 4423 3290
rect 4435 3238 4487 3290
rect 4499 3238 4551 3290
rect 4563 3238 4615 3290
rect 6032 3238 6084 3290
rect 6096 3238 6148 3290
rect 6160 3238 6212 3290
rect 6224 3238 6276 3290
rect 6288 3238 6340 3290
rect 7757 3238 7809 3290
rect 7821 3238 7873 3290
rect 7885 3238 7937 3290
rect 7949 3238 8001 3290
rect 8013 3238 8065 3290
rect 8392 3136 8444 3188
rect 3332 3111 3384 3120
rect 3332 3077 3341 3111
rect 3341 3077 3375 3111
rect 3375 3077 3384 3111
rect 3332 3068 3384 3077
rect 3792 3068 3844 3120
rect 5816 3068 5868 3120
rect 6460 3111 6512 3120
rect 6460 3077 6469 3111
rect 6469 3077 6503 3111
rect 6503 3077 6512 3111
rect 6460 3068 6512 3077
rect 296 3000 348 3052
rect 1492 3043 1544 3052
rect 1492 3009 1501 3043
rect 1501 3009 1535 3043
rect 1535 3009 1544 3043
rect 1492 3000 1544 3009
rect 4804 3000 4856 3052
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 7564 2932 7616 2984
rect 3240 2864 3292 2916
rect 8576 2864 8628 2916
rect 756 2796 808 2848
rect 5724 2796 5776 2848
rect 6000 2796 6052 2848
rect 1720 2694 1772 2746
rect 1784 2694 1836 2746
rect 1848 2694 1900 2746
rect 1912 2694 1964 2746
rect 1976 2694 2028 2746
rect 3445 2694 3497 2746
rect 3509 2694 3561 2746
rect 3573 2694 3625 2746
rect 3637 2694 3689 2746
rect 3701 2694 3753 2746
rect 5170 2694 5222 2746
rect 5234 2694 5286 2746
rect 5298 2694 5350 2746
rect 5362 2694 5414 2746
rect 5426 2694 5478 2746
rect 6895 2694 6947 2746
rect 6959 2694 7011 2746
rect 7023 2694 7075 2746
rect 7087 2694 7139 2746
rect 7151 2694 7203 2746
rect 3884 2592 3936 2644
rect 5172 2592 5224 2644
rect 6460 2592 6512 2644
rect 6000 2567 6052 2576
rect 6000 2533 6009 2567
rect 6009 2533 6043 2567
rect 6043 2533 6052 2567
rect 6000 2524 6052 2533
rect 2780 2456 2832 2508
rect 5908 2456 5960 2508
rect 7288 2499 7340 2508
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 3240 2388 3292 2440
rect 5632 2388 5684 2440
rect 2136 2252 2188 2304
rect 2582 2150 2634 2202
rect 2646 2150 2698 2202
rect 2710 2150 2762 2202
rect 2774 2150 2826 2202
rect 2838 2150 2890 2202
rect 4307 2150 4359 2202
rect 4371 2150 4423 2202
rect 4435 2150 4487 2202
rect 4499 2150 4551 2202
rect 4563 2150 4615 2202
rect 6032 2150 6084 2202
rect 6096 2150 6148 2202
rect 6160 2150 6212 2202
rect 6224 2150 6276 2202
rect 6288 2150 6340 2202
rect 7757 2150 7809 2202
rect 7821 2150 7873 2202
rect 7885 2150 7937 2202
rect 7949 2150 8001 2202
rect 8013 2150 8065 2202
rect 3148 1980 3200 2032
rect 4160 1980 4212 2032
rect 5172 2023 5224 2032
rect 5172 1989 5181 2023
rect 5181 1989 5215 2023
rect 5215 1989 5224 2023
rect 5172 1980 5224 1989
rect 8116 2048 8168 2100
rect 6552 1980 6604 2032
rect 7288 2023 7340 2032
rect 7288 1989 7297 2023
rect 7297 1989 7331 2023
rect 7331 1989 7340 2023
rect 7288 1980 7340 1989
rect 1492 1844 1544 1896
rect 4988 1912 5040 1964
rect 3792 1844 3844 1896
rect 1720 1606 1772 1658
rect 1784 1606 1836 1658
rect 1848 1606 1900 1658
rect 1912 1606 1964 1658
rect 1976 1606 2028 1658
rect 3445 1606 3497 1658
rect 3509 1606 3561 1658
rect 3573 1606 3625 1658
rect 3637 1606 3689 1658
rect 3701 1606 3753 1658
rect 5170 1606 5222 1658
rect 5234 1606 5286 1658
rect 5298 1606 5350 1658
rect 5362 1606 5414 1658
rect 5426 1606 5478 1658
rect 6895 1606 6947 1658
rect 6959 1606 7011 1658
rect 7023 1606 7075 1658
rect 7087 1606 7139 1658
rect 7151 1606 7203 1658
rect 7196 1504 7248 1556
rect 8208 1504 8260 1556
rect 2780 1368 2832 1420
rect 4160 1411 4212 1420
rect 4160 1377 4169 1411
rect 4169 1377 4203 1411
rect 4203 1377 4212 1411
rect 4160 1368 4212 1377
rect 6828 1300 6880 1352
rect 7288 1343 7340 1352
rect 7288 1309 7297 1343
rect 7297 1309 7331 1343
rect 7331 1309 7340 1343
rect 7288 1300 7340 1309
rect 2228 1232 2280 1284
rect 4988 1232 5040 1284
rect 6644 1232 6696 1284
rect 1216 1164 1268 1216
rect 4804 1164 4856 1216
rect 2582 1062 2634 1114
rect 2646 1062 2698 1114
rect 2710 1062 2762 1114
rect 2774 1062 2826 1114
rect 2838 1062 2890 1114
rect 4307 1062 4359 1114
rect 4371 1062 4423 1114
rect 4435 1062 4487 1114
rect 4499 1062 4551 1114
rect 4563 1062 4615 1114
rect 6032 1062 6084 1114
rect 6096 1062 6148 1114
rect 6160 1062 6212 1114
rect 6224 1062 6276 1114
rect 6288 1062 6340 1114
rect 7757 1062 7809 1114
rect 7821 1062 7873 1114
rect 7885 1062 7937 1114
rect 7949 1062 8001 1114
rect 8013 1062 8065 1114
<< metal2 >>
rect 754 9330 810 10000
rect 754 9302 980 9330
rect 754 9200 810 9302
rect 952 8634 980 9302
rect 1030 9200 1086 10000
rect 1306 9200 1362 10000
rect 1582 9330 1638 10000
rect 1412 9302 1638 9330
rect 940 8628 992 8634
rect 940 8570 992 8576
rect 1044 5914 1072 9200
rect 1320 6798 1348 9200
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1320 6458 1348 6734
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 1032 5908 1084 5914
rect 1032 5850 1084 5856
rect 1412 5642 1440 9302
rect 1582 9200 1638 9302
rect 1858 9330 1914 10000
rect 1858 9302 2084 9330
rect 1858 9200 1914 9302
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1780 8401 1808 8434
rect 1582 8392 1638 8401
rect 1582 8327 1638 8336
rect 1766 8392 1822 8401
rect 1766 8327 1822 8336
rect 1596 7546 1624 8327
rect 1720 8188 2028 8197
rect 1720 8186 1726 8188
rect 1782 8186 1806 8188
rect 1862 8186 1886 8188
rect 1942 8186 1966 8188
rect 2022 8186 2028 8188
rect 1782 8134 1784 8186
rect 1964 8134 1966 8186
rect 1720 8132 1726 8134
rect 1782 8132 1806 8134
rect 1862 8132 1886 8134
rect 1942 8132 1966 8134
rect 2022 8132 2028 8134
rect 1720 8123 2028 8132
rect 2056 8090 2084 9302
rect 2134 9200 2190 10000
rect 2410 9200 2466 10000
rect 2686 9200 2742 10000
rect 2962 9330 3018 10000
rect 2962 9302 3188 9330
rect 2962 9200 3018 9302
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2056 7886 2084 8026
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1492 7268 1544 7274
rect 1492 7210 1544 7216
rect 1504 7041 1532 7210
rect 1720 7100 2028 7109
rect 1720 7098 1726 7100
rect 1782 7098 1806 7100
rect 1862 7098 1886 7100
rect 1942 7098 1966 7100
rect 2022 7098 2028 7100
rect 1782 7046 1784 7098
rect 1964 7046 1966 7098
rect 1720 7044 1726 7046
rect 1782 7044 1806 7046
rect 1862 7044 1886 7046
rect 1942 7044 1966 7046
rect 2022 7044 2028 7046
rect 1490 7032 1546 7041
rect 1720 7035 2028 7044
rect 1490 6967 1546 6976
rect 1720 6012 2028 6021
rect 1720 6010 1726 6012
rect 1782 6010 1806 6012
rect 1862 6010 1886 6012
rect 1942 6010 1966 6012
rect 2022 6010 2028 6012
rect 1782 5958 1784 6010
rect 1964 5958 1966 6010
rect 1720 5956 1726 5958
rect 1782 5956 1806 5958
rect 1862 5956 1886 5958
rect 1942 5956 1966 5958
rect 2022 5956 2028 5958
rect 1720 5947 2028 5956
rect 2148 5710 2176 9200
rect 2424 7886 2452 9200
rect 2700 8922 2728 9200
rect 2516 8894 2728 8922
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2516 5778 2544 8894
rect 2582 8732 2890 8741
rect 2582 8730 2588 8732
rect 2644 8730 2668 8732
rect 2724 8730 2748 8732
rect 2804 8730 2828 8732
rect 2884 8730 2890 8732
rect 2644 8678 2646 8730
rect 2826 8678 2828 8730
rect 2582 8676 2588 8678
rect 2644 8676 2668 8678
rect 2724 8676 2748 8678
rect 2804 8676 2828 8678
rect 2884 8676 2890 8678
rect 2582 8667 2890 8676
rect 3160 7954 3188 9302
rect 3238 9200 3294 10000
rect 3514 9330 3570 10000
rect 3514 9302 3740 9330
rect 3514 9200 3570 9302
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2582 7644 2890 7653
rect 2582 7642 2588 7644
rect 2644 7642 2668 7644
rect 2724 7642 2748 7644
rect 2804 7642 2828 7644
rect 2884 7642 2890 7644
rect 2644 7590 2646 7642
rect 2826 7590 2828 7642
rect 2582 7588 2588 7590
rect 2644 7588 2668 7590
rect 2724 7588 2748 7590
rect 2804 7588 2828 7590
rect 2884 7588 2890 7590
rect 2582 7579 2890 7588
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2582 6556 2890 6565
rect 2582 6554 2588 6556
rect 2644 6554 2668 6556
rect 2724 6554 2748 6556
rect 2804 6554 2828 6556
rect 2884 6554 2890 6556
rect 2644 6502 2646 6554
rect 2826 6502 2828 6554
rect 2582 6500 2588 6502
rect 2644 6500 2668 6502
rect 2724 6500 2748 6502
rect 2804 6500 2828 6502
rect 2884 6500 2890 6502
rect 2582 6491 2890 6500
rect 2962 6352 3018 6361
rect 2962 6287 3018 6296
rect 2976 6254 3004 6287
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 1400 5636 1452 5642
rect 1400 5578 1452 5584
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 1504 3058 1532 5510
rect 1720 4924 2028 4933
rect 1720 4922 1726 4924
rect 1782 4922 1806 4924
rect 1862 4922 1886 4924
rect 1942 4922 1966 4924
rect 2022 4922 2028 4924
rect 1782 4870 1784 4922
rect 1964 4870 1966 4922
rect 1720 4868 1726 4870
rect 1782 4868 1806 4870
rect 1862 4868 1886 4870
rect 1942 4868 1966 4870
rect 2022 4868 2028 4870
rect 1720 4859 2028 4868
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 296 3052 348 3058
rect 296 2994 348 3000
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 308 800 336 2994
rect 756 2848 808 2854
rect 756 2790 808 2796
rect 768 800 796 2790
rect 1492 1896 1544 1902
rect 1492 1838 1544 1844
rect 1504 1601 1532 1838
rect 1490 1592 1546 1601
rect 1490 1527 1546 1536
rect 1596 1442 1624 4422
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1720 3836 2028 3845
rect 1720 3834 1726 3836
rect 1782 3834 1806 3836
rect 1862 3834 1886 3836
rect 1942 3834 1966 3836
rect 2022 3834 2028 3836
rect 1782 3782 1784 3834
rect 1964 3782 1966 3834
rect 1720 3780 1726 3782
rect 1782 3780 1806 3782
rect 1862 3780 1886 3782
rect 1942 3780 1966 3782
rect 2022 3780 2028 3782
rect 1720 3771 2028 3780
rect 2056 3534 2084 3878
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1720 2748 2028 2757
rect 1720 2746 1726 2748
rect 1782 2746 1806 2748
rect 1862 2746 1886 2748
rect 1942 2746 1966 2748
rect 2022 2746 2028 2748
rect 1782 2694 1784 2746
rect 1964 2694 1966 2746
rect 1720 2692 1726 2694
rect 1782 2692 1806 2694
rect 1862 2692 1886 2694
rect 1942 2692 1966 2694
rect 2022 2692 2028 2694
rect 1720 2683 2028 2692
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 1720 1660 2028 1669
rect 1720 1658 1726 1660
rect 1782 1658 1806 1660
rect 1862 1658 1886 1660
rect 1942 1658 1966 1660
rect 2022 1658 2028 1660
rect 1782 1606 1784 1658
rect 1964 1606 1966 1658
rect 1720 1604 1726 1606
rect 1782 1604 1806 1606
rect 1862 1604 1886 1606
rect 1942 1604 1966 1606
rect 2022 1604 2028 1606
rect 1720 1595 2028 1604
rect 1596 1414 1716 1442
rect 1216 1216 1268 1222
rect 1216 1158 1268 1164
rect 1228 800 1256 1158
rect 1688 800 1716 1414
rect 2148 800 2176 2246
rect 2240 1290 2268 5510
rect 2582 5468 2890 5477
rect 2582 5466 2588 5468
rect 2644 5466 2668 5468
rect 2724 5466 2748 5468
rect 2804 5466 2828 5468
rect 2884 5466 2890 5468
rect 2644 5414 2646 5466
rect 2826 5414 2828 5466
rect 2582 5412 2588 5414
rect 2644 5412 2668 5414
rect 2724 5412 2748 5414
rect 2804 5412 2828 5414
rect 2884 5412 2890 5414
rect 2582 5403 2890 5412
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4622 2820 4966
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2582 4380 2890 4389
rect 2582 4378 2588 4380
rect 2644 4378 2668 4380
rect 2724 4378 2748 4380
rect 2804 4378 2828 4380
rect 2884 4378 2890 4380
rect 2644 4326 2646 4378
rect 2826 4326 2828 4378
rect 2582 4324 2588 4326
rect 2644 4324 2668 4326
rect 2724 4324 2748 4326
rect 2804 4324 2828 4326
rect 2884 4324 2890 4326
rect 2582 4315 2890 4324
rect 2976 3641 3004 6054
rect 3068 5681 3096 6598
rect 3054 5672 3110 5681
rect 3054 5607 3110 5616
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3068 5030 3096 5170
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2962 3632 3018 3641
rect 2962 3567 3018 3576
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2228 1284 2280 1290
rect 2228 1226 2280 1232
rect 2516 898 2544 3334
rect 2582 3292 2890 3301
rect 2582 3290 2588 3292
rect 2644 3290 2668 3292
rect 2724 3290 2748 3292
rect 2804 3290 2828 3292
rect 2884 3290 2890 3292
rect 2644 3238 2646 3290
rect 2826 3238 2828 3290
rect 2582 3236 2588 3238
rect 2644 3236 2668 3238
rect 2724 3236 2748 3238
rect 2804 3236 2828 3238
rect 2884 3236 2890 3238
rect 2582 3227 2890 3236
rect 2778 2952 2834 2961
rect 2778 2887 2834 2896
rect 2792 2514 2820 2887
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2582 2204 2890 2213
rect 2582 2202 2588 2204
rect 2644 2202 2668 2204
rect 2724 2202 2748 2204
rect 2804 2202 2828 2204
rect 2884 2202 2890 2204
rect 2644 2150 2646 2202
rect 2826 2150 2828 2202
rect 2582 2148 2588 2150
rect 2644 2148 2668 2150
rect 2724 2148 2748 2150
rect 2804 2148 2828 2150
rect 2884 2148 2890 2150
rect 2582 2139 2890 2148
rect 2778 2000 2834 2009
rect 2778 1935 2834 1944
rect 2792 1426 2820 1935
rect 2780 1420 2832 1426
rect 2780 1362 2832 1368
rect 2582 1116 2890 1125
rect 2582 1114 2588 1116
rect 2644 1114 2668 1116
rect 2724 1114 2748 1116
rect 2804 1114 2828 1116
rect 2884 1114 2890 1116
rect 2644 1062 2646 1114
rect 2826 1062 2828 1114
rect 2582 1060 2588 1062
rect 2644 1060 2668 1062
rect 2724 1060 2748 1062
rect 2804 1060 2828 1062
rect 2884 1060 2890 1062
rect 2582 1051 2890 1060
rect 2976 921 3004 3402
rect 2962 912 3018 921
rect 2516 870 2636 898
rect 2608 800 2636 870
rect 2962 847 3018 856
rect 3068 800 3096 4966
rect 3160 2038 3188 5510
rect 3252 4146 3280 9200
rect 3422 9072 3478 9081
rect 3422 9007 3478 9016
rect 3436 8906 3464 9007
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3712 8634 3740 9302
rect 3790 9200 3846 10000
rect 4066 9330 4122 10000
rect 4342 9330 4398 10000
rect 3988 9302 4122 9330
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3445 8188 3753 8197
rect 3445 8186 3451 8188
rect 3507 8186 3531 8188
rect 3587 8186 3611 8188
rect 3667 8186 3691 8188
rect 3747 8186 3753 8188
rect 3507 8134 3509 8186
rect 3689 8134 3691 8186
rect 3445 8132 3451 8134
rect 3507 8132 3531 8134
rect 3587 8132 3611 8134
rect 3667 8132 3691 8134
rect 3747 8132 3753 8134
rect 3445 8123 3753 8132
rect 3330 7440 3386 7449
rect 3330 7375 3386 7384
rect 3344 6934 3372 7375
rect 3445 7100 3753 7109
rect 3445 7098 3451 7100
rect 3507 7098 3531 7100
rect 3587 7098 3611 7100
rect 3667 7098 3691 7100
rect 3747 7098 3753 7100
rect 3507 7046 3509 7098
rect 3689 7046 3691 7098
rect 3445 7044 3451 7046
rect 3507 7044 3531 7046
rect 3587 7044 3611 7046
rect 3667 7044 3691 7046
rect 3747 7044 3753 7046
rect 3445 7035 3753 7044
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3445 6012 3753 6021
rect 3445 6010 3451 6012
rect 3507 6010 3531 6012
rect 3587 6010 3611 6012
rect 3667 6010 3691 6012
rect 3747 6010 3753 6012
rect 3507 5958 3509 6010
rect 3689 5958 3691 6010
rect 3445 5956 3451 5958
rect 3507 5956 3531 5958
rect 3587 5956 3611 5958
rect 3667 5956 3691 5958
rect 3747 5956 3753 5958
rect 3445 5947 3753 5956
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3252 2922 3280 3946
rect 3344 3126 3372 5578
rect 3445 4924 3753 4933
rect 3445 4922 3451 4924
rect 3507 4922 3531 4924
rect 3587 4922 3611 4924
rect 3667 4922 3691 4924
rect 3747 4922 3753 4924
rect 3507 4870 3509 4922
rect 3689 4870 3691 4922
rect 3445 4868 3451 4870
rect 3507 4868 3531 4870
rect 3587 4868 3611 4870
rect 3667 4868 3691 4870
rect 3747 4868 3753 4870
rect 3445 4859 3753 4868
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3712 4010 3740 4762
rect 3804 4690 3832 9200
rect 3882 8936 3938 8945
rect 3882 8871 3938 8880
rect 3896 6390 3924 8871
rect 3988 7410 4016 9302
rect 4066 9200 4122 9302
rect 4172 9302 4398 9330
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 7546 4108 7822
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 4826 3924 5510
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3882 4720 3938 4729
rect 3792 4684 3844 4690
rect 3882 4655 3938 4664
rect 3792 4626 3844 4632
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3445 3836 3753 3845
rect 3445 3834 3451 3836
rect 3507 3834 3531 3836
rect 3587 3834 3611 3836
rect 3667 3834 3691 3836
rect 3747 3834 3753 3836
rect 3507 3782 3509 3834
rect 3689 3782 3691 3834
rect 3445 3780 3451 3782
rect 3507 3780 3531 3782
rect 3587 3780 3611 3782
rect 3667 3780 3691 3782
rect 3747 3780 3753 3782
rect 3445 3771 3753 3780
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3712 2938 3740 3674
rect 3804 3126 3832 3878
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3240 2916 3292 2922
rect 3712 2910 3832 2938
rect 3240 2858 3292 2864
rect 3252 2446 3280 2858
rect 3445 2748 3753 2757
rect 3445 2746 3451 2748
rect 3507 2746 3531 2748
rect 3587 2746 3611 2748
rect 3667 2746 3691 2748
rect 3747 2746 3753 2748
rect 3507 2694 3509 2746
rect 3689 2694 3691 2746
rect 3445 2692 3451 2694
rect 3507 2692 3531 2694
rect 3587 2692 3611 2694
rect 3667 2692 3691 2694
rect 3747 2692 3753 2694
rect 3445 2683 3753 2692
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3148 2032 3200 2038
rect 3148 1974 3200 1980
rect 294 0 350 800
rect 754 0 810 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3160 762 3188 1974
rect 3804 1902 3832 2910
rect 3896 2650 3924 4655
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 3445 1660 3753 1669
rect 3445 1658 3451 1660
rect 3507 1658 3531 1660
rect 3587 1658 3611 1660
rect 3667 1658 3691 1660
rect 3747 1658 3753 1660
rect 3507 1606 3509 1658
rect 3689 1606 3691 1658
rect 3445 1604 3451 1606
rect 3507 1604 3531 1606
rect 3587 1604 3611 1606
rect 3667 1604 3691 1606
rect 3747 1604 3753 1606
rect 3445 1595 3753 1604
rect 3436 870 3556 898
rect 3436 762 3464 870
rect 3528 800 3556 870
rect 3988 800 4016 4558
rect 4080 4282 4108 7278
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 4080 1850 4108 4111
rect 4172 2038 4200 9302
rect 4342 9200 4398 9302
rect 4618 9330 4674 10000
rect 4618 9302 4844 9330
rect 4618 9200 4674 9302
rect 4307 8732 4615 8741
rect 4307 8730 4313 8732
rect 4369 8730 4393 8732
rect 4449 8730 4473 8732
rect 4529 8730 4553 8732
rect 4609 8730 4615 8732
rect 4369 8678 4371 8730
rect 4551 8678 4553 8730
rect 4307 8676 4313 8678
rect 4369 8676 4393 8678
rect 4449 8676 4473 8678
rect 4529 8676 4553 8678
rect 4609 8676 4615 8678
rect 4307 8667 4615 8676
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4632 7857 4660 8366
rect 4710 7984 4766 7993
rect 4816 7954 4844 9302
rect 4894 9200 4950 10000
rect 5170 9330 5226 10000
rect 5446 9330 5502 10000
rect 5092 9302 5226 9330
rect 4710 7919 4766 7928
rect 4804 7948 4856 7954
rect 4618 7848 4674 7857
rect 4618 7783 4674 7792
rect 4307 7644 4615 7653
rect 4307 7642 4313 7644
rect 4369 7642 4393 7644
rect 4449 7642 4473 7644
rect 4529 7642 4553 7644
rect 4609 7642 4615 7644
rect 4369 7590 4371 7642
rect 4551 7590 4553 7642
rect 4307 7588 4313 7590
rect 4369 7588 4393 7590
rect 4449 7588 4473 7590
rect 4529 7588 4553 7590
rect 4609 7588 4615 7590
rect 4307 7579 4615 7588
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4528 6792 4580 6798
rect 4526 6760 4528 6769
rect 4580 6760 4582 6769
rect 4632 6746 4660 7482
rect 4724 7478 4752 7919
rect 4804 7890 4856 7896
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4632 6718 4752 6746
rect 4526 6695 4582 6704
rect 4307 6556 4615 6565
rect 4307 6554 4313 6556
rect 4369 6554 4393 6556
rect 4449 6554 4473 6556
rect 4529 6554 4553 6556
rect 4609 6554 4615 6556
rect 4369 6502 4371 6554
rect 4551 6502 4553 6554
rect 4307 6500 4313 6502
rect 4369 6500 4393 6502
rect 4449 6500 4473 6502
rect 4529 6500 4553 6502
rect 4609 6500 4615 6502
rect 4307 6491 4615 6500
rect 4307 5468 4615 5477
rect 4307 5466 4313 5468
rect 4369 5466 4393 5468
rect 4449 5466 4473 5468
rect 4529 5466 4553 5468
rect 4609 5466 4615 5468
rect 4369 5414 4371 5466
rect 4551 5414 4553 5466
rect 4307 5412 4313 5414
rect 4369 5412 4393 5414
rect 4449 5412 4473 5414
rect 4529 5412 4553 5414
rect 4609 5412 4615 5414
rect 4307 5403 4615 5412
rect 4724 4826 4752 6718
rect 4816 6225 4844 7754
rect 4802 6216 4858 6225
rect 4802 6151 4858 6160
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4307 4380 4615 4389
rect 4307 4378 4313 4380
rect 4369 4378 4393 4380
rect 4449 4378 4473 4380
rect 4529 4378 4553 4380
rect 4609 4378 4615 4380
rect 4369 4326 4371 4378
rect 4551 4326 4553 4378
rect 4307 4324 4313 4326
rect 4369 4324 4393 4326
rect 4449 4324 4473 4326
rect 4529 4324 4553 4326
rect 4609 4324 4615 4326
rect 4307 4315 4615 4324
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4264 3738 4292 4218
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4307 3292 4615 3301
rect 4307 3290 4313 3292
rect 4369 3290 4393 3292
rect 4449 3290 4473 3292
rect 4529 3290 4553 3292
rect 4609 3290 4615 3292
rect 4369 3238 4371 3290
rect 4551 3238 4553 3290
rect 4307 3236 4313 3238
rect 4369 3236 4393 3238
rect 4449 3236 4473 3238
rect 4529 3236 4553 3238
rect 4609 3236 4615 3238
rect 4307 3227 4615 3236
rect 4307 2204 4615 2213
rect 4307 2202 4313 2204
rect 4369 2202 4393 2204
rect 4449 2202 4473 2204
rect 4529 2202 4553 2204
rect 4609 2202 4615 2204
rect 4369 2150 4371 2202
rect 4551 2150 4553 2202
rect 4307 2148 4313 2150
rect 4369 2148 4393 2150
rect 4449 2148 4473 2150
rect 4529 2148 4553 2150
rect 4609 2148 4615 2150
rect 4307 2139 4615 2148
rect 4160 2032 4212 2038
rect 4160 1974 4212 1980
rect 4080 1822 4200 1850
rect 4172 1426 4200 1822
rect 4160 1420 4212 1426
rect 4160 1362 4212 1368
rect 4307 1116 4615 1125
rect 4307 1114 4313 1116
rect 4369 1114 4393 1116
rect 4449 1114 4473 1116
rect 4529 1114 4553 1116
rect 4609 1114 4615 1116
rect 4369 1062 4371 1114
rect 4551 1062 4553 1114
rect 4307 1060 4313 1062
rect 4369 1060 4393 1062
rect 4449 1060 4473 1062
rect 4529 1060 4553 1062
rect 4609 1060 4615 1062
rect 4307 1051 4615 1060
rect 4448 870 4568 898
rect 4448 800 4476 870
rect 3160 734 3464 762
rect 3514 0 3570 800
rect 3974 0 4030 800
rect 4434 0 4490 800
rect 4540 762 4568 870
rect 4724 762 4752 4150
rect 4816 3754 4844 5578
rect 4908 5302 4936 9200
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4908 4282 4936 5034
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4816 3726 4936 3754
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4816 1222 4844 2994
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4908 800 4936 3726
rect 5000 3602 5028 8230
rect 5092 7546 5120 9302
rect 5170 9200 5226 9302
rect 5276 9302 5502 9330
rect 5276 8294 5304 9302
rect 5446 9200 5502 9302
rect 5722 9200 5778 10000
rect 5998 9330 6054 10000
rect 5828 9302 6054 9330
rect 5448 8424 5500 8430
rect 5630 8392 5686 8401
rect 5500 8372 5580 8378
rect 5448 8366 5580 8372
rect 5460 8350 5580 8366
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5170 8188 5478 8197
rect 5170 8186 5176 8188
rect 5232 8186 5256 8188
rect 5312 8186 5336 8188
rect 5392 8186 5416 8188
rect 5472 8186 5478 8188
rect 5232 8134 5234 8186
rect 5414 8134 5416 8186
rect 5170 8132 5176 8134
rect 5232 8132 5256 8134
rect 5312 8132 5336 8134
rect 5392 8132 5416 8134
rect 5472 8132 5478 8134
rect 5170 8123 5478 8132
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7426 5212 8026
rect 5552 7970 5580 8350
rect 5630 8327 5686 8336
rect 5644 8090 5672 8327
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5460 7942 5580 7970
rect 5632 7948 5684 7954
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5368 7546 5396 7822
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5092 7398 5212 7426
rect 5092 6866 5120 7398
rect 5460 7313 5488 7942
rect 5632 7890 5684 7896
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5446 7304 5502 7313
rect 5446 7239 5502 7248
rect 5170 7100 5478 7109
rect 5170 7098 5176 7100
rect 5232 7098 5256 7100
rect 5312 7098 5336 7100
rect 5392 7098 5416 7100
rect 5472 7098 5478 7100
rect 5232 7046 5234 7098
rect 5414 7046 5416 7098
rect 5170 7044 5176 7046
rect 5232 7044 5256 7046
rect 5312 7044 5336 7046
rect 5392 7044 5416 7046
rect 5472 7044 5478 7046
rect 5170 7035 5478 7044
rect 5552 6914 5580 7686
rect 5460 6886 5580 6914
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5092 3482 5120 6598
rect 5460 6361 5488 6886
rect 5446 6352 5502 6361
rect 5446 6287 5502 6296
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5170 6012 5478 6021
rect 5170 6010 5176 6012
rect 5232 6010 5256 6012
rect 5312 6010 5336 6012
rect 5392 6010 5416 6012
rect 5472 6010 5478 6012
rect 5232 5958 5234 6010
rect 5414 5958 5416 6010
rect 5170 5956 5176 5958
rect 5232 5956 5256 5958
rect 5312 5956 5336 5958
rect 5392 5956 5416 5958
rect 5472 5956 5478 5958
rect 5170 5947 5478 5956
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5184 5302 5212 5850
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5460 5012 5488 5646
rect 5552 5302 5580 6190
rect 5644 5914 5672 7890
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5460 4984 5580 5012
rect 5170 4924 5478 4933
rect 5170 4922 5176 4924
rect 5232 4922 5256 4924
rect 5312 4922 5336 4924
rect 5392 4922 5416 4924
rect 5472 4922 5478 4924
rect 5232 4870 5234 4922
rect 5414 4870 5416 4922
rect 5170 4868 5176 4870
rect 5232 4868 5256 4870
rect 5312 4868 5336 4870
rect 5392 4868 5416 4870
rect 5472 4868 5478 4870
rect 5170 4859 5478 4868
rect 5552 4706 5580 4984
rect 5460 4678 5580 4706
rect 5460 4146 5488 4678
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5170 3836 5478 3845
rect 5170 3834 5176 3836
rect 5232 3834 5256 3836
rect 5312 3834 5336 3836
rect 5392 3834 5416 3836
rect 5472 3834 5478 3836
rect 5232 3782 5234 3834
rect 5414 3782 5416 3834
rect 5170 3780 5176 3782
rect 5232 3780 5256 3782
rect 5312 3780 5336 3782
rect 5392 3780 5416 3782
rect 5472 3780 5478 3782
rect 5170 3771 5478 3780
rect 5000 3454 5120 3482
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5000 1970 5028 3454
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4988 1964 5040 1970
rect 4988 1906 5040 1912
rect 4988 1284 5040 1290
rect 4988 1226 5040 1232
rect 5000 921 5028 1226
rect 4986 912 5042 921
rect 4986 847 5042 856
rect 4540 734 4752 762
rect 4894 0 4950 800
rect 5092 762 5120 3334
rect 5460 2938 5488 3470
rect 5460 2910 5580 2938
rect 5170 2748 5478 2757
rect 5170 2746 5176 2748
rect 5232 2746 5256 2748
rect 5312 2746 5336 2748
rect 5392 2746 5416 2748
rect 5472 2746 5478 2748
rect 5232 2694 5234 2746
rect 5414 2694 5416 2746
rect 5170 2692 5176 2694
rect 5232 2692 5256 2694
rect 5312 2692 5336 2694
rect 5392 2692 5416 2694
rect 5472 2692 5478 2694
rect 5170 2683 5478 2692
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5184 2038 5212 2586
rect 5552 2530 5580 2910
rect 5460 2502 5580 2530
rect 5172 2032 5224 2038
rect 5172 1974 5224 1980
rect 5460 1873 5488 2502
rect 5644 2446 5672 5578
rect 5736 4214 5764 9200
rect 5828 4298 5856 9302
rect 5906 9208 5962 9217
rect 5998 9200 6054 9302
rect 6274 9330 6330 10000
rect 6550 9330 6606 10000
rect 6826 9330 6882 10000
rect 6274 9302 6500 9330
rect 6274 9200 6330 9302
rect 5906 9143 5962 9152
rect 5920 6662 5948 9143
rect 6032 8732 6340 8741
rect 6032 8730 6038 8732
rect 6094 8730 6118 8732
rect 6174 8730 6198 8732
rect 6254 8730 6278 8732
rect 6334 8730 6340 8732
rect 6094 8678 6096 8730
rect 6276 8678 6278 8730
rect 6032 8676 6038 8678
rect 6094 8676 6118 8678
rect 6174 8676 6198 8678
rect 6254 8676 6278 8678
rect 6334 8676 6340 8678
rect 6032 8667 6340 8676
rect 6032 7644 6340 7653
rect 6032 7642 6038 7644
rect 6094 7642 6118 7644
rect 6174 7642 6198 7644
rect 6254 7642 6278 7644
rect 6334 7642 6340 7644
rect 6094 7590 6096 7642
rect 6276 7590 6278 7642
rect 6032 7588 6038 7590
rect 6094 7588 6118 7590
rect 6174 7588 6198 7590
rect 6254 7588 6278 7590
rect 6334 7588 6340 7590
rect 6032 7579 6340 7588
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6032 6556 6340 6565
rect 6032 6554 6038 6556
rect 6094 6554 6118 6556
rect 6174 6554 6198 6556
rect 6254 6554 6278 6556
rect 6334 6554 6340 6556
rect 6094 6502 6096 6554
rect 6276 6502 6278 6554
rect 6032 6500 6038 6502
rect 6094 6500 6118 6502
rect 6174 6500 6198 6502
rect 6254 6500 6278 6502
rect 6334 6500 6340 6502
rect 6032 6491 6340 6500
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5920 6118 5948 6394
rect 6380 6390 6408 6598
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5642 5948 6054
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 6032 5468 6340 5477
rect 6032 5466 6038 5468
rect 6094 5466 6118 5468
rect 6174 5466 6198 5468
rect 6254 5466 6278 5468
rect 6334 5466 6340 5468
rect 6094 5414 6096 5466
rect 6276 5414 6278 5466
rect 6032 5412 6038 5414
rect 6094 5412 6118 5414
rect 6174 5412 6198 5414
rect 6254 5412 6278 5414
rect 6334 5412 6340 5414
rect 6032 5403 6340 5412
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5920 4486 5948 5170
rect 6288 4570 6316 5306
rect 6380 5114 6408 6326
rect 6472 5370 6500 9302
rect 6550 9302 6684 9330
rect 6550 9200 6606 9302
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6564 5545 6592 7754
rect 6550 5536 6606 5545
rect 6550 5471 6606 5480
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6380 5086 6592 5114
rect 6288 4542 6500 4570
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6032 4380 6340 4389
rect 6032 4378 6038 4380
rect 6094 4378 6118 4380
rect 6174 4378 6198 4380
rect 6254 4378 6278 4380
rect 6334 4378 6340 4380
rect 6094 4326 6096 4378
rect 6276 4326 6278 4378
rect 6032 4324 6038 4326
rect 6094 4324 6118 4326
rect 6174 4324 6198 4326
rect 6254 4324 6278 4326
rect 6334 4324 6340 4326
rect 6032 4315 6340 4324
rect 5828 4270 5948 4298
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5736 3738 5764 4150
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5736 2854 5764 3470
rect 5828 3398 5856 4082
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5446 1864 5502 1873
rect 5446 1799 5502 1808
rect 5170 1660 5478 1669
rect 5170 1658 5176 1660
rect 5232 1658 5256 1660
rect 5312 1658 5336 1660
rect 5392 1658 5416 1660
rect 5472 1658 5478 1660
rect 5232 1606 5234 1658
rect 5414 1606 5416 1658
rect 5170 1604 5176 1606
rect 5232 1604 5256 1606
rect 5312 1604 5336 1606
rect 5392 1604 5416 1606
rect 5472 1604 5478 1606
rect 5170 1595 5478 1604
rect 5276 870 5396 898
rect 5276 762 5304 870
rect 5368 800 5396 870
rect 5828 800 5856 3062
rect 5920 2514 5948 4270
rect 6032 3292 6340 3301
rect 6032 3290 6038 3292
rect 6094 3290 6118 3292
rect 6174 3290 6198 3292
rect 6254 3290 6278 3292
rect 6334 3290 6340 3292
rect 6094 3238 6096 3290
rect 6276 3238 6278 3290
rect 6032 3236 6038 3238
rect 6094 3236 6118 3238
rect 6174 3236 6198 3238
rect 6254 3236 6278 3238
rect 6334 3236 6340 3238
rect 6032 3227 6340 3236
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6012 2582 6040 2790
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 6032 2204 6340 2213
rect 6032 2202 6038 2204
rect 6094 2202 6118 2204
rect 6174 2202 6198 2204
rect 6254 2202 6278 2204
rect 6334 2202 6340 2204
rect 6094 2150 6096 2202
rect 6276 2150 6278 2202
rect 6032 2148 6038 2150
rect 6094 2148 6118 2150
rect 6174 2148 6198 2150
rect 6254 2148 6278 2150
rect 6334 2148 6340 2150
rect 6032 2139 6340 2148
rect 6032 1116 6340 1125
rect 6032 1114 6038 1116
rect 6094 1114 6118 1116
rect 6174 1114 6198 1116
rect 6254 1114 6278 1116
rect 6334 1114 6340 1116
rect 6094 1062 6096 1114
rect 6276 1062 6278 1114
rect 6032 1060 6038 1062
rect 6094 1060 6118 1062
rect 6174 1060 6198 1062
rect 6254 1060 6278 1062
rect 6334 1060 6340 1062
rect 6032 1051 6340 1060
rect 6380 898 6408 4422
rect 6472 3126 6500 4542
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 6472 2650 6500 3062
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6564 2038 6592 5086
rect 6656 4554 6684 9302
rect 6748 9302 6882 9330
rect 6748 6458 6776 9302
rect 6826 9200 6882 9302
rect 7102 9330 7158 10000
rect 7378 9330 7434 10000
rect 7102 9302 7328 9330
rect 7102 9200 7158 9302
rect 6895 8188 7203 8197
rect 6895 8186 6901 8188
rect 6957 8186 6981 8188
rect 7037 8186 7061 8188
rect 7117 8186 7141 8188
rect 7197 8186 7203 8188
rect 6957 8134 6959 8186
rect 7139 8134 7141 8186
rect 6895 8132 6901 8134
rect 6957 8132 6981 8134
rect 7037 8132 7061 8134
rect 7117 8132 7141 8134
rect 7197 8132 7203 8134
rect 6895 8123 7203 8132
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7410 7144 7686
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6895 7100 7203 7109
rect 6895 7098 6901 7100
rect 6957 7098 6981 7100
rect 7037 7098 7061 7100
rect 7117 7098 7141 7100
rect 7197 7098 7203 7100
rect 6957 7046 6959 7098
rect 7139 7046 7141 7098
rect 6895 7044 6901 7046
rect 6957 7044 6981 7046
rect 7037 7044 7061 7046
rect 7117 7044 7141 7046
rect 7197 7044 7203 7046
rect 6895 7035 7203 7044
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6656 1290 6684 4218
rect 6644 1284 6696 1290
rect 6644 1226 6696 1232
rect 6288 870 6408 898
rect 6288 800 6316 870
rect 6748 800 6776 6258
rect 6895 6012 7203 6021
rect 6895 6010 6901 6012
rect 6957 6010 6981 6012
rect 7037 6010 7061 6012
rect 7117 6010 7141 6012
rect 7197 6010 7203 6012
rect 6957 5958 6959 6010
rect 7139 5958 7141 6010
rect 6895 5956 6901 5958
rect 6957 5956 6981 5958
rect 7037 5956 7061 5958
rect 7117 5956 7141 5958
rect 7197 5956 7203 5958
rect 6895 5947 7203 5956
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7208 5234 7236 5850
rect 7300 5778 7328 9302
rect 7378 9302 7604 9330
rect 7378 9200 7434 9302
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7392 7478 7420 8842
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 6895 4924 7203 4933
rect 6895 4922 6901 4924
rect 6957 4922 6981 4924
rect 7037 4922 7061 4924
rect 7117 4922 7141 4924
rect 7197 4922 7203 4924
rect 6957 4870 6959 4922
rect 7139 4870 7141 4922
rect 6895 4868 6901 4870
rect 6957 4868 6981 4870
rect 7037 4868 7061 4870
rect 7117 4868 7141 4870
rect 7197 4868 7203 4870
rect 6895 4859 7203 4868
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6840 4049 6868 4490
rect 7300 4185 7328 5578
rect 7392 4729 7420 7278
rect 7484 5137 7512 8366
rect 7576 7546 7604 9302
rect 7654 9200 7710 10000
rect 7930 9330 7986 10000
rect 8206 9330 8262 10000
rect 7930 9302 8156 9330
rect 7930 9200 7986 9302
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 6390 7604 7278
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7576 5914 7604 6122
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7470 5128 7526 5137
rect 7470 5063 7526 5072
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7378 4720 7434 4729
rect 7378 4655 7434 4664
rect 7286 4176 7342 4185
rect 7286 4111 7342 4120
rect 7288 4072 7340 4078
rect 6826 4040 6882 4049
rect 7288 4014 7340 4020
rect 6826 3975 6882 3984
rect 6895 3836 7203 3845
rect 6895 3834 6901 3836
rect 6957 3834 6981 3836
rect 7037 3834 7061 3836
rect 7117 3834 7141 3836
rect 7197 3834 7203 3836
rect 6957 3782 6959 3834
rect 7139 3782 7141 3834
rect 6895 3780 6901 3782
rect 6957 3780 6981 3782
rect 7037 3780 7061 3782
rect 7117 3780 7141 3782
rect 7197 3780 7203 3782
rect 6895 3771 7203 3780
rect 7300 3505 7328 4014
rect 7286 3496 7342 3505
rect 7286 3431 7342 3440
rect 7286 3088 7342 3097
rect 7286 3023 7288 3032
rect 7340 3023 7342 3032
rect 7288 2994 7340 3000
rect 7484 2802 7512 4966
rect 7576 2990 7604 5714
rect 7668 3602 7696 9200
rect 7757 8732 8065 8741
rect 7757 8730 7763 8732
rect 7819 8730 7843 8732
rect 7899 8730 7923 8732
rect 7979 8730 8003 8732
rect 8059 8730 8065 8732
rect 7819 8678 7821 8730
rect 8001 8678 8003 8730
rect 7757 8676 7763 8678
rect 7819 8676 7843 8678
rect 7899 8676 7923 8678
rect 7979 8676 8003 8678
rect 8059 8676 8065 8678
rect 7757 8667 8065 8676
rect 7757 7644 8065 7653
rect 7757 7642 7763 7644
rect 7819 7642 7843 7644
rect 7899 7642 7923 7644
rect 7979 7642 8003 7644
rect 8059 7642 8065 7644
rect 7819 7590 7821 7642
rect 8001 7590 8003 7642
rect 7757 7588 7763 7590
rect 7819 7588 7843 7590
rect 7899 7588 7923 7590
rect 7979 7588 8003 7590
rect 8059 7588 8065 7590
rect 7757 7579 8065 7588
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7760 6662 7788 7482
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7757 6556 8065 6565
rect 7757 6554 7763 6556
rect 7819 6554 7843 6556
rect 7899 6554 7923 6556
rect 7979 6554 8003 6556
rect 8059 6554 8065 6556
rect 7819 6502 7821 6554
rect 8001 6502 8003 6554
rect 7757 6500 7763 6502
rect 7819 6500 7843 6502
rect 7899 6500 7923 6502
rect 7979 6500 8003 6502
rect 8059 6500 8065 6502
rect 7757 6491 8065 6500
rect 7757 5468 8065 5477
rect 7757 5466 7763 5468
rect 7819 5466 7843 5468
rect 7899 5466 7923 5468
rect 7979 5466 8003 5468
rect 8059 5466 8065 5468
rect 7819 5414 7821 5466
rect 8001 5414 8003 5466
rect 7757 5412 7763 5414
rect 7819 5412 7843 5414
rect 7899 5412 7923 5414
rect 7979 5412 8003 5414
rect 8059 5412 8065 5414
rect 7757 5403 8065 5412
rect 7757 4380 8065 4389
rect 7757 4378 7763 4380
rect 7819 4378 7843 4380
rect 7899 4378 7923 4380
rect 7979 4378 8003 4380
rect 8059 4378 8065 4380
rect 7819 4326 7821 4378
rect 8001 4326 8003 4378
rect 7757 4324 7763 4326
rect 7819 4324 7843 4326
rect 7899 4324 7923 4326
rect 7979 4324 8003 4326
rect 8059 4324 8065 4326
rect 7757 4315 8065 4324
rect 8128 4282 8156 9302
rect 8206 9302 8432 9330
rect 8206 9200 8262 9302
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7757 3292 8065 3301
rect 7757 3290 7763 3292
rect 7819 3290 7843 3292
rect 7899 3290 7923 3292
rect 7979 3290 8003 3292
rect 8059 3290 8065 3292
rect 7819 3238 7821 3290
rect 8001 3238 8003 3290
rect 7757 3236 7763 3238
rect 7819 3236 7843 3238
rect 7899 3236 7923 3238
rect 7979 3236 8003 3238
rect 8059 3236 8065 3238
rect 7757 3227 8065 3236
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7484 2774 7696 2802
rect 6895 2748 7203 2757
rect 6895 2746 6901 2748
rect 6957 2746 6981 2748
rect 7037 2746 7061 2748
rect 7117 2746 7141 2748
rect 7197 2746 7203 2748
rect 6957 2694 6959 2746
rect 7139 2694 7141 2746
rect 6895 2692 6901 2694
rect 6957 2692 6981 2694
rect 7037 2692 7061 2694
rect 7117 2692 7141 2694
rect 7197 2692 7203 2694
rect 6895 2683 7203 2692
rect 7286 2680 7342 2689
rect 7286 2615 7342 2624
rect 7300 2514 7328 2615
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7286 2408 7342 2417
rect 7286 2343 7342 2352
rect 7300 2038 7328 2343
rect 7288 2032 7340 2038
rect 7288 1974 7340 1980
rect 7286 1864 7342 1873
rect 7286 1799 7342 1808
rect 6895 1660 7203 1669
rect 6895 1658 6901 1660
rect 6957 1658 6981 1660
rect 7037 1658 7061 1660
rect 7117 1658 7141 1660
rect 7197 1658 7203 1660
rect 6957 1606 6959 1658
rect 7139 1606 7141 1658
rect 6895 1604 6901 1606
rect 6957 1604 6981 1606
rect 7037 1604 7061 1606
rect 7117 1604 7141 1606
rect 7197 1604 7203 1606
rect 6895 1595 7203 1604
rect 7196 1556 7248 1562
rect 7196 1498 7248 1504
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 5092 734 5304 762
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 6840 649 6868 1294
rect 7208 800 7236 1498
rect 7300 1358 7328 1799
rect 7288 1352 7340 1358
rect 7288 1294 7340 1300
rect 7668 800 7696 2774
rect 7757 2204 8065 2213
rect 7757 2202 7763 2204
rect 7819 2202 7843 2204
rect 7899 2202 7923 2204
rect 7979 2202 8003 2204
rect 8059 2202 8065 2204
rect 7819 2150 7821 2202
rect 8001 2150 8003 2202
rect 7757 2148 7763 2150
rect 7819 2148 7843 2150
rect 7899 2148 7923 2150
rect 7979 2148 8003 2150
rect 8059 2148 8065 2150
rect 7757 2139 8065 2148
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 7757 1116 8065 1125
rect 7757 1114 7763 1116
rect 7819 1114 7843 1116
rect 7899 1114 7923 1116
rect 7979 1114 8003 1116
rect 8059 1114 8065 1116
rect 7819 1062 7821 1114
rect 8001 1062 8003 1114
rect 7757 1060 7763 1062
rect 7819 1060 7843 1062
rect 7899 1060 7923 1062
rect 7979 1060 8003 1062
rect 8059 1060 8065 1062
rect 7757 1051 8065 1060
rect 8128 800 8156 2042
rect 8220 1562 8248 6666
rect 8404 3194 8432 9302
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8208 1556 8260 1562
rect 8208 1498 8260 1504
rect 8588 800 8616 2858
rect 6826 640 6882 649
rect 6826 575 6882 584
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
<< via2 >>
rect 1582 8336 1638 8392
rect 1766 8336 1822 8392
rect 1726 8186 1782 8188
rect 1806 8186 1862 8188
rect 1886 8186 1942 8188
rect 1966 8186 2022 8188
rect 1726 8134 1772 8186
rect 1772 8134 1782 8186
rect 1806 8134 1836 8186
rect 1836 8134 1848 8186
rect 1848 8134 1862 8186
rect 1886 8134 1900 8186
rect 1900 8134 1912 8186
rect 1912 8134 1942 8186
rect 1966 8134 1976 8186
rect 1976 8134 2022 8186
rect 1726 8132 1782 8134
rect 1806 8132 1862 8134
rect 1886 8132 1942 8134
rect 1966 8132 2022 8134
rect 1726 7098 1782 7100
rect 1806 7098 1862 7100
rect 1886 7098 1942 7100
rect 1966 7098 2022 7100
rect 1726 7046 1772 7098
rect 1772 7046 1782 7098
rect 1806 7046 1836 7098
rect 1836 7046 1848 7098
rect 1848 7046 1862 7098
rect 1886 7046 1900 7098
rect 1900 7046 1912 7098
rect 1912 7046 1942 7098
rect 1966 7046 1976 7098
rect 1976 7046 2022 7098
rect 1726 7044 1782 7046
rect 1806 7044 1862 7046
rect 1886 7044 1942 7046
rect 1966 7044 2022 7046
rect 1490 6976 1546 7032
rect 1726 6010 1782 6012
rect 1806 6010 1862 6012
rect 1886 6010 1942 6012
rect 1966 6010 2022 6012
rect 1726 5958 1772 6010
rect 1772 5958 1782 6010
rect 1806 5958 1836 6010
rect 1836 5958 1848 6010
rect 1848 5958 1862 6010
rect 1886 5958 1900 6010
rect 1900 5958 1912 6010
rect 1912 5958 1942 6010
rect 1966 5958 1976 6010
rect 1976 5958 2022 6010
rect 1726 5956 1782 5958
rect 1806 5956 1862 5958
rect 1886 5956 1942 5958
rect 1966 5956 2022 5958
rect 2588 8730 2644 8732
rect 2668 8730 2724 8732
rect 2748 8730 2804 8732
rect 2828 8730 2884 8732
rect 2588 8678 2634 8730
rect 2634 8678 2644 8730
rect 2668 8678 2698 8730
rect 2698 8678 2710 8730
rect 2710 8678 2724 8730
rect 2748 8678 2762 8730
rect 2762 8678 2774 8730
rect 2774 8678 2804 8730
rect 2828 8678 2838 8730
rect 2838 8678 2884 8730
rect 2588 8676 2644 8678
rect 2668 8676 2724 8678
rect 2748 8676 2804 8678
rect 2828 8676 2884 8678
rect 2588 7642 2644 7644
rect 2668 7642 2724 7644
rect 2748 7642 2804 7644
rect 2828 7642 2884 7644
rect 2588 7590 2634 7642
rect 2634 7590 2644 7642
rect 2668 7590 2698 7642
rect 2698 7590 2710 7642
rect 2710 7590 2724 7642
rect 2748 7590 2762 7642
rect 2762 7590 2774 7642
rect 2774 7590 2804 7642
rect 2828 7590 2838 7642
rect 2838 7590 2884 7642
rect 2588 7588 2644 7590
rect 2668 7588 2724 7590
rect 2748 7588 2804 7590
rect 2828 7588 2884 7590
rect 2588 6554 2644 6556
rect 2668 6554 2724 6556
rect 2748 6554 2804 6556
rect 2828 6554 2884 6556
rect 2588 6502 2634 6554
rect 2634 6502 2644 6554
rect 2668 6502 2698 6554
rect 2698 6502 2710 6554
rect 2710 6502 2724 6554
rect 2748 6502 2762 6554
rect 2762 6502 2774 6554
rect 2774 6502 2804 6554
rect 2828 6502 2838 6554
rect 2838 6502 2884 6554
rect 2588 6500 2644 6502
rect 2668 6500 2724 6502
rect 2748 6500 2804 6502
rect 2828 6500 2884 6502
rect 2962 6296 3018 6352
rect 1726 4922 1782 4924
rect 1806 4922 1862 4924
rect 1886 4922 1942 4924
rect 1966 4922 2022 4924
rect 1726 4870 1772 4922
rect 1772 4870 1782 4922
rect 1806 4870 1836 4922
rect 1836 4870 1848 4922
rect 1848 4870 1862 4922
rect 1886 4870 1900 4922
rect 1900 4870 1912 4922
rect 1912 4870 1942 4922
rect 1966 4870 1976 4922
rect 1976 4870 2022 4922
rect 1726 4868 1782 4870
rect 1806 4868 1862 4870
rect 1886 4868 1942 4870
rect 1966 4868 2022 4870
rect 1490 1536 1546 1592
rect 1726 3834 1782 3836
rect 1806 3834 1862 3836
rect 1886 3834 1942 3836
rect 1966 3834 2022 3836
rect 1726 3782 1772 3834
rect 1772 3782 1782 3834
rect 1806 3782 1836 3834
rect 1836 3782 1848 3834
rect 1848 3782 1862 3834
rect 1886 3782 1900 3834
rect 1900 3782 1912 3834
rect 1912 3782 1942 3834
rect 1966 3782 1976 3834
rect 1976 3782 2022 3834
rect 1726 3780 1782 3782
rect 1806 3780 1862 3782
rect 1886 3780 1942 3782
rect 1966 3780 2022 3782
rect 1726 2746 1782 2748
rect 1806 2746 1862 2748
rect 1886 2746 1942 2748
rect 1966 2746 2022 2748
rect 1726 2694 1772 2746
rect 1772 2694 1782 2746
rect 1806 2694 1836 2746
rect 1836 2694 1848 2746
rect 1848 2694 1862 2746
rect 1886 2694 1900 2746
rect 1900 2694 1912 2746
rect 1912 2694 1942 2746
rect 1966 2694 1976 2746
rect 1976 2694 2022 2746
rect 1726 2692 1782 2694
rect 1806 2692 1862 2694
rect 1886 2692 1942 2694
rect 1966 2692 2022 2694
rect 1726 1658 1782 1660
rect 1806 1658 1862 1660
rect 1886 1658 1942 1660
rect 1966 1658 2022 1660
rect 1726 1606 1772 1658
rect 1772 1606 1782 1658
rect 1806 1606 1836 1658
rect 1836 1606 1848 1658
rect 1848 1606 1862 1658
rect 1886 1606 1900 1658
rect 1900 1606 1912 1658
rect 1912 1606 1942 1658
rect 1966 1606 1976 1658
rect 1976 1606 2022 1658
rect 1726 1604 1782 1606
rect 1806 1604 1862 1606
rect 1886 1604 1942 1606
rect 1966 1604 2022 1606
rect 2588 5466 2644 5468
rect 2668 5466 2724 5468
rect 2748 5466 2804 5468
rect 2828 5466 2884 5468
rect 2588 5414 2634 5466
rect 2634 5414 2644 5466
rect 2668 5414 2698 5466
rect 2698 5414 2710 5466
rect 2710 5414 2724 5466
rect 2748 5414 2762 5466
rect 2762 5414 2774 5466
rect 2774 5414 2804 5466
rect 2828 5414 2838 5466
rect 2838 5414 2884 5466
rect 2588 5412 2644 5414
rect 2668 5412 2724 5414
rect 2748 5412 2804 5414
rect 2828 5412 2884 5414
rect 2588 4378 2644 4380
rect 2668 4378 2724 4380
rect 2748 4378 2804 4380
rect 2828 4378 2884 4380
rect 2588 4326 2634 4378
rect 2634 4326 2644 4378
rect 2668 4326 2698 4378
rect 2698 4326 2710 4378
rect 2710 4326 2724 4378
rect 2748 4326 2762 4378
rect 2762 4326 2774 4378
rect 2774 4326 2804 4378
rect 2828 4326 2838 4378
rect 2838 4326 2884 4378
rect 2588 4324 2644 4326
rect 2668 4324 2724 4326
rect 2748 4324 2804 4326
rect 2828 4324 2884 4326
rect 3054 5616 3110 5672
rect 2962 3576 3018 3632
rect 2588 3290 2644 3292
rect 2668 3290 2724 3292
rect 2748 3290 2804 3292
rect 2828 3290 2884 3292
rect 2588 3238 2634 3290
rect 2634 3238 2644 3290
rect 2668 3238 2698 3290
rect 2698 3238 2710 3290
rect 2710 3238 2724 3290
rect 2748 3238 2762 3290
rect 2762 3238 2774 3290
rect 2774 3238 2804 3290
rect 2828 3238 2838 3290
rect 2838 3238 2884 3290
rect 2588 3236 2644 3238
rect 2668 3236 2724 3238
rect 2748 3236 2804 3238
rect 2828 3236 2884 3238
rect 2778 2896 2834 2952
rect 2588 2202 2644 2204
rect 2668 2202 2724 2204
rect 2748 2202 2804 2204
rect 2828 2202 2884 2204
rect 2588 2150 2634 2202
rect 2634 2150 2644 2202
rect 2668 2150 2698 2202
rect 2698 2150 2710 2202
rect 2710 2150 2724 2202
rect 2748 2150 2762 2202
rect 2762 2150 2774 2202
rect 2774 2150 2804 2202
rect 2828 2150 2838 2202
rect 2838 2150 2884 2202
rect 2588 2148 2644 2150
rect 2668 2148 2724 2150
rect 2748 2148 2804 2150
rect 2828 2148 2884 2150
rect 2778 1944 2834 2000
rect 2588 1114 2644 1116
rect 2668 1114 2724 1116
rect 2748 1114 2804 1116
rect 2828 1114 2884 1116
rect 2588 1062 2634 1114
rect 2634 1062 2644 1114
rect 2668 1062 2698 1114
rect 2698 1062 2710 1114
rect 2710 1062 2724 1114
rect 2748 1062 2762 1114
rect 2762 1062 2774 1114
rect 2774 1062 2804 1114
rect 2828 1062 2838 1114
rect 2838 1062 2884 1114
rect 2588 1060 2644 1062
rect 2668 1060 2724 1062
rect 2748 1060 2804 1062
rect 2828 1060 2884 1062
rect 2962 856 3018 912
rect 3422 9016 3478 9072
rect 3451 8186 3507 8188
rect 3531 8186 3587 8188
rect 3611 8186 3667 8188
rect 3691 8186 3747 8188
rect 3451 8134 3497 8186
rect 3497 8134 3507 8186
rect 3531 8134 3561 8186
rect 3561 8134 3573 8186
rect 3573 8134 3587 8186
rect 3611 8134 3625 8186
rect 3625 8134 3637 8186
rect 3637 8134 3667 8186
rect 3691 8134 3701 8186
rect 3701 8134 3747 8186
rect 3451 8132 3507 8134
rect 3531 8132 3587 8134
rect 3611 8132 3667 8134
rect 3691 8132 3747 8134
rect 3330 7384 3386 7440
rect 3451 7098 3507 7100
rect 3531 7098 3587 7100
rect 3611 7098 3667 7100
rect 3691 7098 3747 7100
rect 3451 7046 3497 7098
rect 3497 7046 3507 7098
rect 3531 7046 3561 7098
rect 3561 7046 3573 7098
rect 3573 7046 3587 7098
rect 3611 7046 3625 7098
rect 3625 7046 3637 7098
rect 3637 7046 3667 7098
rect 3691 7046 3701 7098
rect 3701 7046 3747 7098
rect 3451 7044 3507 7046
rect 3531 7044 3587 7046
rect 3611 7044 3667 7046
rect 3691 7044 3747 7046
rect 3451 6010 3507 6012
rect 3531 6010 3587 6012
rect 3611 6010 3667 6012
rect 3691 6010 3747 6012
rect 3451 5958 3497 6010
rect 3497 5958 3507 6010
rect 3531 5958 3561 6010
rect 3561 5958 3573 6010
rect 3573 5958 3587 6010
rect 3611 5958 3625 6010
rect 3625 5958 3637 6010
rect 3637 5958 3667 6010
rect 3691 5958 3701 6010
rect 3701 5958 3747 6010
rect 3451 5956 3507 5958
rect 3531 5956 3587 5958
rect 3611 5956 3667 5958
rect 3691 5956 3747 5958
rect 3451 4922 3507 4924
rect 3531 4922 3587 4924
rect 3611 4922 3667 4924
rect 3691 4922 3747 4924
rect 3451 4870 3497 4922
rect 3497 4870 3507 4922
rect 3531 4870 3561 4922
rect 3561 4870 3573 4922
rect 3573 4870 3587 4922
rect 3611 4870 3625 4922
rect 3625 4870 3637 4922
rect 3637 4870 3667 4922
rect 3691 4870 3701 4922
rect 3701 4870 3747 4922
rect 3451 4868 3507 4870
rect 3531 4868 3587 4870
rect 3611 4868 3667 4870
rect 3691 4868 3747 4870
rect 3882 8880 3938 8936
rect 3882 4664 3938 4720
rect 3451 3834 3507 3836
rect 3531 3834 3587 3836
rect 3611 3834 3667 3836
rect 3691 3834 3747 3836
rect 3451 3782 3497 3834
rect 3497 3782 3507 3834
rect 3531 3782 3561 3834
rect 3561 3782 3573 3834
rect 3573 3782 3587 3834
rect 3611 3782 3625 3834
rect 3625 3782 3637 3834
rect 3637 3782 3667 3834
rect 3691 3782 3701 3834
rect 3701 3782 3747 3834
rect 3451 3780 3507 3782
rect 3531 3780 3587 3782
rect 3611 3780 3667 3782
rect 3691 3780 3747 3782
rect 3451 2746 3507 2748
rect 3531 2746 3587 2748
rect 3611 2746 3667 2748
rect 3691 2746 3747 2748
rect 3451 2694 3497 2746
rect 3497 2694 3507 2746
rect 3531 2694 3561 2746
rect 3561 2694 3573 2746
rect 3573 2694 3587 2746
rect 3611 2694 3625 2746
rect 3625 2694 3637 2746
rect 3637 2694 3667 2746
rect 3691 2694 3701 2746
rect 3701 2694 3747 2746
rect 3451 2692 3507 2694
rect 3531 2692 3587 2694
rect 3611 2692 3667 2694
rect 3691 2692 3747 2694
rect 3451 1658 3507 1660
rect 3531 1658 3587 1660
rect 3611 1658 3667 1660
rect 3691 1658 3747 1660
rect 3451 1606 3497 1658
rect 3497 1606 3507 1658
rect 3531 1606 3561 1658
rect 3561 1606 3573 1658
rect 3573 1606 3587 1658
rect 3611 1606 3625 1658
rect 3625 1606 3637 1658
rect 3637 1606 3667 1658
rect 3691 1606 3701 1658
rect 3701 1606 3747 1658
rect 3451 1604 3507 1606
rect 3531 1604 3587 1606
rect 3611 1604 3667 1606
rect 3691 1604 3747 1606
rect 4066 4120 4122 4176
rect 4313 8730 4369 8732
rect 4393 8730 4449 8732
rect 4473 8730 4529 8732
rect 4553 8730 4609 8732
rect 4313 8678 4359 8730
rect 4359 8678 4369 8730
rect 4393 8678 4423 8730
rect 4423 8678 4435 8730
rect 4435 8678 4449 8730
rect 4473 8678 4487 8730
rect 4487 8678 4499 8730
rect 4499 8678 4529 8730
rect 4553 8678 4563 8730
rect 4563 8678 4609 8730
rect 4313 8676 4369 8678
rect 4393 8676 4449 8678
rect 4473 8676 4529 8678
rect 4553 8676 4609 8678
rect 4710 7928 4766 7984
rect 4618 7792 4674 7848
rect 4313 7642 4369 7644
rect 4393 7642 4449 7644
rect 4473 7642 4529 7644
rect 4553 7642 4609 7644
rect 4313 7590 4359 7642
rect 4359 7590 4369 7642
rect 4393 7590 4423 7642
rect 4423 7590 4435 7642
rect 4435 7590 4449 7642
rect 4473 7590 4487 7642
rect 4487 7590 4499 7642
rect 4499 7590 4529 7642
rect 4553 7590 4563 7642
rect 4563 7590 4609 7642
rect 4313 7588 4369 7590
rect 4393 7588 4449 7590
rect 4473 7588 4529 7590
rect 4553 7588 4609 7590
rect 4526 6740 4528 6760
rect 4528 6740 4580 6760
rect 4580 6740 4582 6760
rect 4526 6704 4582 6740
rect 4313 6554 4369 6556
rect 4393 6554 4449 6556
rect 4473 6554 4529 6556
rect 4553 6554 4609 6556
rect 4313 6502 4359 6554
rect 4359 6502 4369 6554
rect 4393 6502 4423 6554
rect 4423 6502 4435 6554
rect 4435 6502 4449 6554
rect 4473 6502 4487 6554
rect 4487 6502 4499 6554
rect 4499 6502 4529 6554
rect 4553 6502 4563 6554
rect 4563 6502 4609 6554
rect 4313 6500 4369 6502
rect 4393 6500 4449 6502
rect 4473 6500 4529 6502
rect 4553 6500 4609 6502
rect 4313 5466 4369 5468
rect 4393 5466 4449 5468
rect 4473 5466 4529 5468
rect 4553 5466 4609 5468
rect 4313 5414 4359 5466
rect 4359 5414 4369 5466
rect 4393 5414 4423 5466
rect 4423 5414 4435 5466
rect 4435 5414 4449 5466
rect 4473 5414 4487 5466
rect 4487 5414 4499 5466
rect 4499 5414 4529 5466
rect 4553 5414 4563 5466
rect 4563 5414 4609 5466
rect 4313 5412 4369 5414
rect 4393 5412 4449 5414
rect 4473 5412 4529 5414
rect 4553 5412 4609 5414
rect 4802 6160 4858 6216
rect 4313 4378 4369 4380
rect 4393 4378 4449 4380
rect 4473 4378 4529 4380
rect 4553 4378 4609 4380
rect 4313 4326 4359 4378
rect 4359 4326 4369 4378
rect 4393 4326 4423 4378
rect 4423 4326 4435 4378
rect 4435 4326 4449 4378
rect 4473 4326 4487 4378
rect 4487 4326 4499 4378
rect 4499 4326 4529 4378
rect 4553 4326 4563 4378
rect 4563 4326 4609 4378
rect 4313 4324 4369 4326
rect 4393 4324 4449 4326
rect 4473 4324 4529 4326
rect 4553 4324 4609 4326
rect 4313 3290 4369 3292
rect 4393 3290 4449 3292
rect 4473 3290 4529 3292
rect 4553 3290 4609 3292
rect 4313 3238 4359 3290
rect 4359 3238 4369 3290
rect 4393 3238 4423 3290
rect 4423 3238 4435 3290
rect 4435 3238 4449 3290
rect 4473 3238 4487 3290
rect 4487 3238 4499 3290
rect 4499 3238 4529 3290
rect 4553 3238 4563 3290
rect 4563 3238 4609 3290
rect 4313 3236 4369 3238
rect 4393 3236 4449 3238
rect 4473 3236 4529 3238
rect 4553 3236 4609 3238
rect 4313 2202 4369 2204
rect 4393 2202 4449 2204
rect 4473 2202 4529 2204
rect 4553 2202 4609 2204
rect 4313 2150 4359 2202
rect 4359 2150 4369 2202
rect 4393 2150 4423 2202
rect 4423 2150 4435 2202
rect 4435 2150 4449 2202
rect 4473 2150 4487 2202
rect 4487 2150 4499 2202
rect 4499 2150 4529 2202
rect 4553 2150 4563 2202
rect 4563 2150 4609 2202
rect 4313 2148 4369 2150
rect 4393 2148 4449 2150
rect 4473 2148 4529 2150
rect 4553 2148 4609 2150
rect 4313 1114 4369 1116
rect 4393 1114 4449 1116
rect 4473 1114 4529 1116
rect 4553 1114 4609 1116
rect 4313 1062 4359 1114
rect 4359 1062 4369 1114
rect 4393 1062 4423 1114
rect 4423 1062 4435 1114
rect 4435 1062 4449 1114
rect 4473 1062 4487 1114
rect 4487 1062 4499 1114
rect 4499 1062 4529 1114
rect 4553 1062 4563 1114
rect 4563 1062 4609 1114
rect 4313 1060 4369 1062
rect 4393 1060 4449 1062
rect 4473 1060 4529 1062
rect 4553 1060 4609 1062
rect 5176 8186 5232 8188
rect 5256 8186 5312 8188
rect 5336 8186 5392 8188
rect 5416 8186 5472 8188
rect 5176 8134 5222 8186
rect 5222 8134 5232 8186
rect 5256 8134 5286 8186
rect 5286 8134 5298 8186
rect 5298 8134 5312 8186
rect 5336 8134 5350 8186
rect 5350 8134 5362 8186
rect 5362 8134 5392 8186
rect 5416 8134 5426 8186
rect 5426 8134 5472 8186
rect 5176 8132 5232 8134
rect 5256 8132 5312 8134
rect 5336 8132 5392 8134
rect 5416 8132 5472 8134
rect 5630 8336 5686 8392
rect 5446 7248 5502 7304
rect 5176 7098 5232 7100
rect 5256 7098 5312 7100
rect 5336 7098 5392 7100
rect 5416 7098 5472 7100
rect 5176 7046 5222 7098
rect 5222 7046 5232 7098
rect 5256 7046 5286 7098
rect 5286 7046 5298 7098
rect 5298 7046 5312 7098
rect 5336 7046 5350 7098
rect 5350 7046 5362 7098
rect 5362 7046 5392 7098
rect 5416 7046 5426 7098
rect 5426 7046 5472 7098
rect 5176 7044 5232 7046
rect 5256 7044 5312 7046
rect 5336 7044 5392 7046
rect 5416 7044 5472 7046
rect 5446 6296 5502 6352
rect 5176 6010 5232 6012
rect 5256 6010 5312 6012
rect 5336 6010 5392 6012
rect 5416 6010 5472 6012
rect 5176 5958 5222 6010
rect 5222 5958 5232 6010
rect 5256 5958 5286 6010
rect 5286 5958 5298 6010
rect 5298 5958 5312 6010
rect 5336 5958 5350 6010
rect 5350 5958 5362 6010
rect 5362 5958 5392 6010
rect 5416 5958 5426 6010
rect 5426 5958 5472 6010
rect 5176 5956 5232 5958
rect 5256 5956 5312 5958
rect 5336 5956 5392 5958
rect 5416 5956 5472 5958
rect 5176 4922 5232 4924
rect 5256 4922 5312 4924
rect 5336 4922 5392 4924
rect 5416 4922 5472 4924
rect 5176 4870 5222 4922
rect 5222 4870 5232 4922
rect 5256 4870 5286 4922
rect 5286 4870 5298 4922
rect 5298 4870 5312 4922
rect 5336 4870 5350 4922
rect 5350 4870 5362 4922
rect 5362 4870 5392 4922
rect 5416 4870 5426 4922
rect 5426 4870 5472 4922
rect 5176 4868 5232 4870
rect 5256 4868 5312 4870
rect 5336 4868 5392 4870
rect 5416 4868 5472 4870
rect 5176 3834 5232 3836
rect 5256 3834 5312 3836
rect 5336 3834 5392 3836
rect 5416 3834 5472 3836
rect 5176 3782 5222 3834
rect 5222 3782 5232 3834
rect 5256 3782 5286 3834
rect 5286 3782 5298 3834
rect 5298 3782 5312 3834
rect 5336 3782 5350 3834
rect 5350 3782 5362 3834
rect 5362 3782 5392 3834
rect 5416 3782 5426 3834
rect 5426 3782 5472 3834
rect 5176 3780 5232 3782
rect 5256 3780 5312 3782
rect 5336 3780 5392 3782
rect 5416 3780 5472 3782
rect 4986 856 5042 912
rect 5176 2746 5232 2748
rect 5256 2746 5312 2748
rect 5336 2746 5392 2748
rect 5416 2746 5472 2748
rect 5176 2694 5222 2746
rect 5222 2694 5232 2746
rect 5256 2694 5286 2746
rect 5286 2694 5298 2746
rect 5298 2694 5312 2746
rect 5336 2694 5350 2746
rect 5350 2694 5362 2746
rect 5362 2694 5392 2746
rect 5416 2694 5426 2746
rect 5426 2694 5472 2746
rect 5176 2692 5232 2694
rect 5256 2692 5312 2694
rect 5336 2692 5392 2694
rect 5416 2692 5472 2694
rect 5906 9152 5962 9208
rect 6038 8730 6094 8732
rect 6118 8730 6174 8732
rect 6198 8730 6254 8732
rect 6278 8730 6334 8732
rect 6038 8678 6084 8730
rect 6084 8678 6094 8730
rect 6118 8678 6148 8730
rect 6148 8678 6160 8730
rect 6160 8678 6174 8730
rect 6198 8678 6212 8730
rect 6212 8678 6224 8730
rect 6224 8678 6254 8730
rect 6278 8678 6288 8730
rect 6288 8678 6334 8730
rect 6038 8676 6094 8678
rect 6118 8676 6174 8678
rect 6198 8676 6254 8678
rect 6278 8676 6334 8678
rect 6038 7642 6094 7644
rect 6118 7642 6174 7644
rect 6198 7642 6254 7644
rect 6278 7642 6334 7644
rect 6038 7590 6084 7642
rect 6084 7590 6094 7642
rect 6118 7590 6148 7642
rect 6148 7590 6160 7642
rect 6160 7590 6174 7642
rect 6198 7590 6212 7642
rect 6212 7590 6224 7642
rect 6224 7590 6254 7642
rect 6278 7590 6288 7642
rect 6288 7590 6334 7642
rect 6038 7588 6094 7590
rect 6118 7588 6174 7590
rect 6198 7588 6254 7590
rect 6278 7588 6334 7590
rect 6038 6554 6094 6556
rect 6118 6554 6174 6556
rect 6198 6554 6254 6556
rect 6278 6554 6334 6556
rect 6038 6502 6084 6554
rect 6084 6502 6094 6554
rect 6118 6502 6148 6554
rect 6148 6502 6160 6554
rect 6160 6502 6174 6554
rect 6198 6502 6212 6554
rect 6212 6502 6224 6554
rect 6224 6502 6254 6554
rect 6278 6502 6288 6554
rect 6288 6502 6334 6554
rect 6038 6500 6094 6502
rect 6118 6500 6174 6502
rect 6198 6500 6254 6502
rect 6278 6500 6334 6502
rect 6038 5466 6094 5468
rect 6118 5466 6174 5468
rect 6198 5466 6254 5468
rect 6278 5466 6334 5468
rect 6038 5414 6084 5466
rect 6084 5414 6094 5466
rect 6118 5414 6148 5466
rect 6148 5414 6160 5466
rect 6160 5414 6174 5466
rect 6198 5414 6212 5466
rect 6212 5414 6224 5466
rect 6224 5414 6254 5466
rect 6278 5414 6288 5466
rect 6288 5414 6334 5466
rect 6038 5412 6094 5414
rect 6118 5412 6174 5414
rect 6198 5412 6254 5414
rect 6278 5412 6334 5414
rect 6550 5480 6606 5536
rect 6038 4378 6094 4380
rect 6118 4378 6174 4380
rect 6198 4378 6254 4380
rect 6278 4378 6334 4380
rect 6038 4326 6084 4378
rect 6084 4326 6094 4378
rect 6118 4326 6148 4378
rect 6148 4326 6160 4378
rect 6160 4326 6174 4378
rect 6198 4326 6212 4378
rect 6212 4326 6224 4378
rect 6224 4326 6254 4378
rect 6278 4326 6288 4378
rect 6288 4326 6334 4378
rect 6038 4324 6094 4326
rect 6118 4324 6174 4326
rect 6198 4324 6254 4326
rect 6278 4324 6334 4326
rect 5446 1808 5502 1864
rect 5176 1658 5232 1660
rect 5256 1658 5312 1660
rect 5336 1658 5392 1660
rect 5416 1658 5472 1660
rect 5176 1606 5222 1658
rect 5222 1606 5232 1658
rect 5256 1606 5286 1658
rect 5286 1606 5298 1658
rect 5298 1606 5312 1658
rect 5336 1606 5350 1658
rect 5350 1606 5362 1658
rect 5362 1606 5392 1658
rect 5416 1606 5426 1658
rect 5426 1606 5472 1658
rect 5176 1604 5232 1606
rect 5256 1604 5312 1606
rect 5336 1604 5392 1606
rect 5416 1604 5472 1606
rect 6038 3290 6094 3292
rect 6118 3290 6174 3292
rect 6198 3290 6254 3292
rect 6278 3290 6334 3292
rect 6038 3238 6084 3290
rect 6084 3238 6094 3290
rect 6118 3238 6148 3290
rect 6148 3238 6160 3290
rect 6160 3238 6174 3290
rect 6198 3238 6212 3290
rect 6212 3238 6224 3290
rect 6224 3238 6254 3290
rect 6278 3238 6288 3290
rect 6288 3238 6334 3290
rect 6038 3236 6094 3238
rect 6118 3236 6174 3238
rect 6198 3236 6254 3238
rect 6278 3236 6334 3238
rect 6038 2202 6094 2204
rect 6118 2202 6174 2204
rect 6198 2202 6254 2204
rect 6278 2202 6334 2204
rect 6038 2150 6084 2202
rect 6084 2150 6094 2202
rect 6118 2150 6148 2202
rect 6148 2150 6160 2202
rect 6160 2150 6174 2202
rect 6198 2150 6212 2202
rect 6212 2150 6224 2202
rect 6224 2150 6254 2202
rect 6278 2150 6288 2202
rect 6288 2150 6334 2202
rect 6038 2148 6094 2150
rect 6118 2148 6174 2150
rect 6198 2148 6254 2150
rect 6278 2148 6334 2150
rect 6038 1114 6094 1116
rect 6118 1114 6174 1116
rect 6198 1114 6254 1116
rect 6278 1114 6334 1116
rect 6038 1062 6084 1114
rect 6084 1062 6094 1114
rect 6118 1062 6148 1114
rect 6148 1062 6160 1114
rect 6160 1062 6174 1114
rect 6198 1062 6212 1114
rect 6212 1062 6224 1114
rect 6224 1062 6254 1114
rect 6278 1062 6288 1114
rect 6288 1062 6334 1114
rect 6038 1060 6094 1062
rect 6118 1060 6174 1062
rect 6198 1060 6254 1062
rect 6278 1060 6334 1062
rect 6901 8186 6957 8188
rect 6981 8186 7037 8188
rect 7061 8186 7117 8188
rect 7141 8186 7197 8188
rect 6901 8134 6947 8186
rect 6947 8134 6957 8186
rect 6981 8134 7011 8186
rect 7011 8134 7023 8186
rect 7023 8134 7037 8186
rect 7061 8134 7075 8186
rect 7075 8134 7087 8186
rect 7087 8134 7117 8186
rect 7141 8134 7151 8186
rect 7151 8134 7197 8186
rect 6901 8132 6957 8134
rect 6981 8132 7037 8134
rect 7061 8132 7117 8134
rect 7141 8132 7197 8134
rect 6901 7098 6957 7100
rect 6981 7098 7037 7100
rect 7061 7098 7117 7100
rect 7141 7098 7197 7100
rect 6901 7046 6947 7098
rect 6947 7046 6957 7098
rect 6981 7046 7011 7098
rect 7011 7046 7023 7098
rect 7023 7046 7037 7098
rect 7061 7046 7075 7098
rect 7075 7046 7087 7098
rect 7087 7046 7117 7098
rect 7141 7046 7151 7098
rect 7151 7046 7197 7098
rect 6901 7044 6957 7046
rect 6981 7044 7037 7046
rect 7061 7044 7117 7046
rect 7141 7044 7197 7046
rect 6901 6010 6957 6012
rect 6981 6010 7037 6012
rect 7061 6010 7117 6012
rect 7141 6010 7197 6012
rect 6901 5958 6947 6010
rect 6947 5958 6957 6010
rect 6981 5958 7011 6010
rect 7011 5958 7023 6010
rect 7023 5958 7037 6010
rect 7061 5958 7075 6010
rect 7075 5958 7087 6010
rect 7087 5958 7117 6010
rect 7141 5958 7151 6010
rect 7151 5958 7197 6010
rect 6901 5956 6957 5958
rect 6981 5956 7037 5958
rect 7061 5956 7117 5958
rect 7141 5956 7197 5958
rect 6901 4922 6957 4924
rect 6981 4922 7037 4924
rect 7061 4922 7117 4924
rect 7141 4922 7197 4924
rect 6901 4870 6947 4922
rect 6947 4870 6957 4922
rect 6981 4870 7011 4922
rect 7011 4870 7023 4922
rect 7023 4870 7037 4922
rect 7061 4870 7075 4922
rect 7075 4870 7087 4922
rect 7087 4870 7117 4922
rect 7141 4870 7151 4922
rect 7151 4870 7197 4922
rect 6901 4868 6957 4870
rect 6981 4868 7037 4870
rect 7061 4868 7117 4870
rect 7141 4868 7197 4870
rect 7470 5072 7526 5128
rect 7378 4664 7434 4720
rect 7286 4120 7342 4176
rect 6826 3984 6882 4040
rect 6901 3834 6957 3836
rect 6981 3834 7037 3836
rect 7061 3834 7117 3836
rect 7141 3834 7197 3836
rect 6901 3782 6947 3834
rect 6947 3782 6957 3834
rect 6981 3782 7011 3834
rect 7011 3782 7023 3834
rect 7023 3782 7037 3834
rect 7061 3782 7075 3834
rect 7075 3782 7087 3834
rect 7087 3782 7117 3834
rect 7141 3782 7151 3834
rect 7151 3782 7197 3834
rect 6901 3780 6957 3782
rect 6981 3780 7037 3782
rect 7061 3780 7117 3782
rect 7141 3780 7197 3782
rect 7286 3440 7342 3496
rect 7286 3052 7342 3088
rect 7286 3032 7288 3052
rect 7288 3032 7340 3052
rect 7340 3032 7342 3052
rect 7763 8730 7819 8732
rect 7843 8730 7899 8732
rect 7923 8730 7979 8732
rect 8003 8730 8059 8732
rect 7763 8678 7809 8730
rect 7809 8678 7819 8730
rect 7843 8678 7873 8730
rect 7873 8678 7885 8730
rect 7885 8678 7899 8730
rect 7923 8678 7937 8730
rect 7937 8678 7949 8730
rect 7949 8678 7979 8730
rect 8003 8678 8013 8730
rect 8013 8678 8059 8730
rect 7763 8676 7819 8678
rect 7843 8676 7899 8678
rect 7923 8676 7979 8678
rect 8003 8676 8059 8678
rect 7763 7642 7819 7644
rect 7843 7642 7899 7644
rect 7923 7642 7979 7644
rect 8003 7642 8059 7644
rect 7763 7590 7809 7642
rect 7809 7590 7819 7642
rect 7843 7590 7873 7642
rect 7873 7590 7885 7642
rect 7885 7590 7899 7642
rect 7923 7590 7937 7642
rect 7937 7590 7949 7642
rect 7949 7590 7979 7642
rect 8003 7590 8013 7642
rect 8013 7590 8059 7642
rect 7763 7588 7819 7590
rect 7843 7588 7899 7590
rect 7923 7588 7979 7590
rect 8003 7588 8059 7590
rect 7763 6554 7819 6556
rect 7843 6554 7899 6556
rect 7923 6554 7979 6556
rect 8003 6554 8059 6556
rect 7763 6502 7809 6554
rect 7809 6502 7819 6554
rect 7843 6502 7873 6554
rect 7873 6502 7885 6554
rect 7885 6502 7899 6554
rect 7923 6502 7937 6554
rect 7937 6502 7949 6554
rect 7949 6502 7979 6554
rect 8003 6502 8013 6554
rect 8013 6502 8059 6554
rect 7763 6500 7819 6502
rect 7843 6500 7899 6502
rect 7923 6500 7979 6502
rect 8003 6500 8059 6502
rect 7763 5466 7819 5468
rect 7843 5466 7899 5468
rect 7923 5466 7979 5468
rect 8003 5466 8059 5468
rect 7763 5414 7809 5466
rect 7809 5414 7819 5466
rect 7843 5414 7873 5466
rect 7873 5414 7885 5466
rect 7885 5414 7899 5466
rect 7923 5414 7937 5466
rect 7937 5414 7949 5466
rect 7949 5414 7979 5466
rect 8003 5414 8013 5466
rect 8013 5414 8059 5466
rect 7763 5412 7819 5414
rect 7843 5412 7899 5414
rect 7923 5412 7979 5414
rect 8003 5412 8059 5414
rect 7763 4378 7819 4380
rect 7843 4378 7899 4380
rect 7923 4378 7979 4380
rect 8003 4378 8059 4380
rect 7763 4326 7809 4378
rect 7809 4326 7819 4378
rect 7843 4326 7873 4378
rect 7873 4326 7885 4378
rect 7885 4326 7899 4378
rect 7923 4326 7937 4378
rect 7937 4326 7949 4378
rect 7949 4326 7979 4378
rect 8003 4326 8013 4378
rect 8013 4326 8059 4378
rect 7763 4324 7819 4326
rect 7843 4324 7899 4326
rect 7923 4324 7979 4326
rect 8003 4324 8059 4326
rect 7763 3290 7819 3292
rect 7843 3290 7899 3292
rect 7923 3290 7979 3292
rect 8003 3290 8059 3292
rect 7763 3238 7809 3290
rect 7809 3238 7819 3290
rect 7843 3238 7873 3290
rect 7873 3238 7885 3290
rect 7885 3238 7899 3290
rect 7923 3238 7937 3290
rect 7937 3238 7949 3290
rect 7949 3238 7979 3290
rect 8003 3238 8013 3290
rect 8013 3238 8059 3290
rect 7763 3236 7819 3238
rect 7843 3236 7899 3238
rect 7923 3236 7979 3238
rect 8003 3236 8059 3238
rect 6901 2746 6957 2748
rect 6981 2746 7037 2748
rect 7061 2746 7117 2748
rect 7141 2746 7197 2748
rect 6901 2694 6947 2746
rect 6947 2694 6957 2746
rect 6981 2694 7011 2746
rect 7011 2694 7023 2746
rect 7023 2694 7037 2746
rect 7061 2694 7075 2746
rect 7075 2694 7087 2746
rect 7087 2694 7117 2746
rect 7141 2694 7151 2746
rect 7151 2694 7197 2746
rect 6901 2692 6957 2694
rect 6981 2692 7037 2694
rect 7061 2692 7117 2694
rect 7141 2692 7197 2694
rect 7286 2624 7342 2680
rect 7286 2352 7342 2408
rect 7286 1808 7342 1864
rect 6901 1658 6957 1660
rect 6981 1658 7037 1660
rect 7061 1658 7117 1660
rect 7141 1658 7197 1660
rect 6901 1606 6947 1658
rect 6947 1606 6957 1658
rect 6981 1606 7011 1658
rect 7011 1606 7023 1658
rect 7023 1606 7037 1658
rect 7061 1606 7075 1658
rect 7075 1606 7087 1658
rect 7087 1606 7117 1658
rect 7141 1606 7151 1658
rect 7151 1606 7197 1658
rect 6901 1604 6957 1606
rect 6981 1604 7037 1606
rect 7061 1604 7117 1606
rect 7141 1604 7197 1606
rect 7763 2202 7819 2204
rect 7843 2202 7899 2204
rect 7923 2202 7979 2204
rect 8003 2202 8059 2204
rect 7763 2150 7809 2202
rect 7809 2150 7819 2202
rect 7843 2150 7873 2202
rect 7873 2150 7885 2202
rect 7885 2150 7899 2202
rect 7923 2150 7937 2202
rect 7937 2150 7949 2202
rect 7949 2150 7979 2202
rect 8003 2150 8013 2202
rect 8013 2150 8059 2202
rect 7763 2148 7819 2150
rect 7843 2148 7899 2150
rect 7923 2148 7979 2150
rect 8003 2148 8059 2150
rect 7763 1114 7819 1116
rect 7843 1114 7899 1116
rect 7923 1114 7979 1116
rect 8003 1114 8059 1116
rect 7763 1062 7809 1114
rect 7809 1062 7819 1114
rect 7843 1062 7873 1114
rect 7873 1062 7885 1114
rect 7885 1062 7899 1114
rect 7923 1062 7937 1114
rect 7937 1062 7949 1114
rect 7949 1062 7979 1114
rect 8003 1062 8013 1114
rect 8013 1062 8059 1114
rect 7763 1060 7819 1062
rect 7843 1060 7899 1062
rect 7923 1060 7979 1062
rect 8003 1060 8059 1062
rect 6826 584 6882 640
<< metal3 >>
rect 5901 9210 5967 9213
rect 8200 9210 9000 9240
rect 5901 9208 9000 9210
rect 5901 9152 5906 9208
rect 5962 9152 9000 9208
rect 5901 9150 9000 9152
rect 5901 9147 5967 9150
rect 8200 9120 9000 9150
rect 0 9074 800 9104
rect 3417 9074 3483 9077
rect 0 9072 3483 9074
rect 0 9016 3422 9072
rect 3478 9016 3483 9072
rect 0 9014 3483 9016
rect 0 8984 800 9014
rect 3417 9011 3483 9014
rect 3877 8938 3943 8941
rect 3877 8936 8218 8938
rect 3877 8880 3882 8936
rect 3938 8880 8218 8936
rect 3877 8878 8218 8880
rect 3877 8875 3943 8878
rect 8158 8832 8218 8878
rect 8158 8742 9000 8832
rect 2578 8736 2894 8737
rect 2578 8672 2584 8736
rect 2648 8672 2664 8736
rect 2728 8672 2744 8736
rect 2808 8672 2824 8736
rect 2888 8672 2894 8736
rect 2578 8671 2894 8672
rect 4303 8736 4619 8737
rect 4303 8672 4309 8736
rect 4373 8672 4389 8736
rect 4453 8672 4469 8736
rect 4533 8672 4549 8736
rect 4613 8672 4619 8736
rect 4303 8671 4619 8672
rect 6028 8736 6344 8737
rect 6028 8672 6034 8736
rect 6098 8672 6114 8736
rect 6178 8672 6194 8736
rect 6258 8672 6274 8736
rect 6338 8672 6344 8736
rect 6028 8671 6344 8672
rect 7753 8736 8069 8737
rect 7753 8672 7759 8736
rect 7823 8672 7839 8736
rect 7903 8672 7919 8736
rect 7983 8672 7999 8736
rect 8063 8672 8069 8736
rect 8200 8712 9000 8742
rect 7753 8671 8069 8672
rect 0 8394 800 8424
rect 1577 8394 1643 8397
rect 1761 8394 1827 8397
rect 0 8392 1827 8394
rect 0 8336 1582 8392
rect 1638 8336 1766 8392
rect 1822 8336 1827 8392
rect 0 8334 1827 8336
rect 0 8304 800 8334
rect 1577 8331 1643 8334
rect 1761 8331 1827 8334
rect 5625 8394 5691 8397
rect 8200 8394 9000 8424
rect 5625 8392 9000 8394
rect 5625 8336 5630 8392
rect 5686 8336 9000 8392
rect 5625 8334 9000 8336
rect 5625 8331 5691 8334
rect 8200 8304 9000 8334
rect 1716 8192 2032 8193
rect 1716 8128 1722 8192
rect 1786 8128 1802 8192
rect 1866 8128 1882 8192
rect 1946 8128 1962 8192
rect 2026 8128 2032 8192
rect 1716 8127 2032 8128
rect 3441 8192 3757 8193
rect 3441 8128 3447 8192
rect 3511 8128 3527 8192
rect 3591 8128 3607 8192
rect 3671 8128 3687 8192
rect 3751 8128 3757 8192
rect 3441 8127 3757 8128
rect 5166 8192 5482 8193
rect 5166 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5482 8192
rect 5166 8127 5482 8128
rect 6891 8192 7207 8193
rect 6891 8128 6897 8192
rect 6961 8128 6977 8192
rect 7041 8128 7057 8192
rect 7121 8128 7137 8192
rect 7201 8128 7207 8192
rect 6891 8127 7207 8128
rect 4705 7986 4771 7989
rect 8200 7986 9000 8016
rect 4705 7984 9000 7986
rect 4705 7928 4710 7984
rect 4766 7928 9000 7984
rect 4705 7926 9000 7928
rect 4705 7923 4771 7926
rect 8200 7896 9000 7926
rect 4613 7850 4679 7853
rect 4613 7848 8034 7850
rect 4613 7792 4618 7848
rect 4674 7816 8034 7848
rect 4674 7792 8218 7816
rect 4613 7790 8218 7792
rect 4613 7787 4679 7790
rect 7974 7756 8218 7790
rect 0 7714 800 7744
rect 0 7654 2514 7714
rect 0 7624 800 7654
rect 2454 7442 2514 7654
rect 2578 7648 2894 7649
rect 2578 7584 2584 7648
rect 2648 7584 2664 7648
rect 2728 7584 2744 7648
rect 2808 7584 2824 7648
rect 2888 7584 2894 7648
rect 2578 7583 2894 7584
rect 4303 7648 4619 7649
rect 4303 7584 4309 7648
rect 4373 7584 4389 7648
rect 4453 7584 4469 7648
rect 4533 7584 4549 7648
rect 4613 7584 4619 7648
rect 4303 7583 4619 7584
rect 6028 7648 6344 7649
rect 6028 7584 6034 7648
rect 6098 7584 6114 7648
rect 6178 7584 6194 7648
rect 6258 7584 6274 7648
rect 6338 7584 6344 7648
rect 6028 7583 6344 7584
rect 7753 7648 8069 7649
rect 7753 7584 7759 7648
rect 7823 7584 7839 7648
rect 7903 7584 7919 7648
rect 7983 7584 7999 7648
rect 8063 7584 8069 7648
rect 7753 7583 8069 7584
rect 8158 7608 8218 7756
rect 8158 7518 9000 7608
rect 8200 7488 9000 7518
rect 3325 7442 3391 7445
rect 2454 7440 3391 7442
rect 2454 7384 3330 7440
rect 3386 7384 3391 7440
rect 2454 7382 3391 7384
rect 3325 7379 3391 7382
rect 5441 7306 5507 7309
rect 5441 7304 7482 7306
rect 5441 7248 5446 7304
rect 5502 7248 7482 7304
rect 5441 7246 7482 7248
rect 5441 7243 5507 7246
rect 7422 7170 7482 7246
rect 8200 7170 9000 7200
rect 7422 7110 9000 7170
rect 1716 7104 2032 7105
rect 0 7034 800 7064
rect 1716 7040 1722 7104
rect 1786 7040 1802 7104
rect 1866 7040 1882 7104
rect 1946 7040 1962 7104
rect 2026 7040 2032 7104
rect 1716 7039 2032 7040
rect 3441 7104 3757 7105
rect 3441 7040 3447 7104
rect 3511 7040 3527 7104
rect 3591 7040 3607 7104
rect 3671 7040 3687 7104
rect 3751 7040 3757 7104
rect 3441 7039 3757 7040
rect 5166 7104 5482 7105
rect 5166 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5482 7104
rect 5166 7039 5482 7040
rect 6891 7104 7207 7105
rect 6891 7040 6897 7104
rect 6961 7040 6977 7104
rect 7041 7040 7057 7104
rect 7121 7040 7137 7104
rect 7201 7040 7207 7104
rect 8200 7080 9000 7110
rect 6891 7039 7207 7040
rect 1485 7034 1551 7037
rect 0 7032 1551 7034
rect 0 6976 1490 7032
rect 1546 6976 1551 7032
rect 0 6974 1551 6976
rect 0 6944 800 6974
rect 1485 6971 1551 6974
rect 4521 6762 4587 6765
rect 8200 6762 9000 6792
rect 4521 6760 9000 6762
rect 4521 6704 4526 6760
rect 4582 6704 9000 6760
rect 4521 6702 9000 6704
rect 4521 6699 4587 6702
rect 8200 6672 9000 6702
rect 2578 6560 2894 6561
rect 2578 6496 2584 6560
rect 2648 6496 2664 6560
rect 2728 6496 2744 6560
rect 2808 6496 2824 6560
rect 2888 6496 2894 6560
rect 2578 6495 2894 6496
rect 4303 6560 4619 6561
rect 4303 6496 4309 6560
rect 4373 6496 4389 6560
rect 4453 6496 4469 6560
rect 4533 6496 4549 6560
rect 4613 6496 4619 6560
rect 4303 6495 4619 6496
rect 6028 6560 6344 6561
rect 6028 6496 6034 6560
rect 6098 6496 6114 6560
rect 6178 6496 6194 6560
rect 6258 6496 6274 6560
rect 6338 6496 6344 6560
rect 6028 6495 6344 6496
rect 7753 6560 8069 6561
rect 7753 6496 7759 6560
rect 7823 6496 7839 6560
rect 7903 6496 7919 6560
rect 7983 6496 7999 6560
rect 8063 6496 8069 6560
rect 7753 6495 8069 6496
rect 0 6354 800 6384
rect 2957 6354 3023 6357
rect 0 6352 3023 6354
rect 0 6296 2962 6352
rect 3018 6296 3023 6352
rect 0 6294 3023 6296
rect 0 6264 800 6294
rect 2957 6291 3023 6294
rect 5441 6354 5507 6357
rect 8200 6354 9000 6384
rect 5441 6352 9000 6354
rect 5441 6296 5446 6352
rect 5502 6296 9000 6352
rect 5441 6294 9000 6296
rect 5441 6291 5507 6294
rect 8200 6264 9000 6294
rect 4797 6218 4863 6221
rect 4797 6216 7666 6218
rect 4797 6160 4802 6216
rect 4858 6160 7666 6216
rect 4797 6158 7666 6160
rect 4797 6155 4863 6158
rect 1716 6016 2032 6017
rect 1716 5952 1722 6016
rect 1786 5952 1802 6016
rect 1866 5952 1882 6016
rect 1946 5952 1962 6016
rect 2026 5952 2032 6016
rect 1716 5951 2032 5952
rect 3441 6016 3757 6017
rect 3441 5952 3447 6016
rect 3511 5952 3527 6016
rect 3591 5952 3607 6016
rect 3671 5952 3687 6016
rect 3751 5952 3757 6016
rect 3441 5951 3757 5952
rect 5166 6016 5482 6017
rect 5166 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5482 6016
rect 5166 5951 5482 5952
rect 6891 6016 7207 6017
rect 6891 5952 6897 6016
rect 6961 5952 6977 6016
rect 7041 5952 7057 6016
rect 7121 5952 7137 6016
rect 7201 5952 7207 6016
rect 6891 5951 7207 5952
rect 7606 5946 7666 6158
rect 8200 5946 9000 5976
rect 7606 5886 9000 5946
rect 8200 5856 9000 5886
rect 0 5674 800 5704
rect 3049 5674 3115 5677
rect 0 5672 3115 5674
rect 0 5616 3054 5672
rect 3110 5616 3115 5672
rect 0 5614 3115 5616
rect 0 5584 800 5614
rect 3049 5611 3115 5614
rect 7606 5614 8218 5674
rect 6545 5538 6611 5541
rect 7606 5538 7666 5614
rect 6545 5536 7666 5538
rect 6545 5480 6550 5536
rect 6606 5480 7666 5536
rect 6545 5478 7666 5480
rect 8158 5568 8218 5614
rect 8158 5478 9000 5568
rect 6545 5475 6611 5478
rect 2578 5472 2894 5473
rect 2578 5408 2584 5472
rect 2648 5408 2664 5472
rect 2728 5408 2744 5472
rect 2808 5408 2824 5472
rect 2888 5408 2894 5472
rect 2578 5407 2894 5408
rect 4303 5472 4619 5473
rect 4303 5408 4309 5472
rect 4373 5408 4389 5472
rect 4453 5408 4469 5472
rect 4533 5408 4549 5472
rect 4613 5408 4619 5472
rect 4303 5407 4619 5408
rect 6028 5472 6344 5473
rect 6028 5408 6034 5472
rect 6098 5408 6114 5472
rect 6178 5408 6194 5472
rect 6258 5408 6274 5472
rect 6338 5408 6344 5472
rect 6028 5407 6344 5408
rect 7753 5472 8069 5473
rect 7753 5408 7759 5472
rect 7823 5408 7839 5472
rect 7903 5408 7919 5472
rect 7983 5408 7999 5472
rect 8063 5408 8069 5472
rect 8200 5448 9000 5478
rect 7753 5407 8069 5408
rect 7465 5130 7531 5133
rect 8200 5130 9000 5160
rect 7465 5128 9000 5130
rect 7465 5072 7470 5128
rect 7526 5072 9000 5128
rect 7465 5070 9000 5072
rect 7465 5067 7531 5070
rect 8200 5040 9000 5070
rect 0 4994 800 5024
rect 0 4934 1594 4994
rect 0 4904 800 4934
rect 1534 4722 1594 4934
rect 1716 4928 2032 4929
rect 1716 4864 1722 4928
rect 1786 4864 1802 4928
rect 1866 4864 1882 4928
rect 1946 4864 1962 4928
rect 2026 4864 2032 4928
rect 1716 4863 2032 4864
rect 3441 4928 3757 4929
rect 3441 4864 3447 4928
rect 3511 4864 3527 4928
rect 3591 4864 3607 4928
rect 3671 4864 3687 4928
rect 3751 4864 3757 4928
rect 3441 4863 3757 4864
rect 5166 4928 5482 4929
rect 5166 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5482 4928
rect 5166 4863 5482 4864
rect 6891 4928 7207 4929
rect 6891 4864 6897 4928
rect 6961 4864 6977 4928
rect 7041 4864 7057 4928
rect 7121 4864 7137 4928
rect 7201 4864 7207 4928
rect 6891 4863 7207 4864
rect 3877 4722 3943 4725
rect 1534 4720 3943 4722
rect 1534 4664 3882 4720
rect 3938 4664 3943 4720
rect 1534 4662 3943 4664
rect 3877 4659 3943 4662
rect 7373 4722 7439 4725
rect 8200 4722 9000 4752
rect 7373 4720 9000 4722
rect 7373 4664 7378 4720
rect 7434 4664 9000 4720
rect 7373 4662 9000 4664
rect 7373 4659 7439 4662
rect 8200 4632 9000 4662
rect 2578 4384 2894 4385
rect 0 4314 800 4344
rect 2578 4320 2584 4384
rect 2648 4320 2664 4384
rect 2728 4320 2744 4384
rect 2808 4320 2824 4384
rect 2888 4320 2894 4384
rect 2578 4319 2894 4320
rect 4303 4384 4619 4385
rect 4303 4320 4309 4384
rect 4373 4320 4389 4384
rect 4453 4320 4469 4384
rect 4533 4320 4549 4384
rect 4613 4320 4619 4384
rect 4303 4319 4619 4320
rect 6028 4384 6344 4385
rect 6028 4320 6034 4384
rect 6098 4320 6114 4384
rect 6178 4320 6194 4384
rect 6258 4320 6274 4384
rect 6338 4320 6344 4384
rect 6028 4319 6344 4320
rect 7753 4384 8069 4385
rect 7753 4320 7759 4384
rect 7823 4320 7839 4384
rect 7903 4320 7919 4384
rect 7983 4320 7999 4384
rect 8063 4320 8069 4384
rect 7753 4319 8069 4320
rect 8200 4314 9000 4344
rect 0 4254 2146 4314
rect 0 4224 800 4254
rect 2086 4178 2146 4254
rect 8158 4224 9000 4314
rect 4061 4178 4127 4181
rect 2086 4176 4127 4178
rect 2086 4120 4066 4176
rect 4122 4120 4127 4176
rect 2086 4118 4127 4120
rect 4061 4115 4127 4118
rect 7281 4178 7347 4181
rect 8158 4178 8218 4224
rect 7281 4176 8218 4178
rect 7281 4120 7286 4176
rect 7342 4120 8218 4176
rect 7281 4118 8218 4120
rect 7281 4115 7347 4118
rect 6821 4042 6887 4045
rect 6821 4040 7482 4042
rect 6821 3984 6826 4040
rect 6882 3984 7482 4040
rect 6821 3982 7482 3984
rect 6821 3979 6887 3982
rect 7422 3906 7482 3982
rect 8200 3906 9000 3936
rect 7422 3846 9000 3906
rect 1716 3840 2032 3841
rect 1716 3776 1722 3840
rect 1786 3776 1802 3840
rect 1866 3776 1882 3840
rect 1946 3776 1962 3840
rect 2026 3776 2032 3840
rect 1716 3775 2032 3776
rect 3441 3840 3757 3841
rect 3441 3776 3447 3840
rect 3511 3776 3527 3840
rect 3591 3776 3607 3840
rect 3671 3776 3687 3840
rect 3751 3776 3757 3840
rect 3441 3775 3757 3776
rect 5166 3840 5482 3841
rect 5166 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5482 3840
rect 5166 3775 5482 3776
rect 6891 3840 7207 3841
rect 6891 3776 6897 3840
rect 6961 3776 6977 3840
rect 7041 3776 7057 3840
rect 7121 3776 7137 3840
rect 7201 3776 7207 3840
rect 8200 3816 9000 3846
rect 6891 3775 7207 3776
rect 0 3634 800 3664
rect 2957 3634 3023 3637
rect 0 3632 3023 3634
rect 0 3576 2962 3632
rect 3018 3576 3023 3632
rect 0 3574 3023 3576
rect 0 3544 800 3574
rect 2957 3571 3023 3574
rect 7281 3498 7347 3501
rect 8200 3498 9000 3528
rect 7281 3496 9000 3498
rect 7281 3440 7286 3496
rect 7342 3440 9000 3496
rect 7281 3438 9000 3440
rect 7281 3435 7347 3438
rect 8200 3408 9000 3438
rect 2578 3296 2894 3297
rect 2578 3232 2584 3296
rect 2648 3232 2664 3296
rect 2728 3232 2744 3296
rect 2808 3232 2824 3296
rect 2888 3232 2894 3296
rect 2578 3231 2894 3232
rect 4303 3296 4619 3297
rect 4303 3232 4309 3296
rect 4373 3232 4389 3296
rect 4453 3232 4469 3296
rect 4533 3232 4549 3296
rect 4613 3232 4619 3296
rect 4303 3231 4619 3232
rect 6028 3296 6344 3297
rect 6028 3232 6034 3296
rect 6098 3232 6114 3296
rect 6178 3232 6194 3296
rect 6258 3232 6274 3296
rect 6338 3232 6344 3296
rect 6028 3231 6344 3232
rect 7753 3296 8069 3297
rect 7753 3232 7759 3296
rect 7823 3232 7839 3296
rect 7903 3232 7919 3296
rect 7983 3232 7999 3296
rect 8063 3232 8069 3296
rect 7753 3231 8069 3232
rect 7281 3090 7347 3093
rect 8200 3090 9000 3120
rect 7281 3088 9000 3090
rect 7281 3032 7286 3088
rect 7342 3032 9000 3088
rect 7281 3030 9000 3032
rect 7281 3027 7347 3030
rect 8200 3000 9000 3030
rect 0 2954 800 2984
rect 2773 2954 2839 2957
rect 0 2952 2839 2954
rect 0 2896 2778 2952
rect 2834 2896 2839 2952
rect 0 2894 2839 2896
rect 0 2864 800 2894
rect 2773 2891 2839 2894
rect 1716 2752 2032 2753
rect 1716 2688 1722 2752
rect 1786 2688 1802 2752
rect 1866 2688 1882 2752
rect 1946 2688 1962 2752
rect 2026 2688 2032 2752
rect 1716 2687 2032 2688
rect 3441 2752 3757 2753
rect 3441 2688 3447 2752
rect 3511 2688 3527 2752
rect 3591 2688 3607 2752
rect 3671 2688 3687 2752
rect 3751 2688 3757 2752
rect 3441 2687 3757 2688
rect 5166 2752 5482 2753
rect 5166 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5482 2752
rect 5166 2687 5482 2688
rect 6891 2752 7207 2753
rect 6891 2688 6897 2752
rect 6961 2688 6977 2752
rect 7041 2688 7057 2752
rect 7121 2688 7137 2752
rect 7201 2688 7207 2752
rect 6891 2687 7207 2688
rect 7281 2682 7347 2685
rect 8200 2682 9000 2712
rect 7281 2680 9000 2682
rect 7281 2624 7286 2680
rect 7342 2624 9000 2680
rect 7281 2622 9000 2624
rect 7281 2619 7347 2622
rect 8200 2592 9000 2622
rect 7281 2410 7347 2413
rect 7281 2408 8218 2410
rect 7281 2352 7286 2408
rect 7342 2352 8218 2408
rect 7281 2350 8218 2352
rect 7281 2347 7347 2350
rect 8158 2304 8218 2350
rect 0 2274 800 2304
rect 0 2214 1410 2274
rect 8158 2214 9000 2304
rect 0 2184 800 2214
rect 1350 2002 1410 2214
rect 2578 2208 2894 2209
rect 2578 2144 2584 2208
rect 2648 2144 2664 2208
rect 2728 2144 2744 2208
rect 2808 2144 2824 2208
rect 2888 2144 2894 2208
rect 2578 2143 2894 2144
rect 4303 2208 4619 2209
rect 4303 2144 4309 2208
rect 4373 2144 4389 2208
rect 4453 2144 4469 2208
rect 4533 2144 4549 2208
rect 4613 2144 4619 2208
rect 4303 2143 4619 2144
rect 6028 2208 6344 2209
rect 6028 2144 6034 2208
rect 6098 2144 6114 2208
rect 6178 2144 6194 2208
rect 6258 2144 6274 2208
rect 6338 2144 6344 2208
rect 6028 2143 6344 2144
rect 7753 2208 8069 2209
rect 7753 2144 7759 2208
rect 7823 2144 7839 2208
rect 7903 2144 7919 2208
rect 7983 2144 7999 2208
rect 8063 2144 8069 2208
rect 8200 2184 9000 2214
rect 7753 2143 8069 2144
rect 2773 2002 2839 2005
rect 1350 2000 2839 2002
rect 1350 1944 2778 2000
rect 2834 1944 2839 2000
rect 1350 1942 2839 1944
rect 2773 1939 2839 1942
rect 5441 1866 5507 1869
rect 7281 1866 7347 1869
rect 8200 1866 9000 1896
rect 5441 1864 5642 1866
rect 5441 1808 5446 1864
rect 5502 1808 5642 1864
rect 5441 1806 5642 1808
rect 5441 1803 5507 1806
rect 1716 1664 2032 1665
rect 0 1594 800 1624
rect 1716 1600 1722 1664
rect 1786 1600 1802 1664
rect 1866 1600 1882 1664
rect 1946 1600 1962 1664
rect 2026 1600 2032 1664
rect 1716 1599 2032 1600
rect 3441 1664 3757 1665
rect 3441 1600 3447 1664
rect 3511 1600 3527 1664
rect 3591 1600 3607 1664
rect 3671 1600 3687 1664
rect 3751 1600 3757 1664
rect 3441 1599 3757 1600
rect 5166 1664 5482 1665
rect 5166 1600 5172 1664
rect 5236 1600 5252 1664
rect 5316 1600 5332 1664
rect 5396 1600 5412 1664
rect 5476 1600 5482 1664
rect 5166 1599 5482 1600
rect 1485 1594 1551 1597
rect 0 1592 1551 1594
rect 0 1536 1490 1592
rect 1546 1536 1551 1592
rect 0 1534 1551 1536
rect 0 1504 800 1534
rect 1485 1531 1551 1534
rect 5582 1458 5642 1806
rect 7281 1864 9000 1866
rect 7281 1808 7286 1864
rect 7342 1808 9000 1864
rect 7281 1806 9000 1808
rect 7281 1803 7347 1806
rect 8200 1776 9000 1806
rect 6891 1664 7207 1665
rect 6891 1600 6897 1664
rect 6961 1600 6977 1664
rect 7041 1600 7057 1664
rect 7121 1600 7137 1664
rect 7201 1600 7207 1664
rect 6891 1599 7207 1600
rect 8200 1458 9000 1488
rect 5582 1398 9000 1458
rect 8200 1368 9000 1398
rect 2578 1120 2894 1121
rect 2578 1056 2584 1120
rect 2648 1056 2664 1120
rect 2728 1056 2744 1120
rect 2808 1056 2824 1120
rect 2888 1056 2894 1120
rect 2578 1055 2894 1056
rect 4303 1120 4619 1121
rect 4303 1056 4309 1120
rect 4373 1056 4389 1120
rect 4453 1056 4469 1120
rect 4533 1056 4549 1120
rect 4613 1056 4619 1120
rect 4303 1055 4619 1056
rect 6028 1120 6344 1121
rect 6028 1056 6034 1120
rect 6098 1056 6114 1120
rect 6178 1056 6194 1120
rect 6258 1056 6274 1120
rect 6338 1056 6344 1120
rect 6028 1055 6344 1056
rect 7753 1120 8069 1121
rect 7753 1056 7759 1120
rect 7823 1056 7839 1120
rect 7903 1056 7919 1120
rect 7983 1056 7999 1120
rect 8063 1056 8069 1120
rect 7753 1055 8069 1056
rect 8200 1050 9000 1080
rect 8158 960 9000 1050
rect 0 914 800 944
rect 2957 914 3023 917
rect 0 912 3023 914
rect 0 856 2962 912
rect 3018 856 3023 912
rect 0 854 3023 856
rect 0 824 800 854
rect 2957 851 3023 854
rect 4981 914 5047 917
rect 8158 914 8218 960
rect 4981 912 8218 914
rect 4981 856 4986 912
rect 5042 856 8218 912
rect 4981 854 8218 856
rect 4981 851 5047 854
rect 6821 642 6887 645
rect 8200 642 9000 672
rect 6821 640 9000 642
rect 6821 584 6826 640
rect 6882 584 9000 640
rect 6821 582 9000 584
rect 6821 579 6887 582
rect 8200 552 9000 582
<< via3 >>
rect 2584 8732 2648 8736
rect 2584 8676 2588 8732
rect 2588 8676 2644 8732
rect 2644 8676 2648 8732
rect 2584 8672 2648 8676
rect 2664 8732 2728 8736
rect 2664 8676 2668 8732
rect 2668 8676 2724 8732
rect 2724 8676 2728 8732
rect 2664 8672 2728 8676
rect 2744 8732 2808 8736
rect 2744 8676 2748 8732
rect 2748 8676 2804 8732
rect 2804 8676 2808 8732
rect 2744 8672 2808 8676
rect 2824 8732 2888 8736
rect 2824 8676 2828 8732
rect 2828 8676 2884 8732
rect 2884 8676 2888 8732
rect 2824 8672 2888 8676
rect 4309 8732 4373 8736
rect 4309 8676 4313 8732
rect 4313 8676 4369 8732
rect 4369 8676 4373 8732
rect 4309 8672 4373 8676
rect 4389 8732 4453 8736
rect 4389 8676 4393 8732
rect 4393 8676 4449 8732
rect 4449 8676 4453 8732
rect 4389 8672 4453 8676
rect 4469 8732 4533 8736
rect 4469 8676 4473 8732
rect 4473 8676 4529 8732
rect 4529 8676 4533 8732
rect 4469 8672 4533 8676
rect 4549 8732 4613 8736
rect 4549 8676 4553 8732
rect 4553 8676 4609 8732
rect 4609 8676 4613 8732
rect 4549 8672 4613 8676
rect 6034 8732 6098 8736
rect 6034 8676 6038 8732
rect 6038 8676 6094 8732
rect 6094 8676 6098 8732
rect 6034 8672 6098 8676
rect 6114 8732 6178 8736
rect 6114 8676 6118 8732
rect 6118 8676 6174 8732
rect 6174 8676 6178 8732
rect 6114 8672 6178 8676
rect 6194 8732 6258 8736
rect 6194 8676 6198 8732
rect 6198 8676 6254 8732
rect 6254 8676 6258 8732
rect 6194 8672 6258 8676
rect 6274 8732 6338 8736
rect 6274 8676 6278 8732
rect 6278 8676 6334 8732
rect 6334 8676 6338 8732
rect 6274 8672 6338 8676
rect 7759 8732 7823 8736
rect 7759 8676 7763 8732
rect 7763 8676 7819 8732
rect 7819 8676 7823 8732
rect 7759 8672 7823 8676
rect 7839 8732 7903 8736
rect 7839 8676 7843 8732
rect 7843 8676 7899 8732
rect 7899 8676 7903 8732
rect 7839 8672 7903 8676
rect 7919 8732 7983 8736
rect 7919 8676 7923 8732
rect 7923 8676 7979 8732
rect 7979 8676 7983 8732
rect 7919 8672 7983 8676
rect 7999 8732 8063 8736
rect 7999 8676 8003 8732
rect 8003 8676 8059 8732
rect 8059 8676 8063 8732
rect 7999 8672 8063 8676
rect 1722 8188 1786 8192
rect 1722 8132 1726 8188
rect 1726 8132 1782 8188
rect 1782 8132 1786 8188
rect 1722 8128 1786 8132
rect 1802 8188 1866 8192
rect 1802 8132 1806 8188
rect 1806 8132 1862 8188
rect 1862 8132 1866 8188
rect 1802 8128 1866 8132
rect 1882 8188 1946 8192
rect 1882 8132 1886 8188
rect 1886 8132 1942 8188
rect 1942 8132 1946 8188
rect 1882 8128 1946 8132
rect 1962 8188 2026 8192
rect 1962 8132 1966 8188
rect 1966 8132 2022 8188
rect 2022 8132 2026 8188
rect 1962 8128 2026 8132
rect 3447 8188 3511 8192
rect 3447 8132 3451 8188
rect 3451 8132 3507 8188
rect 3507 8132 3511 8188
rect 3447 8128 3511 8132
rect 3527 8188 3591 8192
rect 3527 8132 3531 8188
rect 3531 8132 3587 8188
rect 3587 8132 3591 8188
rect 3527 8128 3591 8132
rect 3607 8188 3671 8192
rect 3607 8132 3611 8188
rect 3611 8132 3667 8188
rect 3667 8132 3671 8188
rect 3607 8128 3671 8132
rect 3687 8188 3751 8192
rect 3687 8132 3691 8188
rect 3691 8132 3747 8188
rect 3747 8132 3751 8188
rect 3687 8128 3751 8132
rect 5172 8188 5236 8192
rect 5172 8132 5176 8188
rect 5176 8132 5232 8188
rect 5232 8132 5236 8188
rect 5172 8128 5236 8132
rect 5252 8188 5316 8192
rect 5252 8132 5256 8188
rect 5256 8132 5312 8188
rect 5312 8132 5316 8188
rect 5252 8128 5316 8132
rect 5332 8188 5396 8192
rect 5332 8132 5336 8188
rect 5336 8132 5392 8188
rect 5392 8132 5396 8188
rect 5332 8128 5396 8132
rect 5412 8188 5476 8192
rect 5412 8132 5416 8188
rect 5416 8132 5472 8188
rect 5472 8132 5476 8188
rect 5412 8128 5476 8132
rect 6897 8188 6961 8192
rect 6897 8132 6901 8188
rect 6901 8132 6957 8188
rect 6957 8132 6961 8188
rect 6897 8128 6961 8132
rect 6977 8188 7041 8192
rect 6977 8132 6981 8188
rect 6981 8132 7037 8188
rect 7037 8132 7041 8188
rect 6977 8128 7041 8132
rect 7057 8188 7121 8192
rect 7057 8132 7061 8188
rect 7061 8132 7117 8188
rect 7117 8132 7121 8188
rect 7057 8128 7121 8132
rect 7137 8188 7201 8192
rect 7137 8132 7141 8188
rect 7141 8132 7197 8188
rect 7197 8132 7201 8188
rect 7137 8128 7201 8132
rect 2584 7644 2648 7648
rect 2584 7588 2588 7644
rect 2588 7588 2644 7644
rect 2644 7588 2648 7644
rect 2584 7584 2648 7588
rect 2664 7644 2728 7648
rect 2664 7588 2668 7644
rect 2668 7588 2724 7644
rect 2724 7588 2728 7644
rect 2664 7584 2728 7588
rect 2744 7644 2808 7648
rect 2744 7588 2748 7644
rect 2748 7588 2804 7644
rect 2804 7588 2808 7644
rect 2744 7584 2808 7588
rect 2824 7644 2888 7648
rect 2824 7588 2828 7644
rect 2828 7588 2884 7644
rect 2884 7588 2888 7644
rect 2824 7584 2888 7588
rect 4309 7644 4373 7648
rect 4309 7588 4313 7644
rect 4313 7588 4369 7644
rect 4369 7588 4373 7644
rect 4309 7584 4373 7588
rect 4389 7644 4453 7648
rect 4389 7588 4393 7644
rect 4393 7588 4449 7644
rect 4449 7588 4453 7644
rect 4389 7584 4453 7588
rect 4469 7644 4533 7648
rect 4469 7588 4473 7644
rect 4473 7588 4529 7644
rect 4529 7588 4533 7644
rect 4469 7584 4533 7588
rect 4549 7644 4613 7648
rect 4549 7588 4553 7644
rect 4553 7588 4609 7644
rect 4609 7588 4613 7644
rect 4549 7584 4613 7588
rect 6034 7644 6098 7648
rect 6034 7588 6038 7644
rect 6038 7588 6094 7644
rect 6094 7588 6098 7644
rect 6034 7584 6098 7588
rect 6114 7644 6178 7648
rect 6114 7588 6118 7644
rect 6118 7588 6174 7644
rect 6174 7588 6178 7644
rect 6114 7584 6178 7588
rect 6194 7644 6258 7648
rect 6194 7588 6198 7644
rect 6198 7588 6254 7644
rect 6254 7588 6258 7644
rect 6194 7584 6258 7588
rect 6274 7644 6338 7648
rect 6274 7588 6278 7644
rect 6278 7588 6334 7644
rect 6334 7588 6338 7644
rect 6274 7584 6338 7588
rect 7759 7644 7823 7648
rect 7759 7588 7763 7644
rect 7763 7588 7819 7644
rect 7819 7588 7823 7644
rect 7759 7584 7823 7588
rect 7839 7644 7903 7648
rect 7839 7588 7843 7644
rect 7843 7588 7899 7644
rect 7899 7588 7903 7644
rect 7839 7584 7903 7588
rect 7919 7644 7983 7648
rect 7919 7588 7923 7644
rect 7923 7588 7979 7644
rect 7979 7588 7983 7644
rect 7919 7584 7983 7588
rect 7999 7644 8063 7648
rect 7999 7588 8003 7644
rect 8003 7588 8059 7644
rect 8059 7588 8063 7644
rect 7999 7584 8063 7588
rect 1722 7100 1786 7104
rect 1722 7044 1726 7100
rect 1726 7044 1782 7100
rect 1782 7044 1786 7100
rect 1722 7040 1786 7044
rect 1802 7100 1866 7104
rect 1802 7044 1806 7100
rect 1806 7044 1862 7100
rect 1862 7044 1866 7100
rect 1802 7040 1866 7044
rect 1882 7100 1946 7104
rect 1882 7044 1886 7100
rect 1886 7044 1942 7100
rect 1942 7044 1946 7100
rect 1882 7040 1946 7044
rect 1962 7100 2026 7104
rect 1962 7044 1966 7100
rect 1966 7044 2022 7100
rect 2022 7044 2026 7100
rect 1962 7040 2026 7044
rect 3447 7100 3511 7104
rect 3447 7044 3451 7100
rect 3451 7044 3507 7100
rect 3507 7044 3511 7100
rect 3447 7040 3511 7044
rect 3527 7100 3591 7104
rect 3527 7044 3531 7100
rect 3531 7044 3587 7100
rect 3587 7044 3591 7100
rect 3527 7040 3591 7044
rect 3607 7100 3671 7104
rect 3607 7044 3611 7100
rect 3611 7044 3667 7100
rect 3667 7044 3671 7100
rect 3607 7040 3671 7044
rect 3687 7100 3751 7104
rect 3687 7044 3691 7100
rect 3691 7044 3747 7100
rect 3747 7044 3751 7100
rect 3687 7040 3751 7044
rect 5172 7100 5236 7104
rect 5172 7044 5176 7100
rect 5176 7044 5232 7100
rect 5232 7044 5236 7100
rect 5172 7040 5236 7044
rect 5252 7100 5316 7104
rect 5252 7044 5256 7100
rect 5256 7044 5312 7100
rect 5312 7044 5316 7100
rect 5252 7040 5316 7044
rect 5332 7100 5396 7104
rect 5332 7044 5336 7100
rect 5336 7044 5392 7100
rect 5392 7044 5396 7100
rect 5332 7040 5396 7044
rect 5412 7100 5476 7104
rect 5412 7044 5416 7100
rect 5416 7044 5472 7100
rect 5472 7044 5476 7100
rect 5412 7040 5476 7044
rect 6897 7100 6961 7104
rect 6897 7044 6901 7100
rect 6901 7044 6957 7100
rect 6957 7044 6961 7100
rect 6897 7040 6961 7044
rect 6977 7100 7041 7104
rect 6977 7044 6981 7100
rect 6981 7044 7037 7100
rect 7037 7044 7041 7100
rect 6977 7040 7041 7044
rect 7057 7100 7121 7104
rect 7057 7044 7061 7100
rect 7061 7044 7117 7100
rect 7117 7044 7121 7100
rect 7057 7040 7121 7044
rect 7137 7100 7201 7104
rect 7137 7044 7141 7100
rect 7141 7044 7197 7100
rect 7197 7044 7201 7100
rect 7137 7040 7201 7044
rect 2584 6556 2648 6560
rect 2584 6500 2588 6556
rect 2588 6500 2644 6556
rect 2644 6500 2648 6556
rect 2584 6496 2648 6500
rect 2664 6556 2728 6560
rect 2664 6500 2668 6556
rect 2668 6500 2724 6556
rect 2724 6500 2728 6556
rect 2664 6496 2728 6500
rect 2744 6556 2808 6560
rect 2744 6500 2748 6556
rect 2748 6500 2804 6556
rect 2804 6500 2808 6556
rect 2744 6496 2808 6500
rect 2824 6556 2888 6560
rect 2824 6500 2828 6556
rect 2828 6500 2884 6556
rect 2884 6500 2888 6556
rect 2824 6496 2888 6500
rect 4309 6556 4373 6560
rect 4309 6500 4313 6556
rect 4313 6500 4369 6556
rect 4369 6500 4373 6556
rect 4309 6496 4373 6500
rect 4389 6556 4453 6560
rect 4389 6500 4393 6556
rect 4393 6500 4449 6556
rect 4449 6500 4453 6556
rect 4389 6496 4453 6500
rect 4469 6556 4533 6560
rect 4469 6500 4473 6556
rect 4473 6500 4529 6556
rect 4529 6500 4533 6556
rect 4469 6496 4533 6500
rect 4549 6556 4613 6560
rect 4549 6500 4553 6556
rect 4553 6500 4609 6556
rect 4609 6500 4613 6556
rect 4549 6496 4613 6500
rect 6034 6556 6098 6560
rect 6034 6500 6038 6556
rect 6038 6500 6094 6556
rect 6094 6500 6098 6556
rect 6034 6496 6098 6500
rect 6114 6556 6178 6560
rect 6114 6500 6118 6556
rect 6118 6500 6174 6556
rect 6174 6500 6178 6556
rect 6114 6496 6178 6500
rect 6194 6556 6258 6560
rect 6194 6500 6198 6556
rect 6198 6500 6254 6556
rect 6254 6500 6258 6556
rect 6194 6496 6258 6500
rect 6274 6556 6338 6560
rect 6274 6500 6278 6556
rect 6278 6500 6334 6556
rect 6334 6500 6338 6556
rect 6274 6496 6338 6500
rect 7759 6556 7823 6560
rect 7759 6500 7763 6556
rect 7763 6500 7819 6556
rect 7819 6500 7823 6556
rect 7759 6496 7823 6500
rect 7839 6556 7903 6560
rect 7839 6500 7843 6556
rect 7843 6500 7899 6556
rect 7899 6500 7903 6556
rect 7839 6496 7903 6500
rect 7919 6556 7983 6560
rect 7919 6500 7923 6556
rect 7923 6500 7979 6556
rect 7979 6500 7983 6556
rect 7919 6496 7983 6500
rect 7999 6556 8063 6560
rect 7999 6500 8003 6556
rect 8003 6500 8059 6556
rect 8059 6500 8063 6556
rect 7999 6496 8063 6500
rect 1722 6012 1786 6016
rect 1722 5956 1726 6012
rect 1726 5956 1782 6012
rect 1782 5956 1786 6012
rect 1722 5952 1786 5956
rect 1802 6012 1866 6016
rect 1802 5956 1806 6012
rect 1806 5956 1862 6012
rect 1862 5956 1866 6012
rect 1802 5952 1866 5956
rect 1882 6012 1946 6016
rect 1882 5956 1886 6012
rect 1886 5956 1942 6012
rect 1942 5956 1946 6012
rect 1882 5952 1946 5956
rect 1962 6012 2026 6016
rect 1962 5956 1966 6012
rect 1966 5956 2022 6012
rect 2022 5956 2026 6012
rect 1962 5952 2026 5956
rect 3447 6012 3511 6016
rect 3447 5956 3451 6012
rect 3451 5956 3507 6012
rect 3507 5956 3511 6012
rect 3447 5952 3511 5956
rect 3527 6012 3591 6016
rect 3527 5956 3531 6012
rect 3531 5956 3587 6012
rect 3587 5956 3591 6012
rect 3527 5952 3591 5956
rect 3607 6012 3671 6016
rect 3607 5956 3611 6012
rect 3611 5956 3667 6012
rect 3667 5956 3671 6012
rect 3607 5952 3671 5956
rect 3687 6012 3751 6016
rect 3687 5956 3691 6012
rect 3691 5956 3747 6012
rect 3747 5956 3751 6012
rect 3687 5952 3751 5956
rect 5172 6012 5236 6016
rect 5172 5956 5176 6012
rect 5176 5956 5232 6012
rect 5232 5956 5236 6012
rect 5172 5952 5236 5956
rect 5252 6012 5316 6016
rect 5252 5956 5256 6012
rect 5256 5956 5312 6012
rect 5312 5956 5316 6012
rect 5252 5952 5316 5956
rect 5332 6012 5396 6016
rect 5332 5956 5336 6012
rect 5336 5956 5392 6012
rect 5392 5956 5396 6012
rect 5332 5952 5396 5956
rect 5412 6012 5476 6016
rect 5412 5956 5416 6012
rect 5416 5956 5472 6012
rect 5472 5956 5476 6012
rect 5412 5952 5476 5956
rect 6897 6012 6961 6016
rect 6897 5956 6901 6012
rect 6901 5956 6957 6012
rect 6957 5956 6961 6012
rect 6897 5952 6961 5956
rect 6977 6012 7041 6016
rect 6977 5956 6981 6012
rect 6981 5956 7037 6012
rect 7037 5956 7041 6012
rect 6977 5952 7041 5956
rect 7057 6012 7121 6016
rect 7057 5956 7061 6012
rect 7061 5956 7117 6012
rect 7117 5956 7121 6012
rect 7057 5952 7121 5956
rect 7137 6012 7201 6016
rect 7137 5956 7141 6012
rect 7141 5956 7197 6012
rect 7197 5956 7201 6012
rect 7137 5952 7201 5956
rect 2584 5468 2648 5472
rect 2584 5412 2588 5468
rect 2588 5412 2644 5468
rect 2644 5412 2648 5468
rect 2584 5408 2648 5412
rect 2664 5468 2728 5472
rect 2664 5412 2668 5468
rect 2668 5412 2724 5468
rect 2724 5412 2728 5468
rect 2664 5408 2728 5412
rect 2744 5468 2808 5472
rect 2744 5412 2748 5468
rect 2748 5412 2804 5468
rect 2804 5412 2808 5468
rect 2744 5408 2808 5412
rect 2824 5468 2888 5472
rect 2824 5412 2828 5468
rect 2828 5412 2884 5468
rect 2884 5412 2888 5468
rect 2824 5408 2888 5412
rect 4309 5468 4373 5472
rect 4309 5412 4313 5468
rect 4313 5412 4369 5468
rect 4369 5412 4373 5468
rect 4309 5408 4373 5412
rect 4389 5468 4453 5472
rect 4389 5412 4393 5468
rect 4393 5412 4449 5468
rect 4449 5412 4453 5468
rect 4389 5408 4453 5412
rect 4469 5468 4533 5472
rect 4469 5412 4473 5468
rect 4473 5412 4529 5468
rect 4529 5412 4533 5468
rect 4469 5408 4533 5412
rect 4549 5468 4613 5472
rect 4549 5412 4553 5468
rect 4553 5412 4609 5468
rect 4609 5412 4613 5468
rect 4549 5408 4613 5412
rect 6034 5468 6098 5472
rect 6034 5412 6038 5468
rect 6038 5412 6094 5468
rect 6094 5412 6098 5468
rect 6034 5408 6098 5412
rect 6114 5468 6178 5472
rect 6114 5412 6118 5468
rect 6118 5412 6174 5468
rect 6174 5412 6178 5468
rect 6114 5408 6178 5412
rect 6194 5468 6258 5472
rect 6194 5412 6198 5468
rect 6198 5412 6254 5468
rect 6254 5412 6258 5468
rect 6194 5408 6258 5412
rect 6274 5468 6338 5472
rect 6274 5412 6278 5468
rect 6278 5412 6334 5468
rect 6334 5412 6338 5468
rect 6274 5408 6338 5412
rect 7759 5468 7823 5472
rect 7759 5412 7763 5468
rect 7763 5412 7819 5468
rect 7819 5412 7823 5468
rect 7759 5408 7823 5412
rect 7839 5468 7903 5472
rect 7839 5412 7843 5468
rect 7843 5412 7899 5468
rect 7899 5412 7903 5468
rect 7839 5408 7903 5412
rect 7919 5468 7983 5472
rect 7919 5412 7923 5468
rect 7923 5412 7979 5468
rect 7979 5412 7983 5468
rect 7919 5408 7983 5412
rect 7999 5468 8063 5472
rect 7999 5412 8003 5468
rect 8003 5412 8059 5468
rect 8059 5412 8063 5468
rect 7999 5408 8063 5412
rect 1722 4924 1786 4928
rect 1722 4868 1726 4924
rect 1726 4868 1782 4924
rect 1782 4868 1786 4924
rect 1722 4864 1786 4868
rect 1802 4924 1866 4928
rect 1802 4868 1806 4924
rect 1806 4868 1862 4924
rect 1862 4868 1866 4924
rect 1802 4864 1866 4868
rect 1882 4924 1946 4928
rect 1882 4868 1886 4924
rect 1886 4868 1942 4924
rect 1942 4868 1946 4924
rect 1882 4864 1946 4868
rect 1962 4924 2026 4928
rect 1962 4868 1966 4924
rect 1966 4868 2022 4924
rect 2022 4868 2026 4924
rect 1962 4864 2026 4868
rect 3447 4924 3511 4928
rect 3447 4868 3451 4924
rect 3451 4868 3507 4924
rect 3507 4868 3511 4924
rect 3447 4864 3511 4868
rect 3527 4924 3591 4928
rect 3527 4868 3531 4924
rect 3531 4868 3587 4924
rect 3587 4868 3591 4924
rect 3527 4864 3591 4868
rect 3607 4924 3671 4928
rect 3607 4868 3611 4924
rect 3611 4868 3667 4924
rect 3667 4868 3671 4924
rect 3607 4864 3671 4868
rect 3687 4924 3751 4928
rect 3687 4868 3691 4924
rect 3691 4868 3747 4924
rect 3747 4868 3751 4924
rect 3687 4864 3751 4868
rect 5172 4924 5236 4928
rect 5172 4868 5176 4924
rect 5176 4868 5232 4924
rect 5232 4868 5236 4924
rect 5172 4864 5236 4868
rect 5252 4924 5316 4928
rect 5252 4868 5256 4924
rect 5256 4868 5312 4924
rect 5312 4868 5316 4924
rect 5252 4864 5316 4868
rect 5332 4924 5396 4928
rect 5332 4868 5336 4924
rect 5336 4868 5392 4924
rect 5392 4868 5396 4924
rect 5332 4864 5396 4868
rect 5412 4924 5476 4928
rect 5412 4868 5416 4924
rect 5416 4868 5472 4924
rect 5472 4868 5476 4924
rect 5412 4864 5476 4868
rect 6897 4924 6961 4928
rect 6897 4868 6901 4924
rect 6901 4868 6957 4924
rect 6957 4868 6961 4924
rect 6897 4864 6961 4868
rect 6977 4924 7041 4928
rect 6977 4868 6981 4924
rect 6981 4868 7037 4924
rect 7037 4868 7041 4924
rect 6977 4864 7041 4868
rect 7057 4924 7121 4928
rect 7057 4868 7061 4924
rect 7061 4868 7117 4924
rect 7117 4868 7121 4924
rect 7057 4864 7121 4868
rect 7137 4924 7201 4928
rect 7137 4868 7141 4924
rect 7141 4868 7197 4924
rect 7197 4868 7201 4924
rect 7137 4864 7201 4868
rect 2584 4380 2648 4384
rect 2584 4324 2588 4380
rect 2588 4324 2644 4380
rect 2644 4324 2648 4380
rect 2584 4320 2648 4324
rect 2664 4380 2728 4384
rect 2664 4324 2668 4380
rect 2668 4324 2724 4380
rect 2724 4324 2728 4380
rect 2664 4320 2728 4324
rect 2744 4380 2808 4384
rect 2744 4324 2748 4380
rect 2748 4324 2804 4380
rect 2804 4324 2808 4380
rect 2744 4320 2808 4324
rect 2824 4380 2888 4384
rect 2824 4324 2828 4380
rect 2828 4324 2884 4380
rect 2884 4324 2888 4380
rect 2824 4320 2888 4324
rect 4309 4380 4373 4384
rect 4309 4324 4313 4380
rect 4313 4324 4369 4380
rect 4369 4324 4373 4380
rect 4309 4320 4373 4324
rect 4389 4380 4453 4384
rect 4389 4324 4393 4380
rect 4393 4324 4449 4380
rect 4449 4324 4453 4380
rect 4389 4320 4453 4324
rect 4469 4380 4533 4384
rect 4469 4324 4473 4380
rect 4473 4324 4529 4380
rect 4529 4324 4533 4380
rect 4469 4320 4533 4324
rect 4549 4380 4613 4384
rect 4549 4324 4553 4380
rect 4553 4324 4609 4380
rect 4609 4324 4613 4380
rect 4549 4320 4613 4324
rect 6034 4380 6098 4384
rect 6034 4324 6038 4380
rect 6038 4324 6094 4380
rect 6094 4324 6098 4380
rect 6034 4320 6098 4324
rect 6114 4380 6178 4384
rect 6114 4324 6118 4380
rect 6118 4324 6174 4380
rect 6174 4324 6178 4380
rect 6114 4320 6178 4324
rect 6194 4380 6258 4384
rect 6194 4324 6198 4380
rect 6198 4324 6254 4380
rect 6254 4324 6258 4380
rect 6194 4320 6258 4324
rect 6274 4380 6338 4384
rect 6274 4324 6278 4380
rect 6278 4324 6334 4380
rect 6334 4324 6338 4380
rect 6274 4320 6338 4324
rect 7759 4380 7823 4384
rect 7759 4324 7763 4380
rect 7763 4324 7819 4380
rect 7819 4324 7823 4380
rect 7759 4320 7823 4324
rect 7839 4380 7903 4384
rect 7839 4324 7843 4380
rect 7843 4324 7899 4380
rect 7899 4324 7903 4380
rect 7839 4320 7903 4324
rect 7919 4380 7983 4384
rect 7919 4324 7923 4380
rect 7923 4324 7979 4380
rect 7979 4324 7983 4380
rect 7919 4320 7983 4324
rect 7999 4380 8063 4384
rect 7999 4324 8003 4380
rect 8003 4324 8059 4380
rect 8059 4324 8063 4380
rect 7999 4320 8063 4324
rect 1722 3836 1786 3840
rect 1722 3780 1726 3836
rect 1726 3780 1782 3836
rect 1782 3780 1786 3836
rect 1722 3776 1786 3780
rect 1802 3836 1866 3840
rect 1802 3780 1806 3836
rect 1806 3780 1862 3836
rect 1862 3780 1866 3836
rect 1802 3776 1866 3780
rect 1882 3836 1946 3840
rect 1882 3780 1886 3836
rect 1886 3780 1942 3836
rect 1942 3780 1946 3836
rect 1882 3776 1946 3780
rect 1962 3836 2026 3840
rect 1962 3780 1966 3836
rect 1966 3780 2022 3836
rect 2022 3780 2026 3836
rect 1962 3776 2026 3780
rect 3447 3836 3511 3840
rect 3447 3780 3451 3836
rect 3451 3780 3507 3836
rect 3507 3780 3511 3836
rect 3447 3776 3511 3780
rect 3527 3836 3591 3840
rect 3527 3780 3531 3836
rect 3531 3780 3587 3836
rect 3587 3780 3591 3836
rect 3527 3776 3591 3780
rect 3607 3836 3671 3840
rect 3607 3780 3611 3836
rect 3611 3780 3667 3836
rect 3667 3780 3671 3836
rect 3607 3776 3671 3780
rect 3687 3836 3751 3840
rect 3687 3780 3691 3836
rect 3691 3780 3747 3836
rect 3747 3780 3751 3836
rect 3687 3776 3751 3780
rect 5172 3836 5236 3840
rect 5172 3780 5176 3836
rect 5176 3780 5232 3836
rect 5232 3780 5236 3836
rect 5172 3776 5236 3780
rect 5252 3836 5316 3840
rect 5252 3780 5256 3836
rect 5256 3780 5312 3836
rect 5312 3780 5316 3836
rect 5252 3776 5316 3780
rect 5332 3836 5396 3840
rect 5332 3780 5336 3836
rect 5336 3780 5392 3836
rect 5392 3780 5396 3836
rect 5332 3776 5396 3780
rect 5412 3836 5476 3840
rect 5412 3780 5416 3836
rect 5416 3780 5472 3836
rect 5472 3780 5476 3836
rect 5412 3776 5476 3780
rect 6897 3836 6961 3840
rect 6897 3780 6901 3836
rect 6901 3780 6957 3836
rect 6957 3780 6961 3836
rect 6897 3776 6961 3780
rect 6977 3836 7041 3840
rect 6977 3780 6981 3836
rect 6981 3780 7037 3836
rect 7037 3780 7041 3836
rect 6977 3776 7041 3780
rect 7057 3836 7121 3840
rect 7057 3780 7061 3836
rect 7061 3780 7117 3836
rect 7117 3780 7121 3836
rect 7057 3776 7121 3780
rect 7137 3836 7201 3840
rect 7137 3780 7141 3836
rect 7141 3780 7197 3836
rect 7197 3780 7201 3836
rect 7137 3776 7201 3780
rect 2584 3292 2648 3296
rect 2584 3236 2588 3292
rect 2588 3236 2644 3292
rect 2644 3236 2648 3292
rect 2584 3232 2648 3236
rect 2664 3292 2728 3296
rect 2664 3236 2668 3292
rect 2668 3236 2724 3292
rect 2724 3236 2728 3292
rect 2664 3232 2728 3236
rect 2744 3292 2808 3296
rect 2744 3236 2748 3292
rect 2748 3236 2804 3292
rect 2804 3236 2808 3292
rect 2744 3232 2808 3236
rect 2824 3292 2888 3296
rect 2824 3236 2828 3292
rect 2828 3236 2884 3292
rect 2884 3236 2888 3292
rect 2824 3232 2888 3236
rect 4309 3292 4373 3296
rect 4309 3236 4313 3292
rect 4313 3236 4369 3292
rect 4369 3236 4373 3292
rect 4309 3232 4373 3236
rect 4389 3292 4453 3296
rect 4389 3236 4393 3292
rect 4393 3236 4449 3292
rect 4449 3236 4453 3292
rect 4389 3232 4453 3236
rect 4469 3292 4533 3296
rect 4469 3236 4473 3292
rect 4473 3236 4529 3292
rect 4529 3236 4533 3292
rect 4469 3232 4533 3236
rect 4549 3292 4613 3296
rect 4549 3236 4553 3292
rect 4553 3236 4609 3292
rect 4609 3236 4613 3292
rect 4549 3232 4613 3236
rect 6034 3292 6098 3296
rect 6034 3236 6038 3292
rect 6038 3236 6094 3292
rect 6094 3236 6098 3292
rect 6034 3232 6098 3236
rect 6114 3292 6178 3296
rect 6114 3236 6118 3292
rect 6118 3236 6174 3292
rect 6174 3236 6178 3292
rect 6114 3232 6178 3236
rect 6194 3292 6258 3296
rect 6194 3236 6198 3292
rect 6198 3236 6254 3292
rect 6254 3236 6258 3292
rect 6194 3232 6258 3236
rect 6274 3292 6338 3296
rect 6274 3236 6278 3292
rect 6278 3236 6334 3292
rect 6334 3236 6338 3292
rect 6274 3232 6338 3236
rect 7759 3292 7823 3296
rect 7759 3236 7763 3292
rect 7763 3236 7819 3292
rect 7819 3236 7823 3292
rect 7759 3232 7823 3236
rect 7839 3292 7903 3296
rect 7839 3236 7843 3292
rect 7843 3236 7899 3292
rect 7899 3236 7903 3292
rect 7839 3232 7903 3236
rect 7919 3292 7983 3296
rect 7919 3236 7923 3292
rect 7923 3236 7979 3292
rect 7979 3236 7983 3292
rect 7919 3232 7983 3236
rect 7999 3292 8063 3296
rect 7999 3236 8003 3292
rect 8003 3236 8059 3292
rect 8059 3236 8063 3292
rect 7999 3232 8063 3236
rect 1722 2748 1786 2752
rect 1722 2692 1726 2748
rect 1726 2692 1782 2748
rect 1782 2692 1786 2748
rect 1722 2688 1786 2692
rect 1802 2748 1866 2752
rect 1802 2692 1806 2748
rect 1806 2692 1862 2748
rect 1862 2692 1866 2748
rect 1802 2688 1866 2692
rect 1882 2748 1946 2752
rect 1882 2692 1886 2748
rect 1886 2692 1942 2748
rect 1942 2692 1946 2748
rect 1882 2688 1946 2692
rect 1962 2748 2026 2752
rect 1962 2692 1966 2748
rect 1966 2692 2022 2748
rect 2022 2692 2026 2748
rect 1962 2688 2026 2692
rect 3447 2748 3511 2752
rect 3447 2692 3451 2748
rect 3451 2692 3507 2748
rect 3507 2692 3511 2748
rect 3447 2688 3511 2692
rect 3527 2748 3591 2752
rect 3527 2692 3531 2748
rect 3531 2692 3587 2748
rect 3587 2692 3591 2748
rect 3527 2688 3591 2692
rect 3607 2748 3671 2752
rect 3607 2692 3611 2748
rect 3611 2692 3667 2748
rect 3667 2692 3671 2748
rect 3607 2688 3671 2692
rect 3687 2748 3751 2752
rect 3687 2692 3691 2748
rect 3691 2692 3747 2748
rect 3747 2692 3751 2748
rect 3687 2688 3751 2692
rect 5172 2748 5236 2752
rect 5172 2692 5176 2748
rect 5176 2692 5232 2748
rect 5232 2692 5236 2748
rect 5172 2688 5236 2692
rect 5252 2748 5316 2752
rect 5252 2692 5256 2748
rect 5256 2692 5312 2748
rect 5312 2692 5316 2748
rect 5252 2688 5316 2692
rect 5332 2748 5396 2752
rect 5332 2692 5336 2748
rect 5336 2692 5392 2748
rect 5392 2692 5396 2748
rect 5332 2688 5396 2692
rect 5412 2748 5476 2752
rect 5412 2692 5416 2748
rect 5416 2692 5472 2748
rect 5472 2692 5476 2748
rect 5412 2688 5476 2692
rect 6897 2748 6961 2752
rect 6897 2692 6901 2748
rect 6901 2692 6957 2748
rect 6957 2692 6961 2748
rect 6897 2688 6961 2692
rect 6977 2748 7041 2752
rect 6977 2692 6981 2748
rect 6981 2692 7037 2748
rect 7037 2692 7041 2748
rect 6977 2688 7041 2692
rect 7057 2748 7121 2752
rect 7057 2692 7061 2748
rect 7061 2692 7117 2748
rect 7117 2692 7121 2748
rect 7057 2688 7121 2692
rect 7137 2748 7201 2752
rect 7137 2692 7141 2748
rect 7141 2692 7197 2748
rect 7197 2692 7201 2748
rect 7137 2688 7201 2692
rect 2584 2204 2648 2208
rect 2584 2148 2588 2204
rect 2588 2148 2644 2204
rect 2644 2148 2648 2204
rect 2584 2144 2648 2148
rect 2664 2204 2728 2208
rect 2664 2148 2668 2204
rect 2668 2148 2724 2204
rect 2724 2148 2728 2204
rect 2664 2144 2728 2148
rect 2744 2204 2808 2208
rect 2744 2148 2748 2204
rect 2748 2148 2804 2204
rect 2804 2148 2808 2204
rect 2744 2144 2808 2148
rect 2824 2204 2888 2208
rect 2824 2148 2828 2204
rect 2828 2148 2884 2204
rect 2884 2148 2888 2204
rect 2824 2144 2888 2148
rect 4309 2204 4373 2208
rect 4309 2148 4313 2204
rect 4313 2148 4369 2204
rect 4369 2148 4373 2204
rect 4309 2144 4373 2148
rect 4389 2204 4453 2208
rect 4389 2148 4393 2204
rect 4393 2148 4449 2204
rect 4449 2148 4453 2204
rect 4389 2144 4453 2148
rect 4469 2204 4533 2208
rect 4469 2148 4473 2204
rect 4473 2148 4529 2204
rect 4529 2148 4533 2204
rect 4469 2144 4533 2148
rect 4549 2204 4613 2208
rect 4549 2148 4553 2204
rect 4553 2148 4609 2204
rect 4609 2148 4613 2204
rect 4549 2144 4613 2148
rect 6034 2204 6098 2208
rect 6034 2148 6038 2204
rect 6038 2148 6094 2204
rect 6094 2148 6098 2204
rect 6034 2144 6098 2148
rect 6114 2204 6178 2208
rect 6114 2148 6118 2204
rect 6118 2148 6174 2204
rect 6174 2148 6178 2204
rect 6114 2144 6178 2148
rect 6194 2204 6258 2208
rect 6194 2148 6198 2204
rect 6198 2148 6254 2204
rect 6254 2148 6258 2204
rect 6194 2144 6258 2148
rect 6274 2204 6338 2208
rect 6274 2148 6278 2204
rect 6278 2148 6334 2204
rect 6334 2148 6338 2204
rect 6274 2144 6338 2148
rect 7759 2204 7823 2208
rect 7759 2148 7763 2204
rect 7763 2148 7819 2204
rect 7819 2148 7823 2204
rect 7759 2144 7823 2148
rect 7839 2204 7903 2208
rect 7839 2148 7843 2204
rect 7843 2148 7899 2204
rect 7899 2148 7903 2204
rect 7839 2144 7903 2148
rect 7919 2204 7983 2208
rect 7919 2148 7923 2204
rect 7923 2148 7979 2204
rect 7979 2148 7983 2204
rect 7919 2144 7983 2148
rect 7999 2204 8063 2208
rect 7999 2148 8003 2204
rect 8003 2148 8059 2204
rect 8059 2148 8063 2204
rect 7999 2144 8063 2148
rect 1722 1660 1786 1664
rect 1722 1604 1726 1660
rect 1726 1604 1782 1660
rect 1782 1604 1786 1660
rect 1722 1600 1786 1604
rect 1802 1660 1866 1664
rect 1802 1604 1806 1660
rect 1806 1604 1862 1660
rect 1862 1604 1866 1660
rect 1802 1600 1866 1604
rect 1882 1660 1946 1664
rect 1882 1604 1886 1660
rect 1886 1604 1942 1660
rect 1942 1604 1946 1660
rect 1882 1600 1946 1604
rect 1962 1660 2026 1664
rect 1962 1604 1966 1660
rect 1966 1604 2022 1660
rect 2022 1604 2026 1660
rect 1962 1600 2026 1604
rect 3447 1660 3511 1664
rect 3447 1604 3451 1660
rect 3451 1604 3507 1660
rect 3507 1604 3511 1660
rect 3447 1600 3511 1604
rect 3527 1660 3591 1664
rect 3527 1604 3531 1660
rect 3531 1604 3587 1660
rect 3587 1604 3591 1660
rect 3527 1600 3591 1604
rect 3607 1660 3671 1664
rect 3607 1604 3611 1660
rect 3611 1604 3667 1660
rect 3667 1604 3671 1660
rect 3607 1600 3671 1604
rect 3687 1660 3751 1664
rect 3687 1604 3691 1660
rect 3691 1604 3747 1660
rect 3747 1604 3751 1660
rect 3687 1600 3751 1604
rect 5172 1660 5236 1664
rect 5172 1604 5176 1660
rect 5176 1604 5232 1660
rect 5232 1604 5236 1660
rect 5172 1600 5236 1604
rect 5252 1660 5316 1664
rect 5252 1604 5256 1660
rect 5256 1604 5312 1660
rect 5312 1604 5316 1660
rect 5252 1600 5316 1604
rect 5332 1660 5396 1664
rect 5332 1604 5336 1660
rect 5336 1604 5392 1660
rect 5392 1604 5396 1660
rect 5332 1600 5396 1604
rect 5412 1660 5476 1664
rect 5412 1604 5416 1660
rect 5416 1604 5472 1660
rect 5472 1604 5476 1660
rect 5412 1600 5476 1604
rect 6897 1660 6961 1664
rect 6897 1604 6901 1660
rect 6901 1604 6957 1660
rect 6957 1604 6961 1660
rect 6897 1600 6961 1604
rect 6977 1660 7041 1664
rect 6977 1604 6981 1660
rect 6981 1604 7037 1660
rect 7037 1604 7041 1660
rect 6977 1600 7041 1604
rect 7057 1660 7121 1664
rect 7057 1604 7061 1660
rect 7061 1604 7117 1660
rect 7117 1604 7121 1660
rect 7057 1600 7121 1604
rect 7137 1660 7201 1664
rect 7137 1604 7141 1660
rect 7141 1604 7197 1660
rect 7197 1604 7201 1660
rect 7137 1600 7201 1604
rect 2584 1116 2648 1120
rect 2584 1060 2588 1116
rect 2588 1060 2644 1116
rect 2644 1060 2648 1116
rect 2584 1056 2648 1060
rect 2664 1116 2728 1120
rect 2664 1060 2668 1116
rect 2668 1060 2724 1116
rect 2724 1060 2728 1116
rect 2664 1056 2728 1060
rect 2744 1116 2808 1120
rect 2744 1060 2748 1116
rect 2748 1060 2804 1116
rect 2804 1060 2808 1116
rect 2744 1056 2808 1060
rect 2824 1116 2888 1120
rect 2824 1060 2828 1116
rect 2828 1060 2884 1116
rect 2884 1060 2888 1116
rect 2824 1056 2888 1060
rect 4309 1116 4373 1120
rect 4309 1060 4313 1116
rect 4313 1060 4369 1116
rect 4369 1060 4373 1116
rect 4309 1056 4373 1060
rect 4389 1116 4453 1120
rect 4389 1060 4393 1116
rect 4393 1060 4449 1116
rect 4449 1060 4453 1116
rect 4389 1056 4453 1060
rect 4469 1116 4533 1120
rect 4469 1060 4473 1116
rect 4473 1060 4529 1116
rect 4529 1060 4533 1116
rect 4469 1056 4533 1060
rect 4549 1116 4613 1120
rect 4549 1060 4553 1116
rect 4553 1060 4609 1116
rect 4609 1060 4613 1116
rect 4549 1056 4613 1060
rect 6034 1116 6098 1120
rect 6034 1060 6038 1116
rect 6038 1060 6094 1116
rect 6094 1060 6098 1116
rect 6034 1056 6098 1060
rect 6114 1116 6178 1120
rect 6114 1060 6118 1116
rect 6118 1060 6174 1116
rect 6174 1060 6178 1116
rect 6114 1056 6178 1060
rect 6194 1116 6258 1120
rect 6194 1060 6198 1116
rect 6198 1060 6254 1116
rect 6254 1060 6258 1116
rect 6194 1056 6258 1060
rect 6274 1116 6338 1120
rect 6274 1060 6278 1116
rect 6278 1060 6334 1116
rect 6334 1060 6338 1116
rect 6274 1056 6338 1060
rect 7759 1116 7823 1120
rect 7759 1060 7763 1116
rect 7763 1060 7819 1116
rect 7819 1060 7823 1116
rect 7759 1056 7823 1060
rect 7839 1116 7903 1120
rect 7839 1060 7843 1116
rect 7843 1060 7899 1116
rect 7899 1060 7903 1116
rect 7839 1056 7903 1060
rect 7919 1116 7983 1120
rect 7919 1060 7923 1116
rect 7923 1060 7979 1116
rect 7979 1060 7983 1116
rect 7919 1056 7983 1060
rect 7999 1116 8063 1120
rect 7999 1060 8003 1116
rect 8003 1060 8059 1116
rect 8059 1060 8063 1116
rect 7999 1056 8063 1060
<< metal4 >>
rect 1714 8192 2034 8752
rect 1714 8128 1722 8192
rect 1786 8128 1802 8192
rect 1866 8128 1882 8192
rect 1946 8128 1962 8192
rect 2026 8128 2034 8192
rect 1714 7104 2034 8128
rect 1714 7040 1722 7104
rect 1786 7040 1802 7104
rect 1866 7040 1882 7104
rect 1946 7040 1962 7104
rect 2026 7040 2034 7104
rect 1714 6016 2034 7040
rect 1714 5952 1722 6016
rect 1786 5952 1802 6016
rect 1866 5952 1882 6016
rect 1946 5952 1962 6016
rect 2026 5952 2034 6016
rect 1714 4928 2034 5952
rect 1714 4864 1722 4928
rect 1786 4864 1802 4928
rect 1866 4864 1882 4928
rect 1946 4864 1962 4928
rect 2026 4864 2034 4928
rect 1714 3840 2034 4864
rect 1714 3776 1722 3840
rect 1786 3776 1802 3840
rect 1866 3776 1882 3840
rect 1946 3776 1962 3840
rect 2026 3776 2034 3840
rect 1714 2752 2034 3776
rect 1714 2688 1722 2752
rect 1786 2688 1802 2752
rect 1866 2688 1882 2752
rect 1946 2688 1962 2752
rect 2026 2688 2034 2752
rect 1714 1664 2034 2688
rect 1714 1600 1722 1664
rect 1786 1600 1802 1664
rect 1866 1600 1882 1664
rect 1946 1600 1962 1664
rect 2026 1600 2034 1664
rect 1714 1040 2034 1600
rect 2576 8736 2896 8752
rect 2576 8672 2584 8736
rect 2648 8672 2664 8736
rect 2728 8672 2744 8736
rect 2808 8672 2824 8736
rect 2888 8672 2896 8736
rect 2576 7648 2896 8672
rect 2576 7584 2584 7648
rect 2648 7584 2664 7648
rect 2728 7584 2744 7648
rect 2808 7584 2824 7648
rect 2888 7584 2896 7648
rect 2576 6560 2896 7584
rect 2576 6496 2584 6560
rect 2648 6496 2664 6560
rect 2728 6496 2744 6560
rect 2808 6496 2824 6560
rect 2888 6496 2896 6560
rect 2576 5472 2896 6496
rect 2576 5408 2584 5472
rect 2648 5408 2664 5472
rect 2728 5408 2744 5472
rect 2808 5408 2824 5472
rect 2888 5408 2896 5472
rect 2576 4384 2896 5408
rect 2576 4320 2584 4384
rect 2648 4320 2664 4384
rect 2728 4320 2744 4384
rect 2808 4320 2824 4384
rect 2888 4320 2896 4384
rect 2576 3296 2896 4320
rect 2576 3232 2584 3296
rect 2648 3232 2664 3296
rect 2728 3232 2744 3296
rect 2808 3232 2824 3296
rect 2888 3232 2896 3296
rect 2576 2208 2896 3232
rect 2576 2144 2584 2208
rect 2648 2144 2664 2208
rect 2728 2144 2744 2208
rect 2808 2144 2824 2208
rect 2888 2144 2896 2208
rect 2576 1120 2896 2144
rect 2576 1056 2584 1120
rect 2648 1056 2664 1120
rect 2728 1056 2744 1120
rect 2808 1056 2824 1120
rect 2888 1056 2896 1120
rect 2576 1040 2896 1056
rect 3439 8192 3759 8752
rect 3439 8128 3447 8192
rect 3511 8128 3527 8192
rect 3591 8128 3607 8192
rect 3671 8128 3687 8192
rect 3751 8128 3759 8192
rect 3439 7104 3759 8128
rect 3439 7040 3447 7104
rect 3511 7040 3527 7104
rect 3591 7040 3607 7104
rect 3671 7040 3687 7104
rect 3751 7040 3759 7104
rect 3439 6016 3759 7040
rect 3439 5952 3447 6016
rect 3511 5952 3527 6016
rect 3591 5952 3607 6016
rect 3671 5952 3687 6016
rect 3751 5952 3759 6016
rect 3439 4928 3759 5952
rect 3439 4864 3447 4928
rect 3511 4864 3527 4928
rect 3591 4864 3607 4928
rect 3671 4864 3687 4928
rect 3751 4864 3759 4928
rect 3439 3840 3759 4864
rect 3439 3776 3447 3840
rect 3511 3776 3527 3840
rect 3591 3776 3607 3840
rect 3671 3776 3687 3840
rect 3751 3776 3759 3840
rect 3439 2752 3759 3776
rect 3439 2688 3447 2752
rect 3511 2688 3527 2752
rect 3591 2688 3607 2752
rect 3671 2688 3687 2752
rect 3751 2688 3759 2752
rect 3439 1664 3759 2688
rect 3439 1600 3447 1664
rect 3511 1600 3527 1664
rect 3591 1600 3607 1664
rect 3671 1600 3687 1664
rect 3751 1600 3759 1664
rect 3439 1040 3759 1600
rect 4301 8736 4621 8752
rect 4301 8672 4309 8736
rect 4373 8672 4389 8736
rect 4453 8672 4469 8736
rect 4533 8672 4549 8736
rect 4613 8672 4621 8736
rect 4301 7648 4621 8672
rect 4301 7584 4309 7648
rect 4373 7584 4389 7648
rect 4453 7584 4469 7648
rect 4533 7584 4549 7648
rect 4613 7584 4621 7648
rect 4301 6560 4621 7584
rect 4301 6496 4309 6560
rect 4373 6496 4389 6560
rect 4453 6496 4469 6560
rect 4533 6496 4549 6560
rect 4613 6496 4621 6560
rect 4301 5472 4621 6496
rect 4301 5408 4309 5472
rect 4373 5408 4389 5472
rect 4453 5408 4469 5472
rect 4533 5408 4549 5472
rect 4613 5408 4621 5472
rect 4301 4384 4621 5408
rect 4301 4320 4309 4384
rect 4373 4320 4389 4384
rect 4453 4320 4469 4384
rect 4533 4320 4549 4384
rect 4613 4320 4621 4384
rect 4301 3296 4621 4320
rect 4301 3232 4309 3296
rect 4373 3232 4389 3296
rect 4453 3232 4469 3296
rect 4533 3232 4549 3296
rect 4613 3232 4621 3296
rect 4301 2208 4621 3232
rect 4301 2144 4309 2208
rect 4373 2144 4389 2208
rect 4453 2144 4469 2208
rect 4533 2144 4549 2208
rect 4613 2144 4621 2208
rect 4301 1120 4621 2144
rect 4301 1056 4309 1120
rect 4373 1056 4389 1120
rect 4453 1056 4469 1120
rect 4533 1056 4549 1120
rect 4613 1056 4621 1120
rect 4301 1040 4621 1056
rect 5164 8192 5484 8752
rect 5164 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5484 8192
rect 5164 7104 5484 8128
rect 5164 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5484 7104
rect 5164 6016 5484 7040
rect 5164 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5484 6016
rect 5164 4928 5484 5952
rect 5164 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5484 4928
rect 5164 3840 5484 4864
rect 5164 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5484 3840
rect 5164 2752 5484 3776
rect 5164 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5484 2752
rect 5164 1664 5484 2688
rect 5164 1600 5172 1664
rect 5236 1600 5252 1664
rect 5316 1600 5332 1664
rect 5396 1600 5412 1664
rect 5476 1600 5484 1664
rect 5164 1040 5484 1600
rect 6026 8736 6346 8752
rect 6026 8672 6034 8736
rect 6098 8672 6114 8736
rect 6178 8672 6194 8736
rect 6258 8672 6274 8736
rect 6338 8672 6346 8736
rect 6026 7648 6346 8672
rect 6026 7584 6034 7648
rect 6098 7584 6114 7648
rect 6178 7584 6194 7648
rect 6258 7584 6274 7648
rect 6338 7584 6346 7648
rect 6026 6560 6346 7584
rect 6026 6496 6034 6560
rect 6098 6496 6114 6560
rect 6178 6496 6194 6560
rect 6258 6496 6274 6560
rect 6338 6496 6346 6560
rect 6026 5472 6346 6496
rect 6026 5408 6034 5472
rect 6098 5408 6114 5472
rect 6178 5408 6194 5472
rect 6258 5408 6274 5472
rect 6338 5408 6346 5472
rect 6026 4384 6346 5408
rect 6026 4320 6034 4384
rect 6098 4320 6114 4384
rect 6178 4320 6194 4384
rect 6258 4320 6274 4384
rect 6338 4320 6346 4384
rect 6026 3296 6346 4320
rect 6026 3232 6034 3296
rect 6098 3232 6114 3296
rect 6178 3232 6194 3296
rect 6258 3232 6274 3296
rect 6338 3232 6346 3296
rect 6026 2208 6346 3232
rect 6026 2144 6034 2208
rect 6098 2144 6114 2208
rect 6178 2144 6194 2208
rect 6258 2144 6274 2208
rect 6338 2144 6346 2208
rect 6026 1120 6346 2144
rect 6026 1056 6034 1120
rect 6098 1056 6114 1120
rect 6178 1056 6194 1120
rect 6258 1056 6274 1120
rect 6338 1056 6346 1120
rect 6026 1040 6346 1056
rect 6889 8192 7209 8752
rect 6889 8128 6897 8192
rect 6961 8128 6977 8192
rect 7041 8128 7057 8192
rect 7121 8128 7137 8192
rect 7201 8128 7209 8192
rect 6889 7104 7209 8128
rect 6889 7040 6897 7104
rect 6961 7040 6977 7104
rect 7041 7040 7057 7104
rect 7121 7040 7137 7104
rect 7201 7040 7209 7104
rect 6889 6016 7209 7040
rect 6889 5952 6897 6016
rect 6961 5952 6977 6016
rect 7041 5952 7057 6016
rect 7121 5952 7137 6016
rect 7201 5952 7209 6016
rect 6889 4928 7209 5952
rect 6889 4864 6897 4928
rect 6961 4864 6977 4928
rect 7041 4864 7057 4928
rect 7121 4864 7137 4928
rect 7201 4864 7209 4928
rect 6889 3840 7209 4864
rect 6889 3776 6897 3840
rect 6961 3776 6977 3840
rect 7041 3776 7057 3840
rect 7121 3776 7137 3840
rect 7201 3776 7209 3840
rect 6889 2752 7209 3776
rect 6889 2688 6897 2752
rect 6961 2688 6977 2752
rect 7041 2688 7057 2752
rect 7121 2688 7137 2752
rect 7201 2688 7209 2752
rect 6889 1664 7209 2688
rect 6889 1600 6897 1664
rect 6961 1600 6977 1664
rect 7041 1600 7057 1664
rect 7121 1600 7137 1664
rect 7201 1600 7209 1664
rect 6889 1040 7209 1600
rect 7751 8736 8071 8752
rect 7751 8672 7759 8736
rect 7823 8672 7839 8736
rect 7903 8672 7919 8736
rect 7983 8672 7999 8736
rect 8063 8672 8071 8736
rect 7751 7648 8071 8672
rect 7751 7584 7759 7648
rect 7823 7584 7839 7648
rect 7903 7584 7919 7648
rect 7983 7584 7999 7648
rect 8063 7584 8071 7648
rect 7751 6560 8071 7584
rect 7751 6496 7759 6560
rect 7823 6496 7839 6560
rect 7903 6496 7919 6560
rect 7983 6496 7999 6560
rect 8063 6496 8071 6560
rect 7751 5472 8071 6496
rect 7751 5408 7759 5472
rect 7823 5408 7839 5472
rect 7903 5408 7919 5472
rect 7983 5408 7999 5472
rect 8063 5408 8071 5472
rect 7751 4384 8071 5408
rect 7751 4320 7759 4384
rect 7823 4320 7839 4384
rect 7903 4320 7919 4384
rect 7983 4320 7999 4384
rect 8063 4320 8071 4384
rect 7751 3296 8071 4320
rect 7751 3232 7759 3296
rect 7823 3232 7839 3296
rect 7903 3232 7919 3296
rect 7983 3232 7999 3296
rect 8063 3232 8071 3296
rect 7751 2208 8071 3232
rect 7751 2144 7759 2208
rect 7823 2144 7839 2208
rect 7903 2144 7919 2208
rect 7983 2144 7999 2208
rect 8063 2144 8071 2208
rect 7751 1120 8071 2144
rect 7751 1056 7759 1120
rect 7823 1056 7839 1120
rect 7903 1056 7919 1120
rect 7983 1056 7999 1120
rect 8063 1056 8071 1120
rect 7751 1040 8071 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[0\]_A swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[1\]_A
timestamp 1673029049
transform 1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[2\]_A
timestamp 1673029049
transform -1 0 5520 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[3\]_A
timestamp 1673029049
transform -1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[4\]_A
timestamp 1673029049
transform -1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[5\]_A
timestamp 1673029049
transform -1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[6\]_A
timestamp 1673029049
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[7\]_A
timestamp 1673029049
transform -1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[8\]_A
timestamp 1673029049
transform -1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[9\]_A
timestamp 1673029049
transform -1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[10\]_A
timestamp 1673029049
transform -1 0 5428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[11\]_A
timestamp 1673029049
transform -1 0 6072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[12\]_A
timestamp 1673029049
transform -1 0 2576 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[13\]_A
timestamp 1673029049
transform 1 0 5888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[14\]_A
timestamp 1673029049
transform -1 0 5980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[15\]_A
timestamp 1673029049
transform -1 0 6072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[16\]_A
timestamp 1673029049
transform -1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[17\]_A
timestamp 1673029049
transform -1 0 1840 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[18\]_A
timestamp 1673029049
transform -1 0 3404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[19\]_A
timestamp 1673029049
transform -1 0 2024 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[20\]_A
timestamp 1673029049
transform -1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[21\]_A
timestamp 1673029049
transform -1 0 2024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[22\]_A
timestamp 1673029049
transform -1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[23\]_A
timestamp 1673029049
transform -1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[24\]_A
timestamp 1673029049
transform -1 0 4876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[25\]_A
timestamp 1673029049
transform -1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[26\]_A
timestamp 1673029049
transform -1 0 5520 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[27\]_A
timestamp 1673029049
transform 1 0 5336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[28\]_A
timestamp 1673029049
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[29\]_A
timestamp 1673029049
transform -1 0 7268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[30\]_A
timestamp 1673029049
transform -1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[31\]_A
timestamp 1673029049
transform -1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[32\]_A
timestamp 1673029049
transform -1 0 4232 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[33\]_A
timestamp 1673029049
transform -1 0 1840 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[34\]_A
timestamp 1673029049
transform -1 0 1840 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[35\]_A
timestamp 1673029049
transform -1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[36\]_A
timestamp 1673029049
transform -1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[37\]_A
timestamp 1673029049
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[38\]_A
timestamp 1673029049
transform -1 0 3404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[39\]_A
timestamp 1673029049
transform 1 0 2208 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[40\]_A
timestamp 1673029049
transform -1 0 4784 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[0\] swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1472 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[1\]
timestamp 1673029049
transform 1 0 6440 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[2\]
timestamp 1673029049
transform 1 0 4600 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[3\]
timestamp 1673029049
transform 1 0 3864 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[4\]
timestamp 1673029049
transform 1 0 3864 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[5\]
timestamp 1673029049
transform 1 0 3864 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[6\]
timestamp 1673029049
transform 1 0 3588 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[7\]
timestamp 1673029049
transform 1 0 3588 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[8\]
timestamp 1673029049
transform 1 0 2392 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[9\]
timestamp 1673029049
transform -1 0 4508 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[10\]
timestamp 1673029049
transform -1 0 4876 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[11\]
timestamp 1673029049
transform -1 0 5888 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[12\]
timestamp 1673029049
transform -1 0 4232 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[13\]
timestamp 1673029049
transform -1 0 5980 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[14\]
timestamp 1673029049
transform 1 0 6440 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[15\]
timestamp 1673029049
transform -1 0 7452 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[16\]
timestamp 1673029049
transform -1 0 7452 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[17\]
timestamp 1673029049
transform -1 0 5980 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[18\]
timestamp 1673029049
transform -1 0 3404 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[19\]
timestamp 1673029049
transform -1 0 4968 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[20\]
timestamp 1673029049
transform -1 0 3404 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[21\]
timestamp 1673029049
transform -1 0 3404 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[22\]
timestamp 1673029049
transform 1 0 6440 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[23\]
timestamp 1673029049
transform 1 0 6440 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[24\]
timestamp 1673029049
transform 1 0 6440 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[25\]
timestamp 1673029049
transform 1 0 6440 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[26\]
timestamp 1673029049
transform 1 0 6440 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[27\]
timestamp 1673029049
transform 1 0 6440 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[28\]
timestamp 1673029049
transform 1 0 6440 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[29\]
timestamp 1673029049
transform 1 0 6440 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[30\]
timestamp 1673029049
transform 1 0 6440 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[31\]
timestamp 1673029049
transform 1 0 5704 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[32\]
timestamp 1673029049
transform 1 0 3864 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[33\]
timestamp 1673029049
transform 1 0 2208 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[34\]
timestamp 1673029049
transform 1 0 1840 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[35\]
timestamp 1673029049
transform 1 0 3864 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[36\]
timestamp 1673029049
transform 1 0 1748 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[37\]
timestamp 1673029049
transform 1 0 2668 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[38\]
timestamp 1673029049
transform 1 0 4048 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[39\]
timestamp 1673029049
transform 1 0 2760 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[40\]
timestamp 1673029049
transform 1 0 2208 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1288 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2024 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3404 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3680 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43
timestamp 1673029049
transform 1 0 4968 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1673029049
transform 1 0 5520 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6072 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1673029049
transform 1 0 6256 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1673029049
transform 1 0 7452 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1673029049
transform 1 0 1288 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1673029049
transform 1 0 1840 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1673029049
transform 1 0 3220 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1673029049
transform 1 0 4600 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1673029049
transform 1 0 5980 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1673029049
transform 1 0 6256 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 1673029049
transform 1 0 7452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1673029049
transform 1 0 1288 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1673029049
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1673029049
transform 1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1673029049
transform 1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1673029049
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46
timestamp 1673029049
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_49
timestamp 1673029049
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1673029049
transform 1 0 6072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 1673029049
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1673029049
transform 1 0 1288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_16 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1673029049
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1673029049
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1673029049
transform 1 0 6256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1673029049
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1673029049
transform 1 0 1288 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1673029049
transform 1 0 2024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1673029049
transform 1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1673029049
transform 1 0 3680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_42
timestamp 1673029049
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_46
timestamp 1673029049
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_49
timestamp 1673029049
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_55
timestamp 1673029049
transform 1 0 6072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1673029049
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1673029049
transform 1 0 1288 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1673029049
transform 1 0 2024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1673029049
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1673029049
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1673029049
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1673029049
transform 1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1673029049
transform 1 0 6256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_70
timestamp 1673029049
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1673029049
transform 1 0 1288 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1673029049
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1673029049
transform 1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1673029049
transform 1 0 3680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1673029049
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1673029049
transform 1 0 5244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_49
timestamp 1673029049
transform 1 0 5520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1673029049
transform 1 0 6072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_70
timestamp 1673029049
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1673029049
transform 1 0 1288 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1673029049
transform 1 0 1840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1673029049
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1673029049
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 1673029049
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1673029049
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1673029049
transform 1 0 5980 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1673029049
transform 1 0 6256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_70
timestamp 1673029049
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1673029049
transform 1 0 1288 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1673029049
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp 1673029049
transform 1 0 2024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1673029049
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_20
timestamp 1673029049
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1673029049
transform 1 0 3404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1673029049
transform 1 0 3680 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_42
timestamp 1673029049
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1673029049
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_52
timestamp 1673029049
transform 1 0 5796 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_55
timestamp 1673029049
transform 1 0 6072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp 1673029049
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1673029049
transform 1 0 1288 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1673029049
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1673029049
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1673029049
transform 1 0 3772 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_36
timestamp 1673029049
transform 1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_42
timestamp 1673029049
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_48
timestamp 1673029049
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1673029049
transform 1 0 5980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1673029049
transform 1 0 6256 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1673029049
transform 1 0 7452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1673029049
transform 1 0 1288 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_20
timestamp 1673029049
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1673029049
transform 1 0 3404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1673029049
transform 1 0 3680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_44
timestamp 1673029049
transform 1 0 5060 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_52
timestamp 1673029049
transform 1 0 5796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 1673029049
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1673029049
transform 1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1673029049
transform 1 0 1288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_8
timestamp 1673029049
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1673029049
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_29
timestamp 1673029049
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1673029049
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_41
timestamp 1673029049
transform 1 0 4784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1673029049
transform 1 0 5704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1673029049
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1673029049
transform 1 0 6256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1673029049
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1673029049
transform 1 0 1288 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1673029049
transform 1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1673029049
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1673029049
transform 1 0 3680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_42
timestamp 1673029049
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_50
timestamp 1673029049
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1673029049
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_68
timestamp 1673029049
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1673029049
transform 1 0 1288 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1673029049
transform 1 0 1656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1673029049
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_23
timestamp 1673029049
transform 1 0 3128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1673029049
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1673029049
transform 1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_42
timestamp 1673029049
transform 1 0 4876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1673029049
transform 1 0 5612 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1673029049
transform 1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1673029049
transform 1 0 6256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1673029049
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 1012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 1012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 7912 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 1012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 1012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 1012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1673029049
transform 1 0 1012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1673029049
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1673029049
transform 1 0 1012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1673029049
transform -1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1673029049
transform 1 0 1012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1673029049
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1673029049
transform 1 0 1012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1673029049
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1673029049
transform 1 0 1012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1673029049
transform -1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1673029049
transform 1 0 1012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1673029049
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1673029049
transform 1 0 1012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1673029049
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1673029049
transform 1 0 1012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1673029049
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1673029049
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1673029049
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1673029049
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1673029049
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1673029049
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1673029049
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1673029049
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1673029049
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1673029049
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1673029049
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1673029049
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1673029049
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1673029049
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1673029049
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1673029049
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 2576 1040 2896 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4301 1040 4621 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6026 1040 6346 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7751 1040 8071 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1714 1040 2034 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3439 1040 3759 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5164 1040 5484 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6889 1040 7209 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 7930 9200 7986 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[0]
port 2 nsew signal input
flabel metal2 s 2410 9200 2466 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[10]
port 3 nsew signal input
flabel metal2 s 1858 9200 1914 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[11]
port 4 nsew signal input
flabel metal2 s 1306 9200 1362 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[12]
port 5 nsew signal input
flabel metal2 s 754 9200 810 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[13]
port 6 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 mgmt_gpio_in[14]
port 7 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 mgmt_gpio_in[15]
port 8 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 mgmt_gpio_in[16]
port 9 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 mgmt_gpio_in[17]
port 10 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 mgmt_gpio_in[18]
port 11 nsew signal input
flabel metal2 s 7378 9200 7434 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[1]
port 12 nsew signal input
flabel metal2 s 6826 9200 6882 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[2]
port 13 nsew signal input
flabel metal2 s 6274 9200 6330 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[3]
port 14 nsew signal input
flabel metal2 s 5722 9200 5778 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[4]
port 15 nsew signal input
flabel metal2 s 5170 9200 5226 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[5]
port 16 nsew signal input
flabel metal2 s 4618 9200 4674 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[6]
port 17 nsew signal input
flabel metal2 s 4066 9200 4122 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[7]
port 18 nsew signal input
flabel metal2 s 3514 9200 3570 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[8]
port 19 nsew signal input
flabel metal2 s 2962 9200 3018 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[9]
port 20 nsew signal input
flabel metal3 s 8200 1776 9000 1896 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[0]
port 21 nsew signal tristate
flabel metal3 s 8200 5856 9000 5976 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[10]
port 22 nsew signal tristate
flabel metal3 s 8200 6264 9000 6384 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[11]
port 23 nsew signal tristate
flabel metal3 s 8200 6672 9000 6792 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[12]
port 24 nsew signal tristate
flabel metal3 s 8200 7080 9000 7200 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[13]
port 25 nsew signal tristate
flabel metal3 s 8200 7488 9000 7608 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[14]
port 26 nsew signal tristate
flabel metal3 s 8200 7896 9000 8016 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[15]
port 27 nsew signal tristate
flabel metal3 s 8200 8304 9000 8424 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[16]
port 28 nsew signal tristate
flabel metal3 s 8200 8712 9000 8832 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[17]
port 29 nsew signal tristate
flabel metal3 s 8200 9120 9000 9240 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[18]
port 30 nsew signal tristate
flabel metal3 s 8200 2184 9000 2304 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[1]
port 31 nsew signal tristate
flabel metal3 s 8200 2592 9000 2712 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[2]
port 32 nsew signal tristate
flabel metal3 s 8200 3000 9000 3120 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[3]
port 33 nsew signal tristate
flabel metal3 s 8200 3408 9000 3528 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[4]
port 34 nsew signal tristate
flabel metal3 s 8200 3816 9000 3936 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[5]
port 35 nsew signal tristate
flabel metal3 s 8200 4224 9000 4344 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[6]
port 36 nsew signal tristate
flabel metal3 s 8200 4632 9000 4752 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[7]
port 37 nsew signal tristate
flabel metal3 s 8200 5040 9000 5160 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[8]
port 38 nsew signal tristate
flabel metal3 s 8200 5448 9000 5568 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[9]
port 39 nsew signal tristate
flabel metal3 s 8200 552 9000 672 0 FreeSans 480 0 0 0 mgmt_gpio_oeb[0]
port 40 nsew signal input
flabel metal3 s 8200 960 9000 1080 0 FreeSans 480 0 0 0 mgmt_gpio_oeb[1]
port 41 nsew signal input
flabel metal3 s 8200 1368 9000 1488 0 FreeSans 480 0 0 0 mgmt_gpio_oeb[2]
port 42 nsew signal input
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 mgmt_gpio_oeb_buf[0]
port 43 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 mgmt_gpio_oeb_buf[1]
port 44 nsew signal tristate
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 mgmt_gpio_oeb_buf[2]
port 45 nsew signal tristate
flabel metal2 s 294 0 350 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[0]
port 46 nsew signal input
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[10]
port 47 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[11]
port 48 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[12]
port 49 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[13]
port 50 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[14]
port 51 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[15]
port 52 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[16]
port 53 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[17]
port 54 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[18]
port 55 nsew signal input
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[1]
port 56 nsew signal input
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[2]
port 57 nsew signal input
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[3]
port 58 nsew signal input
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[4]
port 59 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[5]
port 60 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[6]
port 61 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[7]
port 62 nsew signal input
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[8]
port 63 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[9]
port 64 nsew signal input
flabel metal2 s 8206 9200 8262 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[0]
port 65 nsew signal tristate
flabel metal2 s 2686 9200 2742 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[10]
port 66 nsew signal tristate
flabel metal2 s 2134 9200 2190 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[11]
port 67 nsew signal tristate
flabel metal2 s 1582 9200 1638 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[12]
port 68 nsew signal tristate
flabel metal2 s 1030 9200 1086 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[13]
port 69 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[14]
port 70 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[15]
port 71 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[16]
port 72 nsew signal tristate
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[17]
port 73 nsew signal tristate
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[18]
port 74 nsew signal tristate
flabel metal2 s 7654 9200 7710 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[1]
port 75 nsew signal tristate
flabel metal2 s 7102 9200 7158 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[2]
port 76 nsew signal tristate
flabel metal2 s 6550 9200 6606 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[3]
port 77 nsew signal tristate
flabel metal2 s 5998 9200 6054 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[4]
port 78 nsew signal tristate
flabel metal2 s 5446 9200 5502 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[5]
port 79 nsew signal tristate
flabel metal2 s 4894 9200 4950 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[6]
port 80 nsew signal tristate
flabel metal2 s 4342 9200 4398 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[7]
port 81 nsew signal tristate
flabel metal2 s 3790 9200 3846 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[8]
port 82 nsew signal tristate
flabel metal2 s 3238 9200 3294 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[9]
port 83 nsew signal tristate
rlabel via1 4541 8704 4541 8704 0 VGND
rlabel metal1 4462 8160 4462 8160 0 VPWR
rlabel metal2 4922 4658 4922 4658 0 mgmt_gpio_in[0]
rlabel metal1 3174 7854 3174 7854 0 mgmt_gpio_in[10]
rlabel metal1 1932 8058 1932 8058 0 mgmt_gpio_in[11]
rlabel metal1 1610 6766 1610 6766 0 mgmt_gpio_in[12]
rlabel metal1 2116 8602 2116 8602 0 mgmt_gpio_in[13]
rlabel metal2 1794 8415 1794 8415 0 mgmt_gpio_in[14]
rlabel metal1 1840 7242 1840 7242 0 mgmt_gpio_in[15]
rlabel metal1 3174 6630 3174 6630 0 mgmt_gpio_in[16]
rlabel metal1 2668 6086 2668 6086 0 mgmt_gpio_in[17]
rlabel metal1 2254 1904 2254 1904 0 mgmt_gpio_in[18]
rlabel metal2 6394 5865 6394 5865 0 mgmt_gpio_in[1]
rlabel metal1 5382 6086 5382 6086 0 mgmt_gpio_in[2]
rlabel metal2 6486 3825 6486 3825 0 mgmt_gpio_in[3]
rlabel metal1 6118 4182 6118 4182 0 mgmt_gpio_in[4]
rlabel metal1 5060 4794 5060 4794 0 mgmt_gpio_in[5]
rlabel metal1 5796 5882 5796 5882 0 mgmt_gpio_in[6]
rlabel metal1 5244 7378 5244 7378 0 mgmt_gpio_in[7]
rlabel metal1 4784 8602 4784 8602 0 mgmt_gpio_in[8]
rlabel metal1 5244 7854 5244 7854 0 mgmt_gpio_in[9]
rlabel metal2 7314 1581 7314 1581 0 mgmt_gpio_in_buf[0]
rlabel metal1 4784 7786 4784 7786 0 mgmt_gpio_in_buf[10]
rlabel metal2 5474 6612 5474 6612 0 mgmt_gpio_in_buf[11]
rlabel via2 4554 6749 4554 6749 0 mgmt_gpio_in_buf[12]
rlabel metal2 5474 7616 5474 7616 0 mgmt_gpio_in_buf[13]
rlabel metal2 4646 8109 4646 8109 0 mgmt_gpio_in_buf[14]
rlabel metal1 4140 7446 4140 7446 0 mgmt_gpio_in_buf[15]
rlabel metal1 5014 6834 5014 6834 0 mgmt_gpio_in_buf[16]
rlabel metal1 3772 6358 3772 6358 0 mgmt_gpio_in_buf[17]
rlabel metal1 4048 1938 4048 1938 0 mgmt_gpio_in_buf[18]
rlabel metal2 7314 2193 7314 2193 0 mgmt_gpio_in_buf[1]
rlabel metal2 7314 2567 7314 2567 0 mgmt_gpio_in_buf[2]
rlabel via2 7314 3043 7314 3043 0 mgmt_gpio_in_buf[3]
rlabel metal2 7314 3757 7314 3757 0 mgmt_gpio_in_buf[4]
rlabel metal2 6854 4267 6854 4267 0 mgmt_gpio_in_buf[5]
rlabel metal2 7314 4879 7314 4879 0 mgmt_gpio_in_buf[6]
rlabel metal3 7874 4692 7874 4692 0 mgmt_gpio_in_buf[7]
rlabel metal3 7920 5100 7920 5100 0 mgmt_gpio_in_buf[8]
rlabel metal2 6578 6647 6578 6647 0 mgmt_gpio_in_buf[9]
rlabel metal1 3450 1326 3450 1326 0 mgmt_gpio_oeb[0]
rlabel metal1 2806 1258 2806 1258 0 mgmt_gpio_oeb[1]
rlabel metal1 4416 3502 4416 3502 0 mgmt_gpio_oeb[2]
rlabel metal3 1395 4284 1395 4284 0 mgmt_gpio_oeb_buf[0]
rlabel metal3 1027 2244 1027 2244 0 mgmt_gpio_oeb_buf[1]
rlabel metal3 1832 884 1832 884 0 mgmt_gpio_oeb_buf[2]
rlabel metal1 920 3026 920 3026 0 mgmt_gpio_out[0]
rlabel metal2 4830 4675 4830 4675 0 mgmt_gpio_out[10]
rlabel metal1 5566 3366 5566 3366 0 mgmt_gpio_out[11]
rlabel metal1 5014 3094 5014 3094 0 mgmt_gpio_out[12]
rlabel metal1 6210 4454 6210 4454 0 mgmt_gpio_out[13]
rlabel metal1 6624 6290 6624 6290 0 mgmt_gpio_out[14]
rlabel metal2 8234 4114 8234 4114 0 mgmt_gpio_out[15]
rlabel metal1 7452 5202 7452 5202 0 mgmt_gpio_out[16]
rlabel metal1 5934 2040 5934 2040 0 mgmt_gpio_out[17]
rlabel metal1 3312 2414 3312 2414 0 mgmt_gpio_out[18]
rlabel metal2 6026 2686 6026 2686 0 mgmt_gpio_out[1]
rlabel metal1 3312 1190 3312 1190 0 mgmt_gpio_out[2]
rlabel metal1 1748 4454 1748 4454 0 mgmt_gpio_out[3]
rlabel metal1 2070 2278 2070 2278 0 mgmt_gpio_out[4]
rlabel metal1 2254 3366 2254 3366 0 mgmt_gpio_out[5]
rlabel metal2 3082 2880 3082 2880 0 mgmt_gpio_out[6]
rlabel metal1 3404 2006 3404 2006 0 mgmt_gpio_out[7]
rlabel metal1 3220 4590 3220 4590 0 mgmt_gpio_out[8]
rlabel metal1 4600 4182 4600 4182 0 mgmt_gpio_out[9]
rlabel metal1 2346 3128 2346 3128 0 mgmt_gpio_out_buf[0]
rlabel metal1 3266 5746 3266 5746 0 mgmt_gpio_out_buf[10]
rlabel metal1 3818 5678 3818 5678 0 mgmt_gpio_out_buf[11]
rlabel metal1 2392 5610 2392 5610 0 mgmt_gpio_out_buf[12]
rlabel metal1 3128 5882 3128 5882 0 mgmt_gpio_out_buf[13]
rlabel metal3 2062 9044 2062 9044 0 mgmt_gpio_out_buf[14]
rlabel metal3 1579 7684 1579 7684 0 mgmt_gpio_out_buf[15]
rlabel metal3 1832 6324 1832 6324 0 mgmt_gpio_out_buf[16]
rlabel metal3 1119 4964 1119 4964 0 mgmt_gpio_out_buf[17]
rlabel metal3 1740 2924 1740 2924 0 mgmt_gpio_out_buf[18]
rlabel metal1 7498 3570 7498 3570 0 mgmt_gpio_out_buf[1]
rlabel metal2 7590 4352 7590 4352 0 mgmt_gpio_out_buf[2]
rlabel metal1 5704 4522 5704 4522 0 mgmt_gpio_out_buf[3]
rlabel metal1 5336 2482 5336 2482 0 mgmt_gpio_out_buf[4]
rlabel metal1 4876 3570 4876 3570 0 mgmt_gpio_out_buf[5]
rlabel metal1 4692 5270 4692 5270 0 mgmt_gpio_out_buf[6]
rlabel metal1 4278 2006 4278 2006 0 mgmt_gpio_out_buf[7]
rlabel metal1 3542 4658 3542 4658 0 mgmt_gpio_out_buf[8]
rlabel metal1 3450 4114 3450 4114 0 mgmt_gpio_out_buf[9]
<< properties >>
string FIXED_BBOX 0 0 9000 10000
<< end >>
