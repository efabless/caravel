VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_core
  CLASS BLOCK ;
  FOREIGN caravel_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 3165.000 BY 4767.000 ;
  PIN clock_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.135 -2.000 725.415 4.000 ;
    END
  END clock_core
  PIN flash_clk_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.335 -2.000 1597.615 4.000 ;
    END
  END flash_clk_frame
  PIN flash_clk_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.975 -2.000 1613.255 4.000 ;
    END
  END flash_clk_oeb
  PIN flash_csb_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.335 -2.000 1323.615 4.000 ;
    END
  END flash_csb_frame
  PIN flash_csb_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.975 -2.000 1339.255 4.000 ;
    END
  END flash_csb_oeb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.135 -2.000 1816.415 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.335 -2.000 1871.615 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.715 -2.000 1849.995 4.000 ;
    END
  END flash_io0_ieb
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.975 -2.000 1887.255 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.135 -2.000 2090.415 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.335 -2.000 2145.615 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2123.715 -2.000 2123.995 4.000 ;
    END
  END flash_io1_ieb
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.975 -2.000 2161.255 4.000 ;
    END
  END flash_io1_oeb
  PIN gpio_in_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.135 -2.000 2364.415 4.000 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2397.715 -2.000 2397.995 4.000 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2391.735 -2.000 2392.015 4.000 ;
    END
  END gpio_mode0_core
  PIN gpio_mode1_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.355 -2.000 2413.635 4.000 ;
    END
  END gpio_mode1_core
  PIN gpio_out_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.335 -2.000 2419.615 4.000 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.975 -2.000 2435.255 4.000 ;
    END
  END gpio_outenb_core
  PIN mprj_analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2545.395 3167.185 2545.995 ;
    END
  END mprj_analog_io[0]
  PIN mprj_analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.165 4763.000 2215.445 4768.935 ;
    END
  END mprj_analog_io[10]
  PIN mprj_analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.165 4763.000 1770.445 4768.935 ;
    END
  END mprj_analog_io[11]
  PIN mprj_analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.165 4763.000 1261.445 4768.935 ;
    END
  END mprj_analog_io[12]
  PIN mprj_analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.165 4763.000 1003.445 4768.935 ;
    END
  END mprj_analog_io[13]
  PIN mprj_analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.165 4763.000 746.445 4768.935 ;
    END
  END mprj_analog_io[14]
  PIN mprj_analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.165 4763.000 489.445 4768.935 ;
    END
  END mprj_analog_io[15]
  PIN mprj_analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.165 4763.000 232.445 4768.935 ;
    END
  END mprj_analog_io[16]
  PIN mprj_analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4623.005 4.000 4623.605 ;
    END
  END mprj_analog_io[17]
  PIN mprj_analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3774.005 4.000 3774.605 ;
    END
  END mprj_analog_io[18]
  PIN mprj_analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3558.005 4.000 3558.605 ;
    END
  END mprj_analog_io[19]
  PIN mprj_analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2771.395 3167.185 2771.995 ;
    END
  END mprj_analog_io[1]
  PIN mprj_analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3342.005 4.000 3342.605 ;
    END
  END mprj_analog_io[20]
  PIN mprj_analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3126.005 4.000 3126.605 ;
    END
  END mprj_analog_io[21]
  PIN mprj_analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2910.005 4.000 2910.605 ;
    END
  END mprj_analog_io[22]
  PIN mprj_analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2694.005 4.000 2694.605 ;
    END
  END mprj_analog_io[23]
  PIN mprj_analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2478.005 4.000 2478.605 ;
    END
  END mprj_analog_io[24]
  PIN mprj_analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1840.005 4.000 1840.605 ;
    END
  END mprj_analog_io[25]
  PIN mprj_analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1624.005 4.000 1624.605 ;
    END
  END mprj_analog_io[26]
  PIN mprj_analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1408.005 4.000 1408.605 ;
    END
  END mprj_analog_io[27]
  PIN mprj_analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1192.005 4.000 1192.605 ;
    END
  END mprj_analog_io[28]
  PIN mprj_analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2996.395 3167.185 2996.995 ;
    END
  END mprj_analog_io[2]
  PIN mprj_analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3222.395 3167.185 3222.995 ;
    END
  END mprj_analog_io[3]
  PIN mprj_analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3447.395 3167.185 3447.995 ;
    END
  END mprj_analog_io[4]
  PIN mprj_analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3672.395 3167.185 3672.995 ;
    END
  END mprj_analog_io[5]
  PIN mprj_analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4118.395 3167.185 4118.995 ;
    END
  END mprj_analog_io[6]
  PIN mprj_analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4564.395 3167.185 4564.995 ;
    END
  END mprj_analog_io[7]
  PIN mprj_analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2981.165 4763.000 2981.445 4768.935 ;
    END
  END mprj_analog_io[8]
  PIN mprj_analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.165 4763.000 2472.445 4768.935 ;
    END
  END mprj_analog_io[9]
  PIN mprj_io_analog_en[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 318.355 3167.185 318.955 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_en[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3234.355 3167.185 3234.955 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_en[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3459.355 3167.185 3459.955 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_en[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3684.355 3167.185 3684.955 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_en[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4130.355 3167.185 4130.955 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_en[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4576.355 3167.185 4576.955 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_en[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2969.205 4763.000 2969.485 4768.935 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_en[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.205 4763.000 2460.485 4768.935 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_en[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.205 4763.000 2203.485 4768.935 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_en[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.205 4763.000 1758.485 4768.935 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_en[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.205 4763.000 1249.485 4768.935 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_en[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 544.355 3167.185 544.955 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_en[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.205 4763.000 991.485 4768.935 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_en[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.205 4763.000 734.485 4768.935 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_en[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.205 4763.000 477.485 4768.935 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_en[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.205 4763.000 220.485 4768.935 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_en[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4611.045 4.000 4611.645 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_en[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3762.045 4.000 3762.645 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_en[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3546.045 4.000 3546.645 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_en[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3330.045 4.000 3330.645 ;
    END
  END mprj_io_analog_en[27]
  PIN mprj_io_analog_en[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3114.045 4.290 3114.645 ;
    END
  END mprj_io_analog_en[28]
  PIN mprj_io_analog_en[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2898.045 4.000 2898.645 ;
    END
  END mprj_io_analog_en[29]
  PIN mprj_io_analog_en[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 769.355 3167.185 769.955 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_en[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2682.045 4.000 2682.645 ;
    END
  END mprj_io_analog_en[30]
  PIN mprj_io_analog_en[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2466.045 4.000 2466.645 ;
    END
  END mprj_io_analog_en[31]
  PIN mprj_io_analog_en[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1828.045 4.000 1828.645 ;
    END
  END mprj_io_analog_en[32]
  PIN mprj_io_analog_en[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1612.045 4.000 1612.645 ;
    END
  END mprj_io_analog_en[33]
  PIN mprj_io_analog_en[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1396.045 4.000 1396.645 ;
    END
  END mprj_io_analog_en[34]
  PIN mprj_io_analog_en[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1180.045 4.000 1180.645 ;
    END
  END mprj_io_analog_en[35]
  PIN mprj_io_analog_en[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 964.045 4.000 964.645 ;
    END
  END mprj_io_analog_en[36]
  PIN mprj_io_analog_en[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 748.045 4.000 748.645 ;
    END
  END mprj_io_analog_en[37]
  PIN mprj_io_analog_en[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 995.355 3167.185 995.955 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_en[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1220.355 3167.185 1220.955 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_en[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1445.355 3167.185 1445.955 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_en[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1671.355 3167.185 1671.955 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_en[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2557.355 3167.185 2557.955 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_en[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2783.355 3167.185 2783.955 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_en[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3008.355 3167.185 3008.955 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 324.795 3167.185 325.395 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_pol[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3240.795 3167.185 3241.395 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_pol[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3465.795 3167.185 3466.395 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_pol[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3690.795 3167.185 3691.395 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_pol[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4136.795 3167.185 4137.395 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_pol[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4582.795 3167.185 4583.395 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_pol[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2962.765 4763.000 2963.045 4768.935 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_pol[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.765 4763.000 2454.045 4768.935 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_pol[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.765 4763.000 2197.045 4768.935 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_pol[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.765 4763.000 1752.045 4768.935 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_pol[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.765 4763.000 1243.045 4768.935 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_pol[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 550.795 3167.185 551.395 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_pol[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.765 4763.000 985.045 4768.935 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_pol[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.765 4763.000 728.045 4768.935 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_pol[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.765 4763.000 471.045 4768.935 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_pol[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.765 4763.000 214.045 4768.935 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_pol[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4604.605 4.000 4605.205 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_pol[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3755.605 4.000 3756.205 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_pol[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3539.605 4.000 3540.205 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_pol[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3323.605 4.000 3324.205 ;
    END
  END mprj_io_analog_pol[27]
  PIN mprj_io_analog_pol[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3107.605 4.000 3108.205 ;
    END
  END mprj_io_analog_pol[28]
  PIN mprj_io_analog_pol[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2891.605 4.000 2892.205 ;
    END
  END mprj_io_analog_pol[29]
  PIN mprj_io_analog_pol[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 775.795 3167.185 776.395 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_pol[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2675.605 4.000 2676.205 ;
    END
  END mprj_io_analog_pol[30]
  PIN mprj_io_analog_pol[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2459.605 4.000 2460.205 ;
    END
  END mprj_io_analog_pol[31]
  PIN mprj_io_analog_pol[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1821.605 4.000 1822.205 ;
    END
  END mprj_io_analog_pol[32]
  PIN mprj_io_analog_pol[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1605.605 4.000 1606.205 ;
    END
  END mprj_io_analog_pol[33]
  PIN mprj_io_analog_pol[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1389.605 4.000 1390.205 ;
    END
  END mprj_io_analog_pol[34]
  PIN mprj_io_analog_pol[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1173.605 4.000 1174.205 ;
    END
  END mprj_io_analog_pol[35]
  PIN mprj_io_analog_pol[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 957.605 4.000 958.205 ;
    END
  END mprj_io_analog_pol[36]
  PIN mprj_io_analog_pol[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 741.605 4.000 742.205 ;
    END
  END mprj_io_analog_pol[37]
  PIN mprj_io_analog_pol[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1001.795 3167.185 1002.395 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_pol[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1226.795 3167.185 1227.395 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_pol[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1451.795 3167.185 1452.395 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_pol[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1677.795 3167.185 1678.395 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_pol[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2563.795 3167.185 2564.395 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_pol[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2789.795 3167.185 2790.395 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_pol[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3014.795 3167.185 3015.395 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 339.975 3167.185 340.575 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_analog_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3255.975 3167.185 3256.575 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_analog_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3480.975 3167.185 3481.575 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_analog_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3705.975 3167.185 3706.575 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_analog_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4151.975 3167.185 4152.575 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_analog_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4597.975 3167.185 4598.575 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_analog_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2947.585 4763.000 2947.865 4768.935 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_analog_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2438.585 4763.000 2438.865 4768.935 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_analog_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2181.585 4763.000 2181.865 4768.935 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_analog_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.585 4763.000 1736.865 4768.935 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_analog_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.585 4763.000 1227.865 4768.935 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_analog_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 565.975 3167.185 566.575 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_analog_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.585 4763.000 969.865 4768.935 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_analog_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.585 4763.000 712.865 4768.935 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_analog_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.585 4763.000 455.865 4768.935 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_analog_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.585 4763.000 198.865 4768.935 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_analog_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4589.425 4.000 4590.025 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_analog_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3740.425 4.000 3741.025 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_analog_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3524.425 4.000 3525.025 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_analog_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3308.425 4.000 3309.025 ;
    END
  END mprj_io_analog_sel[27]
  PIN mprj_io_analog_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3092.425 4.000 3093.025 ;
    END
  END mprj_io_analog_sel[28]
  PIN mprj_io_analog_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2876.425 4.000 2877.025 ;
    END
  END mprj_io_analog_sel[29]
  PIN mprj_io_analog_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 790.975 3167.185 791.575 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_analog_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2660.425 4.000 2661.025 ;
    END
  END mprj_io_analog_sel[30]
  PIN mprj_io_analog_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2444.425 4.000 2445.025 ;
    END
  END mprj_io_analog_sel[31]
  PIN mprj_io_analog_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1806.425 4.000 1807.025 ;
    END
  END mprj_io_analog_sel[32]
  PIN mprj_io_analog_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1590.425 4.000 1591.025 ;
    END
  END mprj_io_analog_sel[33]
  PIN mprj_io_analog_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1374.425 4.000 1375.025 ;
    END
  END mprj_io_analog_sel[34]
  PIN mprj_io_analog_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1158.425 4.000 1159.025 ;
    END
  END mprj_io_analog_sel[35]
  PIN mprj_io_analog_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 942.425 4.000 943.025 ;
    END
  END mprj_io_analog_sel[36]
  PIN mprj_io_analog_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 726.425 4.000 727.025 ;
    END
  END mprj_io_analog_sel[37]
  PIN mprj_io_analog_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1016.975 3167.185 1017.575 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_analog_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1241.975 3167.185 1242.575 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_analog_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1466.975 3167.185 1467.575 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_analog_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1692.975 3167.185 1693.575 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_analog_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2578.975 3167.185 2579.575 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_analog_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2804.975 3167.185 2805.575 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_analog_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3029.975 3167.185 3030.575 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 321.575 3167.185 322.175 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1618.025 4.000 1618.625 ;
    END
  END mprj_io_dm[100]
  PIN mprj_io_dm[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1587.205 4.000 1587.805 ;
    END
  END mprj_io_dm[101]
  PIN mprj_io_dm[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1392.825 4.000 1393.425 ;
    END
  END mprj_io_dm[102]
  PIN mprj_io_dm[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1402.025 4.000 1402.625 ;
    END
  END mprj_io_dm[103]
  PIN mprj_io_dm[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1371.205 4.000 1371.805 ;
    END
  END mprj_io_dm[104]
  PIN mprj_io_dm[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1176.825 4.290 1177.425 ;
    END
  END mprj_io_dm[105]
  PIN mprj_io_dm[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1186.025 4.000 1186.625 ;
    END
  END mprj_io_dm[106]
  PIN mprj_io_dm[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1155.205 4.000 1155.805 ;
    END
  END mprj_io_dm[107]
  PIN mprj_io_dm[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 960.825 4.000 961.425 ;
    END
  END mprj_io_dm[108]
  PIN mprj_io_dm[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 970.025 4.000 970.625 ;
    END
  END mprj_io_dm[109]
  PIN mprj_io_dm[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 989.375 3167.185 989.975 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 939.205 4.000 939.805 ;
    END
  END mprj_io_dm[110]
  PIN mprj_io_dm[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 744.825 4.000 745.425 ;
    END
  END mprj_io_dm[111]
  PIN mprj_io_dm[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 754.025 4.000 754.625 ;
    END
  END mprj_io_dm[112]
  PIN mprj_io_dm[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 723.205 4.000 723.805 ;
    END
  END mprj_io_dm[113]
  PIN mprj_io_dm[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1020.195 3167.185 1020.795 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1223.575 3167.185 1224.175 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1214.375 3167.185 1214.975 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1245.195 3167.185 1245.795 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_dm[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1448.575 3167.185 1449.175 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1439.375 3167.185 1439.975 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1470.195 3167.185 1470.795 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_dm[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1674.575 3167.185 1675.175 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1665.375 3167.185 1665.975 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 312.375 3167.185 312.975 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1696.195 3167.185 1696.795 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_dm[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2560.575 3167.185 2561.175 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2551.375 3167.185 2551.975 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2582.195 3167.185 2582.795 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_dm[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2786.575 3167.185 2787.175 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2777.375 3167.185 2777.975 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2808.195 3167.185 2808.795 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_dm[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3011.575 3167.185 3012.175 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3002.375 3167.185 3002.975 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3033.195 3167.185 3033.795 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_dm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 343.195 3167.185 343.795 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_dm[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3237.575 3167.185 3238.175 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3228.375 3167.185 3228.975 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3259.195 3167.185 3259.795 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_dm[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3462.575 3167.185 3463.175 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3453.375 3167.185 3453.975 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3484.195 3167.185 3484.795 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_dm[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3687.575 3167.185 3688.175 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3678.375 3167.185 3678.975 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3709.195 3167.185 3709.795 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_dm[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4133.575 3167.185 4134.175 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 547.575 3167.185 548.175 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4124.375 3167.185 4124.975 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4155.195 3167.185 4155.795 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_dm[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4579.575 3167.185 4580.175 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4570.375 3167.185 4570.975 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4601.195 3167.185 4601.795 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_dm[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2965.985 4763.000 2966.265 4768.935 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2975.185 4763.000 2975.465 4768.935 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2944.365 4763.000 2944.645 4768.935 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_dm[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.985 4763.000 2457.265 4768.935 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.185 4763.000 2466.465 4768.935 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 538.375 3167.185 538.975 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2435.365 4763.000 2435.645 4768.935 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_dm[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.985 4763.000 2200.265 4768.935 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.185 4763.000 2209.465 4768.935 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.365 4763.000 2178.645 4768.935 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_dm[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.985 4763.000 1755.265 4768.935 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.185 4763.000 1764.465 4768.935 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.365 4763.000 1733.645 4768.935 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_dm[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.985 4763.000 1246.265 4768.935 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.185 4763.000 1255.465 4768.935 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.365 4763.000 1224.645 4768.935 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_dm[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 569.195 3167.185 569.795 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_dm[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.985 4763.000 988.265 4768.935 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.185 4763.000 997.465 4768.935 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.365 4763.000 966.645 4768.935 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_dm[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.985 4763.000 731.265 4768.935 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.185 4763.000 740.465 4768.935 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.365 4763.000 709.645 4768.935 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_dm[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.985 4763.000 474.265 4768.935 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.185 4763.000 483.465 4768.935 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.365 4763.000 452.645 4768.935 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_dm[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.985 4763.000 217.265 4768.935 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 772.575 3167.185 773.175 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.185 4763.000 226.465 4768.935 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.365 4763.000 195.645 4768.935 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_dm[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4607.825 4.000 4608.425 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4617.025 4.000 4617.625 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4586.205 4.000 4586.805 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_dm[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3758.825 4.000 3759.425 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3768.025 4.000 3768.625 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3737.205 4.000 3737.805 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_dm[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3542.825 4.000 3543.425 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3552.025 4.000 3552.625 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 763.375 3167.185 763.975 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3521.205 4.000 3521.805 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_dm[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3326.825 4.000 3327.425 ;
    END
  END mprj_io_dm[81]
  PIN mprj_io_dm[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3336.025 4.000 3336.625 ;
    END
  END mprj_io_dm[82]
  PIN mprj_io_dm[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3305.205 4.000 3305.805 ;
    END
  END mprj_io_dm[83]
  PIN mprj_io_dm[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3110.825 4.000 3111.425 ;
    END
  END mprj_io_dm[84]
  PIN mprj_io_dm[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3120.025 4.000 3120.625 ;
    END
  END mprj_io_dm[85]
  PIN mprj_io_dm[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3089.205 4.000 3089.805 ;
    END
  END mprj_io_dm[86]
  PIN mprj_io_dm[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2894.825 4.000 2895.425 ;
    END
  END mprj_io_dm[87]
  PIN mprj_io_dm[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2904.025 4.000 2904.625 ;
    END
  END mprj_io_dm[88]
  PIN mprj_io_dm[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2873.205 4.000 2873.805 ;
    END
  END mprj_io_dm[89]
  PIN mprj_io_dm[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 794.195 3167.185 794.795 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_dm[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2678.825 4.000 2679.425 ;
    END
  END mprj_io_dm[90]
  PIN mprj_io_dm[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2688.025 4.000 2688.625 ;
    END
  END mprj_io_dm[91]
  PIN mprj_io_dm[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2657.205 4.000 2657.805 ;
    END
  END mprj_io_dm[92]
  PIN mprj_io_dm[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2462.825 4.000 2463.425 ;
    END
  END mprj_io_dm[93]
  PIN mprj_io_dm[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2472.025 4.000 2472.625 ;
    END
  END mprj_io_dm[94]
  PIN mprj_io_dm[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2441.205 4.000 2441.805 ;
    END
  END mprj_io_dm[95]
  PIN mprj_io_dm[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1824.825 4.000 1825.425 ;
    END
  END mprj_io_dm[96]
  PIN mprj_io_dm[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1834.025 4.000 1834.625 ;
    END
  END mprj_io_dm[97]
  PIN mprj_io_dm[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1803.205 4.000 1803.805 ;
    END
  END mprj_io_dm[98]
  PIN mprj_io_dm[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1608.825 4.000 1609.425 ;
    END
  END mprj_io_dm[99]
  PIN mprj_io_dm[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 998.575 3167.185 999.175 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 346.415 3167.185 347.015 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_holdover[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3262.415 3167.185 3263.015 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_holdover[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3487.415 3167.185 3488.015 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_holdover[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3712.415 3167.185 3713.015 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_holdover[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4158.415 3167.185 4159.015 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_holdover[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4604.415 3167.185 4605.015 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_holdover[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2941.145 4763.000 2941.425 4768.935 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_holdover[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2432.145 4763.000 2432.425 4768.935 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_holdover[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.145 4763.000 2175.425 4768.935 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_holdover[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.145 4763.000 1730.425 4768.935 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_holdover[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.145 4763.000 1221.425 4768.935 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_holdover[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 572.415 3167.185 573.015 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_holdover[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.145 4763.000 963.425 4768.935 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_holdover[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.145 4763.000 706.425 4768.935 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_holdover[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.145 4763.000 449.425 4768.935 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_holdover[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.145 4763.000 192.425 4768.935 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_holdover[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4582.985 4.000 4583.585 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_holdover[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3733.985 4.000 3734.585 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_holdover[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3517.985 4.000 3518.585 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_holdover[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3301.985 4.000 3302.585 ;
    END
  END mprj_io_holdover[27]
  PIN mprj_io_holdover[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3085.985 4.000 3086.585 ;
    END
  END mprj_io_holdover[28]
  PIN mprj_io_holdover[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2869.985 4.000 2870.585 ;
    END
  END mprj_io_holdover[29]
  PIN mprj_io_holdover[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 797.415 3167.185 798.015 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_holdover[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2653.985 4.000 2654.585 ;
    END
  END mprj_io_holdover[30]
  PIN mprj_io_holdover[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2437.985 4.000 2438.585 ;
    END
  END mprj_io_holdover[31]
  PIN mprj_io_holdover[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1799.985 4.000 1800.585 ;
    END
  END mprj_io_holdover[32]
  PIN mprj_io_holdover[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1583.985 4.000 1584.585 ;
    END
  END mprj_io_holdover[33]
  PIN mprj_io_holdover[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1367.985 4.000 1368.585 ;
    END
  END mprj_io_holdover[34]
  PIN mprj_io_holdover[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1151.985 4.000 1152.585 ;
    END
  END mprj_io_holdover[35]
  PIN mprj_io_holdover[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 935.985 4.000 936.585 ;
    END
  END mprj_io_holdover[36]
  PIN mprj_io_holdover[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 719.985 4.000 720.585 ;
    END
  END mprj_io_holdover[37]
  PIN mprj_io_holdover[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1023.415 3167.185 1024.015 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_holdover[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1248.415 3167.185 1249.015 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_holdover[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1473.415 3167.185 1474.015 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_holdover[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1699.415 3167.185 1700.015 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_holdover[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2585.415 3167.185 2586.015 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_holdover[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2811.415 3167.185 2812.015 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_holdover[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3036.415 3167.185 3037.015 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 361.595 3167.185 362.195 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3277.595 3167.185 3278.195 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3502.595 3167.185 3503.195 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3727.595 3167.185 3728.195 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4173.595 3167.185 4174.195 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4619.595 3167.185 4620.195 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2925.965 4763.000 2926.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.965 4763.000 2417.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2159.965 4763.000 2160.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.965 4763.000 1715.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.965 4763.000 1206.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 587.595 3167.185 588.195 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.965 4763.000 948.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.965 4763.000 691.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.965 4763.000 434.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.965 4763.000 177.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4567.805 4.000 4568.405 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3718.805 4.000 3719.405 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3502.805 4.000 3503.405 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_ib_mode_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3286.805 4.000 3287.405 ;
    END
  END mprj_io_ib_mode_sel[27]
  PIN mprj_io_ib_mode_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3070.805 4.000 3071.405 ;
    END
  END mprj_io_ib_mode_sel[28]
  PIN mprj_io_ib_mode_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2854.805 4.000 2855.405 ;
    END
  END mprj_io_ib_mode_sel[29]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 812.595 3167.185 813.195 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_ib_mode_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2638.805 4.000 2639.405 ;
    END
  END mprj_io_ib_mode_sel[30]
  PIN mprj_io_ib_mode_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2422.805 4.000 2423.405 ;
    END
  END mprj_io_ib_mode_sel[31]
  PIN mprj_io_ib_mode_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1784.805 4.000 1785.405 ;
    END
  END mprj_io_ib_mode_sel[32]
  PIN mprj_io_ib_mode_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1568.805 4.000 1569.405 ;
    END
  END mprj_io_ib_mode_sel[33]
  PIN mprj_io_ib_mode_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1352.805 4.000 1353.405 ;
    END
  END mprj_io_ib_mode_sel[34]
  PIN mprj_io_ib_mode_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1136.805 4.000 1137.405 ;
    END
  END mprj_io_ib_mode_sel[35]
  PIN mprj_io_ib_mode_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 920.805 4.000 921.405 ;
    END
  END mprj_io_ib_mode_sel[36]
  PIN mprj_io_ib_mode_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 704.805 4.000 705.405 ;
    END
  END mprj_io_ib_mode_sel[37]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1038.595 3167.185 1039.195 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1263.595 3167.185 1264.195 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1488.595 3167.185 1489.195 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1714.595 3167.185 1715.195 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2600.595 3167.185 2601.195 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2826.595 3167.185 2827.195 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3051.595 3167.185 3052.195 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 293.975 3167.185 294.575 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3209.975 3167.185 3210.575 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3434.975 3167.185 3435.575 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3659.975 3167.185 3660.575 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4105.975 3167.185 4106.575 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4551.975 3167.185 4552.575 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2993.585 4763.000 2993.865 4768.935 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2484.585 4763.000 2484.865 4768.935 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2227.585 4763.000 2227.865 4768.935 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.585 4763.000 1782.865 4768.935 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.585 4763.000 1273.865 4768.935 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 519.975 3167.185 520.575 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.585 4763.000 1015.865 4768.935 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.585 4763.000 758.865 4768.935 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.585 4763.000 501.865 4768.935 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.585 4763.000 244.865 4768.935 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4635.425 4.000 4636.025 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3786.425 4.000 3787.025 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3570.425 4.000 3571.025 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3354.425 4.000 3355.025 ;
    END
  END mprj_io_in[27]
  PIN mprj_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3138.425 4.000 3139.025 ;
    END
  END mprj_io_in[28]
  PIN mprj_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2922.425 4.000 2923.025 ;
    END
  END mprj_io_in[29]
  PIN mprj_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 744.975 3167.185 745.575 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2706.425 4.000 2707.025 ;
    END
  END mprj_io_in[30]
  PIN mprj_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2490.425 4.000 2491.025 ;
    END
  END mprj_io_in[31]
  PIN mprj_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1852.425 4.000 1853.025 ;
    END
  END mprj_io_in[32]
  PIN mprj_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1636.425 4.000 1637.025 ;
    END
  END mprj_io_in[33]
  PIN mprj_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1420.425 4.000 1421.025 ;
    END
  END mprj_io_in[34]
  PIN mprj_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1204.425 4.000 1205.025 ;
    END
  END mprj_io_in[35]
  PIN mprj_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 988.425 4.000 989.025 ;
    END
  END mprj_io_in[36]
  PIN mprj_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 772.425 4.000 773.025 ;
    END
  END mprj_io_in[37]
  PIN mprj_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 970.975 3167.185 971.575 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1195.975 3167.185 1196.575 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1420.975 3167.185 1421.575 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1646.975 3167.185 1647.575 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2532.975 3167.185 2533.575 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2758.975 3167.185 2759.575 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2983.975 3167.185 2984.575 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_inp_dis[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 327.555 3167.185 328.155 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_inp_dis[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3243.555 3167.185 3244.155 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_inp_dis[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3468.555 3167.185 3469.155 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_inp_dis[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3693.555 3167.185 3694.155 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_inp_dis[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4139.555 3167.185 4140.155 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_inp_dis[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4585.555 3167.185 4586.155 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_inp_dis[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2960.005 4763.000 2960.285 4768.935 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_inp_dis[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2451.005 4763.000 2451.285 4768.935 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_inp_dis[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.005 4763.000 2194.285 4768.935 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_inp_dis[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.005 4763.000 1749.285 4768.935 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_inp_dis[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.005 4763.000 1240.285 4768.935 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_inp_dis[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 553.555 3167.185 554.155 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_inp_dis[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.005 4763.000 982.285 4768.935 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_inp_dis[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.005 4763.000 725.285 4768.935 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_inp_dis[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.005 4763.000 468.285 4768.935 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_inp_dis[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.005 4763.000 211.285 4768.935 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_inp_dis[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4601.845 4.000 4602.445 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_inp_dis[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3752.845 4.000 3753.445 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_inp_dis[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3536.845 4.000 3537.445 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_inp_dis[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3320.845 4.000 3321.445 ;
    END
  END mprj_io_inp_dis[27]
  PIN mprj_io_inp_dis[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3104.845 4.000 3105.445 ;
    END
  END mprj_io_inp_dis[28]
  PIN mprj_io_inp_dis[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2888.845 4.000 2889.445 ;
    END
  END mprj_io_inp_dis[29]
  PIN mprj_io_inp_dis[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 778.555 3167.185 779.155 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_inp_dis[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2672.845 4.000 2673.445 ;
    END
  END mprj_io_inp_dis[30]
  PIN mprj_io_inp_dis[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2456.845 4.000 2457.445 ;
    END
  END mprj_io_inp_dis[31]
  PIN mprj_io_inp_dis[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1818.845 4.000 1819.445 ;
    END
  END mprj_io_inp_dis[32]
  PIN mprj_io_inp_dis[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1602.845 4.000 1603.445 ;
    END
  END mprj_io_inp_dis[33]
  PIN mprj_io_inp_dis[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1386.845 4.000 1387.445 ;
    END
  END mprj_io_inp_dis[34]
  PIN mprj_io_inp_dis[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1170.845 4.000 1171.445 ;
    END
  END mprj_io_inp_dis[35]
  PIN mprj_io_inp_dis[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 954.845 4.000 955.445 ;
    END
  END mprj_io_inp_dis[36]
  PIN mprj_io_inp_dis[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 738.845 4.000 739.445 ;
    END
  END mprj_io_inp_dis[37]
  PIN mprj_io_inp_dis[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1004.555 3167.185 1005.155 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_inp_dis[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1229.555 3167.185 1230.155 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_inp_dis[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1454.555 3167.185 1455.155 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_inp_dis[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1680.555 3167.185 1681.155 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_inp_dis[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2566.555 3167.185 2567.155 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_inp_dis[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2792.555 3167.185 2793.155 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_inp_dis[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3017.555 3167.185 3018.155 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 364.815 3167.185 365.415 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3280.815 3167.185 3281.415 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3505.815 3167.185 3506.415 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3730.815 3167.185 3731.415 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4176.815 3167.185 4177.415 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4622.815 3167.185 4623.415 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2922.745 4763.000 2923.025 4768.935 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.745 4763.000 2414.025 4768.935 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.745 4763.000 2157.025 4768.935 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.745 4763.000 1712.025 4768.935 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.745 4763.000 1203.025 4768.935 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 590.815 3167.185 591.415 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.745 4763.000 945.025 4768.935 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.745 4763.000 688.025 4768.935 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.745 4763.000 431.025 4768.935 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.745 4763.000 174.025 4768.935 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4564.585 4.000 4565.185 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3715.585 4.000 3716.185 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3499.585 4.000 3500.185 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3283.585 4.000 3284.185 ;
    END
  END mprj_io_oeb[27]
  PIN mprj_io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3067.585 4.000 3068.185 ;
    END
  END mprj_io_oeb[28]
  PIN mprj_io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2851.585 4.000 2852.185 ;
    END
  END mprj_io_oeb[29]
  PIN mprj_io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 815.815 3167.185 816.415 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2635.585 4.000 2636.185 ;
    END
  END mprj_io_oeb[30]
  PIN mprj_io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2419.585 4.000 2420.185 ;
    END
  END mprj_io_oeb[31]
  PIN mprj_io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1781.585 4.000 1782.185 ;
    END
  END mprj_io_oeb[32]
  PIN mprj_io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1565.585 4.000 1566.185 ;
    END
  END mprj_io_oeb[33]
  PIN mprj_io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1349.585 4.000 1350.185 ;
    END
  END mprj_io_oeb[34]
  PIN mprj_io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1133.585 4.000 1134.185 ;
    END
  END mprj_io_oeb[35]
  PIN mprj_io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 917.585 4.000 918.185 ;
    END
  END mprj_io_oeb[36]
  PIN mprj_io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 701.585 4.000 702.185 ;
    END
  END mprj_io_oeb[37]
  PIN mprj_io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1041.815 3167.185 1042.415 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1266.815 3167.185 1267.415 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1491.815 3167.185 1492.415 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1717.815 3167.185 1718.415 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2603.815 3167.185 2604.415 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2829.815 3167.185 2830.415 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3054.815 3167.185 3055.415 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_one[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 299.955 3167.185 300.555 ;
    END
  END mprj_io_one[0]
  PIN mprj_io_one[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3215.955 3167.185 3216.555 ;
    END
  END mprj_io_one[10]
  PIN mprj_io_one[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3440.955 3167.185 3441.555 ;
    END
  END mprj_io_one[11]
  PIN mprj_io_one[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3665.955 3167.185 3666.555 ;
    END
  END mprj_io_one[12]
  PIN mprj_io_one[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4111.955 3167.185 4112.555 ;
    END
  END mprj_io_one[13]
  PIN mprj_io_one[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4557.955 3167.185 4558.555 ;
    END
  END mprj_io_one[14]
  PIN mprj_io_one[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2987.605 4763.000 2987.885 4768.935 ;
    END
  END mprj_io_one[15]
  PIN mprj_io_one[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2478.605 4763.000 2478.885 4768.935 ;
    END
  END mprj_io_one[16]
  PIN mprj_io_one[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.605 4763.000 2221.885 4768.935 ;
    END
  END mprj_io_one[17]
  PIN mprj_io_one[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.605 4763.000 1776.885 4768.935 ;
    END
  END mprj_io_one[18]
  PIN mprj_io_one[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.605 4763.000 1267.885 4768.935 ;
    END
  END mprj_io_one[19]
  PIN mprj_io_one[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 525.955 3167.185 526.555 ;
    END
  END mprj_io_one[1]
  PIN mprj_io_one[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.605 4763.000 1009.885 4768.935 ;
    END
  END mprj_io_one[20]
  PIN mprj_io_one[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.605 4763.000 752.885 4768.935 ;
    END
  END mprj_io_one[21]
  PIN mprj_io_one[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.605 4763.000 495.885 4768.935 ;
    END
  END mprj_io_one[22]
  PIN mprj_io_one[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.605 4763.000 238.885 4768.935 ;
    END
  END mprj_io_one[23]
  PIN mprj_io_one[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4629.445 4.000 4630.045 ;
    END
  END mprj_io_one[24]
  PIN mprj_io_one[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3780.445 4.000 3781.045 ;
    END
  END mprj_io_one[25]
  PIN mprj_io_one[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3564.445 4.000 3565.045 ;
    END
  END mprj_io_one[26]
  PIN mprj_io_one[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3348.445 4.000 3349.045 ;
    END
  END mprj_io_one[27]
  PIN mprj_io_one[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3132.445 4.000 3133.045 ;
    END
  END mprj_io_one[28]
  PIN mprj_io_one[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2916.445 4.000 2917.045 ;
    END
  END mprj_io_one[29]
  PIN mprj_io_one[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 750.955 3167.185 751.555 ;
    END
  END mprj_io_one[2]
  PIN mprj_io_one[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2700.445 4.000 2701.045 ;
    END
  END mprj_io_one[30]
  PIN mprj_io_one[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2484.445 4.000 2485.045 ;
    END
  END mprj_io_one[31]
  PIN mprj_io_one[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1846.445 4.000 1847.045 ;
    END
  END mprj_io_one[32]
  PIN mprj_io_one[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1630.445 4.000 1631.045 ;
    END
  END mprj_io_one[33]
  PIN mprj_io_one[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1414.445 4.000 1415.045 ;
    END
  END mprj_io_one[34]
  PIN mprj_io_one[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1198.445 4.290 1199.045 ;
    END
  END mprj_io_one[35]
  PIN mprj_io_one[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 982.445 4.000 983.045 ;
    END
  END mprj_io_one[36]
  PIN mprj_io_one[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 766.445 4.000 767.045 ;
    END
  END mprj_io_one[37]
  PIN mprj_io_one[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 976.955 3167.185 977.555 ;
    END
  END mprj_io_one[3]
  PIN mprj_io_one[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1201.955 3167.185 1202.555 ;
    END
  END mprj_io_one[4]
  PIN mprj_io_one[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1426.955 3167.185 1427.555 ;
    END
  END mprj_io_one[5]
  PIN mprj_io_one[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1652.955 3167.185 1653.555 ;
    END
  END mprj_io_one[6]
  PIN mprj_io_one[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2538.955 3167.185 2539.555 ;
    END
  END mprj_io_one[7]
  PIN mprj_io_one[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2764.955 3167.185 2765.555 ;
    END
  END mprj_io_one[8]
  PIN mprj_io_one[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2989.955 3167.185 2990.555 ;
    END
  END mprj_io_one[9]
  PIN mprj_io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 349.175 3167.185 349.775 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3265.175 3167.185 3265.775 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3490.175 3167.185 3490.775 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3715.175 3167.185 3715.775 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4161.175 3167.185 4161.775 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4607.175 3167.185 4607.775 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2938.385 4763.000 2938.665 4768.935 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2429.385 4763.000 2429.665 4768.935 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.385 4763.000 2172.665 4768.935 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.385 4763.000 1727.665 4768.935 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.385 4763.000 1218.665 4768.935 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 575.175 3167.185 575.775 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.385 4763.000 960.665 4768.935 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.385 4763.000 703.665 4768.935 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.385 4763.000 446.665 4768.935 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.385 4763.000 189.665 4768.935 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4580.225 4.000 4580.825 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3731.225 4.000 3731.825 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3515.225 4.000 3515.825 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3299.225 4.000 3299.825 ;
    END
  END mprj_io_out[27]
  PIN mprj_io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3083.225 4.000 3083.825 ;
    END
  END mprj_io_out[28]
  PIN mprj_io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2867.225 4.000 2867.825 ;
    END
  END mprj_io_out[29]
  PIN mprj_io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 800.175 3167.185 800.775 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2651.225 4.000 2651.825 ;
    END
  END mprj_io_out[30]
  PIN mprj_io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2435.225 4.000 2435.825 ;
    END
  END mprj_io_out[31]
  PIN mprj_io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1797.225 4.000 1797.825 ;
    END
  END mprj_io_out[32]
  PIN mprj_io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1581.225 4.000 1581.825 ;
    END
  END mprj_io_out[33]
  PIN mprj_io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1365.225 4.000 1365.825 ;
    END
  END mprj_io_out[34]
  PIN mprj_io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1149.225 4.000 1149.825 ;
    END
  END mprj_io_out[35]
  PIN mprj_io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 933.225 4.000 933.825 ;
    END
  END mprj_io_out[36]
  PIN mprj_io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 717.225 4.000 717.825 ;
    END
  END mprj_io_out[37]
  PIN mprj_io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1026.175 3167.185 1026.775 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1251.175 3167.185 1251.775 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1476.175 3167.185 1476.775 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1702.175 3167.185 1702.775 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2588.175 3167.185 2588.775 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2814.175 3167.185 2814.775 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3039.175 3167.185 3039.775 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 303.175 3167.185 303.775 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_slow_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3219.175 3167.185 3219.775 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_slow_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3444.175 3167.185 3444.775 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_slow_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3669.175 3167.185 3669.775 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_slow_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4115.175 3167.185 4115.775 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_slow_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4561.175 3167.185 4561.775 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_slow_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2984.385 4763.000 2984.665 4768.935 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_slow_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2475.385 4763.000 2475.665 4768.935 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_slow_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.385 4763.000 2218.665 4768.935 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_slow_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.385 4763.000 1773.665 4768.935 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_slow_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.385 4763.000 1264.665 4768.935 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_slow_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 529.175 3167.185 529.775 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_slow_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.385 4763.000 1006.665 4768.935 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_slow_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.385 4763.000 749.665 4768.935 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_slow_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.385 4763.000 492.665 4768.935 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_slow_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.385 4763.000 235.665 4768.935 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_slow_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4626.225 4.000 4626.825 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_slow_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3777.225 4.000 3777.825 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_slow_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3561.225 4.000 3561.825 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_slow_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3345.225 4.000 3345.825 ;
    END
  END mprj_io_slow_sel[27]
  PIN mprj_io_slow_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3129.225 4.000 3129.825 ;
    END
  END mprj_io_slow_sel[28]
  PIN mprj_io_slow_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2913.225 4.000 2913.825 ;
    END
  END mprj_io_slow_sel[29]
  PIN mprj_io_slow_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 754.175 3167.185 754.775 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_slow_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2697.225 4.000 2697.825 ;
    END
  END mprj_io_slow_sel[30]
  PIN mprj_io_slow_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2481.225 4.000 2481.825 ;
    END
  END mprj_io_slow_sel[31]
  PIN mprj_io_slow_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1843.225 4.000 1843.825 ;
    END
  END mprj_io_slow_sel[32]
  PIN mprj_io_slow_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1627.225 4.000 1627.825 ;
    END
  END mprj_io_slow_sel[33]
  PIN mprj_io_slow_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1411.225 4.000 1411.825 ;
    END
  END mprj_io_slow_sel[34]
  PIN mprj_io_slow_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1195.225 4.000 1195.825 ;
    END
  END mprj_io_slow_sel[35]
  PIN mprj_io_slow_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 979.225 4.000 979.825 ;
    END
  END mprj_io_slow_sel[36]
  PIN mprj_io_slow_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 763.225 4.000 763.825 ;
    END
  END mprj_io_slow_sel[37]
  PIN mprj_io_slow_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 980.175 3167.185 980.775 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_slow_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1205.175 3167.185 1205.775 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_slow_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1430.175 3167.185 1430.775 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_slow_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1656.175 3167.185 1656.775 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_slow_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2542.175 3167.185 2542.775 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_slow_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2768.175 3167.185 2768.775 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_slow_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2993.175 3167.185 2993.775 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 358.375 3167.185 358.975 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3274.375 3167.185 3274.975 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3499.375 3167.185 3499.975 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3724.375 3167.185 3724.975 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4170.375 3167.185 4170.975 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4616.375 3167.185 4616.975 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2929.185 4763.000 2929.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.185 4763.000 2420.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.185 4763.000 2163.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.185 4763.000 1718.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.185 4763.000 1209.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 584.375 3167.185 584.975 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.185 4763.000 951.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.185 4763.000 694.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.185 4763.000 437.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.185 4763.000 180.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4571.025 4.000 4571.625 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3722.025 4.000 3722.625 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3506.025 4.000 3506.625 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_vtrip_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3290.025 4.000 3290.625 ;
    END
  END mprj_io_vtrip_sel[27]
  PIN mprj_io_vtrip_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3074.025 4.000 3074.625 ;
    END
  END mprj_io_vtrip_sel[28]
  PIN mprj_io_vtrip_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2858.025 4.000 2858.625 ;
    END
  END mprj_io_vtrip_sel[29]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 809.375 3167.185 809.975 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_vtrip_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2642.025 4.000 2642.625 ;
    END
  END mprj_io_vtrip_sel[30]
  PIN mprj_io_vtrip_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2426.025 4.000 2426.625 ;
    END
  END mprj_io_vtrip_sel[31]
  PIN mprj_io_vtrip_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1788.025 4.000 1788.625 ;
    END
  END mprj_io_vtrip_sel[32]
  PIN mprj_io_vtrip_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1572.025 4.000 1572.625 ;
    END
  END mprj_io_vtrip_sel[33]
  PIN mprj_io_vtrip_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1356.025 4.000 1356.625 ;
    END
  END mprj_io_vtrip_sel[34]
  PIN mprj_io_vtrip_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1140.025 4.000 1140.625 ;
    END
  END mprj_io_vtrip_sel[35]
  PIN mprj_io_vtrip_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 924.025 4.000 924.625 ;
    END
  END mprj_io_vtrip_sel[36]
  PIN mprj_io_vtrip_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 708.025 4.000 708.625 ;
    END
  END mprj_io_vtrip_sel[37]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1035.375 3167.185 1035.975 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1260.375 3167.185 1260.975 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1485.375 3167.185 1485.975 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1711.375 3167.185 1711.975 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2597.375 3167.185 2597.975 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2823.375 3167.185 2823.975 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3048.375 3167.185 3048.975 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN por_l
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.715 -2.000 758.995 4.000 ;
    END
  END por_l
  PIN porb_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.775 -2.000 1330.055 4.000 ;
    END
  END porb_h
  PIN rstb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.835 -10.525 497.115 4.000 ;
    END
  END rstb_h
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.920 10.640 15.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3147.180 10.640 3152.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 10.880 3154.920 20.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4735.060 3154.920 4748.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.920 10.640 72.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3087.180 10.640 3089.180 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 10.640 130.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 4596.300 130.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.920 10.640 230.320 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.920 620.365 230.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.920 4596.300 230.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.920 10.640 330.320 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.920 620.365 330.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.920 4596.300 330.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.920 10.640 430.320 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.920 620.365 430.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.920 4596.300 430.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.920 10.640 530.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.920 4596.300 530.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.920 10.640 630.320 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.920 620.365 630.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.920 4596.300 630.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.920 10.640 730.320 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.920 620.365 730.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.920 4596.300 730.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.920 10.640 830.320 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.920 620.365 830.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.920 4596.300 830.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.920 10.640 930.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.920 4596.300 930.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.920 34.080 1030.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.920 4596.300 1030.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1123.920 10.640 1130.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1123.920 4596.300 1130.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.920 10.640 1230.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.920 4596.300 1230.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.920 10.640 1330.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.920 4596.300 1330.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1423.920 10.640 1430.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1423.920 4596.300 1430.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.920 10.640 1530.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.920 4596.300 1530.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.920 10.640 1630.320 177.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.920 284.020 1630.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.920 4596.300 1630.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1723.920 10.640 1730.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1723.920 4596.300 1730.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.920 10.640 1830.320 123.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.920 570.365 1830.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.920 4596.300 1830.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.920 10.640 1930.320 123.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.920 570.365 1930.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.920 4596.300 1930.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.920 10.640 2030.320 123.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.920 570.365 2030.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.920 4596.300 2030.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.920 10.640 2130.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.920 4596.300 2130.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.920 10.640 2230.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.920 4596.300 2230.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2323.920 10.640 2330.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2323.920 4596.300 2330.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.920 10.640 2430.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.920 4596.300 2430.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.920 10.640 2530.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.920 4596.300 2530.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2623.920 10.640 2630.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2623.920 4596.300 2630.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.920 10.640 2730.320 193.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.920 733.285 2730.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.920 4596.300 2730.320 4603.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.920 10.640 2830.320 192.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.920 737.100 2830.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.920 4596.300 2830.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2923.920 10.640 2930.320 193.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2923.920 733.285 2930.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2923.920 4596.300 2930.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3023.920 10.640 3030.320 193.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 3023.920 733.285 3030.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3023.920 4596.300 3030.320 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 308.680 3154.920 315.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 428.680 3154.920 435.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 548.680 3154.920 555.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 668.680 3154.920 675.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 788.680 3154.920 795.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 908.680 3154.920 915.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1028.680 75.920 1035.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1148.680 75.920 1155.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1268.680 75.920 1275.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1388.680 75.920 1395.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1508.680 75.920 1515.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1628.680 75.920 1635.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1748.680 75.920 1755.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1868.680 75.920 1875.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2108.680 75.920 2115.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2348.680 75.920 2355.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2468.680 75.920 2475.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2588.680 75.920 2595.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2708.680 75.920 2715.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2828.680 75.920 2835.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2948.680 75.920 2955.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3068.680 75.920 3075.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3188.680 75.920 3195.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3308.680 75.920 3315.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3428.680 75.920 3435.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3548.680 75.920 3555.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3668.680 75.920 3675.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3788.680 75.920 3795.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3908.680 75.920 3915.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4028.680 75.920 4035.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4148.680 75.920 4155.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4268.680 75.920 4275.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4508.680 75.920 4515.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 28.000 188.680 3154.920 195.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1028.680 3154.920 1035.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1148.680 3154.920 1155.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1268.680 3154.920 1275.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1388.680 3154.920 1395.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1508.680 3154.920 1515.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1628.680 3154.920 1635.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1748.680 3154.920 1755.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1988.680 3154.920 1995.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2228.680 3154.920 2235.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2468.680 3154.920 2475.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2588.680 3154.920 2595.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2708.680 3154.920 2715.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2828.680 3154.920 2835.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2948.680 3154.920 2955.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3068.680 3154.920 3075.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3188.680 3154.920 3195.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3308.680 3154.920 3315.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3428.680 3154.920 3435.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3548.680 3154.920 3555.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3668.680 3154.920 3675.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3788.680 3154.920 3795.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4028.680 3154.920 4035.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4148.680 3154.920 4155.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4268.680 3154.920 4275.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4508.680 3154.920 4515.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 242.680 3154.920 257.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 362.680 3154.920 377.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 482.680 3154.920 497.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 602.680 3154.920 617.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 722.680 3154.920 737.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 953.000 3154.920 967.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2650.320 4640.080 2655.320 4692.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 2623.920 4597.700 2837.920 4599.300 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.920 10.640 27.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3135.180 10.640 3140.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 34.080 3154.920 44.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4705.860 3154.920 4718.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 815.480 3154.920 820.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.720 10.640 1280.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.720 10.640 1380.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 10.640 1480.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 4596.300 1480.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.640 4596.300 270.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.640 10.640 570.040 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.640 4596.300 570.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1163.640 10.640 1170.040 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1163.640 4596.300 1170.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.640 10.640 1470.040 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.640 4596.300 1470.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.640 10.640 1770.040 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.640 4596.300 1770.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2063.640 4596.300 2070.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.640 10.640 2370.040 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.640 4596.300 2370.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2763.640 4596.300 2770.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 963.640 4596.300 970.040 4754.800 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 64.920 10.640 69.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3093.180 10.640 3098.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 115.280 3154.920 125.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4603.660 3154.920 4616.660 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 831.480 3154.920 836.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 850.720 620.365 855.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 900.720 10.640 905.520 989.000 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 52.920 10.640 57.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3105.180 10.640 3110.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 92.080 3154.920 102.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4632.860 3154.920 4645.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 847.480 3154.920 852.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1843.720 570.365 1848.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1883.720 570.365 1888.520 989.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 40.920 10.640 45.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3117.180 10.640 3122.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 68.880 3154.920 78.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4662.060 3154.920 4675.060 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 863.480 3154.920 868.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1859.720 570.365 1864.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1899.720 570.365 1904.520 989.000 ;
    END
  END vdda2
  PIN vddio
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 650.000 145.380 1082.115 150.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 650.000 159.380 1082.115 164.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.720 10.640 659.520 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 1040.720 34.080 1045.520 189.000 ;
    END
  END vddio
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.920 10.640 51.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3111.180 10.640 3116.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 80.480 3154.920 90.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4647.460 3154.920 4660.460 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 855.480 3154.920 860.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1851.720 570.365 1856.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.720 570.365 1896.520 989.000 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.920 10.640 39.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3123.180 10.640 3128.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 57.280 3154.920 67.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4676.660 3154.920 4689.660 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 871.480 3154.920 876.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1867.720 570.365 1872.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1907.720 570.365 1912.520 989.000 ;
    END
  END vssa2
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.920 10.640 21.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3141.180 10.640 3146.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 22.480 3154.920 32.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4720.460 3154.920 4733.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.920 10.640 75.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3090.180 10.640 3092.180 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.520 10.640 137.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.520 4596.300 137.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.520 10.640 237.920 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.520 620.365 237.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.520 4596.300 237.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.520 10.640 337.920 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.520 620.365 337.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.520 4596.300 337.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 431.520 10.640 437.920 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 431.520 620.365 437.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 431.520 4596.300 437.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.520 10.640 537.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.520 4596.300 537.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.520 10.640 637.920 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.520 620.365 637.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.520 4596.300 637.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 731.520 10.640 737.920 169.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 731.520 620.365 737.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 731.520 4596.300 737.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.520 10.640 837.920 173.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.520 620.365 837.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.520 4596.300 837.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.520 10.640 937.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.520 4596.300 937.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1031.520 34.080 1037.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1031.520 4596.300 1037.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.520 10.640 1137.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.520 4596.300 1137.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.520 10.640 1237.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.520 4596.300 1237.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1331.520 10.640 1337.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1331.520 4596.300 1337.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1431.520 10.640 1437.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1431.520 4596.300 1437.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1531.520 10.640 1537.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1531.520 4596.300 1537.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1631.520 10.640 1637.920 177.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1631.520 284.020 1637.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1631.520 4596.300 1637.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1731.520 10.640 1737.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1731.520 4596.300 1737.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.520 10.640 1837.920 123.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.520 570.365 1837.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.520 4596.300 1837.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.520 10.640 1937.920 123.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.520 570.365 1937.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.520 4596.300 1937.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2031.520 10.640 2037.920 119.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2031.520 570.365 2037.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2031.520 4596.300 2037.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2131.520 10.640 2137.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2131.520 4596.300 2137.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.520 10.640 2237.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.520 4596.300 2237.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2331.520 10.640 2337.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2331.520 4596.300 2337.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2431.520 10.640 2437.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2431.520 4596.300 2437.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2531.520 10.640 2537.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2531.520 4596.300 2537.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2631.520 10.640 2637.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2631.520 4596.300 2637.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.520 10.640 2737.920 193.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.520 733.285 2737.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.520 4596.300 2737.920 4603.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.520 10.640 2837.920 193.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.520 733.285 2837.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.520 4596.300 2837.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.520 10.640 2937.920 193.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.520 733.285 2937.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.520 4596.300 2937.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3031.520 10.640 3037.920 193.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 3031.520 733.285 3037.920 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3031.520 4596.300 3037.920 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 317.480 3154.920 323.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 437.480 3154.920 443.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 557.480 3154.920 563.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 677.480 3154.920 683.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 797.480 3154.920 803.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 917.480 3154.920 923.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1037.480 75.920 1043.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1157.480 75.920 1163.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1277.480 75.920 1283.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1397.480 75.920 1403.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1517.480 75.920 1523.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1637.480 75.920 1643.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1757.480 75.920 1763.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1877.480 75.920 1883.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2117.480 75.920 2123.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2357.480 75.920 2363.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2477.480 75.920 2483.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2597.480 75.920 2603.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2717.480 75.920 2723.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2837.480 75.920 2843.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2957.480 75.920 2963.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3077.480 75.920 3083.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3197.480 75.920 3203.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3317.480 75.920 3323.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3437.480 75.920 3443.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3557.480 75.920 3563.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3677.480 75.920 3683.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3797.480 75.920 3803.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3917.480 75.920 3923.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4037.480 75.920 4043.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4157.480 75.920 4163.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4277.480 75.920 4283.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4517.480 75.920 4523.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 28.000 197.480 3154.920 203.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1037.480 3154.920 1043.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1157.480 3154.920 1163.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1277.480 3154.920 1283.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1397.480 3154.920 1403.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1517.480 3154.920 1523.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1637.480 3154.920 1643.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1757.480 3154.920 1763.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1997.480 3154.920 2003.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2237.480 3154.920 2243.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2477.480 3154.920 2483.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2597.480 3154.920 2603.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2717.480 3154.920 2723.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2837.480 3154.920 2843.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2957.480 3154.920 2963.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3077.480 3154.920 3083.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3197.480 3154.920 3203.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3317.480 3154.920 3323.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3437.480 3154.920 3443.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3557.480 3154.920 3563.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3677.480 3154.920 3683.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3797.480 3154.920 3803.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4037.480 3154.920 4043.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4157.480 3154.920 4163.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4277.480 3154.920 4283.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4517.480 3154.920 4523.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 259.480 3154.920 273.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 379.480 3154.920 393.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 499.480 3154.920 513.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 619.480 3154.920 633.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 739.480 3154.920 753.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 969.800 3154.920 984.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.760 4640.080 2661.760 4692.240 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.920 10.640 33.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3129.180 10.640 3134.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 45.680 3154.920 55.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4691.260 3154.920 4704.260 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 823.480 3154.920 828.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.720 10.640 1288.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1383.720 10.640 1388.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1483.720 10.640 1488.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.040 4596.300 262.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 556.040 10.640 562.440 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 556.040 4596.300 562.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.040 10.640 1162.440 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.040 4596.300 1162.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1456.040 10.640 1462.440 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1456.040 4596.300 1462.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.040 10.640 1762.440 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.040 4596.300 1762.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.040 4596.300 2062.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.040 10.640 2362.440 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.040 4596.300 2362.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2756.040 4596.300 2762.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.040 10.640 962.440 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.040 4596.300 962.440 4754.800 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 58.920 10.640 63.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3099.180 10.640 3104.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 103.680 3154.920 113.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4618.260 3154.920 4631.260 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 839.480 3154.920 844.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.720 620.365 863.520 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.720 10.640 913.520 989.000 ;
    END
  END vssd2
  PIN vssio
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 650.000 152.380 1082.115 157.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 650.000 166.380 1082.115 171.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.520 10.640 666.320 169.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1047.520 34.080 1052.320 189.000 ;
    END
  END vssio
  OBS
      LAYER li1 ;
        RECT 10.120 10.795 3154.680 4754.645 ;
      LAYER met1 ;
        RECT 4.670 10.240 3159.210 4762.680 ;
      LAYER met2 ;
        RECT 4.690 4762.720 173.465 4763.810 ;
        RECT 174.305 4762.720 176.685 4763.810 ;
        RECT 177.525 4762.720 179.905 4763.810 ;
        RECT 180.745 4762.720 189.105 4763.810 ;
        RECT 189.945 4762.720 191.865 4763.810 ;
        RECT 192.705 4762.720 195.085 4763.810 ;
        RECT 195.925 4762.720 198.305 4763.810 ;
        RECT 199.145 4762.720 210.725 4763.810 ;
        RECT 211.565 4762.720 213.485 4763.810 ;
        RECT 214.325 4762.720 216.705 4763.810 ;
        RECT 217.545 4762.720 219.925 4763.810 ;
        RECT 220.765 4762.720 225.905 4763.810 ;
        RECT 226.745 4762.720 231.885 4763.810 ;
        RECT 232.725 4762.720 235.105 4763.810 ;
        RECT 235.945 4762.720 238.325 4763.810 ;
        RECT 239.165 4762.720 244.305 4763.810 ;
        RECT 245.145 4762.720 430.465 4763.810 ;
        RECT 431.305 4762.720 433.685 4763.810 ;
        RECT 434.525 4762.720 436.905 4763.810 ;
        RECT 437.745 4762.720 446.105 4763.810 ;
        RECT 446.945 4762.720 448.865 4763.810 ;
        RECT 449.705 4762.720 452.085 4763.810 ;
        RECT 452.925 4762.720 455.305 4763.810 ;
        RECT 456.145 4762.720 467.725 4763.810 ;
        RECT 468.565 4762.720 470.485 4763.810 ;
        RECT 471.325 4762.720 473.705 4763.810 ;
        RECT 474.545 4762.720 476.925 4763.810 ;
        RECT 477.765 4762.720 482.905 4763.810 ;
        RECT 483.745 4762.720 488.885 4763.810 ;
        RECT 489.725 4762.720 492.105 4763.810 ;
        RECT 492.945 4762.720 495.325 4763.810 ;
        RECT 496.165 4762.720 501.305 4763.810 ;
        RECT 502.145 4762.720 687.465 4763.810 ;
        RECT 688.305 4762.720 690.685 4763.810 ;
        RECT 691.525 4762.720 693.905 4763.810 ;
        RECT 694.745 4762.720 703.105 4763.810 ;
        RECT 703.945 4762.720 705.865 4763.810 ;
        RECT 706.705 4762.720 709.085 4763.810 ;
        RECT 709.925 4762.720 712.305 4763.810 ;
        RECT 713.145 4762.720 724.725 4763.810 ;
        RECT 725.565 4762.720 727.485 4763.810 ;
        RECT 728.325 4762.720 730.705 4763.810 ;
        RECT 731.545 4762.720 733.925 4763.810 ;
        RECT 734.765 4762.720 739.905 4763.810 ;
        RECT 740.745 4762.720 745.885 4763.810 ;
        RECT 746.725 4762.720 749.105 4763.810 ;
        RECT 749.945 4762.720 752.325 4763.810 ;
        RECT 753.165 4762.720 758.305 4763.810 ;
        RECT 759.145 4762.720 944.465 4763.810 ;
        RECT 945.305 4762.720 947.685 4763.810 ;
        RECT 948.525 4762.720 950.905 4763.810 ;
        RECT 951.745 4762.720 960.105 4763.810 ;
        RECT 960.945 4762.720 962.865 4763.810 ;
        RECT 963.705 4762.720 966.085 4763.810 ;
        RECT 966.925 4762.720 969.305 4763.810 ;
        RECT 970.145 4762.720 981.725 4763.810 ;
        RECT 982.565 4762.720 984.485 4763.810 ;
        RECT 985.325 4762.720 987.705 4763.810 ;
        RECT 988.545 4762.720 990.925 4763.810 ;
        RECT 991.765 4762.720 996.905 4763.810 ;
        RECT 997.745 4762.720 1002.885 4763.810 ;
        RECT 1003.725 4762.720 1006.105 4763.810 ;
        RECT 1006.945 4762.720 1009.325 4763.810 ;
        RECT 1010.165 4762.720 1015.305 4763.810 ;
        RECT 1016.145 4762.720 1202.465 4763.810 ;
        RECT 1203.305 4762.720 1205.685 4763.810 ;
        RECT 1206.525 4762.720 1208.905 4763.810 ;
        RECT 1209.745 4762.720 1218.105 4763.810 ;
        RECT 1218.945 4762.720 1220.865 4763.810 ;
        RECT 1221.705 4762.720 1224.085 4763.810 ;
        RECT 1224.925 4762.720 1227.305 4763.810 ;
        RECT 1228.145 4762.720 1239.725 4763.810 ;
        RECT 1240.565 4762.720 1242.485 4763.810 ;
        RECT 1243.325 4762.720 1245.705 4763.810 ;
        RECT 1246.545 4762.720 1248.925 4763.810 ;
        RECT 1249.765 4762.720 1254.905 4763.810 ;
        RECT 1255.745 4762.720 1260.885 4763.810 ;
        RECT 1261.725 4762.720 1264.105 4763.810 ;
        RECT 1264.945 4762.720 1267.325 4763.810 ;
        RECT 1268.165 4762.720 1273.305 4763.810 ;
        RECT 1274.145 4762.720 1711.465 4763.810 ;
        RECT 1712.305 4762.720 1714.685 4763.810 ;
        RECT 1715.525 4762.720 1717.905 4763.810 ;
        RECT 1718.745 4762.720 1727.105 4763.810 ;
        RECT 1727.945 4762.720 1729.865 4763.810 ;
        RECT 1730.705 4762.720 1733.085 4763.810 ;
        RECT 1733.925 4762.720 1736.305 4763.810 ;
        RECT 1737.145 4762.720 1748.725 4763.810 ;
        RECT 1749.565 4762.720 1751.485 4763.810 ;
        RECT 1752.325 4762.720 1754.705 4763.810 ;
        RECT 1755.545 4762.720 1757.925 4763.810 ;
        RECT 1758.765 4762.720 1763.905 4763.810 ;
        RECT 1764.745 4762.720 1769.885 4763.810 ;
        RECT 1770.725 4762.720 1773.105 4763.810 ;
        RECT 1773.945 4762.720 1776.325 4763.810 ;
        RECT 1777.165 4762.720 1782.305 4763.810 ;
        RECT 1783.145 4762.720 2156.465 4763.810 ;
        RECT 2157.305 4762.720 2159.685 4763.810 ;
        RECT 2160.525 4762.720 2162.905 4763.810 ;
        RECT 2163.745 4762.720 2172.105 4763.810 ;
        RECT 2172.945 4762.720 2174.865 4763.810 ;
        RECT 2175.705 4762.720 2178.085 4763.810 ;
        RECT 2178.925 4762.720 2181.305 4763.810 ;
        RECT 2182.145 4762.720 2193.725 4763.810 ;
        RECT 2194.565 4762.720 2196.485 4763.810 ;
        RECT 2197.325 4762.720 2199.705 4763.810 ;
        RECT 2200.545 4762.720 2202.925 4763.810 ;
        RECT 2203.765 4762.720 2208.905 4763.810 ;
        RECT 2209.745 4762.720 2214.885 4763.810 ;
        RECT 2215.725 4762.720 2218.105 4763.810 ;
        RECT 2218.945 4762.720 2221.325 4763.810 ;
        RECT 2222.165 4762.720 2227.305 4763.810 ;
        RECT 2228.145 4762.720 2413.465 4763.810 ;
        RECT 2414.305 4762.720 2416.685 4763.810 ;
        RECT 2417.525 4762.720 2419.905 4763.810 ;
        RECT 2420.745 4762.720 2429.105 4763.810 ;
        RECT 2429.945 4762.720 2431.865 4763.810 ;
        RECT 2432.705 4762.720 2435.085 4763.810 ;
        RECT 2435.925 4762.720 2438.305 4763.810 ;
        RECT 2439.145 4762.720 2450.725 4763.810 ;
        RECT 2451.565 4762.720 2453.485 4763.810 ;
        RECT 2454.325 4762.720 2456.705 4763.810 ;
        RECT 2457.545 4762.720 2459.925 4763.810 ;
        RECT 2460.765 4762.720 2465.905 4763.810 ;
        RECT 2466.745 4762.720 2471.885 4763.810 ;
        RECT 2472.725 4762.720 2475.105 4763.810 ;
        RECT 2475.945 4762.720 2478.325 4763.810 ;
        RECT 2479.165 4762.720 2484.305 4763.810 ;
        RECT 2485.145 4762.720 2922.465 4763.810 ;
        RECT 2923.305 4762.720 2925.685 4763.810 ;
        RECT 2926.525 4762.720 2928.905 4763.810 ;
        RECT 2929.745 4762.720 2938.105 4763.810 ;
        RECT 2938.945 4762.720 2940.865 4763.810 ;
        RECT 2941.705 4762.720 2944.085 4763.810 ;
        RECT 2944.925 4762.720 2947.305 4763.810 ;
        RECT 2948.145 4762.720 2959.725 4763.810 ;
        RECT 2960.565 4762.720 2962.485 4763.810 ;
        RECT 2963.325 4762.720 2965.705 4763.810 ;
        RECT 2966.545 4762.720 2968.925 4763.810 ;
        RECT 2969.765 4762.720 2974.905 4763.810 ;
        RECT 2975.745 4762.720 2980.885 4763.810 ;
        RECT 2981.725 4762.720 2984.105 4763.810 ;
        RECT 2984.945 4762.720 2987.325 4763.810 ;
        RECT 2988.165 4762.720 2993.305 4763.810 ;
        RECT 2994.145 4762.720 3159.190 4763.810 ;
        RECT 4.690 4.280 3159.190 4762.720 ;
        RECT 4.690 3.670 496.555 4.280 ;
        RECT 497.395 3.670 724.855 4.280 ;
        RECT 725.695 3.670 758.435 4.280 ;
        RECT 759.275 3.670 1323.055 4.280 ;
        RECT 1323.895 3.670 1329.495 4.280 ;
        RECT 1330.335 3.670 1338.695 4.280 ;
        RECT 1339.535 3.670 1597.055 4.280 ;
        RECT 1597.895 3.670 1612.695 4.280 ;
        RECT 1613.535 3.670 1815.855 4.280 ;
        RECT 1816.695 3.670 1849.435 4.280 ;
        RECT 1850.275 3.670 1871.055 4.280 ;
        RECT 1871.895 3.670 1886.695 4.280 ;
        RECT 1887.535 3.670 2089.855 4.280 ;
        RECT 2090.695 3.670 2123.435 4.280 ;
        RECT 2124.275 3.670 2145.055 4.280 ;
        RECT 2145.895 3.670 2160.695 4.280 ;
        RECT 2161.535 3.670 2363.855 4.280 ;
        RECT 2364.695 3.670 2391.455 4.280 ;
        RECT 2392.295 3.670 2397.435 4.280 ;
        RECT 2398.275 3.670 2413.075 4.280 ;
        RECT 2413.915 3.670 2419.055 4.280 ;
        RECT 2419.895 3.670 2434.695 4.280 ;
        RECT 2435.535 3.670 3159.190 4.280 ;
      LAYER met3 ;
        RECT 0.000 4763.400 2666.935 4767.000 ;
      LAYER met3 ;
        RECT 2666.935 4763.400 2690.965 4777.980 ;
      LAYER met3 ;
        RECT 2690.965 4763.400 2716.840 4767.000 ;
      LAYER met3 ;
        RECT 2716.840 4763.400 2740.870 4777.980 ;
      LAYER met3 ;
        RECT 2740.870 4763.400 3165.000 4767.000 ;
        RECT 0.000 4636.425 3165.000 4763.400 ;
        RECT 4.400 4635.025 3165.000 4636.425 ;
        RECT 0.000 4630.445 3165.000 4635.025 ;
        RECT 4.400 4629.045 3165.000 4630.445 ;
        RECT 0.000 4627.225 3165.000 4629.045 ;
        RECT 4.400 4625.825 3165.000 4627.225 ;
        RECT 0.000 4624.005 3165.000 4625.825 ;
        RECT 4.400 4623.815 3165.000 4624.005 ;
        RECT 4.400 4622.605 3160.600 4623.815 ;
        RECT 0.000 4622.415 3160.600 4622.605 ;
        RECT 0.000 4620.595 3165.000 4622.415 ;
        RECT 0.000 4619.195 3160.600 4620.595 ;
        RECT 0.000 4618.025 3165.000 4619.195 ;
        RECT 4.400 4617.375 3165.000 4618.025 ;
        RECT 4.400 4616.625 3160.600 4617.375 ;
        RECT 0.000 4615.975 3160.600 4616.625 ;
        RECT 0.000 4612.045 3165.000 4615.975 ;
        RECT 4.400 4610.645 3165.000 4612.045 ;
        RECT 0.000 4608.825 3165.000 4610.645 ;
        RECT 4.400 4608.175 3165.000 4608.825 ;
        RECT 4.400 4607.425 3160.600 4608.175 ;
        RECT 0.000 4606.775 3160.600 4607.425 ;
        RECT 0.000 4605.605 3165.000 4606.775 ;
        RECT 4.400 4605.415 3165.000 4605.605 ;
        RECT 4.400 4604.205 3160.600 4605.415 ;
        RECT 0.000 4604.015 3160.600 4604.205 ;
        RECT 0.000 4602.845 3165.000 4604.015 ;
        RECT 4.400 4602.195 3165.000 4602.845 ;
        RECT 4.400 4601.445 3160.600 4602.195 ;
        RECT 0.000 4600.795 3160.600 4601.445 ;
        RECT 0.000 4598.975 3165.000 4600.795 ;
        RECT 0.000 4597.575 3160.600 4598.975 ;
        RECT 0.000 4590.425 3165.000 4597.575 ;
        RECT 4.400 4589.025 3165.000 4590.425 ;
        RECT 0.000 4587.205 3165.000 4589.025 ;
        RECT 4.400 4586.555 3165.000 4587.205 ;
        RECT 4.400 4585.805 3160.600 4586.555 ;
        RECT 0.000 4585.155 3160.600 4585.805 ;
        RECT 0.000 4583.985 3165.000 4585.155 ;
        RECT 4.400 4583.795 3165.000 4583.985 ;
        RECT 4.400 4582.585 3160.600 4583.795 ;
        RECT 0.000 4582.395 3160.600 4582.585 ;
        RECT 0.000 4581.225 3165.000 4582.395 ;
        RECT 4.400 4580.575 3165.000 4581.225 ;
        RECT 4.400 4579.825 3160.600 4580.575 ;
        RECT 0.000 4579.175 3160.600 4579.825 ;
        RECT 0.000 4577.355 3165.000 4579.175 ;
        RECT 0.000 4575.955 3160.600 4577.355 ;
        RECT 0.000 4572.025 3165.000 4575.955 ;
        RECT 4.400 4571.375 3165.000 4572.025 ;
        RECT 4.400 4570.625 3160.600 4571.375 ;
        RECT 0.000 4569.975 3160.600 4570.625 ;
        RECT 0.000 4568.805 3165.000 4569.975 ;
        RECT 4.400 4567.405 3165.000 4568.805 ;
        RECT 0.000 4565.585 3165.000 4567.405 ;
        RECT 4.400 4565.395 3165.000 4565.585 ;
        RECT 4.400 4564.185 3160.600 4565.395 ;
        RECT 0.000 4563.995 3160.600 4564.185 ;
        RECT 0.000 4562.175 3165.000 4563.995 ;
        RECT 0.000 4560.775 3160.600 4562.175 ;
        RECT 0.000 4558.955 3165.000 4560.775 ;
        RECT 0.000 4557.555 3160.600 4558.955 ;
        RECT 0.000 4552.975 3165.000 4557.555 ;
        RECT 0.000 4551.575 3160.600 4552.975 ;
        RECT 0.000 4424.200 3165.000 4551.575 ;
      LAYER met3 ;
        RECT -16.080 4400.255 5.910 4424.200 ;
      LAYER met3 ;
        RECT 5.910 4402.000 3165.000 4424.200 ;
        RECT 5.910 4400.255 3156.030 4402.000 ;
        RECT 0.000 4398.650 3156.030 4400.255 ;
      LAYER met3 ;
        RECT -11.000 4375.600 5.910 4398.650 ;
      LAYER met3 ;
        RECT 5.910 4378.055 3156.030 4398.650 ;
      LAYER met3 ;
        RECT 3156.030 4378.055 3178.020 4402.000 ;
      LAYER met3 ;
        RECT 5.910 4376.450 3165.000 4378.055 ;
        RECT 5.910 4375.600 3156.030 4376.450 ;
        RECT 0.000 4374.000 3156.030 4375.600 ;
      LAYER met3 ;
        RECT -16.080 4350.055 5.910 4374.000 ;
      LAYER met3 ;
        RECT 5.910 4353.345 3156.030 4374.000 ;
      LAYER met3 ;
        RECT 3156.030 4353.345 3176.020 4376.450 ;
      LAYER met3 ;
        RECT 5.910 4351.745 3165.000 4353.345 ;
        RECT 5.910 4350.055 3156.030 4351.745 ;
        RECT 0.000 4327.800 3156.030 4350.055 ;
      LAYER met3 ;
        RECT 3156.030 4327.800 3178.020 4351.745 ;
      LAYER met3 ;
        RECT 0.000 4177.815 3165.000 4327.800 ;
        RECT 0.000 4176.415 3160.600 4177.815 ;
        RECT 0.000 4174.595 3165.000 4176.415 ;
        RECT 0.000 4173.195 3160.600 4174.595 ;
        RECT 0.000 4171.375 3165.000 4173.195 ;
        RECT 0.000 4169.975 3160.600 4171.375 ;
        RECT 0.000 4162.175 3165.000 4169.975 ;
        RECT 0.000 4160.775 3160.600 4162.175 ;
        RECT 0.000 4159.415 3165.000 4160.775 ;
        RECT 0.000 4158.015 3160.600 4159.415 ;
        RECT 0.000 4156.195 3165.000 4158.015 ;
        RECT 0.000 4154.795 3160.600 4156.195 ;
        RECT 0.000 4152.975 3165.000 4154.795 ;
        RECT 0.000 4151.575 3160.600 4152.975 ;
        RECT 0.000 4140.555 3165.000 4151.575 ;
        RECT 0.000 4139.155 3160.600 4140.555 ;
        RECT 0.000 4137.795 3165.000 4139.155 ;
        RECT 0.000 4136.395 3160.600 4137.795 ;
        RECT 0.000 4134.575 3165.000 4136.395 ;
        RECT 0.000 4133.175 3160.600 4134.575 ;
        RECT 0.000 4131.355 3165.000 4133.175 ;
        RECT 0.000 4129.955 3160.600 4131.355 ;
        RECT 0.000 4125.375 3165.000 4129.955 ;
        RECT 0.000 4123.975 3160.600 4125.375 ;
        RECT 0.000 4119.395 3165.000 4123.975 ;
        RECT 0.000 4117.995 3160.600 4119.395 ;
        RECT 0.000 4116.175 3165.000 4117.995 ;
        RECT 0.000 4114.775 3160.600 4116.175 ;
        RECT 0.000 4112.955 3165.000 4114.775 ;
        RECT 0.000 4111.555 3160.600 4112.955 ;
        RECT 0.000 4106.975 3165.000 4111.555 ;
        RECT 0.000 4105.575 3160.600 4106.975 ;
        RECT 0.000 4001.790 3165.000 4105.575 ;
      LAYER met3 ;
        RECT -16.080 3977.845 5.910 4001.790 ;
      LAYER met3 ;
        RECT 5.910 3977.845 3165.000 4001.790 ;
        RECT 0.000 3956.005 3165.000 3977.845 ;
        RECT 0.000 3951.895 3156.030 3956.005 ;
      LAYER met3 ;
        RECT -16.080 3927.950 5.910 3951.895 ;
      LAYER met3 ;
        RECT 5.910 3932.060 3156.030 3951.895 ;
      LAYER met3 ;
        RECT 3156.030 3932.060 3178.020 3956.005 ;
      LAYER met3 ;
        RECT 5.910 3927.950 3165.000 3932.060 ;
        RECT 0.000 3906.090 3165.000 3927.950 ;
        RECT 0.000 3882.145 3156.030 3906.090 ;
      LAYER met3 ;
        RECT 3156.030 3882.145 3178.020 3906.090 ;
      LAYER met3 ;
        RECT 0.000 3787.425 3165.000 3882.145 ;
        RECT 4.400 3786.025 3165.000 3787.425 ;
        RECT 0.000 3781.445 3165.000 3786.025 ;
        RECT 4.400 3780.045 3165.000 3781.445 ;
        RECT 0.000 3778.225 3165.000 3780.045 ;
        RECT 4.400 3776.825 3165.000 3778.225 ;
        RECT 0.000 3775.005 3165.000 3776.825 ;
        RECT 4.400 3773.605 3165.000 3775.005 ;
        RECT 0.000 3769.025 3165.000 3773.605 ;
        RECT 4.400 3767.625 3165.000 3769.025 ;
        RECT 0.000 3763.045 3165.000 3767.625 ;
        RECT 4.400 3761.645 3165.000 3763.045 ;
        RECT 0.000 3759.825 3165.000 3761.645 ;
        RECT 4.400 3758.425 3165.000 3759.825 ;
        RECT 0.000 3756.605 3165.000 3758.425 ;
        RECT 4.400 3755.205 3165.000 3756.605 ;
        RECT 0.000 3753.845 3165.000 3755.205 ;
        RECT 4.400 3752.445 3165.000 3753.845 ;
        RECT 0.000 3741.425 3165.000 3752.445 ;
        RECT 4.400 3740.025 3165.000 3741.425 ;
        RECT 0.000 3738.205 3165.000 3740.025 ;
        RECT 4.400 3736.805 3165.000 3738.205 ;
        RECT 0.000 3734.985 3165.000 3736.805 ;
        RECT 4.400 3733.585 3165.000 3734.985 ;
        RECT 0.000 3732.225 3165.000 3733.585 ;
        RECT 4.400 3731.815 3165.000 3732.225 ;
        RECT 4.400 3730.825 3160.600 3731.815 ;
        RECT 0.000 3730.415 3160.600 3730.825 ;
        RECT 0.000 3728.595 3165.000 3730.415 ;
        RECT 0.000 3727.195 3160.600 3728.595 ;
        RECT 0.000 3725.375 3165.000 3727.195 ;
        RECT 0.000 3723.975 3160.600 3725.375 ;
        RECT 0.000 3723.025 3165.000 3723.975 ;
        RECT 4.400 3721.625 3165.000 3723.025 ;
        RECT 0.000 3719.805 3165.000 3721.625 ;
        RECT 4.400 3718.405 3165.000 3719.805 ;
        RECT 0.000 3716.585 3165.000 3718.405 ;
        RECT 4.400 3716.175 3165.000 3716.585 ;
        RECT 4.400 3715.185 3160.600 3716.175 ;
        RECT 0.000 3714.775 3160.600 3715.185 ;
        RECT 0.000 3713.415 3165.000 3714.775 ;
        RECT 0.000 3712.015 3160.600 3713.415 ;
        RECT 0.000 3710.195 3165.000 3712.015 ;
        RECT 0.000 3708.795 3160.600 3710.195 ;
        RECT 0.000 3706.975 3165.000 3708.795 ;
        RECT 0.000 3705.575 3160.600 3706.975 ;
        RECT 0.000 3694.555 3165.000 3705.575 ;
        RECT 0.000 3693.155 3160.600 3694.555 ;
        RECT 0.000 3691.795 3165.000 3693.155 ;
        RECT 0.000 3690.395 3160.600 3691.795 ;
        RECT 0.000 3688.575 3165.000 3690.395 ;
        RECT 0.000 3687.175 3160.600 3688.575 ;
        RECT 0.000 3685.355 3165.000 3687.175 ;
        RECT 0.000 3683.955 3160.600 3685.355 ;
        RECT 0.000 3679.375 3165.000 3683.955 ;
        RECT 0.000 3677.975 3160.600 3679.375 ;
        RECT 0.000 3673.395 3165.000 3677.975 ;
        RECT 0.000 3671.995 3160.600 3673.395 ;
        RECT 0.000 3670.175 3165.000 3671.995 ;
        RECT 0.000 3668.775 3160.600 3670.175 ;
        RECT 0.000 3666.955 3165.000 3668.775 ;
        RECT 0.000 3665.555 3160.600 3666.955 ;
        RECT 0.000 3660.975 3165.000 3665.555 ;
        RECT 0.000 3659.575 3160.600 3660.975 ;
        RECT 0.000 3571.425 3165.000 3659.575 ;
        RECT 4.400 3570.025 3165.000 3571.425 ;
        RECT 0.000 3565.445 3165.000 3570.025 ;
        RECT 4.400 3564.045 3165.000 3565.445 ;
        RECT 0.000 3562.225 3165.000 3564.045 ;
        RECT 4.400 3560.825 3165.000 3562.225 ;
        RECT 0.000 3559.005 3165.000 3560.825 ;
        RECT 4.400 3557.605 3165.000 3559.005 ;
        RECT 0.000 3553.025 3165.000 3557.605 ;
        RECT 4.400 3551.625 3165.000 3553.025 ;
        RECT 0.000 3547.045 3165.000 3551.625 ;
        RECT 4.400 3545.645 3165.000 3547.045 ;
        RECT 0.000 3543.825 3165.000 3545.645 ;
        RECT 4.400 3542.425 3165.000 3543.825 ;
        RECT 0.000 3540.605 3165.000 3542.425 ;
        RECT 4.400 3539.205 3165.000 3540.605 ;
        RECT 0.000 3537.845 3165.000 3539.205 ;
        RECT 4.400 3536.445 3165.000 3537.845 ;
        RECT 0.000 3525.425 3165.000 3536.445 ;
        RECT 4.400 3524.025 3165.000 3525.425 ;
        RECT 0.000 3522.205 3165.000 3524.025 ;
        RECT 4.400 3520.805 3165.000 3522.205 ;
        RECT 0.000 3518.985 3165.000 3520.805 ;
        RECT 4.400 3517.585 3165.000 3518.985 ;
        RECT 0.000 3516.225 3165.000 3517.585 ;
        RECT 4.400 3514.825 3165.000 3516.225 ;
        RECT 0.000 3507.025 3165.000 3514.825 ;
        RECT 4.400 3506.815 3165.000 3507.025 ;
        RECT 4.400 3505.625 3160.600 3506.815 ;
        RECT 0.000 3505.415 3160.600 3505.625 ;
        RECT 0.000 3503.805 3165.000 3505.415 ;
        RECT 4.400 3503.595 3165.000 3503.805 ;
        RECT 4.400 3502.405 3160.600 3503.595 ;
        RECT 0.000 3502.195 3160.600 3502.405 ;
        RECT 0.000 3500.585 3165.000 3502.195 ;
        RECT 4.400 3500.375 3165.000 3500.585 ;
        RECT 4.400 3499.185 3160.600 3500.375 ;
        RECT 0.000 3498.975 3160.600 3499.185 ;
        RECT 0.000 3491.175 3165.000 3498.975 ;
        RECT 0.000 3489.775 3160.600 3491.175 ;
        RECT 0.000 3488.415 3165.000 3489.775 ;
        RECT 0.000 3487.015 3160.600 3488.415 ;
        RECT 0.000 3485.195 3165.000 3487.015 ;
        RECT 0.000 3483.795 3160.600 3485.195 ;
        RECT 0.000 3481.975 3165.000 3483.795 ;
        RECT 0.000 3480.575 3160.600 3481.975 ;
        RECT 0.000 3469.555 3165.000 3480.575 ;
        RECT 0.000 3468.155 3160.600 3469.555 ;
        RECT 0.000 3466.795 3165.000 3468.155 ;
        RECT 0.000 3465.395 3160.600 3466.795 ;
        RECT 0.000 3463.575 3165.000 3465.395 ;
        RECT 0.000 3462.175 3160.600 3463.575 ;
        RECT 0.000 3460.355 3165.000 3462.175 ;
        RECT 0.000 3458.955 3160.600 3460.355 ;
        RECT 0.000 3454.375 3165.000 3458.955 ;
        RECT 0.000 3452.975 3160.600 3454.375 ;
        RECT 0.000 3448.395 3165.000 3452.975 ;
        RECT 0.000 3446.995 3160.600 3448.395 ;
        RECT 0.000 3445.175 3165.000 3446.995 ;
        RECT 0.000 3443.775 3160.600 3445.175 ;
        RECT 0.000 3441.955 3165.000 3443.775 ;
        RECT 0.000 3440.555 3160.600 3441.955 ;
        RECT 0.000 3435.975 3165.000 3440.555 ;
        RECT 0.000 3434.575 3160.600 3435.975 ;
        RECT 0.000 3355.425 3165.000 3434.575 ;
        RECT 4.400 3354.025 3165.000 3355.425 ;
        RECT 0.000 3349.445 3165.000 3354.025 ;
        RECT 4.400 3348.045 3165.000 3349.445 ;
        RECT 0.000 3346.225 3165.000 3348.045 ;
        RECT 4.400 3344.825 3165.000 3346.225 ;
        RECT 0.000 3343.005 3165.000 3344.825 ;
        RECT 4.400 3341.605 3165.000 3343.005 ;
        RECT 0.000 3337.025 3165.000 3341.605 ;
        RECT 4.400 3335.625 3165.000 3337.025 ;
        RECT 0.000 3331.045 3165.000 3335.625 ;
        RECT 4.400 3329.645 3165.000 3331.045 ;
        RECT 0.000 3327.825 3165.000 3329.645 ;
        RECT 4.400 3326.425 3165.000 3327.825 ;
        RECT 0.000 3324.605 3165.000 3326.425 ;
        RECT 4.400 3323.205 3165.000 3324.605 ;
        RECT 0.000 3321.845 3165.000 3323.205 ;
        RECT 4.400 3320.445 3165.000 3321.845 ;
        RECT 0.000 3309.425 3165.000 3320.445 ;
        RECT 4.400 3308.025 3165.000 3309.425 ;
        RECT 0.000 3306.205 3165.000 3308.025 ;
        RECT 4.400 3304.805 3165.000 3306.205 ;
        RECT 0.000 3302.985 3165.000 3304.805 ;
        RECT 4.400 3301.585 3165.000 3302.985 ;
        RECT 0.000 3300.225 3165.000 3301.585 ;
        RECT 4.400 3298.825 3165.000 3300.225 ;
        RECT 0.000 3291.025 3165.000 3298.825 ;
        RECT 4.400 3289.625 3165.000 3291.025 ;
        RECT 0.000 3287.805 3165.000 3289.625 ;
        RECT 4.400 3286.405 3165.000 3287.805 ;
        RECT 0.000 3284.585 3165.000 3286.405 ;
        RECT 4.400 3283.185 3165.000 3284.585 ;
        RECT 0.000 3281.815 3165.000 3283.185 ;
        RECT 0.000 3280.415 3160.600 3281.815 ;
        RECT 0.000 3278.595 3165.000 3280.415 ;
        RECT 0.000 3277.195 3160.600 3278.595 ;
        RECT 0.000 3275.375 3165.000 3277.195 ;
        RECT 0.000 3273.975 3160.600 3275.375 ;
        RECT 0.000 3266.175 3165.000 3273.975 ;
        RECT 0.000 3264.775 3160.600 3266.175 ;
        RECT 0.000 3263.415 3165.000 3264.775 ;
        RECT 0.000 3262.015 3160.600 3263.415 ;
        RECT 0.000 3260.195 3165.000 3262.015 ;
        RECT 0.000 3258.795 3160.600 3260.195 ;
        RECT 0.000 3256.975 3165.000 3258.795 ;
        RECT 0.000 3255.575 3160.600 3256.975 ;
        RECT 0.000 3244.555 3165.000 3255.575 ;
        RECT 0.000 3243.155 3160.600 3244.555 ;
        RECT 0.000 3241.795 3165.000 3243.155 ;
        RECT 0.000 3240.395 3160.600 3241.795 ;
        RECT 0.000 3238.575 3165.000 3240.395 ;
        RECT 0.000 3237.175 3160.600 3238.575 ;
        RECT 0.000 3235.355 3165.000 3237.175 ;
        RECT 0.000 3233.955 3160.600 3235.355 ;
        RECT 0.000 3229.375 3165.000 3233.955 ;
        RECT 0.000 3227.975 3160.600 3229.375 ;
        RECT 0.000 3223.395 3165.000 3227.975 ;
        RECT 0.000 3221.995 3160.600 3223.395 ;
        RECT 0.000 3220.175 3165.000 3221.995 ;
        RECT 0.000 3218.775 3160.600 3220.175 ;
        RECT 0.000 3216.955 3165.000 3218.775 ;
        RECT 0.000 3215.555 3160.600 3216.955 ;
        RECT 0.000 3210.975 3165.000 3215.555 ;
        RECT 0.000 3209.575 3160.600 3210.975 ;
        RECT 0.000 3139.425 3165.000 3209.575 ;
        RECT 4.400 3138.025 3165.000 3139.425 ;
        RECT 0.000 3133.445 3165.000 3138.025 ;
        RECT 4.400 3132.045 3165.000 3133.445 ;
        RECT 0.000 3130.225 3165.000 3132.045 ;
        RECT 4.400 3128.825 3165.000 3130.225 ;
        RECT 0.000 3127.005 3165.000 3128.825 ;
        RECT 4.400 3125.605 3165.000 3127.005 ;
        RECT 0.000 3121.025 3165.000 3125.605 ;
        RECT 4.400 3119.625 3165.000 3121.025 ;
        RECT 0.000 3115.045 3165.000 3119.625 ;
        RECT 4.690 3113.645 3165.000 3115.045 ;
        RECT 0.000 3111.825 3165.000 3113.645 ;
        RECT 4.400 3110.425 3165.000 3111.825 ;
        RECT 0.000 3108.605 3165.000 3110.425 ;
        RECT 4.400 3107.205 3165.000 3108.605 ;
        RECT 0.000 3105.845 3165.000 3107.205 ;
        RECT 4.400 3104.445 3165.000 3105.845 ;
        RECT 0.000 3093.425 3165.000 3104.445 ;
        RECT 4.400 3092.025 3165.000 3093.425 ;
        RECT 0.000 3090.205 3165.000 3092.025 ;
        RECT 4.400 3088.805 3165.000 3090.205 ;
        RECT 0.000 3086.985 3165.000 3088.805 ;
        RECT 4.400 3085.585 3165.000 3086.985 ;
        RECT 0.000 3084.225 3165.000 3085.585 ;
        RECT 4.400 3082.825 3165.000 3084.225 ;
        RECT 0.000 3075.025 3165.000 3082.825 ;
        RECT 4.400 3073.625 3165.000 3075.025 ;
        RECT 0.000 3071.805 3165.000 3073.625 ;
        RECT 4.400 3070.405 3165.000 3071.805 ;
        RECT 0.000 3068.585 3165.000 3070.405 ;
        RECT 4.400 3067.185 3165.000 3068.585 ;
        RECT 0.000 3055.815 3165.000 3067.185 ;
        RECT 0.000 3054.415 3160.600 3055.815 ;
        RECT 0.000 3052.595 3165.000 3054.415 ;
        RECT 0.000 3051.195 3160.600 3052.595 ;
        RECT 0.000 3049.375 3165.000 3051.195 ;
        RECT 0.000 3047.975 3160.600 3049.375 ;
        RECT 0.000 3040.175 3165.000 3047.975 ;
        RECT 0.000 3038.775 3160.600 3040.175 ;
        RECT 0.000 3037.415 3165.000 3038.775 ;
        RECT 0.000 3036.015 3160.600 3037.415 ;
        RECT 0.000 3034.195 3165.000 3036.015 ;
        RECT 0.000 3032.795 3160.600 3034.195 ;
        RECT 0.000 3030.975 3165.000 3032.795 ;
        RECT 0.000 3029.575 3160.600 3030.975 ;
        RECT 0.000 3018.555 3165.000 3029.575 ;
        RECT 0.000 3017.155 3160.600 3018.555 ;
        RECT 0.000 3015.795 3165.000 3017.155 ;
        RECT 0.000 3014.395 3160.600 3015.795 ;
        RECT 0.000 3012.575 3165.000 3014.395 ;
        RECT 0.000 3011.175 3160.600 3012.575 ;
        RECT 0.000 3009.355 3165.000 3011.175 ;
        RECT 0.000 3007.955 3160.600 3009.355 ;
        RECT 0.000 3003.375 3165.000 3007.955 ;
        RECT 0.000 3001.975 3160.600 3003.375 ;
        RECT 0.000 2997.395 3165.000 3001.975 ;
        RECT 0.000 2995.995 3160.600 2997.395 ;
        RECT 0.000 2994.175 3165.000 2995.995 ;
        RECT 0.000 2992.775 3160.600 2994.175 ;
        RECT 0.000 2990.955 3165.000 2992.775 ;
        RECT 0.000 2989.555 3160.600 2990.955 ;
        RECT 0.000 2984.975 3165.000 2989.555 ;
        RECT 0.000 2983.575 3160.600 2984.975 ;
        RECT 0.000 2923.425 3165.000 2983.575 ;
        RECT 4.400 2922.025 3165.000 2923.425 ;
        RECT 0.000 2917.445 3165.000 2922.025 ;
        RECT 4.400 2916.045 3165.000 2917.445 ;
        RECT 0.000 2914.225 3165.000 2916.045 ;
        RECT 4.400 2912.825 3165.000 2914.225 ;
        RECT 0.000 2911.005 3165.000 2912.825 ;
        RECT 4.400 2909.605 3165.000 2911.005 ;
        RECT 0.000 2905.025 3165.000 2909.605 ;
        RECT 4.400 2903.625 3165.000 2905.025 ;
        RECT 0.000 2899.045 3165.000 2903.625 ;
        RECT 4.400 2897.645 3165.000 2899.045 ;
        RECT 0.000 2895.825 3165.000 2897.645 ;
        RECT 4.400 2894.425 3165.000 2895.825 ;
        RECT 0.000 2892.605 3165.000 2894.425 ;
        RECT 4.400 2891.205 3165.000 2892.605 ;
        RECT 0.000 2889.845 3165.000 2891.205 ;
        RECT 4.400 2888.445 3165.000 2889.845 ;
        RECT 0.000 2877.425 3165.000 2888.445 ;
        RECT 4.400 2876.025 3165.000 2877.425 ;
        RECT 0.000 2874.205 3165.000 2876.025 ;
        RECT 4.400 2872.805 3165.000 2874.205 ;
        RECT 0.000 2870.985 3165.000 2872.805 ;
        RECT 4.400 2869.585 3165.000 2870.985 ;
        RECT 0.000 2868.225 3165.000 2869.585 ;
        RECT 4.400 2866.825 3165.000 2868.225 ;
        RECT 0.000 2859.025 3165.000 2866.825 ;
        RECT 4.400 2857.625 3165.000 2859.025 ;
        RECT 0.000 2855.805 3165.000 2857.625 ;
        RECT 4.400 2854.405 3165.000 2855.805 ;
        RECT 0.000 2852.585 3165.000 2854.405 ;
        RECT 4.400 2851.185 3165.000 2852.585 ;
        RECT 0.000 2830.815 3165.000 2851.185 ;
        RECT 0.000 2829.415 3160.600 2830.815 ;
        RECT 0.000 2827.595 3165.000 2829.415 ;
        RECT 0.000 2826.195 3160.600 2827.595 ;
        RECT 0.000 2824.375 3165.000 2826.195 ;
        RECT 0.000 2822.975 3160.600 2824.375 ;
        RECT 0.000 2815.175 3165.000 2822.975 ;
        RECT 0.000 2813.775 3160.600 2815.175 ;
        RECT 0.000 2812.415 3165.000 2813.775 ;
        RECT 0.000 2811.015 3160.600 2812.415 ;
        RECT 0.000 2809.195 3165.000 2811.015 ;
        RECT 0.000 2807.795 3160.600 2809.195 ;
        RECT 0.000 2805.975 3165.000 2807.795 ;
        RECT 0.000 2804.575 3160.600 2805.975 ;
        RECT 0.000 2793.555 3165.000 2804.575 ;
        RECT 0.000 2792.155 3160.600 2793.555 ;
        RECT 0.000 2790.795 3165.000 2792.155 ;
        RECT 0.000 2789.395 3160.600 2790.795 ;
        RECT 0.000 2787.575 3165.000 2789.395 ;
        RECT 0.000 2786.175 3160.600 2787.575 ;
        RECT 0.000 2784.355 3165.000 2786.175 ;
        RECT 0.000 2782.955 3160.600 2784.355 ;
        RECT 0.000 2778.375 3165.000 2782.955 ;
        RECT 0.000 2776.975 3160.600 2778.375 ;
        RECT 0.000 2772.395 3165.000 2776.975 ;
        RECT 0.000 2770.995 3160.600 2772.395 ;
        RECT 0.000 2769.175 3165.000 2770.995 ;
        RECT 0.000 2767.775 3160.600 2769.175 ;
        RECT 0.000 2765.955 3165.000 2767.775 ;
        RECT 0.000 2764.555 3160.600 2765.955 ;
        RECT 0.000 2759.975 3165.000 2764.555 ;
        RECT 0.000 2758.575 3160.600 2759.975 ;
        RECT 0.000 2707.425 3165.000 2758.575 ;
        RECT 4.400 2706.025 3165.000 2707.425 ;
        RECT 0.000 2701.445 3165.000 2706.025 ;
        RECT 4.400 2700.045 3165.000 2701.445 ;
        RECT 0.000 2698.225 3165.000 2700.045 ;
        RECT 4.400 2696.825 3165.000 2698.225 ;
        RECT 0.000 2695.005 3165.000 2696.825 ;
        RECT 4.400 2693.605 3165.000 2695.005 ;
        RECT 0.000 2689.025 3165.000 2693.605 ;
        RECT 4.400 2687.625 3165.000 2689.025 ;
        RECT 0.000 2683.045 3165.000 2687.625 ;
        RECT 4.400 2681.645 3165.000 2683.045 ;
        RECT 0.000 2679.825 3165.000 2681.645 ;
        RECT 4.400 2678.425 3165.000 2679.825 ;
        RECT 0.000 2676.605 3165.000 2678.425 ;
        RECT 4.400 2675.205 3165.000 2676.605 ;
        RECT 0.000 2673.845 3165.000 2675.205 ;
        RECT 4.400 2672.445 3165.000 2673.845 ;
        RECT 0.000 2661.425 3165.000 2672.445 ;
        RECT 4.400 2660.025 3165.000 2661.425 ;
        RECT 0.000 2658.205 3165.000 2660.025 ;
        RECT 4.400 2656.805 3165.000 2658.205 ;
        RECT 0.000 2654.985 3165.000 2656.805 ;
        RECT 4.400 2653.585 3165.000 2654.985 ;
        RECT 0.000 2652.225 3165.000 2653.585 ;
        RECT 4.400 2650.825 3165.000 2652.225 ;
        RECT 0.000 2643.025 3165.000 2650.825 ;
        RECT 4.400 2641.625 3165.000 2643.025 ;
        RECT 0.000 2639.805 3165.000 2641.625 ;
        RECT 4.400 2638.405 3165.000 2639.805 ;
        RECT 0.000 2636.585 3165.000 2638.405 ;
        RECT 4.400 2635.185 3165.000 2636.585 ;
        RECT 0.000 2604.815 3165.000 2635.185 ;
        RECT 0.000 2603.415 3160.600 2604.815 ;
        RECT 0.000 2601.595 3165.000 2603.415 ;
        RECT 0.000 2600.195 3160.600 2601.595 ;
        RECT 0.000 2598.375 3165.000 2600.195 ;
        RECT 0.000 2596.975 3160.600 2598.375 ;
        RECT 0.000 2589.175 3165.000 2596.975 ;
        RECT 0.000 2587.775 3160.600 2589.175 ;
        RECT 0.000 2586.415 3165.000 2587.775 ;
        RECT 0.000 2585.015 3160.600 2586.415 ;
        RECT 0.000 2583.195 3165.000 2585.015 ;
        RECT 0.000 2581.795 3160.600 2583.195 ;
        RECT 0.000 2579.975 3165.000 2581.795 ;
        RECT 0.000 2578.575 3160.600 2579.975 ;
        RECT 0.000 2567.555 3165.000 2578.575 ;
        RECT 0.000 2566.155 3160.600 2567.555 ;
        RECT 0.000 2564.795 3165.000 2566.155 ;
        RECT 0.000 2563.395 3160.600 2564.795 ;
        RECT 0.000 2561.575 3165.000 2563.395 ;
        RECT 0.000 2560.175 3160.600 2561.575 ;
        RECT 0.000 2558.355 3165.000 2560.175 ;
        RECT 0.000 2556.955 3160.600 2558.355 ;
        RECT 0.000 2552.375 3165.000 2556.955 ;
        RECT 0.000 2550.975 3160.600 2552.375 ;
        RECT 0.000 2546.395 3165.000 2550.975 ;
        RECT 0.000 2544.995 3160.600 2546.395 ;
        RECT 0.000 2543.175 3165.000 2544.995 ;
        RECT 0.000 2541.775 3160.600 2543.175 ;
        RECT 0.000 2539.955 3165.000 2541.775 ;
        RECT 0.000 2538.555 3160.600 2539.955 ;
        RECT 0.000 2533.975 3165.000 2538.555 ;
        RECT 0.000 2532.575 3160.600 2533.975 ;
        RECT 0.000 2491.425 3165.000 2532.575 ;
        RECT 4.400 2490.025 3165.000 2491.425 ;
        RECT 0.000 2485.445 3165.000 2490.025 ;
        RECT 4.400 2484.045 3165.000 2485.445 ;
        RECT 0.000 2482.225 3165.000 2484.045 ;
        RECT 4.400 2480.825 3165.000 2482.225 ;
        RECT 0.000 2479.005 3165.000 2480.825 ;
        RECT 4.400 2477.605 3165.000 2479.005 ;
        RECT 0.000 2473.025 3165.000 2477.605 ;
        RECT 4.400 2471.625 3165.000 2473.025 ;
        RECT 0.000 2467.045 3165.000 2471.625 ;
        RECT 4.400 2465.645 3165.000 2467.045 ;
        RECT 0.000 2463.825 3165.000 2465.645 ;
        RECT 4.400 2462.425 3165.000 2463.825 ;
        RECT 0.000 2460.605 3165.000 2462.425 ;
        RECT 4.400 2459.205 3165.000 2460.605 ;
        RECT 0.000 2457.845 3165.000 2459.205 ;
        RECT 4.400 2456.445 3165.000 2457.845 ;
        RECT 0.000 2445.425 3165.000 2456.445 ;
        RECT 4.400 2444.025 3165.000 2445.425 ;
        RECT 0.000 2442.205 3165.000 2444.025 ;
        RECT 4.400 2440.805 3165.000 2442.205 ;
        RECT 0.000 2438.985 3165.000 2440.805 ;
        RECT 4.400 2437.585 3165.000 2438.985 ;
        RECT 0.000 2436.225 3165.000 2437.585 ;
        RECT 4.400 2434.825 3165.000 2436.225 ;
        RECT 0.000 2427.025 3165.000 2434.825 ;
        RECT 4.400 2425.625 3165.000 2427.025 ;
        RECT 0.000 2423.805 3165.000 2425.625 ;
        RECT 4.400 2422.405 3165.000 2423.805 ;
        RECT 0.000 2420.585 3165.000 2422.405 ;
        RECT 4.400 2419.185 3165.000 2420.585 ;
        RECT 0.000 2383.005 3165.000 2419.185 ;
        RECT 0.000 2359.060 3156.030 2383.005 ;
      LAYER met3 ;
        RECT 3156.030 2359.060 3178.020 2383.005 ;
      LAYER met3 ;
        RECT 0.000 2333.090 3165.000 2359.060 ;
        RECT 0.000 2309.145 3156.030 2333.090 ;
      LAYER met3 ;
        RECT 3156.030 2309.145 3178.020 2333.090 ;
      LAYER met3 ;
        RECT 0.000 2278.790 3165.000 2309.145 ;
      LAYER met3 ;
        RECT -16.080 2254.845 5.910 2278.790 ;
      LAYER met3 ;
        RECT 5.910 2254.845 3165.000 2278.790 ;
        RECT 0.000 2228.895 3165.000 2254.845 ;
      LAYER met3 ;
        RECT -16.080 2204.950 5.910 2228.895 ;
      LAYER met3 ;
        RECT 5.910 2204.950 3165.000 2228.895 ;
        RECT 0.000 2163.000 3165.000 2204.950 ;
        RECT 0.000 2139.055 3156.030 2163.000 ;
      LAYER met3 ;
        RECT 3156.030 2139.055 3178.020 2163.000 ;
      LAYER met3 ;
        RECT 0.000 2137.450 3165.000 2139.055 ;
        RECT 0.000 2114.345 3156.030 2137.450 ;
      LAYER met3 ;
        RECT 3156.030 2114.345 3176.020 2137.450 ;
      LAYER met3 ;
        RECT 0.000 2112.745 3165.000 2114.345 ;
        RECT 0.000 2088.800 3156.030 2112.745 ;
      LAYER met3 ;
        RECT 3156.030 2088.800 3178.020 2112.745 ;
      LAYER met3 ;
        RECT 0.000 2068.200 3165.000 2088.800 ;
      LAYER met3 ;
        RECT -16.080 2044.255 5.910 2068.200 ;
      LAYER met3 ;
        RECT 5.910 2044.255 3165.000 2068.200 ;
        RECT 0.000 2042.650 3165.000 2044.255 ;
      LAYER met3 ;
        RECT -11.080 2019.600 5.910 2042.650 ;
      LAYER met3 ;
        RECT 5.910 2019.600 3165.000 2042.650 ;
        RECT 0.000 2018.000 3165.000 2019.600 ;
      LAYER met3 ;
        RECT -16.080 1994.055 5.910 2018.000 ;
      LAYER met3 ;
        RECT 5.910 1994.055 3165.000 2018.000 ;
        RECT 0.000 1942.045 3165.000 1994.055 ;
        RECT 0.000 1918.100 3156.030 1942.045 ;
      LAYER met3 ;
        RECT 3156.030 1918.100 3178.020 1942.045 ;
      LAYER met3 ;
        RECT 0.000 1892.130 3165.000 1918.100 ;
        RECT 0.000 1868.185 3156.030 1892.130 ;
      LAYER met3 ;
        RECT 3156.030 1868.185 3178.020 1892.130 ;
      LAYER met3 ;
        RECT 0.000 1853.425 3165.000 1868.185 ;
        RECT 4.400 1852.025 3165.000 1853.425 ;
        RECT 0.000 1847.445 3165.000 1852.025 ;
        RECT 4.400 1846.045 3165.000 1847.445 ;
        RECT 0.000 1844.225 3165.000 1846.045 ;
        RECT 4.400 1842.825 3165.000 1844.225 ;
        RECT 0.000 1841.005 3165.000 1842.825 ;
        RECT 4.400 1839.605 3165.000 1841.005 ;
        RECT 0.000 1835.025 3165.000 1839.605 ;
        RECT 4.400 1833.625 3165.000 1835.025 ;
        RECT 0.000 1829.045 3165.000 1833.625 ;
        RECT 4.400 1827.645 3165.000 1829.045 ;
        RECT 0.000 1825.825 3165.000 1827.645 ;
        RECT 4.400 1824.425 3165.000 1825.825 ;
        RECT 0.000 1822.605 3165.000 1824.425 ;
        RECT 4.400 1821.205 3165.000 1822.605 ;
        RECT 0.000 1819.845 3165.000 1821.205 ;
        RECT 4.400 1818.445 3165.000 1819.845 ;
        RECT 0.000 1807.425 3165.000 1818.445 ;
        RECT 4.400 1806.025 3165.000 1807.425 ;
        RECT 0.000 1804.205 3165.000 1806.025 ;
        RECT 4.400 1802.805 3165.000 1804.205 ;
        RECT 0.000 1800.985 3165.000 1802.805 ;
        RECT 4.400 1799.585 3165.000 1800.985 ;
        RECT 0.000 1798.225 3165.000 1799.585 ;
        RECT 4.400 1796.825 3165.000 1798.225 ;
        RECT 0.000 1789.025 3165.000 1796.825 ;
        RECT 4.400 1787.625 3165.000 1789.025 ;
        RECT 0.000 1785.805 3165.000 1787.625 ;
        RECT 4.400 1784.405 3165.000 1785.805 ;
        RECT 0.000 1782.585 3165.000 1784.405 ;
        RECT 4.400 1781.185 3165.000 1782.585 ;
        RECT 0.000 1718.815 3165.000 1781.185 ;
        RECT 0.000 1717.415 3160.600 1718.815 ;
        RECT 0.000 1715.595 3165.000 1717.415 ;
        RECT 0.000 1714.195 3160.600 1715.595 ;
        RECT 0.000 1712.375 3165.000 1714.195 ;
        RECT 0.000 1710.975 3160.600 1712.375 ;
        RECT 0.000 1703.175 3165.000 1710.975 ;
        RECT 0.000 1701.775 3160.600 1703.175 ;
        RECT 0.000 1700.415 3165.000 1701.775 ;
        RECT 0.000 1699.015 3160.600 1700.415 ;
        RECT 0.000 1697.195 3165.000 1699.015 ;
        RECT 0.000 1695.795 3160.600 1697.195 ;
        RECT 0.000 1693.975 3165.000 1695.795 ;
        RECT 0.000 1692.575 3160.600 1693.975 ;
        RECT 0.000 1681.555 3165.000 1692.575 ;
        RECT 0.000 1680.155 3160.600 1681.555 ;
        RECT 0.000 1678.795 3165.000 1680.155 ;
        RECT 0.000 1677.395 3160.600 1678.795 ;
        RECT 0.000 1675.575 3165.000 1677.395 ;
        RECT 0.000 1674.175 3160.600 1675.575 ;
        RECT 0.000 1672.355 3165.000 1674.175 ;
        RECT 0.000 1670.955 3160.600 1672.355 ;
        RECT 0.000 1666.375 3165.000 1670.955 ;
        RECT 0.000 1664.975 3160.600 1666.375 ;
        RECT 0.000 1657.175 3165.000 1664.975 ;
        RECT 0.000 1655.775 3160.600 1657.175 ;
        RECT 0.000 1653.955 3165.000 1655.775 ;
        RECT 0.000 1652.555 3160.600 1653.955 ;
        RECT 0.000 1647.975 3165.000 1652.555 ;
        RECT 0.000 1646.575 3160.600 1647.975 ;
        RECT 0.000 1637.425 3165.000 1646.575 ;
        RECT 4.400 1636.025 3165.000 1637.425 ;
        RECT 0.000 1631.445 3165.000 1636.025 ;
        RECT 4.400 1630.045 3165.000 1631.445 ;
        RECT 0.000 1628.225 3165.000 1630.045 ;
        RECT 4.400 1626.825 3165.000 1628.225 ;
        RECT 0.000 1625.005 3165.000 1626.825 ;
        RECT 4.400 1623.605 3165.000 1625.005 ;
        RECT 0.000 1619.025 3165.000 1623.605 ;
        RECT 4.400 1617.625 3165.000 1619.025 ;
        RECT 0.000 1613.045 3165.000 1617.625 ;
        RECT 4.400 1611.645 3165.000 1613.045 ;
        RECT 0.000 1609.825 3165.000 1611.645 ;
        RECT 4.400 1608.425 3165.000 1609.825 ;
        RECT 0.000 1606.605 3165.000 1608.425 ;
        RECT 4.400 1605.205 3165.000 1606.605 ;
        RECT 0.000 1603.845 3165.000 1605.205 ;
        RECT 4.400 1602.445 3165.000 1603.845 ;
        RECT 0.000 1591.425 3165.000 1602.445 ;
        RECT 4.400 1590.025 3165.000 1591.425 ;
        RECT 0.000 1588.205 3165.000 1590.025 ;
        RECT 4.400 1586.805 3165.000 1588.205 ;
        RECT 0.000 1584.985 3165.000 1586.805 ;
        RECT 4.400 1583.585 3165.000 1584.985 ;
        RECT 0.000 1582.225 3165.000 1583.585 ;
        RECT 4.400 1580.825 3165.000 1582.225 ;
        RECT 0.000 1573.025 3165.000 1580.825 ;
        RECT 4.400 1571.625 3165.000 1573.025 ;
        RECT 0.000 1569.805 3165.000 1571.625 ;
        RECT 4.400 1568.405 3165.000 1569.805 ;
        RECT 0.000 1566.585 3165.000 1568.405 ;
        RECT 4.400 1565.185 3165.000 1566.585 ;
        RECT 0.000 1492.815 3165.000 1565.185 ;
        RECT 0.000 1491.415 3160.600 1492.815 ;
        RECT 0.000 1489.595 3165.000 1491.415 ;
        RECT 0.000 1488.195 3160.600 1489.595 ;
        RECT 0.000 1486.375 3165.000 1488.195 ;
        RECT 0.000 1484.975 3160.600 1486.375 ;
        RECT 0.000 1477.175 3165.000 1484.975 ;
        RECT 0.000 1475.775 3160.600 1477.175 ;
        RECT 0.000 1474.415 3165.000 1475.775 ;
        RECT 0.000 1473.015 3160.600 1474.415 ;
        RECT 0.000 1471.195 3165.000 1473.015 ;
        RECT 0.000 1469.795 3160.600 1471.195 ;
        RECT 0.000 1467.975 3165.000 1469.795 ;
        RECT 0.000 1466.575 3160.600 1467.975 ;
        RECT 0.000 1455.555 3165.000 1466.575 ;
        RECT 0.000 1454.155 3160.600 1455.555 ;
        RECT 0.000 1452.795 3165.000 1454.155 ;
        RECT 0.000 1451.395 3160.600 1452.795 ;
        RECT 0.000 1449.575 3165.000 1451.395 ;
        RECT 0.000 1448.175 3160.600 1449.575 ;
        RECT 0.000 1446.355 3165.000 1448.175 ;
        RECT 0.000 1444.955 3160.600 1446.355 ;
        RECT 0.000 1440.375 3165.000 1444.955 ;
        RECT 0.000 1438.975 3160.600 1440.375 ;
        RECT 0.000 1431.175 3165.000 1438.975 ;
        RECT 0.000 1429.775 3160.600 1431.175 ;
        RECT 0.000 1427.955 3165.000 1429.775 ;
        RECT 0.000 1426.555 3160.600 1427.955 ;
        RECT 0.000 1421.975 3165.000 1426.555 ;
        RECT 0.000 1421.425 3160.600 1421.975 ;
        RECT 4.400 1420.575 3160.600 1421.425 ;
        RECT 4.400 1420.025 3165.000 1420.575 ;
        RECT 0.000 1415.445 3165.000 1420.025 ;
        RECT 4.400 1414.045 3165.000 1415.445 ;
        RECT 0.000 1412.225 3165.000 1414.045 ;
        RECT 4.400 1410.825 3165.000 1412.225 ;
        RECT 0.000 1409.005 3165.000 1410.825 ;
        RECT 4.400 1407.605 3165.000 1409.005 ;
        RECT 0.000 1403.025 3165.000 1407.605 ;
        RECT 4.400 1401.625 3165.000 1403.025 ;
        RECT 0.000 1397.045 3165.000 1401.625 ;
        RECT 4.400 1395.645 3165.000 1397.045 ;
        RECT 0.000 1393.825 3165.000 1395.645 ;
        RECT 4.400 1392.425 3165.000 1393.825 ;
        RECT 0.000 1390.605 3165.000 1392.425 ;
        RECT 4.400 1389.205 3165.000 1390.605 ;
        RECT 0.000 1387.845 3165.000 1389.205 ;
        RECT 4.400 1386.445 3165.000 1387.845 ;
        RECT 0.000 1375.425 3165.000 1386.445 ;
        RECT 4.400 1374.025 3165.000 1375.425 ;
        RECT 0.000 1372.205 3165.000 1374.025 ;
        RECT 4.400 1370.805 3165.000 1372.205 ;
        RECT 0.000 1368.985 3165.000 1370.805 ;
        RECT 4.400 1367.585 3165.000 1368.985 ;
        RECT 0.000 1366.225 3165.000 1367.585 ;
        RECT 4.400 1364.825 3165.000 1366.225 ;
        RECT 0.000 1357.025 3165.000 1364.825 ;
        RECT 4.400 1355.625 3165.000 1357.025 ;
        RECT 0.000 1353.805 3165.000 1355.625 ;
        RECT 4.400 1352.405 3165.000 1353.805 ;
        RECT 0.000 1350.585 3165.000 1352.405 ;
        RECT 4.400 1349.185 3165.000 1350.585 ;
        RECT 0.000 1267.815 3165.000 1349.185 ;
        RECT 0.000 1266.415 3160.600 1267.815 ;
        RECT 0.000 1264.595 3165.000 1266.415 ;
        RECT 0.000 1263.195 3160.600 1264.595 ;
        RECT 0.000 1261.375 3165.000 1263.195 ;
        RECT 0.000 1259.975 3160.600 1261.375 ;
        RECT 0.000 1252.175 3165.000 1259.975 ;
        RECT 0.000 1250.775 3160.600 1252.175 ;
        RECT 0.000 1249.415 3165.000 1250.775 ;
        RECT 0.000 1248.015 3160.600 1249.415 ;
        RECT 0.000 1246.195 3165.000 1248.015 ;
        RECT 0.000 1244.795 3160.600 1246.195 ;
        RECT 0.000 1242.975 3165.000 1244.795 ;
        RECT 0.000 1241.575 3160.600 1242.975 ;
        RECT 0.000 1230.555 3165.000 1241.575 ;
        RECT 0.000 1229.155 3160.600 1230.555 ;
        RECT 0.000 1227.795 3165.000 1229.155 ;
        RECT 0.000 1226.395 3160.600 1227.795 ;
        RECT 0.000 1224.575 3165.000 1226.395 ;
        RECT 0.000 1223.175 3160.600 1224.575 ;
        RECT 0.000 1221.355 3165.000 1223.175 ;
        RECT 0.000 1219.955 3160.600 1221.355 ;
        RECT 0.000 1215.375 3165.000 1219.955 ;
        RECT 0.000 1213.975 3160.600 1215.375 ;
        RECT 0.000 1206.175 3165.000 1213.975 ;
        RECT 0.000 1205.425 3160.600 1206.175 ;
        RECT 4.400 1204.775 3160.600 1205.425 ;
        RECT 4.400 1204.025 3165.000 1204.775 ;
        RECT 0.000 1202.955 3165.000 1204.025 ;
        RECT 0.000 1201.555 3160.600 1202.955 ;
        RECT 0.000 1199.445 3165.000 1201.555 ;
        RECT 4.690 1198.045 3165.000 1199.445 ;
        RECT 0.000 1196.975 3165.000 1198.045 ;
        RECT 0.000 1196.225 3160.600 1196.975 ;
        RECT 4.400 1195.575 3160.600 1196.225 ;
        RECT 4.400 1194.825 3165.000 1195.575 ;
        RECT 0.000 1193.005 3165.000 1194.825 ;
        RECT 4.400 1191.605 3165.000 1193.005 ;
        RECT 0.000 1187.025 3165.000 1191.605 ;
        RECT 4.400 1185.625 3165.000 1187.025 ;
        RECT 0.000 1181.045 3165.000 1185.625 ;
        RECT 4.400 1179.645 3165.000 1181.045 ;
        RECT 0.000 1177.825 3165.000 1179.645 ;
        RECT 4.690 1176.425 3165.000 1177.825 ;
        RECT 0.000 1174.605 3165.000 1176.425 ;
        RECT 4.400 1173.205 3165.000 1174.605 ;
        RECT 0.000 1171.845 3165.000 1173.205 ;
        RECT 4.400 1170.445 3165.000 1171.845 ;
        RECT 0.000 1159.425 3165.000 1170.445 ;
        RECT 4.400 1158.025 3165.000 1159.425 ;
        RECT 0.000 1156.205 3165.000 1158.025 ;
        RECT 4.400 1154.805 3165.000 1156.205 ;
        RECT 0.000 1152.985 3165.000 1154.805 ;
        RECT 4.400 1151.585 3165.000 1152.985 ;
        RECT 0.000 1150.225 3165.000 1151.585 ;
        RECT 4.400 1148.825 3165.000 1150.225 ;
        RECT 0.000 1141.025 3165.000 1148.825 ;
        RECT 4.400 1139.625 3165.000 1141.025 ;
        RECT 0.000 1137.805 3165.000 1139.625 ;
        RECT 4.400 1136.405 3165.000 1137.805 ;
        RECT 0.000 1134.585 3165.000 1136.405 ;
        RECT 4.400 1133.185 3165.000 1134.585 ;
        RECT 0.000 1042.815 3165.000 1133.185 ;
        RECT 0.000 1041.415 3160.600 1042.815 ;
        RECT 0.000 1039.595 3165.000 1041.415 ;
        RECT 0.000 1038.195 3160.600 1039.595 ;
        RECT 0.000 1036.375 3165.000 1038.195 ;
        RECT 0.000 1034.975 3160.600 1036.375 ;
        RECT 0.000 1027.175 3165.000 1034.975 ;
        RECT 0.000 1025.775 3160.600 1027.175 ;
        RECT 0.000 1024.415 3165.000 1025.775 ;
        RECT 0.000 1023.015 3160.600 1024.415 ;
        RECT 0.000 1021.195 3165.000 1023.015 ;
        RECT 0.000 1019.795 3160.600 1021.195 ;
        RECT 0.000 1017.975 3165.000 1019.795 ;
        RECT 0.000 1016.575 3160.600 1017.975 ;
        RECT 0.000 1005.555 3165.000 1016.575 ;
        RECT 0.000 1004.155 3160.600 1005.555 ;
        RECT 0.000 1002.795 3165.000 1004.155 ;
        RECT 0.000 1001.395 3160.600 1002.795 ;
        RECT 0.000 999.575 3165.000 1001.395 ;
        RECT 0.000 998.175 3160.600 999.575 ;
        RECT 0.000 996.355 3165.000 998.175 ;
        RECT 0.000 994.955 3160.600 996.355 ;
        RECT 0.000 990.375 3165.000 994.955 ;
        RECT 0.000 989.425 3160.600 990.375 ;
        RECT 4.400 988.975 3160.600 989.425 ;
        RECT 4.400 988.025 3165.000 988.975 ;
        RECT 0.000 983.445 3165.000 988.025 ;
        RECT 4.400 982.045 3165.000 983.445 ;
        RECT 0.000 981.175 3165.000 982.045 ;
        RECT 0.000 980.225 3160.600 981.175 ;
        RECT 4.400 979.775 3160.600 980.225 ;
        RECT 4.400 978.825 3165.000 979.775 ;
        RECT 0.000 977.955 3165.000 978.825 ;
        RECT 0.000 976.555 3160.600 977.955 ;
        RECT 0.000 971.975 3165.000 976.555 ;
        RECT 0.000 971.025 3160.600 971.975 ;
        RECT 4.400 970.575 3160.600 971.025 ;
        RECT 4.400 969.625 3165.000 970.575 ;
        RECT 0.000 965.045 3165.000 969.625 ;
        RECT 4.400 963.645 3165.000 965.045 ;
        RECT 0.000 961.825 3165.000 963.645 ;
        RECT 4.400 960.425 3165.000 961.825 ;
        RECT 0.000 958.605 3165.000 960.425 ;
        RECT 4.400 957.205 3165.000 958.605 ;
        RECT 0.000 955.845 3165.000 957.205 ;
        RECT 4.400 954.445 3165.000 955.845 ;
        RECT 0.000 943.425 3165.000 954.445 ;
        RECT 4.400 942.025 3165.000 943.425 ;
        RECT 0.000 940.205 3165.000 942.025 ;
        RECT 4.400 938.805 3165.000 940.205 ;
        RECT 0.000 936.985 3165.000 938.805 ;
        RECT 4.400 935.585 3165.000 936.985 ;
        RECT 0.000 934.225 3165.000 935.585 ;
        RECT 4.400 932.825 3165.000 934.225 ;
        RECT 0.000 925.025 3165.000 932.825 ;
        RECT 4.400 923.625 3165.000 925.025 ;
        RECT 0.000 921.805 3165.000 923.625 ;
        RECT 4.400 920.405 3165.000 921.805 ;
        RECT 0.000 918.585 3165.000 920.405 ;
        RECT 4.400 917.185 3165.000 918.585 ;
        RECT 0.000 816.815 3165.000 917.185 ;
        RECT 0.000 815.415 3160.600 816.815 ;
        RECT 0.000 813.595 3165.000 815.415 ;
        RECT 0.000 812.195 3160.600 813.595 ;
        RECT 0.000 810.375 3165.000 812.195 ;
        RECT 0.000 808.975 3160.600 810.375 ;
        RECT 0.000 801.175 3165.000 808.975 ;
        RECT 0.000 799.775 3160.600 801.175 ;
        RECT 0.000 798.415 3165.000 799.775 ;
        RECT 0.000 797.015 3160.600 798.415 ;
        RECT 0.000 795.195 3165.000 797.015 ;
        RECT 0.000 793.795 3160.600 795.195 ;
        RECT 0.000 791.975 3165.000 793.795 ;
        RECT 0.000 790.575 3160.600 791.975 ;
        RECT 0.000 779.555 3165.000 790.575 ;
        RECT 0.000 778.155 3160.600 779.555 ;
        RECT 0.000 776.795 3165.000 778.155 ;
        RECT 0.000 775.395 3160.600 776.795 ;
        RECT 0.000 773.575 3165.000 775.395 ;
        RECT 0.000 773.425 3160.600 773.575 ;
        RECT 4.400 772.175 3160.600 773.425 ;
        RECT 4.400 772.025 3165.000 772.175 ;
        RECT 0.000 770.355 3165.000 772.025 ;
        RECT 0.000 768.955 3160.600 770.355 ;
        RECT 0.000 767.445 3165.000 768.955 ;
        RECT 4.400 766.045 3165.000 767.445 ;
        RECT 0.000 764.375 3165.000 766.045 ;
        RECT 0.000 764.225 3160.600 764.375 ;
        RECT 4.400 762.975 3160.600 764.225 ;
        RECT 4.400 762.825 3165.000 762.975 ;
        RECT 0.000 755.175 3165.000 762.825 ;
        RECT 0.000 755.025 3160.600 755.175 ;
        RECT 4.400 753.775 3160.600 755.025 ;
        RECT 4.400 753.625 3165.000 753.775 ;
        RECT 0.000 751.955 3165.000 753.625 ;
        RECT 0.000 750.555 3160.600 751.955 ;
        RECT 0.000 749.045 3165.000 750.555 ;
        RECT 4.400 747.645 3165.000 749.045 ;
        RECT 0.000 745.975 3165.000 747.645 ;
        RECT 0.000 745.825 3160.600 745.975 ;
        RECT 4.400 744.575 3160.600 745.825 ;
        RECT 4.400 744.425 3165.000 744.575 ;
        RECT 0.000 742.605 3165.000 744.425 ;
        RECT 4.400 741.205 3165.000 742.605 ;
        RECT 0.000 739.845 3165.000 741.205 ;
        RECT 4.400 738.445 3165.000 739.845 ;
        RECT 0.000 727.425 3165.000 738.445 ;
        RECT 4.400 726.025 3165.000 727.425 ;
        RECT 0.000 724.205 3165.000 726.025 ;
        RECT 4.400 722.805 3165.000 724.205 ;
        RECT 0.000 720.985 3165.000 722.805 ;
        RECT 4.400 719.585 3165.000 720.985 ;
        RECT 0.000 718.225 3165.000 719.585 ;
        RECT 4.400 716.825 3165.000 718.225 ;
        RECT 0.000 709.025 3165.000 716.825 ;
        RECT 4.400 707.625 3165.000 709.025 ;
        RECT 0.000 705.805 3165.000 707.625 ;
        RECT 4.400 704.405 3165.000 705.805 ;
        RECT 0.000 702.585 3165.000 704.405 ;
        RECT 4.400 701.185 3165.000 702.585 ;
        RECT 0.000 591.815 3165.000 701.185 ;
        RECT 0.000 590.415 3160.600 591.815 ;
        RECT 0.000 588.595 3165.000 590.415 ;
        RECT 0.000 587.195 3160.600 588.595 ;
        RECT 0.000 585.375 3165.000 587.195 ;
        RECT 0.000 583.975 3160.600 585.375 ;
        RECT 0.000 576.175 3165.000 583.975 ;
        RECT 0.000 574.775 3160.600 576.175 ;
        RECT 0.000 573.415 3165.000 574.775 ;
        RECT 0.000 572.015 3160.600 573.415 ;
        RECT 0.000 570.195 3165.000 572.015 ;
        RECT 0.000 568.795 3160.600 570.195 ;
        RECT 0.000 566.975 3165.000 568.795 ;
        RECT 0.000 565.575 3160.600 566.975 ;
        RECT 0.000 554.555 3165.000 565.575 ;
        RECT 0.000 553.155 3160.600 554.555 ;
        RECT 0.000 551.795 3165.000 553.155 ;
        RECT 0.000 550.395 3160.600 551.795 ;
        RECT 0.000 548.575 3165.000 550.395 ;
        RECT 0.000 547.175 3160.600 548.575 ;
        RECT 0.000 545.355 3165.000 547.175 ;
        RECT 0.000 543.955 3160.600 545.355 ;
        RECT 0.000 539.375 3165.000 543.955 ;
        RECT 0.000 537.975 3160.600 539.375 ;
        RECT 0.000 530.175 3165.000 537.975 ;
        RECT 0.000 528.775 3160.600 530.175 ;
        RECT 0.000 526.955 3165.000 528.775 ;
        RECT 0.000 525.555 3160.600 526.955 ;
        RECT 0.000 520.975 3165.000 525.555 ;
        RECT 0.000 519.575 3160.600 520.975 ;
        RECT 0.000 365.815 3165.000 519.575 ;
        RECT 0.000 364.415 3160.600 365.815 ;
        RECT 0.000 362.595 3165.000 364.415 ;
        RECT 0.000 361.195 3160.600 362.595 ;
        RECT 0.000 359.375 3165.000 361.195 ;
        RECT 0.000 357.975 3160.600 359.375 ;
        RECT 0.000 350.175 3165.000 357.975 ;
        RECT 0.000 348.775 3160.600 350.175 ;
        RECT 0.000 347.415 3165.000 348.775 ;
        RECT 0.000 346.015 3160.600 347.415 ;
        RECT 0.000 344.195 3165.000 346.015 ;
        RECT 0.000 342.795 3160.600 344.195 ;
        RECT 0.000 340.975 3165.000 342.795 ;
        RECT 0.000 339.575 3160.600 340.975 ;
        RECT 0.000 328.555 3165.000 339.575 ;
        RECT 0.000 327.155 3160.600 328.555 ;
        RECT 0.000 325.795 3165.000 327.155 ;
        RECT 0.000 324.395 3160.600 325.795 ;
        RECT 0.000 322.575 3165.000 324.395 ;
        RECT 0.000 321.175 3160.600 322.575 ;
        RECT 0.000 319.355 3165.000 321.175 ;
        RECT 0.000 317.955 3160.600 319.355 ;
        RECT 0.000 313.375 3165.000 317.955 ;
        RECT 0.000 311.975 3160.600 313.375 ;
        RECT 0.000 304.175 3165.000 311.975 ;
        RECT 0.000 302.775 3160.600 304.175 ;
        RECT 0.000 300.955 3165.000 302.775 ;
        RECT 0.000 299.555 3160.600 300.955 ;
        RECT 0.000 294.975 3165.000 299.555 ;
        RECT 0.000 293.575 3160.600 294.975 ;
        RECT 0.000 204.200 3165.000 293.575 ;
      LAYER met3 ;
        RECT -16.080 180.255 5.910 204.200 ;
      LAYER met3 ;
        RECT 5.910 180.255 3165.000 204.200 ;
        RECT 0.000 154.000 3165.000 180.255 ;
      LAYER met3 ;
        RECT -16.080 130.055 5.910 154.000 ;
      LAYER met3 ;
        RECT 5.910 130.055 3165.000 154.000 ;
        RECT 0.000 0.000 3165.000 130.055 ;
      LAYER met3 ;
        RECT 858.500 -31.255 876.510 -0.675 ;
        RECT 966.025 -40.985 979.745 -0.675 ;
        RECT 994.715 -14.690 1018.745 -0.110 ;
        RECT 1044.970 -14.690 1069.000 -0.110 ;
      LAYER met4 ;
        RECT 2666.935 4767.000 2690.965 4772.410 ;
        RECT 2716.840 4767.000 2740.870 4772.410 ;
      LAYER met4 ;
        RECT 0.000 4755.200 3165.000 4767.000 ;
      LAYER met4 ;
        RECT -9.290 4400.255 0.000 4424.200 ;
        RECT -9.290 4375.600 0.000 4398.650 ;
        RECT -9.290 4350.055 0.000 4374.000 ;
        RECT -9.290 3977.845 0.000 4001.790 ;
        RECT -9.290 3927.945 0.000 3951.590 ;
        RECT -9.290 2254.845 0.000 2278.790 ;
        RECT -9.290 2204.945 0.000 2228.590 ;
        RECT -9.290 2044.255 0.000 2068.200 ;
        RECT -9.290 2019.600 0.000 2042.650 ;
        RECT -9.290 1994.055 0.000 2018.000 ;
        RECT -9.290 180.255 0.000 204.200 ;
        RECT -9.290 130.055 0.000 154.000 ;
      LAYER met4 ;
        RECT 0.000 10.240 10.520 4755.200 ;
        RECT 16.320 10.240 16.520 4755.200 ;
        RECT 22.320 10.240 22.520 4755.200 ;
        RECT 28.320 10.240 28.520 4755.200 ;
        RECT 34.320 10.240 34.520 4755.200 ;
        RECT 40.320 10.240 40.520 4755.200 ;
        RECT 46.320 10.240 46.520 4755.200 ;
        RECT 52.320 10.240 52.520 4755.200 ;
        RECT 58.320 10.240 58.520 4755.200 ;
        RECT 64.320 10.240 64.520 4755.200 ;
        RECT 70.320 10.240 70.520 4755.200 ;
        RECT 73.320 10.240 73.520 4755.200 ;
        RECT 76.320 4595.900 123.520 4755.200 ;
        RECT 130.720 4595.900 131.120 4755.200 ;
        RECT 138.320 4595.900 223.520 4755.200 ;
        RECT 230.720 4595.900 231.120 4755.200 ;
        RECT 238.320 4595.900 255.640 4755.200 ;
        RECT 262.840 4595.900 263.240 4755.200 ;
        RECT 270.440 4595.900 323.520 4755.200 ;
        RECT 330.720 4595.900 331.120 4755.200 ;
        RECT 338.320 4595.900 423.520 4755.200 ;
        RECT 430.720 4595.900 431.120 4755.200 ;
        RECT 438.320 4595.900 523.520 4755.200 ;
        RECT 530.720 4595.900 531.120 4755.200 ;
        RECT 538.320 4595.900 555.640 4755.200 ;
        RECT 562.840 4595.900 563.240 4755.200 ;
        RECT 570.440 4595.900 623.520 4755.200 ;
        RECT 630.720 4595.900 631.120 4755.200 ;
        RECT 638.320 4595.900 723.520 4755.200 ;
        RECT 730.720 4595.900 731.120 4755.200 ;
        RECT 738.320 4595.900 823.520 4755.200 ;
        RECT 830.720 4595.900 831.120 4755.200 ;
        RECT 838.320 4595.900 923.520 4755.200 ;
        RECT 930.720 4595.900 931.120 4755.200 ;
        RECT 938.320 4595.900 955.640 4755.200 ;
        RECT 962.840 4595.900 963.240 4755.200 ;
        RECT 970.440 4595.900 1023.520 4755.200 ;
        RECT 1030.720 4595.900 1031.120 4755.200 ;
        RECT 1038.320 4595.900 1123.520 4755.200 ;
        RECT 1130.720 4595.900 1131.120 4755.200 ;
        RECT 1138.320 4595.900 1155.640 4755.200 ;
        RECT 1162.840 4595.900 1163.240 4755.200 ;
        RECT 1170.440 4595.900 1223.520 4755.200 ;
        RECT 1230.720 4595.900 1231.120 4755.200 ;
        RECT 1238.320 4595.900 1323.520 4755.200 ;
        RECT 1330.720 4595.900 1331.120 4755.200 ;
        RECT 1338.320 4595.900 1423.520 4755.200 ;
        RECT 1430.720 4595.900 1431.120 4755.200 ;
        RECT 1438.320 4595.900 1455.640 4755.200 ;
        RECT 1462.840 4595.900 1463.240 4755.200 ;
        RECT 1470.440 4595.900 1475.320 4755.200 ;
        RECT 1480.920 4595.900 1523.520 4755.200 ;
        RECT 1530.720 4595.900 1531.120 4755.200 ;
        RECT 1538.320 4595.900 1623.520 4755.200 ;
        RECT 1630.720 4595.900 1631.120 4755.200 ;
        RECT 1638.320 4595.900 1723.520 4755.200 ;
        RECT 1730.720 4595.900 1731.120 4755.200 ;
        RECT 1738.320 4595.900 1755.640 4755.200 ;
        RECT 1762.840 4595.900 1763.240 4755.200 ;
        RECT 1770.440 4595.900 1823.520 4755.200 ;
        RECT 1830.720 4595.900 1831.120 4755.200 ;
        RECT 1838.320 4595.900 1923.520 4755.200 ;
        RECT 1930.720 4595.900 1931.120 4755.200 ;
        RECT 1938.320 4595.900 2023.520 4755.200 ;
        RECT 2030.720 4595.900 2031.120 4755.200 ;
        RECT 2038.320 4595.900 2055.640 4755.200 ;
        RECT 2062.840 4595.900 2063.240 4755.200 ;
        RECT 2070.440 4595.900 2123.520 4755.200 ;
        RECT 2130.720 4595.900 2131.120 4755.200 ;
        RECT 2138.320 4595.900 2223.520 4755.200 ;
        RECT 2230.720 4595.900 2231.120 4755.200 ;
        RECT 2238.320 4595.900 2323.520 4755.200 ;
        RECT 2330.720 4595.900 2331.120 4755.200 ;
        RECT 2338.320 4595.900 2355.640 4755.200 ;
        RECT 2362.840 4595.900 2363.240 4755.200 ;
        RECT 2370.440 4595.900 2423.520 4755.200 ;
        RECT 2430.720 4595.900 2431.120 4755.200 ;
        RECT 2438.320 4595.900 2523.520 4755.200 ;
        RECT 2530.720 4595.900 2531.120 4755.200 ;
        RECT 2538.320 4595.900 2623.520 4755.200 ;
        RECT 2630.720 4595.900 2631.120 4755.200 ;
        RECT 2638.320 4692.640 2755.640 4755.200 ;
        RECT 2638.320 4639.680 2649.920 4692.640 ;
        RECT 2655.720 4639.680 2656.360 4692.640 ;
        RECT 2662.160 4639.680 2755.640 4692.640 ;
        RECT 2638.320 4603.400 2755.640 4639.680 ;
        RECT 2638.320 4595.900 2723.520 4603.400 ;
        RECT 2730.720 4595.900 2731.120 4603.400 ;
        RECT 2738.320 4595.900 2755.640 4603.400 ;
        RECT 2762.840 4595.900 2763.240 4755.200 ;
        RECT 2770.440 4595.900 2823.520 4755.200 ;
        RECT 2830.720 4595.900 2831.120 4755.200 ;
        RECT 2838.320 4595.900 2923.520 4755.200 ;
        RECT 2930.720 4595.900 2931.120 4755.200 ;
        RECT 2938.320 4595.900 3023.520 4755.200 ;
        RECT 3030.720 4595.900 3031.120 4755.200 ;
        RECT 3038.320 4595.900 3086.780 4755.200 ;
        RECT 76.320 989.400 3086.780 4595.900 ;
        RECT 76.320 10.240 123.520 989.400 ;
        RECT 130.720 10.240 131.120 989.400 ;
        RECT 138.320 619.965 223.520 989.400 ;
        RECT 230.720 619.965 231.120 989.400 ;
        RECT 238.320 619.965 323.520 989.400 ;
        RECT 330.720 619.965 331.120 989.400 ;
        RECT 338.320 619.965 423.520 989.400 ;
        RECT 430.720 619.965 431.120 989.400 ;
        RECT 438.320 619.965 523.520 989.400 ;
        RECT 138.320 174.075 523.520 619.965 ;
        RECT 138.320 10.240 223.520 174.075 ;
        RECT 230.720 10.240 231.120 174.075 ;
        RECT 238.320 10.240 323.520 174.075 ;
        RECT 330.720 10.240 331.120 174.075 ;
        RECT 338.320 10.240 423.520 174.075 ;
        RECT 430.720 10.240 431.120 174.075 ;
        RECT 438.320 10.240 523.520 174.075 ;
        RECT 530.720 10.240 531.120 989.400 ;
        RECT 538.320 10.240 555.640 989.400 ;
        RECT 562.840 10.240 563.240 989.400 ;
        RECT 570.440 619.965 623.520 989.400 ;
        RECT 630.720 619.965 631.120 989.400 ;
        RECT 638.320 619.965 723.520 989.400 ;
        RECT 730.720 619.965 731.120 989.400 ;
        RECT 738.320 619.965 823.520 989.400 ;
        RECT 830.720 619.965 831.120 989.400 ;
        RECT 838.320 619.965 850.320 989.400 ;
        RECT 855.920 619.965 858.320 989.400 ;
        RECT 863.920 619.965 900.320 989.400 ;
        RECT 570.440 174.075 900.320 619.965 ;
        RECT 570.440 10.240 623.520 174.075 ;
        RECT 630.720 10.240 631.120 174.075 ;
        RECT 638.320 10.240 654.320 174.075 ;
        RECT 659.920 169.580 723.520 174.075 ;
        RECT 659.920 10.240 661.120 169.580 ;
        RECT 666.720 10.240 723.520 169.580 ;
        RECT 730.720 169.580 823.520 174.075 ;
        RECT 730.720 10.240 731.120 169.580 ;
        RECT 738.320 10.240 823.520 169.580 ;
        RECT 830.720 10.240 831.120 174.075 ;
        RECT 838.320 10.240 900.320 174.075 ;
        RECT 905.920 10.240 908.320 989.400 ;
        RECT 913.920 10.240 923.520 989.400 ;
        RECT 930.720 10.240 931.120 989.400 ;
        RECT 938.320 10.240 955.640 989.400 ;
        RECT 962.840 33.680 1023.520 989.400 ;
        RECT 1030.720 33.680 1031.120 989.400 ;
        RECT 1038.320 189.400 1123.520 989.400 ;
        RECT 1038.320 33.680 1040.320 189.400 ;
        RECT 1045.920 33.680 1047.120 189.400 ;
        RECT 1052.720 33.680 1123.520 189.400 ;
        RECT 962.840 10.240 1123.520 33.680 ;
        RECT 1130.720 10.240 1131.120 989.400 ;
        RECT 1138.320 10.240 1155.640 989.400 ;
        RECT 1162.840 10.240 1163.240 989.400 ;
        RECT 1170.440 10.240 1223.520 989.400 ;
        RECT 1230.720 10.240 1231.120 989.400 ;
        RECT 1238.320 10.240 1275.320 989.400 ;
        RECT 1280.920 10.240 1283.320 989.400 ;
        RECT 1288.920 10.240 1323.520 989.400 ;
        RECT 1330.720 10.240 1331.120 989.400 ;
        RECT 1338.320 10.240 1375.320 989.400 ;
        RECT 1380.920 10.240 1383.320 989.400 ;
        RECT 1388.920 10.240 1423.520 989.400 ;
        RECT 1430.720 10.240 1431.120 989.400 ;
        RECT 1438.320 10.240 1455.640 989.400 ;
        RECT 1462.840 10.240 1463.240 989.400 ;
        RECT 1470.440 10.240 1475.320 989.400 ;
        RECT 1480.920 10.240 1483.320 989.400 ;
        RECT 1488.920 10.240 1523.520 989.400 ;
        RECT 1530.720 10.240 1531.120 989.400 ;
        RECT 1538.320 283.620 1623.520 989.400 ;
        RECT 1630.720 283.620 1631.120 989.400 ;
        RECT 1638.320 283.620 1723.520 989.400 ;
        RECT 1538.320 177.580 1723.520 283.620 ;
        RECT 1538.320 10.240 1623.520 177.580 ;
        RECT 1630.720 10.240 1631.120 177.580 ;
        RECT 1638.320 10.240 1723.520 177.580 ;
        RECT 1730.720 10.240 1731.120 989.400 ;
        RECT 1738.320 10.240 1755.640 989.400 ;
        RECT 1762.840 10.240 1763.240 989.400 ;
        RECT 1770.440 569.965 1823.520 989.400 ;
        RECT 1830.720 569.965 1831.120 989.400 ;
        RECT 1838.320 569.965 1843.320 989.400 ;
        RECT 1848.920 569.965 1851.320 989.400 ;
        RECT 1856.920 569.965 1859.320 989.400 ;
        RECT 1864.920 569.965 1867.320 989.400 ;
        RECT 1872.920 569.965 1883.320 989.400 ;
        RECT 1888.920 569.965 1891.320 989.400 ;
        RECT 1896.920 569.965 1899.320 989.400 ;
        RECT 1904.920 569.965 1907.320 989.400 ;
        RECT 1912.920 569.965 1923.520 989.400 ;
        RECT 1930.720 569.965 1931.120 989.400 ;
        RECT 1938.320 569.965 2023.520 989.400 ;
        RECT 2030.720 569.965 2031.120 989.400 ;
        RECT 2038.320 569.965 2123.520 989.400 ;
        RECT 1770.440 124.075 2123.520 569.965 ;
        RECT 1770.440 10.240 1823.520 124.075 ;
        RECT 1830.720 10.240 1831.120 124.075 ;
        RECT 1838.320 10.240 1923.520 124.075 ;
        RECT 1930.720 10.240 1931.120 124.075 ;
        RECT 1938.320 10.240 2023.520 124.075 ;
        RECT 2030.720 119.580 2123.520 124.075 ;
        RECT 2030.720 10.240 2031.120 119.580 ;
        RECT 2038.320 10.240 2123.520 119.580 ;
        RECT 2130.720 10.240 2131.120 989.400 ;
        RECT 2138.320 10.240 2223.520 989.400 ;
        RECT 2230.720 10.240 2231.120 989.400 ;
        RECT 2238.320 10.240 2323.520 989.400 ;
        RECT 2330.720 10.240 2331.120 989.400 ;
        RECT 2338.320 10.240 2355.640 989.400 ;
        RECT 2362.840 10.240 2363.240 989.400 ;
        RECT 2370.440 10.240 2423.520 989.400 ;
        RECT 2430.720 10.240 2431.120 989.400 ;
        RECT 2438.320 10.240 2523.520 989.400 ;
        RECT 2530.720 10.240 2531.120 989.400 ;
        RECT 2538.320 10.240 2623.520 989.400 ;
        RECT 2630.720 10.240 2631.120 989.400 ;
        RECT 2638.320 732.885 2723.520 989.400 ;
        RECT 2730.720 732.885 2731.120 989.400 ;
        RECT 2738.320 736.700 2823.520 989.400 ;
        RECT 2830.720 736.700 2831.120 989.400 ;
        RECT 2738.320 732.885 2831.120 736.700 ;
        RECT 2838.320 732.885 2923.520 989.400 ;
        RECT 2930.720 732.885 2931.120 989.400 ;
        RECT 2938.320 732.885 3023.520 989.400 ;
        RECT 3030.720 732.885 3031.120 989.400 ;
        RECT 3038.320 732.885 3086.780 989.400 ;
        RECT 2638.320 193.835 3086.780 732.885 ;
        RECT 2638.320 10.240 2723.520 193.835 ;
        RECT 2730.720 10.240 2731.120 193.835 ;
        RECT 2738.320 192.740 2831.120 193.835 ;
        RECT 2738.320 10.240 2823.520 192.740 ;
        RECT 2830.720 10.240 2831.120 192.740 ;
        RECT 2838.320 10.240 2923.520 193.835 ;
        RECT 2930.720 10.240 2931.120 193.835 ;
        RECT 2938.320 10.240 3023.520 193.835 ;
        RECT 3030.720 10.240 3031.120 193.835 ;
        RECT 3038.320 10.240 3086.780 193.835 ;
        RECT 3089.580 10.240 3089.780 4755.200 ;
        RECT 3092.580 10.240 3092.780 4755.200 ;
        RECT 3098.580 10.240 3098.780 4755.200 ;
        RECT 3104.580 10.240 3104.780 4755.200 ;
        RECT 3110.580 10.240 3110.780 4755.200 ;
        RECT 3116.580 10.240 3116.780 4755.200 ;
        RECT 3122.580 10.240 3122.780 4755.200 ;
        RECT 3128.580 10.240 3128.780 4755.200 ;
        RECT 3134.580 10.240 3134.780 4755.200 ;
        RECT 3140.580 10.240 3140.780 4755.200 ;
        RECT 3146.580 10.240 3146.780 4755.200 ;
        RECT 3152.580 10.240 3165.000 4755.200 ;
      LAYER met4 ;
        RECT 3165.000 4378.055 3171.230 4402.000 ;
        RECT 3165.000 4353.345 3171.230 4376.450 ;
        RECT 3165.000 4327.800 3171.230 4351.745 ;
        RECT 3165.000 3932.060 3171.230 3956.005 ;
        RECT 3165.000 3882.145 3171.230 3906.090 ;
        RECT 3165.000 2359.060 3171.230 2383.005 ;
        RECT 3165.000 2309.145 3171.230 2333.090 ;
        RECT 3165.000 2139.055 3171.230 2163.000 ;
        RECT 3165.000 2114.345 3171.230 2137.450 ;
        RECT 3165.000 2088.800 3171.230 2112.745 ;
        RECT 3165.000 1918.100 3171.230 1942.045 ;
        RECT 3165.000 1868.185 3171.230 1892.130 ;
      LAYER met4 ;
        RECT 0.000 0.000 3165.000 10.240 ;
      LAYER met4 ;
        RECT 858.500 -9.685 876.510 0.000 ;
        RECT 966.025 -9.685 979.745 0.000 ;
        RECT 994.715 -9.120 1018.745 0.000 ;
        RECT 1044.970 -9.120 1069.000 0.000 ;
        RECT 966.540 -40.630 978.860 -36.710 ;
      LAYER met5 ;
        RECT 0.000 4525.480 3165.000 4594.950 ;
        RECT 0.000 4507.080 8.280 4525.480 ;
        RECT 77.520 4507.080 3085.580 4525.480 ;
        RECT 3156.520 4507.080 3165.000 4525.480 ;
      LAYER met5 ;
        RECT -9.290 4400.250 0.000 4424.200 ;
        RECT -9.290 4375.600 0.000 4398.650 ;
        RECT -9.290 4350.050 0.000 4374.000 ;
      LAYER met5 ;
        RECT 0.000 4285.480 3165.000 4507.080 ;
      LAYER met5 ;
        RECT 3165.000 4378.050 3171.230 4402.000 ;
        RECT 3165.000 4353.345 3171.230 4376.450 ;
        RECT 3165.000 4327.795 3171.230 4351.745 ;
      LAYER met5 ;
        RECT 0.000 4267.080 8.280 4285.480 ;
        RECT 77.520 4267.080 3085.580 4285.480 ;
        RECT 3156.520 4267.080 3165.000 4285.480 ;
        RECT 0.000 4165.480 3165.000 4267.080 ;
        RECT 0.000 4147.080 8.280 4165.480 ;
        RECT 77.520 4147.080 3085.580 4165.480 ;
        RECT 3156.520 4147.080 3165.000 4165.480 ;
        RECT 0.000 4045.480 3165.000 4147.080 ;
        RECT 0.000 4027.080 8.280 4045.480 ;
        RECT 77.520 4027.080 3085.580 4045.480 ;
        RECT 3156.520 4027.080 3165.000 4045.480 ;
      LAYER met5 ;
        RECT -9.290 3977.840 0.000 4001.790 ;
        RECT -9.290 3927.945 0.000 3951.895 ;
      LAYER met5 ;
        RECT 0.000 3925.480 3165.000 4027.080 ;
      LAYER met5 ;
        RECT 3165.000 3932.055 3171.230 3956.005 ;
      LAYER met5 ;
        RECT 0.000 3907.080 8.280 3925.480 ;
        RECT 77.520 3907.080 3165.000 3925.480 ;
        RECT 0.000 3805.480 3165.000 3907.080 ;
      LAYER met5 ;
        RECT 3165.000 3882.140 3171.230 3906.090 ;
      LAYER met5 ;
        RECT 0.000 3787.080 8.280 3805.480 ;
        RECT 77.520 3787.080 3085.580 3805.480 ;
        RECT 3156.520 3787.080 3165.000 3805.480 ;
        RECT 0.000 3685.480 3165.000 3787.080 ;
        RECT 0.000 3667.080 8.280 3685.480 ;
        RECT 77.520 3667.080 3085.580 3685.480 ;
        RECT 3156.520 3667.080 3165.000 3685.480 ;
        RECT 0.000 3565.480 3165.000 3667.080 ;
        RECT 0.000 3547.080 8.280 3565.480 ;
        RECT 77.520 3547.080 3085.580 3565.480 ;
        RECT 3156.520 3547.080 3165.000 3565.480 ;
        RECT 0.000 3445.480 3165.000 3547.080 ;
        RECT 0.000 3427.080 8.280 3445.480 ;
        RECT 77.520 3427.080 3085.580 3445.480 ;
        RECT 3156.520 3427.080 3165.000 3445.480 ;
        RECT 0.000 3325.480 3165.000 3427.080 ;
        RECT 0.000 3307.080 8.280 3325.480 ;
        RECT 77.520 3307.080 3085.580 3325.480 ;
        RECT 3156.520 3307.080 3165.000 3325.480 ;
        RECT 0.000 3205.480 3165.000 3307.080 ;
        RECT 0.000 3187.080 8.280 3205.480 ;
        RECT 77.520 3187.080 3085.580 3205.480 ;
        RECT 3156.520 3187.080 3165.000 3205.480 ;
        RECT 0.000 3085.480 3165.000 3187.080 ;
        RECT 0.000 3067.080 8.280 3085.480 ;
        RECT 77.520 3067.080 3085.580 3085.480 ;
        RECT 3156.520 3067.080 3165.000 3085.480 ;
        RECT 0.000 2965.480 3165.000 3067.080 ;
        RECT 0.000 2947.080 8.280 2965.480 ;
        RECT 77.520 2947.080 3085.580 2965.480 ;
        RECT 3156.520 2947.080 3165.000 2965.480 ;
        RECT 0.000 2845.480 3165.000 2947.080 ;
        RECT 0.000 2827.080 8.280 2845.480 ;
        RECT 77.520 2827.080 3085.580 2845.480 ;
        RECT 3156.520 2827.080 3165.000 2845.480 ;
        RECT 0.000 2725.480 3165.000 2827.080 ;
        RECT 0.000 2707.080 8.280 2725.480 ;
        RECT 77.520 2707.080 3085.580 2725.480 ;
        RECT 3156.520 2707.080 3165.000 2725.480 ;
        RECT 0.000 2605.480 3165.000 2707.080 ;
        RECT 0.000 2587.080 8.280 2605.480 ;
        RECT 77.520 2587.080 3085.580 2605.480 ;
        RECT 3156.520 2587.080 3165.000 2605.480 ;
        RECT 0.000 2485.480 3165.000 2587.080 ;
        RECT 0.000 2467.080 8.280 2485.480 ;
        RECT 77.520 2467.080 3085.580 2485.480 ;
        RECT 3156.520 2467.080 3165.000 2485.480 ;
        RECT 0.000 2365.480 3165.000 2467.080 ;
        RECT 0.000 2347.080 8.280 2365.480 ;
        RECT 77.520 2347.080 3165.000 2365.480 ;
      LAYER met5 ;
        RECT 3165.000 2359.055 3171.230 2383.005 ;
        RECT -9.290 2254.840 0.000 2278.790 ;
      LAYER met5 ;
        RECT 0.000 2245.480 3165.000 2347.080 ;
      LAYER met5 ;
        RECT 3165.000 2309.140 3171.230 2333.090 ;
        RECT -9.290 2204.945 0.000 2228.895 ;
      LAYER met5 ;
        RECT 0.000 2227.080 3085.580 2245.480 ;
        RECT 3156.520 2227.080 3165.000 2245.480 ;
        RECT 0.000 2125.480 3165.000 2227.080 ;
      LAYER met5 ;
        RECT 3165.000 2139.050 3171.230 2163.000 ;
      LAYER met5 ;
        RECT 0.000 2107.080 8.280 2125.480 ;
        RECT 77.520 2107.080 3165.000 2125.480 ;
      LAYER met5 ;
        RECT 3165.000 2114.345 3171.230 2137.450 ;
        RECT -9.290 2044.250 0.000 2068.200 ;
        RECT -9.290 2019.600 0.000 2042.650 ;
        RECT -9.290 1994.050 0.000 2018.000 ;
      LAYER met5 ;
        RECT 0.000 2005.480 3165.000 2107.080 ;
      LAYER met5 ;
        RECT 3165.000 2088.795 3171.230 2112.745 ;
      LAYER met5 ;
        RECT 0.000 1987.080 3085.580 2005.480 ;
        RECT 3156.520 1987.080 3165.000 2005.480 ;
        RECT 0.000 1885.480 3165.000 1987.080 ;
      LAYER met5 ;
        RECT 3165.000 1918.095 3171.230 1942.045 ;
      LAYER met5 ;
        RECT 0.000 1867.080 8.280 1885.480 ;
        RECT 77.520 1867.080 3165.000 1885.480 ;
      LAYER met5 ;
        RECT 3165.000 1868.180 3171.230 1892.130 ;
      LAYER met5 ;
        RECT 0.000 1765.480 3165.000 1867.080 ;
        RECT 0.000 1747.080 8.280 1765.480 ;
        RECT 77.520 1747.080 3085.580 1765.480 ;
        RECT 3156.520 1747.080 3165.000 1765.480 ;
        RECT 0.000 1645.480 3165.000 1747.080 ;
        RECT 0.000 1627.080 8.280 1645.480 ;
        RECT 77.520 1627.080 3085.580 1645.480 ;
        RECT 3156.520 1627.080 3165.000 1645.480 ;
        RECT 0.000 1525.480 3165.000 1627.080 ;
        RECT 0.000 1507.080 8.280 1525.480 ;
        RECT 77.520 1507.080 3085.580 1525.480 ;
        RECT 3156.520 1507.080 3165.000 1525.480 ;
        RECT 0.000 1405.480 3165.000 1507.080 ;
        RECT 0.000 1387.080 8.280 1405.480 ;
        RECT 77.520 1387.080 3085.580 1405.480 ;
        RECT 3156.520 1387.080 3165.000 1405.480 ;
        RECT 0.000 1285.480 3165.000 1387.080 ;
        RECT 0.000 1267.080 8.280 1285.480 ;
        RECT 77.520 1267.080 3085.580 1285.480 ;
        RECT 3156.520 1267.080 3165.000 1285.480 ;
        RECT 0.000 1165.480 3165.000 1267.080 ;
        RECT 0.000 1147.080 8.280 1165.480 ;
        RECT 77.520 1147.080 3085.580 1165.480 ;
        RECT 3156.520 1147.080 3165.000 1165.480 ;
        RECT 0.000 1045.480 3165.000 1147.080 ;
        RECT 0.000 1027.080 8.280 1045.480 ;
        RECT 77.520 1027.080 3085.580 1045.480 ;
        RECT 3156.520 1027.080 3165.000 1045.480 ;
        RECT 0.000 985.800 3165.000 1027.080 ;
        RECT 0.000 951.400 8.280 985.800 ;
        RECT 3156.520 951.400 3165.000 985.800 ;
        RECT 0.000 925.480 3165.000 951.400 ;
        RECT 0.000 907.080 8.280 925.480 ;
        RECT 3156.520 907.080 3165.000 925.480 ;
        RECT 0.000 877.880 3165.000 907.080 ;
        RECT 0.000 813.880 8.280 877.880 ;
        RECT 3156.520 813.880 3165.000 877.880 ;
        RECT 0.000 805.480 3165.000 813.880 ;
        RECT 0.000 787.080 8.280 805.480 ;
        RECT 3156.520 787.080 3165.000 805.480 ;
        RECT 0.000 755.480 3165.000 787.080 ;
        RECT 0.000 721.080 8.280 755.480 ;
        RECT 3156.520 721.080 3165.000 755.480 ;
        RECT 0.000 685.480 3165.000 721.080 ;
        RECT 0.000 667.080 8.280 685.480 ;
        RECT 3156.520 667.080 3165.000 685.480 ;
        RECT 0.000 635.480 3165.000 667.080 ;
        RECT 0.000 601.080 8.280 635.480 ;
        RECT 3156.520 601.080 3165.000 635.480 ;
        RECT 0.000 565.480 3165.000 601.080 ;
        RECT 0.000 547.080 8.280 565.480 ;
        RECT 3156.520 547.080 3165.000 565.480 ;
        RECT 0.000 515.480 3165.000 547.080 ;
        RECT 0.000 481.080 8.280 515.480 ;
        RECT 3156.520 481.080 3165.000 515.480 ;
        RECT 0.000 445.480 3165.000 481.080 ;
        RECT 0.000 427.080 8.280 445.480 ;
        RECT 3156.520 427.080 3165.000 445.480 ;
        RECT 0.000 395.480 3165.000 427.080 ;
        RECT 0.000 361.080 8.280 395.480 ;
        RECT 3156.520 361.080 3165.000 395.480 ;
        RECT 0.000 325.480 3165.000 361.080 ;
        RECT 0.000 307.080 8.280 325.480 ;
        RECT 3156.520 307.080 3165.000 325.480 ;
        RECT 0.000 275.480 3165.000 307.080 ;
        RECT 0.000 241.080 8.280 275.480 ;
        RECT 3156.520 241.080 3165.000 275.480 ;
        RECT 0.000 205.480 3165.000 241.080 ;
      LAYER met5 ;
        RECT -9.290 180.250 0.000 204.200 ;
      LAYER met5 ;
        RECT 0.000 187.080 26.400 205.480 ;
        RECT 3156.520 187.080 3165.000 205.480 ;
        RECT 0.000 172.980 3165.000 187.080 ;
      LAYER met5 ;
        RECT -9.290 130.050 0.000 154.000 ;
      LAYER met5 ;
        RECT 0.000 143.780 648.400 172.980 ;
        RECT 1083.715 143.780 3165.000 172.980 ;
        RECT 0.000 130.050 3165.000 143.780 ;
  END
END caravel_core
END LIBRARY

