magic
tech sky130A
magscale 1 2
timestamp 1651019166
<< viali >>
rect 658360 47209 658394 47243
<< metal1 >>
rect 655422 896996 655428 897048
rect 655480 897036 655486 897048
rect 676030 897036 676036 897048
rect 655480 897008 676036 897036
rect 655480 896996 655486 897008
rect 676030 896996 676036 897008
rect 676088 896996 676094 897048
rect 673362 894616 673368 894668
rect 673420 894656 673426 894668
rect 675938 894656 675944 894668
rect 673420 894628 675944 894656
rect 673420 894616 673426 894628
rect 675938 894616 675944 894628
rect 675996 894616 676002 894668
rect 655606 894344 655612 894396
rect 655664 894384 655670 894396
rect 676030 894384 676036 894396
rect 655664 894356 676036 894384
rect 655664 894344 655670 894356
rect 676030 894344 676036 894356
rect 676088 894344 676094 894396
rect 655514 894276 655520 894328
rect 655572 894316 655578 894328
rect 676122 894316 676128 894328
rect 655572 894288 676128 894316
rect 655572 894276 655578 894288
rect 676122 894276 676128 894288
rect 676180 894276 676186 894328
rect 673270 892984 673276 893036
rect 673328 893024 673334 893036
rect 676030 893024 676036 893036
rect 673328 892996 676036 893024
rect 673328 892984 673334 892996
rect 676030 892984 676036 892996
rect 676088 892984 676094 893036
rect 674742 891488 674748 891540
rect 674800 891528 674806 891540
rect 676030 891528 676036 891540
rect 674800 891500 676036 891528
rect 674800 891488 674806 891500
rect 676030 891488 676036 891500
rect 676088 891488 676094 891540
rect 674926 890672 674932 890724
rect 674984 890712 674990 890724
rect 676030 890712 676036 890724
rect 674984 890684 676036 890712
rect 674984 890672 674990 890684
rect 676030 890672 676036 890684
rect 676088 890672 676094 890724
rect 675018 889040 675024 889092
rect 675076 889080 675082 889092
rect 676030 889080 676036 889092
rect 675076 889052 676036 889080
rect 675076 889040 675082 889052
rect 676030 889040 676036 889052
rect 676088 889040 676094 889092
rect 675202 888700 675208 888752
rect 675260 888740 675266 888752
rect 676030 888740 676036 888752
rect 675260 888712 676036 888740
rect 675260 888700 675266 888712
rect 676030 888700 676036 888712
rect 676088 888700 676094 888752
rect 673730 887816 673736 887868
rect 673788 887856 673794 887868
rect 676030 887856 676036 887868
rect 673788 887828 676036 887856
rect 673788 887816 673794 887828
rect 676030 887816 676036 887828
rect 676088 887816 676094 887868
rect 674282 887408 674288 887460
rect 674340 887448 674346 887460
rect 676030 887448 676036 887460
rect 674340 887420 676036 887448
rect 674340 887408 674346 887420
rect 676030 887408 676036 887420
rect 676088 887408 676094 887460
rect 674190 885980 674196 886032
rect 674248 886020 674254 886032
rect 676030 886020 676036 886032
rect 674248 885992 676036 886020
rect 674248 885980 674254 885992
rect 676030 885980 676036 885992
rect 676088 885980 676094 886032
rect 671982 884960 671988 885012
rect 672040 885000 672046 885012
rect 678974 885000 678980 885012
rect 672040 884972 678980 885000
rect 672040 884960 672046 884972
rect 678974 884960 678980 884972
rect 679032 884960 679038 885012
rect 655698 883260 655704 883312
rect 655756 883300 655762 883312
rect 675386 883300 675392 883312
rect 655756 883272 675392 883300
rect 655756 883260 655762 883272
rect 675386 883260 675392 883272
rect 675444 883260 675450 883312
rect 674466 880676 674472 880728
rect 674524 880716 674530 880728
rect 675202 880716 675208 880728
rect 674524 880688 675208 880716
rect 674524 880676 674530 880688
rect 675202 880676 675208 880688
rect 675260 880676 675266 880728
rect 674834 880608 674840 880660
rect 674892 880648 674898 880660
rect 680262 880648 680268 880660
rect 674892 880620 680268 880648
rect 674892 880608 674898 880620
rect 680262 880608 680268 880620
rect 680320 880608 680326 880660
rect 675202 880540 675208 880592
rect 675260 880580 675266 880592
rect 679158 880580 679164 880592
rect 675260 880552 679164 880580
rect 675260 880540 675266 880552
rect 679158 880540 679164 880552
rect 679216 880540 679222 880592
rect 675294 880472 675300 880524
rect 675352 880512 675358 880524
rect 679434 880512 679440 880524
rect 675352 880484 679440 880512
rect 675352 880472 675358 880484
rect 679434 880472 679440 880484
rect 679492 880472 679498 880524
rect 675110 878772 675116 878824
rect 675168 878812 675174 878824
rect 679250 878812 679256 878824
rect 675168 878784 679256 878812
rect 675168 878772 675174 878784
rect 679250 878772 679256 878784
rect 679308 878772 679314 878824
rect 674558 878636 674564 878688
rect 674616 878676 674622 878688
rect 679526 878676 679532 878688
rect 674616 878648 679532 878676
rect 674616 878636 674622 878648
rect 679526 878636 679532 878648
rect 679584 878636 679590 878688
rect 674650 878568 674656 878620
rect 674708 878608 674714 878620
rect 679710 878608 679716 878620
rect 674708 878580 679716 878608
rect 674708 878568 674714 878580
rect 679710 878568 679716 878580
rect 679768 878568 679774 878620
rect 674926 878500 674932 878552
rect 674984 878540 674990 878552
rect 679066 878540 679072 878552
rect 674984 878512 679072 878540
rect 674984 878500 674990 878512
rect 679066 878500 679072 878512
rect 679124 878500 679130 878552
rect 674834 877208 674840 877260
rect 674892 877248 674898 877260
rect 675386 877248 675392 877260
rect 674892 877220 675392 877248
rect 674892 877208 674898 877220
rect 675386 877208 675392 877220
rect 675444 877208 675450 877260
rect 674374 875848 674380 875900
rect 674432 875888 674438 875900
rect 674834 875888 674840 875900
rect 674432 875860 674840 875888
rect 674432 875848 674438 875860
rect 674834 875848 674840 875860
rect 674892 875848 674898 875900
rect 674650 874284 674656 874336
rect 674708 874324 674714 874336
rect 675110 874324 675116 874336
rect 674708 874296 675116 874324
rect 674708 874284 674714 874296
rect 675110 874284 675116 874296
rect 675168 874284 675174 874336
rect 673730 874148 673736 874200
rect 673788 874188 673794 874200
rect 674650 874188 674656 874200
rect 673788 874160 674656 874188
rect 673788 874148 673794 874160
rect 674650 874148 674656 874160
rect 674708 874148 674714 874200
rect 674558 873740 674564 873792
rect 674616 873780 674622 873792
rect 675110 873780 675116 873792
rect 674616 873752 675116 873780
rect 674616 873740 674622 873752
rect 675110 873740 675116 873752
rect 675168 873740 675174 873792
rect 675018 872720 675024 872772
rect 675076 872720 675082 872772
rect 675036 872568 675064 872720
rect 675018 872516 675024 872568
rect 675076 872516 675082 872568
rect 674742 872448 674748 872500
rect 674800 872488 674806 872500
rect 675202 872488 675208 872500
rect 674800 872460 675208 872488
rect 674800 872448 674806 872460
rect 675202 872448 675208 872460
rect 675260 872448 675266 872500
rect 655790 872176 655796 872228
rect 655848 872216 655854 872228
rect 675110 872216 675116 872228
rect 655848 872188 675116 872216
rect 655848 872176 655854 872188
rect 675110 872176 675116 872188
rect 675168 872176 675174 872228
rect 674282 869932 674288 869984
rect 674340 869972 674346 869984
rect 675202 869972 675208 869984
rect 674340 869944 675208 869972
rect 674340 869932 674346 869944
rect 675202 869932 675208 869944
rect 675260 869932 675266 869984
rect 674190 869388 674196 869440
rect 674248 869428 674254 869440
rect 675202 869428 675208 869440
rect 674248 869400 675208 869428
rect 674248 869388 674254 869400
rect 675202 869388 675208 869400
rect 675260 869388 675266 869440
rect 674650 869320 674656 869372
rect 674708 869360 674714 869372
rect 675294 869360 675300 869372
rect 674708 869332 675300 869360
rect 674708 869320 674714 869332
rect 675294 869320 675300 869332
rect 675352 869320 675358 869372
rect 674466 867552 674472 867604
rect 674524 867592 674530 867604
rect 675110 867592 675116 867604
rect 674524 867564 675116 867592
rect 674524 867552 674530 867564
rect 675110 867552 675116 867564
rect 675168 867552 675174 867604
rect 674742 865716 674748 865768
rect 674800 865756 674806 865768
rect 675202 865756 675208 865768
rect 674800 865728 675208 865756
rect 674800 865716 674806 865728
rect 675202 865716 675208 865728
rect 675260 865716 675266 865768
rect 656802 863812 656808 863864
rect 656860 863852 656866 863864
rect 675110 863852 675116 863864
rect 656860 863824 675116 863852
rect 656860 863812 656866 863824
rect 675110 863812 675116 863824
rect 675168 863812 675174 863864
rect 41782 817640 41788 817692
rect 41840 817680 41846 817692
rect 50982 817680 50988 817692
rect 41840 817652 50988 817680
rect 41840 817640 41846 817652
rect 50982 817640 50988 817652
rect 51040 817640 51046 817692
rect 41782 817232 41788 817284
rect 41840 817272 41846 817284
rect 48222 817272 48228 817284
rect 41840 817244 48228 817272
rect 41840 817232 41846 817244
rect 48222 817232 48228 817244
rect 48280 817232 48286 817284
rect 41782 816824 41788 816876
rect 41840 816864 41846 816876
rect 45554 816864 45560 816876
rect 41840 816836 45560 816864
rect 41840 816824 41846 816836
rect 45554 816824 45560 816836
rect 45612 816824 45618 816876
rect 41782 815668 41788 815720
rect 41840 815708 41846 815720
rect 43806 815708 43812 815720
rect 41840 815680 43812 815708
rect 41840 815668 41846 815680
rect 43806 815668 43812 815680
rect 43864 815668 43870 815720
rect 41782 814512 41788 814564
rect 41840 814552 41846 814564
rect 43622 814552 43628 814564
rect 41840 814524 43628 814552
rect 41840 814512 41846 814524
rect 43622 814512 43628 814524
rect 43680 814512 43686 814564
rect 41782 814376 41788 814428
rect 41840 814416 41846 814428
rect 43530 814416 43536 814428
rect 41840 814388 43536 814416
rect 41840 814376 41846 814388
rect 43530 814376 43536 814388
rect 43588 814376 43594 814428
rect 41782 813288 41788 813340
rect 41840 813328 41846 813340
rect 43346 813328 43352 813340
rect 41840 813300 43352 813328
rect 41840 813288 41846 813300
rect 43346 813288 43352 813300
rect 43404 813288 43410 813340
rect 41782 812880 41788 812932
rect 41840 812920 41846 812932
rect 42794 812920 42800 812932
rect 41840 812892 42800 812920
rect 41840 812880 41846 812892
rect 42794 812880 42800 812892
rect 42852 812880 42858 812932
rect 41782 812744 41788 812796
rect 41840 812784 41846 812796
rect 42702 812784 42708 812796
rect 41840 812756 42708 812784
rect 41840 812744 41846 812756
rect 42702 812744 42708 812756
rect 42760 812744 42766 812796
rect 41782 811452 41788 811504
rect 41840 811492 41846 811504
rect 43438 811492 43444 811504
rect 41840 811464 43444 811492
rect 41840 811452 41846 811464
rect 43438 811452 43444 811464
rect 43496 811452 43502 811504
rect 41782 810092 41788 810144
rect 41840 810132 41846 810144
rect 43898 810132 43904 810144
rect 41840 810104 43904 810132
rect 41840 810092 41846 810104
rect 43898 810092 43904 810104
rect 43956 810092 43962 810144
rect 41874 808800 41880 808852
rect 41932 808840 41938 808852
rect 44082 808840 44088 808852
rect 41932 808812 44088 808840
rect 41932 808800 41938 808812
rect 44082 808800 44088 808812
rect 44140 808800 44146 808852
rect 41782 808664 41788 808716
rect 41840 808704 41846 808716
rect 43254 808704 43260 808716
rect 41840 808676 43260 808704
rect 41840 808664 41846 808676
rect 43254 808664 43260 808676
rect 43312 808664 43318 808716
rect 41782 807984 41788 808036
rect 41840 808024 41846 808036
rect 43070 808024 43076 808036
rect 41840 807996 43076 808024
rect 41840 807984 41846 807996
rect 43070 807984 43076 807996
rect 43128 807984 43134 808036
rect 41782 806012 41788 806064
rect 41840 806052 41846 806064
rect 42978 806052 42984 806064
rect 41840 806024 42984 806052
rect 41840 806012 41846 806024
rect 42978 806012 42984 806024
rect 43036 806012 43042 806064
rect 42058 805944 42064 805996
rect 42116 805984 42122 805996
rect 45462 805984 45468 805996
rect 42116 805956 45468 805984
rect 42116 805944 42122 805956
rect 45462 805944 45468 805956
rect 45520 805944 45526 805996
rect 41874 803088 41880 803140
rect 41932 803128 41938 803140
rect 42886 803128 42892 803140
rect 41932 803100 42892 803128
rect 41932 803088 41938 803100
rect 42886 803088 42892 803100
rect 42944 803088 42950 803140
rect 41966 803020 41972 803072
rect 42024 803060 42030 803072
rect 43162 803060 43168 803072
rect 42024 803032 43168 803060
rect 42024 803020 42030 803032
rect 43162 803020 43168 803032
rect 43220 803020 43226 803072
rect 42334 800436 42340 800488
rect 42392 800476 42398 800488
rect 58250 800476 58256 800488
rect 42392 800448 58256 800476
rect 42392 800436 42398 800448
rect 58250 800436 58256 800448
rect 58308 800436 58314 800488
rect 42334 798940 42340 798992
rect 42392 798980 42398 798992
rect 42794 798980 42800 798992
rect 42392 798952 42800 798980
rect 42392 798940 42398 798952
rect 42794 798940 42800 798952
rect 42852 798940 42858 798992
rect 42150 798124 42156 798176
rect 42208 798164 42214 798176
rect 42702 798164 42708 798176
rect 42208 798136 42708 798164
rect 42208 798124 42214 798136
rect 42702 798124 42708 798136
rect 42760 798124 42766 798176
rect 42702 797988 42708 798040
rect 42760 798028 42766 798040
rect 43162 798028 43168 798040
rect 42760 798000 43168 798028
rect 42760 797988 42766 798000
rect 43162 797988 43168 798000
rect 43220 797988 43226 798040
rect 43530 797920 43536 797972
rect 43588 797920 43594 797972
rect 43162 797852 43168 797904
rect 43220 797892 43226 797904
rect 43346 797892 43352 797904
rect 43220 797864 43352 797892
rect 43220 797852 43226 797864
rect 43346 797852 43352 797864
rect 43404 797852 43410 797904
rect 43346 797716 43352 797768
rect 43404 797756 43410 797768
rect 43548 797756 43576 797920
rect 43714 797784 43720 797836
rect 43772 797784 43778 797836
rect 43404 797728 43576 797756
rect 43404 797716 43410 797728
rect 43732 797700 43760 797784
rect 43714 797648 43720 797700
rect 43772 797648 43778 797700
rect 42334 796696 42340 796748
rect 42392 796736 42398 796748
rect 43254 796736 43260 796748
rect 42392 796708 43260 796736
rect 42392 796696 42398 796708
rect 43254 796696 43260 796708
rect 43312 796696 43318 796748
rect 42242 795880 42248 795932
rect 42300 795920 42306 795932
rect 43254 795920 43260 795932
rect 42300 795892 43260 795920
rect 42300 795880 42306 795892
rect 43254 795880 43260 795892
rect 43312 795880 43318 795932
rect 42242 794996 42248 795048
rect 42300 795036 42306 795048
rect 42978 795036 42984 795048
rect 42300 795008 42984 795036
rect 42300 794996 42306 795008
rect 42978 794996 42984 795008
rect 43036 794996 43042 795048
rect 42242 794452 42248 794504
rect 42300 794492 42306 794504
rect 42702 794492 42708 794504
rect 42300 794464 42708 794492
rect 42300 794452 42306 794464
rect 42702 794452 42708 794464
rect 42760 794452 42766 794504
rect 43622 794044 43628 794096
rect 43680 794084 43686 794096
rect 43806 794084 43812 794096
rect 43680 794056 43812 794084
rect 43680 794044 43686 794056
rect 43806 794044 43812 794056
rect 43864 794044 43870 794096
rect 42150 793772 42156 793824
rect 42208 793812 42214 793824
rect 43070 793812 43076 793824
rect 42208 793784 43076 793812
rect 42208 793772 42214 793784
rect 43070 793772 43076 793784
rect 43128 793772 43134 793824
rect 42334 792208 42340 792260
rect 42392 792248 42398 792260
rect 42702 792248 42708 792260
rect 42392 792220 42708 792248
rect 42392 792208 42398 792220
rect 42702 792208 42708 792220
rect 42760 792208 42766 792260
rect 655514 792140 655520 792192
rect 655572 792180 655578 792192
rect 675386 792180 675392 792192
rect 655572 792152 675392 792180
rect 655572 792140 655578 792152
rect 675386 792140 675392 792152
rect 675444 792140 675450 792192
rect 42150 790644 42156 790696
rect 42208 790684 42214 790696
rect 42886 790684 42892 790696
rect 42208 790656 42892 790684
rect 42208 790644 42214 790656
rect 42886 790644 42892 790656
rect 42944 790644 42950 790696
rect 42242 789488 42248 789540
rect 42300 789528 42306 789540
rect 43714 789528 43720 789540
rect 42300 789500 43720 789528
rect 42300 789488 42306 789500
rect 43714 789488 43720 789500
rect 43772 789488 43778 789540
rect 42426 789352 42432 789404
rect 42484 789392 42490 789404
rect 58158 789392 58164 789404
rect 42484 789364 58164 789392
rect 42484 789352 42490 789364
rect 58158 789352 58164 789364
rect 58216 789352 58222 789404
rect 42702 789284 42708 789336
rect 42760 789324 42766 789336
rect 58526 789324 58532 789336
rect 42760 789296 58532 789324
rect 42760 789284 42766 789296
rect 58526 789284 58532 789296
rect 58584 789284 58590 789336
rect 42150 789216 42156 789268
rect 42208 789256 42214 789268
rect 44082 789256 44088 789268
rect 42208 789228 44088 789256
rect 42208 789216 42214 789228
rect 44082 789216 44088 789228
rect 44140 789216 44146 789268
rect 45554 789216 45560 789268
rect 45612 789256 45618 789268
rect 58434 789256 58440 789268
rect 45612 789228 58440 789256
rect 45612 789216 45618 789228
rect 58434 789216 58440 789228
rect 58492 789216 58498 789268
rect 42334 789148 42340 789200
rect 42392 789188 42398 789200
rect 43254 789188 43260 789200
rect 42392 789160 43260 789188
rect 42392 789148 42398 789160
rect 43254 789148 43260 789160
rect 43312 789148 43318 789200
rect 48222 786564 48228 786616
rect 48280 786604 48286 786616
rect 58434 786604 58440 786616
rect 48280 786576 58440 786604
rect 48280 786564 48286 786576
rect 58434 786564 58440 786576
rect 58492 786564 58498 786616
rect 50982 786496 50988 786548
rect 51040 786536 51046 786548
rect 58526 786536 58532 786548
rect 51040 786508 58532 786536
rect 51040 786496 51046 786508
rect 58526 786496 58532 786508
rect 58584 786496 58590 786548
rect 42334 786428 42340 786480
rect 42392 786468 42398 786480
rect 43438 786468 43444 786480
rect 42392 786440 43444 786468
rect 42392 786428 42398 786440
rect 43438 786428 43444 786440
rect 43496 786428 43502 786480
rect 42058 786224 42064 786276
rect 42116 786264 42122 786276
rect 43898 786264 43904 786276
rect 42116 786236 43904 786264
rect 42116 786224 42122 786236
rect 43898 786224 43904 786236
rect 43956 786224 43962 786276
rect 673822 784728 673828 784780
rect 673880 784768 673886 784780
rect 675110 784768 675116 784780
rect 673880 784740 675116 784768
rect 673880 784728 673886 784740
rect 675110 784728 675116 784740
rect 675168 784728 675174 784780
rect 656526 783844 656532 783896
rect 656584 783884 656590 783896
rect 675110 783884 675116 783896
rect 656584 783856 675116 783884
rect 656584 783844 656590 783856
rect 675110 783844 675116 783856
rect 675168 783844 675174 783896
rect 674558 780444 674564 780496
rect 674616 780484 674622 780496
rect 675478 780484 675484 780496
rect 674616 780456 675484 780484
rect 674616 780444 674622 780456
rect 675478 780444 675484 780456
rect 675536 780444 675542 780496
rect 674282 779968 674288 780020
rect 674340 780008 674346 780020
rect 675478 780008 675484 780020
rect 674340 779980 675484 780008
rect 674340 779968 674346 779980
rect 675478 779968 675484 779980
rect 675536 779968 675542 780020
rect 673638 779764 673644 779816
rect 673696 779804 673702 779816
rect 675202 779804 675208 779816
rect 673696 779776 675208 779804
rect 673696 779764 673702 779776
rect 675202 779764 675208 779776
rect 675260 779764 675266 779816
rect 673730 778744 673736 778796
rect 673788 778784 673794 778796
rect 675478 778784 675484 778796
rect 673788 778756 675484 778784
rect 673788 778744 673794 778756
rect 675478 778744 675484 778756
rect 675536 778744 675542 778796
rect 674466 778540 674472 778592
rect 674524 778580 674530 778592
rect 675202 778580 675208 778592
rect 674524 778552 675208 778580
rect 674524 778540 674530 778552
rect 675202 778540 675208 778552
rect 675260 778540 675266 778592
rect 674650 777316 674656 777368
rect 674708 777356 674714 777368
rect 675386 777356 675392 777368
rect 674708 777328 675392 777356
rect 674708 777316 674714 777328
rect 675386 777316 675392 777328
rect 675444 777316 675450 777368
rect 675018 776840 675024 776892
rect 675076 776840 675082 776892
rect 675036 776688 675064 776840
rect 675018 776636 675024 776688
rect 675076 776636 675082 776688
rect 654962 775480 654968 775532
rect 655020 775520 655026 775532
rect 675110 775520 675116 775532
rect 655020 775492 675116 775520
rect 655020 775480 655026 775492
rect 675110 775480 675116 775492
rect 675168 775480 675174 775532
rect 41782 774392 41788 774444
rect 41840 774432 41846 774444
rect 50982 774432 50988 774444
rect 41840 774404 50988 774432
rect 41840 774392 41846 774404
rect 50982 774392 50988 774404
rect 51040 774392 51046 774444
rect 41506 774256 41512 774308
rect 41564 774296 41570 774308
rect 43622 774296 43628 774308
rect 41564 774268 43628 774296
rect 41564 774256 41570 774268
rect 43622 774256 43628 774268
rect 43680 774256 43686 774308
rect 41414 773848 41420 773900
rect 41472 773888 41478 773900
rect 48222 773888 48228 773900
rect 41472 773860 48228 773888
rect 41472 773848 41478 773860
rect 48222 773848 48228 773860
rect 48280 773848 48286 773900
rect 41782 773576 41788 773628
rect 41840 773616 41846 773628
rect 45738 773616 45744 773628
rect 41840 773588 45744 773616
rect 41840 773576 41846 773588
rect 45738 773576 45744 773588
rect 45796 773576 45802 773628
rect 675018 773372 675024 773424
rect 675076 773412 675082 773424
rect 675662 773412 675668 773424
rect 675076 773384 675668 773412
rect 675076 773372 675082 773384
rect 675662 773372 675668 773384
rect 675720 773372 675726 773424
rect 674742 773304 674748 773356
rect 674800 773344 674806 773356
rect 675754 773344 675760 773356
rect 674800 773316 675760 773344
rect 674800 773304 674806 773316
rect 675754 773304 675760 773316
rect 675812 773304 675818 773356
rect 41874 772828 41880 772880
rect 41932 772868 41938 772880
rect 44082 772868 44088 772880
rect 41932 772840 44088 772868
rect 41932 772828 41938 772840
rect 44082 772828 44088 772840
rect 44140 772828 44146 772880
rect 41782 772760 41788 772812
rect 41840 772800 41846 772812
rect 43346 772800 43352 772812
rect 41840 772772 43352 772800
rect 41840 772760 41846 772772
rect 43346 772760 43352 772772
rect 43404 772760 43410 772812
rect 41506 772692 41512 772744
rect 41564 772732 41570 772744
rect 43530 772732 43536 772744
rect 41564 772704 43536 772732
rect 41564 772692 41570 772704
rect 43530 772692 43536 772704
rect 43588 772692 43594 772744
rect 41782 771468 41788 771520
rect 41840 771508 41846 771520
rect 43162 771508 43168 771520
rect 41840 771480 43168 771508
rect 41840 771468 41846 771480
rect 43162 771468 43168 771480
rect 43220 771468 43226 771520
rect 41414 770992 41420 771044
rect 41472 771032 41478 771044
rect 43162 771032 43168 771044
rect 41472 771004 43168 771032
rect 41472 770992 41478 771004
rect 43162 770992 43168 771004
rect 43220 770992 43226 771044
rect 41506 770312 41512 770364
rect 41564 770352 41570 770364
rect 42426 770352 42432 770364
rect 41564 770324 42432 770352
rect 41564 770312 41570 770324
rect 42426 770312 42432 770324
rect 42484 770312 42490 770364
rect 41506 769496 41512 769548
rect 41564 769536 41570 769548
rect 43254 769536 43260 769548
rect 41564 769508 43260 769536
rect 41564 769496 41570 769508
rect 43254 769496 43260 769508
rect 43312 769496 43318 769548
rect 41506 769360 41512 769412
rect 41564 769400 41570 769412
rect 43070 769400 43076 769412
rect 41564 769372 43076 769400
rect 41564 769360 41570 769372
rect 43070 769360 43076 769372
rect 43128 769360 43134 769412
rect 41506 768952 41512 769004
rect 41564 768992 41570 769004
rect 43714 768992 43720 769004
rect 41564 768964 43720 768992
rect 41564 768952 41570 768964
rect 43714 768952 43720 768964
rect 43772 768952 43778 769004
rect 41506 768272 41512 768324
rect 41564 768312 41570 768324
rect 43438 768312 43444 768324
rect 41564 768284 43444 768312
rect 41564 768272 41570 768284
rect 43438 768272 43444 768284
rect 43496 768272 43502 768324
rect 41506 768136 41512 768188
rect 41564 768176 41570 768188
rect 43346 768176 43352 768188
rect 41564 768148 43352 768176
rect 41564 768136 41570 768148
rect 43346 768136 43352 768148
rect 43404 768136 43410 768188
rect 41506 767388 41512 767440
rect 41564 767428 41570 767440
rect 43530 767428 43536 767440
rect 41564 767400 43536 767428
rect 41564 767388 41570 767400
rect 43530 767388 43536 767400
rect 43588 767388 43594 767440
rect 42702 767320 42708 767372
rect 42760 767360 42766 767372
rect 45646 767360 45652 767372
rect 42760 767332 45652 767360
rect 42760 767320 42766 767332
rect 45646 767320 45652 767332
rect 45704 767320 45710 767372
rect 674650 767320 674656 767372
rect 674708 767360 674714 767372
rect 674926 767360 674932 767372
rect 674708 767332 674932 767360
rect 674708 767320 674714 767332
rect 674926 767320 674932 767332
rect 674984 767320 674990 767372
rect 43530 766300 43536 766352
rect 43588 766340 43594 766352
rect 43990 766340 43996 766352
rect 43588 766312 43996 766340
rect 43588 766300 43594 766312
rect 43990 766300 43996 766312
rect 44048 766300 44054 766352
rect 41506 766096 41512 766148
rect 41564 766136 41570 766148
rect 42426 766136 42432 766148
rect 41564 766108 42432 766136
rect 41564 766096 41570 766108
rect 42426 766096 42432 766108
rect 42484 766096 42490 766148
rect 43346 765824 43352 765876
rect 43404 765864 43410 765876
rect 43622 765864 43628 765876
rect 43404 765836 43628 765864
rect 43404 765824 43410 765836
rect 43622 765824 43628 765836
rect 43680 765824 43686 765876
rect 41506 765688 41512 765740
rect 41564 765728 41570 765740
rect 43346 765728 43352 765740
rect 41564 765700 43352 765728
rect 41564 765688 41570 765700
rect 43346 765688 43352 765700
rect 43404 765688 43410 765740
rect 41506 764872 41512 764924
rect 41564 764912 41570 764924
rect 43806 764912 43812 764924
rect 41564 764884 43812 764912
rect 41564 764872 41570 764884
rect 43806 764872 43812 764884
rect 43864 764872 43870 764924
rect 41506 764532 41512 764584
rect 41564 764572 41570 764584
rect 42702 764572 42708 764584
rect 41564 764544 42708 764572
rect 41564 764532 41570 764544
rect 42702 764532 42708 764544
rect 42760 764532 42766 764584
rect 41506 762832 41512 762884
rect 41564 762872 41570 762884
rect 45554 762872 45560 762884
rect 41564 762844 45560 762872
rect 41564 762832 41570 762844
rect 45554 762832 45560 762844
rect 45612 762832 45618 762884
rect 41782 761744 41788 761796
rect 41840 761784 41846 761796
rect 42242 761784 42248 761796
rect 41840 761756 42248 761784
rect 41840 761744 41846 761756
rect 42242 761744 42248 761756
rect 42300 761744 42306 761796
rect 42334 760928 42340 760980
rect 42392 760968 42398 760980
rect 43622 760968 43628 760980
rect 42392 760940 43628 760968
rect 42392 760928 42398 760940
rect 43622 760928 43628 760940
rect 43680 760928 43686 760980
rect 42334 760792 42340 760844
rect 42392 760832 42398 760844
rect 43070 760832 43076 760844
rect 42392 760804 43076 760832
rect 42392 760792 42398 760804
rect 43070 760792 43076 760804
rect 43128 760792 43134 760844
rect 42426 760656 42432 760708
rect 42484 760696 42490 760708
rect 43070 760696 43076 760708
rect 42484 760668 43076 760696
rect 42484 760656 42490 760668
rect 43070 760656 43076 760668
rect 43128 760656 43134 760708
rect 41598 759296 41604 759348
rect 41656 759336 41662 759348
rect 43898 759336 43904 759348
rect 41656 759308 43904 759336
rect 41656 759296 41662 759308
rect 43898 759296 43904 759308
rect 43956 759296 43962 759348
rect 41414 759024 41420 759076
rect 41472 759064 41478 759076
rect 44174 759064 44180 759076
rect 41472 759036 44180 759064
rect 41472 759024 41478 759036
rect 44174 759024 44180 759036
rect 44232 759024 44238 759076
rect 43346 757800 43352 757852
rect 43404 757840 43410 757852
rect 43404 757812 43484 757840
rect 43404 757800 43410 757812
rect 43456 757512 43484 757812
rect 43530 757664 43536 757716
rect 43588 757664 43594 757716
rect 43162 757460 43168 757512
rect 43220 757500 43226 757512
rect 43346 757500 43352 757512
rect 43220 757472 43352 757500
rect 43220 757460 43226 757472
rect 43346 757460 43352 757472
rect 43404 757460 43410 757512
rect 43438 757460 43444 757512
rect 43496 757460 43502 757512
rect 43548 757432 43576 757664
rect 674650 757596 674656 757648
rect 674708 757636 674714 757648
rect 675294 757636 675300 757648
rect 674708 757608 675300 757636
rect 674708 757596 674714 757608
rect 675294 757596 675300 757608
rect 675352 757596 675358 757648
rect 43548 757404 43852 757432
rect 43346 757324 43352 757376
rect 43404 757364 43410 757376
rect 43714 757364 43720 757376
rect 43404 757336 43720 757364
rect 43404 757324 43410 757336
rect 43714 757324 43720 757336
rect 43772 757324 43778 757376
rect 43714 757188 43720 757240
rect 43772 757228 43778 757240
rect 43824 757228 43852 757404
rect 43772 757200 43852 757228
rect 43772 757188 43778 757200
rect 42242 756236 42248 756288
rect 42300 756276 42306 756288
rect 59262 756276 59268 756288
rect 42300 756248 59268 756276
rect 42300 756236 42306 756248
rect 59262 756236 59268 756248
rect 59320 756236 59326 756288
rect 42150 754876 42156 754928
rect 42208 754916 42214 754928
rect 42334 754916 42340 754928
rect 42208 754888 42340 754916
rect 42208 754876 42214 754888
rect 42334 754876 42340 754888
rect 42392 754876 42398 754928
rect 42334 754264 42340 754316
rect 42392 754304 42398 754316
rect 42702 754304 42708 754316
rect 42392 754276 42708 754304
rect 42392 754264 42398 754276
rect 42702 754264 42708 754276
rect 42760 754264 42766 754316
rect 42150 753312 42156 753364
rect 42208 753352 42214 753364
rect 42702 753352 42708 753364
rect 42208 753324 42708 753352
rect 42208 753312 42214 753324
rect 42702 753312 42708 753324
rect 42760 753312 42766 753364
rect 42150 753040 42156 753092
rect 42208 753080 42214 753092
rect 43070 753080 43076 753092
rect 42208 753052 43076 753080
rect 42208 753040 42214 753052
rect 43070 753040 43076 753052
rect 43128 753040 43134 753092
rect 42334 751204 42340 751256
rect 42392 751244 42398 751256
rect 43438 751244 43444 751256
rect 42392 751216 43444 751244
rect 42392 751204 42398 751216
rect 43438 751204 43444 751216
rect 43496 751204 43502 751256
rect 43530 751136 43536 751188
rect 43588 751136 43594 751188
rect 43548 750984 43576 751136
rect 43530 750932 43536 750984
rect 43588 750932 43594 750984
rect 42058 750592 42064 750644
rect 42116 750632 42122 750644
rect 43806 750632 43812 750644
rect 42116 750604 43812 750632
rect 42116 750592 42122 750604
rect 43806 750592 43812 750604
rect 43864 750592 43870 750644
rect 42334 750524 42340 750576
rect 42392 750564 42398 750576
rect 43898 750564 43904 750576
rect 42392 750536 43904 750564
rect 42392 750524 42398 750536
rect 43898 750524 43904 750536
rect 43956 750524 43962 750576
rect 42242 750456 42248 750508
rect 42300 750496 42306 750508
rect 43714 750496 43720 750508
rect 42300 750468 43720 750496
rect 42300 750456 42306 750468
rect 43714 750456 43720 750468
rect 43772 750456 43778 750508
rect 43806 750456 43812 750508
rect 43864 750496 43870 750508
rect 44174 750496 44180 750508
rect 43864 750468 44180 750496
rect 43864 750456 43870 750468
rect 44174 750456 44180 750468
rect 44232 750456 44238 750508
rect 42702 750388 42708 750440
rect 42760 750428 42766 750440
rect 43898 750428 43904 750440
rect 42760 750400 43904 750428
rect 42760 750388 42766 750400
rect 43898 750388 43904 750400
rect 43956 750388 43962 750440
rect 43070 750320 43076 750372
rect 43128 750360 43134 750372
rect 43714 750360 43720 750372
rect 43128 750332 43720 750360
rect 43128 750320 43134 750332
rect 43714 750320 43720 750332
rect 43772 750320 43778 750372
rect 655974 747940 655980 747992
rect 656032 747980 656038 747992
rect 675386 747980 675392 747992
rect 656032 747952 675392 747980
rect 656032 747940 656038 747952
rect 675386 747940 675392 747952
rect 675444 747940 675450 747992
rect 43898 747872 43904 747924
rect 43956 747912 43962 747924
rect 58434 747912 58440 747924
rect 43956 747884 58440 747912
rect 43956 747872 43962 747884
rect 58434 747872 58440 747884
rect 58492 747872 58498 747924
rect 42334 746920 42340 746972
rect 42392 746960 42398 746972
rect 43806 746960 43812 746972
rect 42392 746932 43812 746960
rect 42392 746920 42398 746932
rect 43806 746920 43812 746932
rect 43864 746920 43870 746972
rect 42242 745560 42248 745612
rect 42300 745600 42306 745612
rect 43530 745600 43536 745612
rect 42300 745572 43536 745600
rect 42300 745560 42306 745572
rect 43530 745560 43536 745572
rect 43588 745560 43594 745612
rect 42334 745220 42340 745272
rect 42392 745260 42398 745272
rect 58434 745260 58440 745272
rect 42392 745232 58440 745260
rect 42392 745220 42398 745232
rect 58434 745220 58440 745232
rect 58492 745220 58498 745272
rect 45738 745152 45744 745204
rect 45796 745192 45802 745204
rect 58526 745192 58532 745204
rect 45796 745164 58532 745192
rect 45796 745152 45802 745164
rect 58526 745152 58532 745164
rect 58584 745152 58590 745204
rect 42242 745084 42248 745136
rect 42300 745124 42306 745136
rect 43162 745124 43168 745136
rect 42300 745096 43168 745124
rect 42300 745084 42306 745096
rect 43162 745084 43168 745096
rect 43220 745084 43226 745136
rect 673454 744200 673460 744252
rect 673512 744240 673518 744252
rect 675754 744240 675760 744252
rect 673512 744212 675760 744240
rect 673512 744200 673518 744212
rect 675754 744200 675760 744212
rect 675812 744200 675818 744252
rect 673546 744132 673552 744184
rect 673604 744172 673610 744184
rect 675662 744172 675668 744184
rect 673604 744144 675668 744172
rect 673604 744132 673610 744144
rect 675662 744132 675668 744144
rect 675720 744132 675726 744184
rect 42242 743248 42248 743300
rect 42300 743288 42306 743300
rect 43346 743288 43352 743300
rect 42300 743260 43352 743288
rect 42300 743248 42306 743260
rect 43346 743248 43352 743260
rect 43404 743248 43410 743300
rect 42150 743044 42156 743096
rect 42208 743084 42214 743096
rect 43990 743084 43996 743096
rect 42208 743056 43996 743084
rect 42208 743044 42214 743056
rect 43990 743044 43996 743056
rect 44048 743044 44054 743096
rect 48222 742364 48228 742416
rect 48280 742404 48286 742416
rect 58434 742404 58440 742416
rect 48280 742376 58440 742404
rect 48280 742364 48286 742376
rect 58434 742364 58440 742376
rect 58492 742364 58498 742416
rect 50982 742296 50988 742348
rect 51040 742336 51046 742348
rect 57974 742336 57980 742348
rect 51040 742308 57980 742336
rect 51040 742296 51046 742308
rect 57974 742296 57980 742308
rect 58032 742296 58038 742348
rect 673730 738352 673736 738404
rect 673788 738392 673794 738404
rect 674650 738392 674656 738404
rect 673788 738364 674656 738392
rect 673788 738352 673794 738364
rect 674650 738352 674656 738364
rect 674708 738352 674714 738404
rect 654318 736992 654324 737044
rect 654376 737032 654382 737044
rect 675202 737032 675208 737044
rect 654376 737004 675208 737032
rect 654376 736992 654382 737004
rect 675202 736992 675208 737004
rect 675260 736992 675266 737044
rect 656066 736924 656072 736976
rect 656124 736964 656130 736976
rect 675294 736964 675300 736976
rect 656124 736936 675300 736964
rect 656124 736924 656130 736936
rect 675294 736924 675300 736936
rect 675352 736924 675358 736976
rect 674742 735632 674748 735684
rect 674800 735672 674806 735684
rect 675386 735672 675392 735684
rect 674800 735644 675392 735672
rect 674800 735632 674806 735644
rect 675386 735632 675392 735644
rect 675444 735632 675450 735684
rect 674834 734952 674840 735004
rect 674892 734992 674898 735004
rect 675386 734992 675392 735004
rect 674892 734964 675392 734992
rect 674892 734952 674898 734964
rect 675386 734952 675392 734964
rect 675444 734952 675450 735004
rect 674282 734136 674288 734188
rect 674340 734176 674346 734188
rect 675386 734176 675392 734188
rect 674340 734148 675392 734176
rect 674340 734136 674346 734148
rect 675386 734136 675392 734148
rect 675444 734136 675450 734188
rect 675294 733728 675300 733780
rect 675352 733728 675358 733780
rect 675386 733728 675392 733780
rect 675444 733728 675450 733780
rect 675312 733440 675340 733728
rect 675294 733388 675300 733440
rect 675352 733388 675358 733440
rect 675202 733320 675208 733372
rect 675260 733360 675266 733372
rect 675404 733360 675432 733728
rect 675260 733332 675432 733360
rect 675260 733320 675266 733332
rect 673270 732436 673276 732488
rect 673328 732476 673334 732488
rect 673454 732476 673460 732488
rect 673328 732448 673460 732476
rect 673328 732436 673334 732448
rect 673454 732436 673460 732448
rect 673512 732436 673518 732488
rect 673454 732300 673460 732352
rect 673512 732340 673518 732352
rect 675386 732340 675392 732352
rect 673512 732312 675392 732340
rect 673512 732300 673518 732312
rect 675386 732300 675392 732312
rect 675444 732300 675450 732352
rect 675202 732096 675208 732148
rect 675260 732136 675266 732148
rect 675260 732108 675340 732136
rect 675260 732096 675266 732108
rect 674834 731960 674840 732012
rect 674892 732000 674898 732012
rect 675202 732000 675208 732012
rect 674892 731972 675208 732000
rect 674892 731960 674898 731972
rect 675202 731960 675208 731972
rect 675260 731960 675266 732012
rect 674834 731824 674840 731876
rect 674892 731864 674898 731876
rect 675312 731864 675340 732108
rect 674892 731836 675340 731864
rect 674892 731824 674898 731836
rect 41506 731008 41512 731060
rect 41564 731048 41570 731060
rect 50982 731048 50988 731060
rect 41564 731020 50988 731048
rect 41564 731008 41570 731020
rect 50982 731008 50988 731020
rect 51040 731008 51046 731060
rect 41782 730736 41788 730788
rect 41840 730776 41846 730788
rect 43438 730776 43444 730788
rect 41840 730748 43444 730776
rect 41840 730736 41846 730748
rect 43438 730736 43444 730748
rect 43496 730736 43502 730788
rect 41506 730600 41512 730652
rect 41564 730640 41570 730652
rect 48222 730640 48228 730652
rect 41564 730612 48228 730640
rect 41564 730600 41570 730612
rect 48222 730600 48228 730612
rect 48280 730600 48286 730652
rect 41874 730464 41880 730516
rect 41932 730504 41938 730516
rect 44082 730504 44088 730516
rect 41932 730476 44088 730504
rect 41932 730464 41938 730476
rect 44082 730464 44088 730476
rect 44140 730464 44146 730516
rect 41506 730192 41512 730244
rect 41564 730232 41570 730244
rect 45830 730232 45836 730244
rect 41564 730204 45836 730232
rect 41564 730192 41570 730204
rect 45830 730192 45836 730204
rect 45888 730192 45894 730244
rect 41506 729104 41512 729156
rect 41564 729144 41570 729156
rect 43990 729144 43996 729156
rect 41564 729116 43996 729144
rect 41564 729104 41570 729116
rect 43990 729104 43996 729116
rect 44048 729104 44054 729156
rect 673546 728832 673552 728884
rect 673604 728872 673610 728884
rect 673604 728844 675248 728872
rect 673604 728832 673610 728844
rect 675220 728816 675248 728844
rect 673270 728764 673276 728816
rect 673328 728804 673334 728816
rect 673328 728776 674880 728804
rect 673328 728764 673334 728776
rect 674852 728680 674880 728776
rect 675202 728764 675208 728816
rect 675260 728764 675266 728816
rect 674834 728628 674840 728680
rect 674892 728628 674898 728680
rect 675386 728668 675392 728680
rect 674944 728640 675392 728668
rect 41506 728560 41512 728612
rect 41564 728600 41570 728612
rect 43254 728600 43260 728612
rect 41564 728572 43260 728600
rect 41564 728560 41570 728572
rect 43254 728560 43260 728572
rect 43312 728560 43318 728612
rect 673454 728560 673460 728612
rect 673512 728600 673518 728612
rect 673730 728600 673736 728612
rect 673512 728572 673736 728600
rect 673512 728560 673518 728572
rect 673730 728560 673736 728572
rect 673788 728560 673794 728612
rect 674944 728544 674972 728640
rect 675386 728628 675392 728640
rect 675444 728628 675450 728680
rect 674926 728492 674932 728544
rect 674984 728492 674990 728544
rect 41506 727880 41512 727932
rect 41564 727920 41570 727932
rect 43714 727920 43720 727932
rect 41564 727892 43720 727920
rect 41564 727880 41570 727892
rect 43714 727880 43720 727892
rect 43772 727880 43778 727932
rect 41506 726520 41512 726572
rect 41564 726560 41570 726572
rect 43162 726560 43168 726572
rect 41564 726532 43168 726560
rect 41564 726520 41570 726532
rect 43162 726520 43168 726532
rect 43220 726520 43226 726572
rect 41782 726180 41788 726232
rect 41840 726220 41846 726232
rect 43070 726220 43076 726232
rect 41840 726192 43076 726220
rect 41840 726180 41846 726192
rect 43070 726180 43076 726192
rect 43128 726180 43134 726232
rect 41506 726112 41512 726164
rect 41564 726152 41570 726164
rect 43346 726152 43352 726164
rect 41564 726124 43352 726152
rect 41564 726112 41570 726124
rect 43346 726112 43352 726124
rect 43404 726112 43410 726164
rect 41782 725976 41788 726028
rect 41840 726016 41846 726028
rect 43714 726016 43720 726028
rect 41840 725988 43720 726016
rect 41840 725976 41846 725988
rect 43714 725976 43720 725988
rect 43772 725976 43778 726028
rect 674466 724752 674472 724804
rect 674524 724792 674530 724804
rect 675110 724792 675116 724804
rect 674524 724764 675116 724792
rect 674524 724752 674530 724764
rect 675110 724752 675116 724764
rect 675168 724752 675174 724804
rect 41506 724208 41512 724260
rect 41564 724248 41570 724260
rect 43898 724248 43904 724260
rect 41564 724220 43904 724248
rect 41564 724208 41570 724220
rect 43898 724208 43904 724220
rect 43956 724208 43962 724260
rect 41782 723392 41788 723444
rect 41840 723432 41846 723444
rect 44082 723432 44088 723444
rect 41840 723404 44088 723432
rect 41840 723392 41846 723404
rect 44082 723392 44088 723404
rect 44140 723392 44146 723444
rect 41506 723256 41512 723308
rect 41564 723296 41570 723308
rect 43530 723296 43536 723308
rect 41564 723268 43536 723296
rect 41564 723256 41570 723268
rect 43530 723256 43536 723268
rect 43588 723256 43594 723308
rect 673178 723188 673184 723240
rect 673236 723228 673242 723240
rect 679066 723228 679072 723240
rect 673236 723200 679072 723228
rect 673236 723188 673242 723200
rect 679066 723188 679072 723200
rect 679124 723188 679130 723240
rect 41782 723120 41788 723172
rect 41840 723160 41846 723172
rect 42702 723160 42708 723172
rect 41840 723132 42708 723160
rect 41840 723120 41846 723132
rect 42702 723120 42708 723132
rect 42760 723120 42766 723172
rect 673362 723120 673368 723172
rect 673420 723160 673426 723172
rect 678974 723160 678980 723172
rect 673420 723132 678980 723160
rect 673420 723120 673426 723132
rect 678974 723120 678980 723132
rect 679032 723120 679038 723172
rect 41506 722032 41512 722084
rect 41564 722072 41570 722084
rect 43438 722072 43444 722084
rect 41564 722044 43444 722072
rect 41564 722032 41570 722044
rect 43438 722032 43444 722044
rect 43496 722032 43502 722084
rect 41598 720672 41604 720724
rect 41656 720712 41662 720724
rect 43806 720712 43812 720724
rect 41656 720684 43812 720712
rect 41656 720672 41662 720684
rect 43806 720672 43812 720684
rect 43864 720672 43870 720724
rect 41506 720400 41512 720452
rect 41564 720440 41570 720452
rect 43254 720440 43260 720452
rect 41564 720412 43260 720440
rect 41564 720400 41570 720412
rect 43254 720400 43260 720412
rect 43312 720400 43318 720452
rect 41506 719584 41512 719636
rect 41564 719624 41570 719636
rect 45738 719624 45744 719636
rect 41564 719596 45744 719624
rect 41564 719584 41570 719596
rect 45738 719584 45744 719596
rect 45796 719584 45802 719636
rect 30282 716252 30288 716304
rect 30340 716292 30346 716304
rect 43622 716292 43628 716304
rect 30340 716264 43628 716292
rect 30340 716252 30346 716264
rect 43622 716252 43628 716264
rect 43680 716252 43686 716304
rect 655790 715232 655796 715284
rect 655848 715272 655854 715284
rect 675938 715272 675944 715284
rect 655848 715244 675944 715272
rect 655848 715232 655854 715244
rect 675938 715232 675944 715244
rect 675996 715232 676002 715284
rect 655606 715096 655612 715148
rect 655664 715136 655670 715148
rect 676030 715136 676036 715148
rect 655664 715108 676036 715136
rect 655664 715096 655670 715108
rect 676030 715096 676036 715108
rect 676088 715096 676094 715148
rect 655422 714960 655428 715012
rect 655480 715000 655486 715012
rect 675846 715000 675852 715012
rect 655480 714972 675852 715000
rect 655480 714960 655486 714972
rect 675846 714960 675852 714972
rect 675904 714960 675910 715012
rect 41690 714892 41696 714944
rect 41748 714932 41754 714944
rect 44266 714932 44272 714944
rect 41748 714904 44272 714932
rect 41748 714892 41754 714904
rect 44266 714892 44272 714904
rect 44324 714892 44330 714944
rect 673270 714892 673276 714944
rect 673328 714932 673334 714944
rect 676030 714932 676036 714944
rect 673328 714904 676036 714932
rect 673328 714892 673334 714904
rect 676030 714892 676036 714904
rect 676088 714892 676094 714944
rect 42334 714824 42340 714876
rect 42392 714864 42398 714876
rect 59354 714864 59360 714876
rect 42392 714836 59360 714864
rect 42392 714824 42398 714836
rect 59354 714824 59360 714836
rect 59412 714824 59418 714876
rect 674650 714756 674656 714808
rect 674708 714796 674714 714808
rect 676030 714796 676036 714808
rect 674708 714768 676036 714796
rect 674708 714756 674714 714768
rect 676030 714756 676036 714768
rect 676088 714756 676094 714808
rect 674558 714688 674564 714740
rect 674616 714728 674622 714740
rect 675754 714728 675760 714740
rect 674616 714700 675760 714728
rect 674616 714688 674622 714700
rect 675754 714688 675760 714700
rect 675812 714688 675818 714740
rect 673822 714620 673828 714672
rect 673880 714660 673886 714672
rect 675662 714660 675668 714672
rect 673880 714632 675668 714660
rect 673880 714620 673886 714632
rect 675662 714620 675668 714632
rect 675720 714620 675726 714672
rect 673454 714552 673460 714604
rect 673512 714592 673518 714604
rect 676122 714592 676128 714604
rect 673512 714564 676128 714592
rect 673512 714552 673518 714564
rect 676122 714552 676128 714564
rect 676180 714552 676186 714604
rect 673178 714008 673184 714060
rect 673236 714048 673242 714060
rect 675938 714048 675944 714060
rect 673236 714020 675944 714048
rect 673236 714008 673242 714020
rect 675938 714008 675944 714020
rect 675996 714008 676002 714060
rect 41966 713872 41972 713924
rect 42024 713912 42030 713924
rect 44358 713912 44364 713924
rect 42024 713884 44364 713912
rect 42024 713872 42030 713884
rect 44358 713872 44364 713884
rect 44416 713872 44422 713924
rect 41874 713804 41880 713856
rect 41932 713844 41938 713856
rect 41932 713816 42288 713844
rect 41932 713804 41938 713816
rect 42260 712972 42288 713816
rect 673362 713192 673368 713244
rect 673420 713232 673426 713244
rect 675938 713232 675944 713244
rect 673420 713204 675944 713232
rect 673420 713192 673426 713204
rect 675938 713192 675944 713204
rect 675996 713192 676002 713244
rect 42242 712920 42248 712972
rect 42300 712920 42306 712972
rect 673086 712376 673092 712428
rect 673144 712416 673150 712428
rect 675938 712416 675944 712428
rect 673144 712388 675944 712416
rect 673144 712376 673150 712388
rect 675938 712376 675944 712388
rect 675996 712376 676002 712428
rect 44082 712104 44088 712156
rect 44140 712144 44146 712156
rect 59262 712144 59268 712156
rect 44140 712116 59268 712144
rect 44140 712104 44146 712116
rect 59262 712104 59268 712116
rect 59320 712104 59326 712156
rect 675110 712036 675116 712088
rect 675168 712076 675174 712088
rect 675938 712076 675944 712088
rect 675168 712048 675944 712076
rect 675168 712036 675174 712048
rect 675938 712036 675944 712048
rect 675996 712036 676002 712088
rect 675018 711968 675024 712020
rect 675076 712008 675082 712020
rect 675846 712008 675852 712020
rect 675076 711980 675852 712008
rect 675076 711968 675082 711980
rect 675846 711968 675852 711980
rect 675904 711968 675910 712020
rect 42150 711696 42156 711748
rect 42208 711736 42214 711748
rect 43346 711736 43352 711748
rect 42208 711708 43352 711736
rect 42208 711696 42214 711708
rect 43346 711696 43352 711708
rect 43404 711696 43410 711748
rect 42150 710880 42156 710932
rect 42208 710920 42214 710932
rect 42334 710920 42340 710932
rect 42208 710892 42340 710920
rect 42208 710880 42214 710892
rect 42334 710880 42340 710892
rect 42392 710880 42398 710932
rect 673546 710676 673552 710728
rect 673604 710716 673610 710728
rect 674650 710716 674656 710728
rect 673604 710688 674656 710716
rect 673604 710676 673610 710688
rect 674650 710676 674656 710688
rect 674708 710676 674714 710728
rect 42334 710404 42340 710456
rect 42392 710444 42398 710456
rect 42702 710444 42708 710456
rect 42392 710416 42708 710444
rect 42392 710404 42398 710416
rect 42702 710404 42708 710416
rect 42760 710404 42766 710456
rect 42702 710268 42708 710320
rect 42760 710308 42766 710320
rect 43254 710308 43260 710320
rect 42760 710280 43260 710308
rect 42760 710268 42766 710280
rect 43254 710268 43260 710280
rect 43312 710268 43318 710320
rect 43254 710132 43260 710184
rect 43312 710172 43318 710184
rect 43898 710172 43904 710184
rect 43312 710144 43904 710172
rect 43312 710132 43318 710144
rect 43898 710132 43904 710144
rect 43956 710132 43962 710184
rect 43898 709996 43904 710048
rect 43956 710036 43962 710048
rect 44358 710036 44364 710048
rect 43956 710008 44364 710036
rect 43956 709996 43962 710008
rect 44358 709996 44364 710008
rect 44416 709996 44422 710048
rect 42242 709928 42248 709980
rect 42300 709968 42306 709980
rect 42300 709940 42380 709968
rect 42300 709928 42306 709940
rect 42352 709776 42380 709940
rect 42334 709724 42340 709776
rect 42392 709724 42398 709776
rect 44082 709696 44088 709708
rect 42260 709668 44088 709696
rect 42260 709436 42288 709668
rect 44082 709656 44088 709668
rect 44140 709656 44146 709708
rect 42242 709384 42248 709436
rect 42300 709384 42306 709436
rect 44082 709384 44088 709436
rect 44140 709384 44146 709436
rect 43714 709316 43720 709368
rect 43772 709356 43778 709368
rect 44100 709356 44128 709384
rect 43772 709328 44128 709356
rect 43772 709316 43778 709328
rect 675202 709248 675208 709300
rect 675260 709288 675266 709300
rect 676030 709288 676036 709300
rect 675260 709260 676036 709288
rect 675260 709248 675266 709260
rect 676030 709248 676036 709260
rect 676088 709248 676094 709300
rect 674834 709180 674840 709232
rect 674892 709220 674898 709232
rect 675754 709220 675760 709232
rect 674892 709192 675760 709220
rect 674892 709180 674898 709192
rect 675754 709180 675760 709192
rect 675812 709180 675818 709232
rect 673638 708636 673644 708688
rect 673696 708676 673702 708688
rect 676030 708676 676036 708688
rect 673696 708648 676036 708676
rect 673696 708636 673702 708648
rect 676030 708636 676036 708648
rect 676088 708636 676094 708688
rect 42150 708568 42156 708620
rect 42208 708608 42214 708620
rect 43806 708608 43812 708620
rect 42208 708580 43812 708608
rect 42208 708568 42214 708580
rect 43806 708568 43812 708580
rect 43864 708568 43870 708620
rect 42150 708024 42156 708076
rect 42208 708064 42214 708076
rect 42334 708064 42340 708076
rect 42208 708036 42340 708064
rect 42208 708024 42214 708036
rect 42334 708024 42340 708036
rect 42392 708024 42398 708076
rect 42150 707208 42156 707260
rect 42208 707248 42214 707260
rect 42702 707248 42708 707260
rect 42208 707220 42708 707248
rect 42208 707208 42214 707220
rect 42702 707208 42708 707220
rect 42760 707208 42766 707260
rect 42150 706732 42156 706784
rect 42208 706772 42214 706784
rect 43714 706772 43720 706784
rect 42208 706744 43720 706772
rect 42208 706732 42214 706744
rect 43714 706732 43720 706744
rect 43772 706732 43778 706784
rect 672074 705100 672080 705152
rect 672132 705140 672138 705152
rect 676030 705140 676036 705152
rect 672132 705112 676036 705140
rect 672132 705100 672138 705112
rect 676030 705100 676036 705112
rect 676088 705100 676094 705152
rect 42058 704216 42064 704268
rect 42116 704256 42122 704268
rect 43346 704256 43352 704268
rect 42116 704228 43352 704256
rect 42116 704216 42122 704228
rect 43346 704216 43352 704228
rect 43404 704216 43410 704268
rect 655974 703876 655980 703928
rect 656032 703916 656038 703928
rect 675386 703916 675392 703928
rect 656032 703888 675392 703916
rect 656032 703876 656038 703888
rect 675386 703876 675392 703888
rect 675444 703876 675450 703928
rect 42334 703808 42340 703860
rect 42392 703848 42398 703860
rect 58526 703848 58532 703860
rect 42392 703820 58532 703848
rect 42392 703808 42398 703820
rect 58526 703808 58532 703820
rect 58584 703808 58590 703860
rect 42150 703536 42156 703588
rect 42208 703576 42214 703588
rect 44082 703576 44088 703588
rect 42208 703548 44088 703576
rect 42208 703536 42214 703548
rect 44082 703536 44088 703548
rect 44140 703536 44146 703588
rect 42058 703060 42064 703112
rect 42116 703100 42122 703112
rect 43622 703100 43628 703112
rect 42116 703072 43628 703100
rect 42116 703060 42122 703072
rect 43622 703060 43628 703072
rect 43680 703060 43686 703112
rect 42058 702380 42064 702432
rect 42116 702420 42122 702432
rect 43254 702420 43260 702432
rect 42116 702392 43260 702420
rect 42116 702380 42122 702392
rect 43254 702380 43260 702392
rect 43312 702380 43318 702432
rect 45830 700952 45836 701004
rect 45888 700992 45894 701004
rect 58250 700992 58256 701004
rect 45888 700964 58256 700992
rect 45888 700952 45894 700964
rect 58250 700952 58256 700964
rect 58308 700952 58314 701004
rect 50982 700884 50988 700936
rect 51040 700924 51046 700936
rect 58526 700924 58532 700936
rect 51040 700896 58532 700924
rect 51040 700884 51046 700896
rect 58526 700884 58532 700896
rect 58584 700884 58590 700936
rect 42150 700544 42156 700596
rect 42208 700584 42214 700596
rect 43806 700584 43812 700596
rect 42208 700556 43812 700584
rect 42208 700544 42214 700556
rect 43806 700544 43812 700556
rect 43864 700544 43870 700596
rect 42150 700000 42156 700052
rect 42208 700040 42214 700052
rect 43530 700040 43536 700052
rect 42208 700012 43536 700040
rect 42208 700000 42214 700012
rect 43530 700000 43536 700012
rect 43588 700000 43594 700052
rect 48222 698232 48228 698284
rect 48280 698272 48286 698284
rect 58526 698272 58532 698284
rect 48280 698244 58532 698272
rect 48280 698232 48286 698244
rect 58526 698232 58532 698244
rect 58584 698232 58590 698284
rect 654226 692860 654232 692912
rect 654284 692900 654290 692912
rect 675018 692900 675024 692912
rect 654284 692872 675024 692900
rect 654284 692860 654290 692872
rect 675018 692860 675024 692872
rect 675076 692860 675082 692912
rect 654134 690004 654140 690056
rect 654192 690044 654198 690056
rect 675110 690044 675116 690056
rect 654192 690016 675116 690044
rect 654192 690004 654198 690016
rect 675110 690004 675116 690016
rect 675168 690004 675174 690056
rect 673822 689324 673828 689376
rect 673880 689364 673886 689376
rect 675478 689364 675484 689376
rect 673880 689336 675484 689364
rect 673880 689324 673886 689336
rect 675478 689324 675484 689336
rect 675536 689324 675542 689376
rect 675018 688916 675024 688968
rect 675076 688956 675082 688968
rect 675478 688956 675484 688968
rect 675076 688928 675484 688956
rect 675076 688916 675082 688928
rect 675478 688916 675484 688928
rect 675536 688916 675542 688968
rect 675018 688576 675024 688628
rect 675076 688616 675082 688628
rect 675386 688616 675392 688628
rect 675076 688588 675392 688616
rect 675076 688576 675082 688588
rect 675386 688576 675392 688588
rect 675444 688576 675450 688628
rect 41782 688032 41788 688084
rect 41840 688072 41846 688084
rect 50982 688072 50988 688084
rect 41840 688044 50988 688072
rect 41840 688032 41846 688044
rect 50982 688032 50988 688044
rect 51040 688032 51046 688084
rect 41782 687624 41788 687676
rect 41840 687664 41846 687676
rect 48222 687664 48228 687676
rect 41840 687636 48228 687664
rect 41840 687624 41846 687636
rect 48222 687624 48228 687636
rect 48280 687624 48286 687676
rect 41782 687284 41788 687336
rect 41840 687324 41846 687336
rect 45922 687324 45928 687336
rect 41840 687296 45928 687324
rect 41840 687284 41846 687296
rect 45922 687284 45928 687296
rect 45980 687284 45986 687336
rect 674558 687284 674564 687336
rect 674616 687324 674622 687336
rect 675386 687324 675392 687336
rect 674616 687296 675392 687324
rect 674616 687284 674622 687296
rect 675386 687284 675392 687296
rect 675444 687284 675450 687336
rect 41782 687148 41788 687200
rect 41840 687188 41846 687200
rect 43990 687188 43996 687200
rect 41840 687160 43996 687188
rect 41840 687148 41846 687160
rect 43990 687148 43996 687160
rect 44048 687148 44054 687200
rect 675110 687012 675116 687064
rect 675168 687052 675174 687064
rect 675478 687052 675484 687064
rect 675168 687024 675484 687052
rect 675168 687012 675174 687024
rect 675478 687012 675484 687024
rect 675536 687012 675542 687064
rect 41782 686128 41788 686180
rect 41840 686168 41846 686180
rect 43990 686168 43996 686180
rect 41840 686140 43996 686168
rect 41840 686128 41846 686140
rect 43990 686128 43996 686140
rect 44048 686128 44054 686180
rect 41782 685992 41788 686044
rect 41840 686032 41846 686044
rect 43438 686032 43444 686044
rect 41840 686004 43444 686032
rect 41840 685992 41846 686004
rect 43438 685992 43444 686004
rect 43496 685992 43502 686044
rect 675110 685448 675116 685500
rect 675168 685488 675174 685500
rect 675386 685488 675392 685500
rect 675168 685460 675392 685488
rect 675168 685448 675174 685460
rect 675386 685448 675392 685460
rect 675444 685448 675450 685500
rect 41782 684428 41788 684480
rect 41840 684468 41846 684480
rect 43898 684468 43904 684480
rect 41840 684440 43904 684468
rect 41840 684428 41846 684440
rect 43898 684428 43904 684440
rect 43956 684428 43962 684480
rect 41782 683680 41788 683732
rect 41840 683720 41846 683732
rect 43530 683720 43536 683732
rect 41840 683692 43536 683720
rect 41840 683680 41846 683692
rect 43530 683680 43536 683692
rect 43588 683680 43594 683732
rect 675018 683612 675024 683664
rect 675076 683652 675082 683664
rect 675386 683652 675392 683664
rect 675076 683624 675392 683652
rect 675076 683612 675082 683624
rect 675386 683612 675392 683624
rect 675444 683612 675450 683664
rect 41690 682456 41696 682508
rect 41748 682496 41754 682508
rect 43622 682496 43628 682508
rect 41748 682468 43628 682496
rect 41748 682456 41754 682468
rect 43622 682456 43628 682468
rect 43680 682456 43686 682508
rect 41690 682184 41696 682236
rect 41748 682224 41754 682236
rect 43714 682224 43720 682236
rect 41748 682196 43720 682224
rect 41748 682184 41754 682196
rect 43714 682184 43720 682196
rect 43772 682184 43778 682236
rect 41782 681708 41788 681760
rect 41840 681748 41846 681760
rect 43438 681748 43444 681760
rect 41840 681720 43444 681748
rect 41840 681708 41846 681720
rect 43438 681708 43444 681720
rect 43496 681708 43502 681760
rect 673270 681436 673276 681488
rect 673328 681476 673334 681488
rect 679158 681476 679164 681488
rect 673328 681448 679164 681476
rect 673328 681436 673334 681448
rect 679158 681436 679164 681448
rect 679216 681436 679222 681488
rect 673086 680824 673092 680876
rect 673144 680864 673150 680876
rect 679250 680864 679256 680876
rect 673144 680836 679256 680864
rect 673144 680824 673150 680836
rect 679250 680824 679256 680836
rect 679308 680824 679314 680876
rect 673178 680756 673184 680808
rect 673236 680796 673242 680808
rect 679066 680796 679072 680808
rect 673236 680768 679072 680796
rect 673236 680756 673242 680768
rect 679066 680756 679072 680768
rect 679124 680756 679130 680808
rect 41782 680008 41788 680060
rect 41840 680048 41846 680060
rect 43898 680048 43904 680060
rect 41840 680020 43904 680048
rect 41840 680008 41846 680020
rect 43898 680008 43904 680020
rect 43956 680008 43962 680060
rect 41782 679872 41788 679924
rect 41840 679912 41846 679924
rect 43806 679912 43812 679924
rect 41840 679884 43812 679912
rect 41840 679872 41846 679884
rect 43806 679872 43812 679884
rect 43864 679872 43870 679924
rect 41690 679328 41696 679380
rect 41748 679368 41754 679380
rect 44082 679368 44088 679380
rect 41748 679340 44088 679368
rect 41748 679328 41754 679340
rect 44082 679328 44088 679340
rect 44140 679328 44146 679380
rect 41690 676608 41696 676660
rect 41748 676648 41754 676660
rect 43346 676648 43352 676660
rect 41748 676620 43352 676648
rect 41748 676608 41754 676620
rect 43346 676608 43352 676620
rect 43404 676608 43410 676660
rect 41690 676472 41696 676524
rect 41748 676512 41754 676524
rect 45830 676512 45836 676524
rect 41748 676484 45836 676512
rect 41748 676472 41754 676484
rect 45830 676472 45836 676484
rect 45888 676472 45894 676524
rect 41782 676200 41788 676252
rect 41840 676240 41846 676252
rect 42702 676240 42708 676252
rect 41840 676212 42708 676240
rect 41840 676200 41846 676212
rect 42702 676200 42708 676212
rect 42760 676200 42766 676252
rect 674558 673820 674564 673872
rect 674616 673860 674622 673872
rect 674926 673860 674932 673872
rect 674616 673832 674932 673860
rect 674616 673820 674622 673832
rect 674926 673820 674932 673832
rect 674984 673820 674990 673872
rect 30282 672188 30288 672240
rect 30340 672228 30346 672240
rect 43070 672228 43076 672240
rect 30340 672200 43076 672228
rect 30340 672188 30346 672200
rect 43070 672188 43076 672200
rect 43128 672188 43134 672240
rect 27522 672120 27528 672172
rect 27580 672160 27586 672172
rect 43162 672160 43168 672172
rect 27580 672132 43168 672160
rect 27580 672120 27586 672132
rect 43162 672120 43168 672132
rect 43220 672120 43226 672172
rect 27430 672052 27436 672104
rect 27488 672092 27494 672104
rect 43254 672092 43260 672104
rect 27488 672064 43260 672092
rect 27488 672052 27494 672064
rect 43254 672052 43260 672064
rect 43312 672052 43318 672104
rect 655882 670896 655888 670948
rect 655940 670936 655946 670948
rect 676214 670936 676220 670948
rect 655940 670908 676220 670936
rect 655940 670896 655946 670908
rect 676214 670896 676220 670908
rect 676272 670896 676278 670948
rect 42426 670828 42432 670880
rect 42484 670868 42490 670880
rect 60642 670868 60648 670880
rect 42484 670840 60648 670868
rect 42484 670828 42490 670840
rect 60642 670828 60648 670840
rect 60700 670828 60706 670880
rect 655514 670760 655520 670812
rect 655572 670800 655578 670812
rect 676030 670800 676036 670812
rect 655572 670772 676036 670800
rect 655572 670760 655578 670772
rect 676030 670760 676036 670772
rect 676088 670760 676094 670812
rect 42058 670692 42064 670744
rect 42116 670732 42122 670744
rect 43530 670732 43536 670744
rect 42116 670704 43536 670732
rect 42116 670692 42122 670704
rect 43530 670692 43536 670704
rect 43588 670692 43594 670744
rect 43162 670624 43168 670676
rect 43220 670664 43226 670676
rect 43220 670636 43668 670664
rect 43220 670624 43226 670636
rect 43640 670608 43668 670636
rect 43714 670624 43720 670676
rect 43772 670664 43778 670676
rect 44266 670664 44272 670676
rect 43772 670636 44272 670664
rect 43772 670624 43778 670636
rect 44266 670624 44272 670636
rect 44324 670624 44330 670676
rect 43622 670556 43628 670608
rect 43680 670556 43686 670608
rect 43898 670488 43904 670540
rect 43956 670528 43962 670540
rect 44358 670528 44364 670540
rect 43956 670500 44364 670528
rect 43956 670488 43962 670500
rect 44358 670488 44364 670500
rect 44416 670488 44422 670540
rect 42702 670352 42708 670404
rect 42760 670392 42766 670404
rect 43070 670392 43076 670404
rect 42760 670364 43076 670392
rect 42760 670352 42766 670364
rect 43070 670352 43076 670364
rect 43128 670352 43134 670404
rect 42426 670216 42432 670268
rect 42484 670256 42490 670268
rect 42702 670256 42708 670268
rect 42484 670228 42708 670256
rect 42484 670216 42490 670228
rect 42702 670216 42708 670228
rect 42760 670216 42766 670268
rect 42242 669944 42248 669996
rect 42300 669944 42306 669996
rect 42260 669780 42288 669944
rect 42334 669780 42340 669792
rect 42260 669752 42340 669780
rect 42334 669740 42340 669752
rect 42392 669740 42398 669792
rect 673546 668992 673552 669044
rect 673604 669032 673610 669044
rect 676030 669032 676036 669044
rect 673604 669004 676036 669032
rect 673604 668992 673610 669004
rect 676030 668992 676036 669004
rect 676088 668992 676094 669044
rect 673362 668652 673368 668704
rect 673420 668692 673426 668704
rect 676214 668692 676220 668704
rect 673420 668664 676220 668692
rect 673420 668652 673426 668664
rect 676214 668652 676220 668664
rect 676272 668652 676278 668704
rect 655698 668040 655704 668092
rect 655756 668080 655762 668092
rect 678974 668080 678980 668092
rect 655756 668052 678980 668080
rect 655756 668040 655762 668052
rect 678974 668040 678980 668052
rect 679032 668040 679038 668092
rect 674926 667972 674932 668024
rect 674984 668012 674990 668024
rect 676030 668012 676036 668024
rect 674984 667984 676036 668012
rect 674984 667972 674990 667984
rect 676030 667972 676036 667984
rect 676088 667972 676094 668024
rect 42334 667904 42340 667956
rect 42392 667944 42398 667956
rect 42702 667944 42708 667956
rect 42392 667916 42708 667944
rect 42392 667904 42398 667916
rect 42702 667904 42708 667916
rect 42760 667904 42766 667956
rect 674742 667836 674748 667888
rect 674800 667876 674806 667888
rect 676030 667876 676036 667888
rect 674800 667848 676036 667876
rect 674800 667836 674806 667848
rect 676030 667836 676036 667848
rect 676088 667836 676094 667888
rect 42702 667768 42708 667820
rect 42760 667808 42766 667820
rect 44174 667808 44180 667820
rect 42760 667780 44180 667808
rect 42760 667768 42766 667780
rect 44174 667768 44180 667780
rect 44232 667768 44238 667820
rect 42334 667224 42340 667276
rect 42392 667264 42398 667276
rect 43806 667264 43812 667276
rect 42392 667236 43812 667264
rect 42392 667224 42398 667236
rect 43806 667224 43812 667236
rect 43864 667224 43870 667276
rect 43806 667088 43812 667140
rect 43864 667128 43870 667140
rect 44266 667128 44272 667140
rect 43864 667100 44272 667128
rect 43864 667088 43870 667100
rect 44266 667088 44272 667100
rect 44324 667088 44330 667140
rect 42242 665388 42248 665440
rect 42300 665428 42306 665440
rect 43070 665428 43076 665440
rect 42300 665400 43076 665428
rect 42300 665388 42306 665400
rect 43070 665388 43076 665400
rect 43128 665388 43134 665440
rect 42150 665184 42156 665236
rect 42208 665224 42214 665236
rect 43346 665224 43352 665236
rect 42208 665196 43352 665224
rect 42208 665184 42214 665196
rect 43346 665184 43352 665196
rect 43404 665184 43410 665236
rect 675202 665116 675208 665168
rect 675260 665156 675266 665168
rect 676030 665156 676036 665168
rect 675260 665128 676036 665156
rect 675260 665116 675266 665128
rect 676030 665116 676036 665128
rect 676088 665116 676094 665168
rect 43346 665048 43352 665100
rect 43404 665088 43410 665100
rect 44358 665088 44364 665100
rect 43404 665060 44364 665088
rect 43404 665048 43410 665060
rect 44358 665048 44364 665060
rect 44416 665048 44422 665100
rect 674650 664708 674656 664760
rect 674708 664748 674714 664760
rect 676030 664748 676036 664760
rect 674708 664720 676036 664748
rect 674708 664708 674714 664720
rect 676030 664708 676036 664720
rect 676088 664708 676094 664760
rect 42150 664640 42156 664692
rect 42208 664680 42214 664692
rect 42702 664680 42708 664692
rect 42208 664652 42708 664680
rect 42208 664640 42214 664652
rect 42702 664640 42708 664652
rect 42760 664640 42766 664692
rect 42242 663552 42248 663604
rect 42300 663592 42306 663604
rect 43162 663592 43168 663604
rect 42300 663564 43168 663592
rect 42300 663552 42306 663564
rect 43162 663552 43168 663564
rect 43220 663552 43226 663604
rect 674282 663076 674288 663128
rect 674340 663116 674346 663128
rect 676030 663116 676036 663128
rect 674340 663088 676036 663116
rect 674340 663076 674346 663088
rect 676030 663076 676036 663088
rect 676088 663076 676094 663128
rect 42242 663008 42248 663060
rect 42300 663048 42306 663060
rect 43714 663048 43720 663060
rect 42300 663020 43720 663048
rect 42300 663008 42306 663020
rect 43714 663008 43720 663020
rect 43772 663008 43778 663060
rect 673730 662328 673736 662380
rect 673788 662368 673794 662380
rect 676030 662368 676036 662380
rect 673788 662340 676036 662368
rect 673788 662328 673794 662340
rect 676030 662328 676036 662340
rect 676088 662328 676094 662380
rect 42150 661036 42156 661088
rect 42208 661076 42214 661088
rect 43622 661076 43628 661088
rect 42208 661048 43628 661076
rect 42208 661036 42214 661048
rect 43622 661036 43628 661048
rect 43680 661036 43686 661088
rect 42426 659676 42432 659728
rect 42484 659716 42490 659728
rect 58434 659716 58440 659728
rect 42484 659688 58440 659716
rect 42484 659676 42490 659688
rect 58434 659676 58440 659688
rect 58492 659676 58498 659728
rect 672166 659676 672172 659728
rect 672224 659716 672230 659728
rect 678974 659716 678980 659728
rect 672224 659688 678980 659716
rect 672224 659676 672230 659688
rect 678974 659676 678980 659688
rect 679032 659676 679038 659728
rect 42334 659608 42340 659660
rect 42392 659648 42398 659660
rect 58526 659648 58532 659660
rect 42392 659620 58532 659648
rect 42392 659608 42398 659620
rect 58526 659608 58532 659620
rect 58584 659608 58590 659660
rect 45922 659540 45928 659592
rect 45980 659580 45986 659592
rect 58618 659580 58624 659592
rect 45980 659552 58624 659580
rect 45980 659540 45986 659552
rect 58618 659540 58624 659552
rect 58676 659540 58682 659592
rect 42334 659472 42340 659524
rect 42392 659512 42398 659524
rect 43254 659512 43260 659524
rect 42392 659484 43260 659512
rect 42392 659472 42398 659484
rect 43254 659472 43260 659484
rect 43312 659472 43318 659524
rect 42334 659200 42340 659252
rect 42392 659240 42398 659252
rect 43346 659240 43352 659252
rect 42392 659212 43352 659240
rect 42392 659200 42398 659212
rect 43346 659200 43352 659212
rect 43404 659200 43410 659252
rect 42150 658996 42156 659048
rect 42208 659036 42214 659048
rect 43806 659036 43812 659048
rect 42208 659008 43812 659036
rect 42208 658996 42214 659008
rect 43806 658996 43812 659008
rect 43864 658996 43870 659048
rect 42150 657364 42156 657416
rect 42208 657404 42214 657416
rect 43898 657404 43904 657416
rect 42208 657376 43904 657404
rect 42208 657364 42214 657376
rect 43898 657364 43904 657376
rect 43956 657364 43962 657416
rect 655698 656888 655704 656940
rect 655756 656928 655762 656940
rect 675386 656928 675392 656940
rect 655756 656900 675392 656928
rect 655756 656888 655762 656900
rect 675386 656888 675392 656900
rect 675444 656888 675450 656940
rect 48222 656820 48228 656872
rect 48280 656860 48286 656872
rect 58066 656860 58072 656872
rect 48280 656832 58072 656860
rect 48280 656820 48286 656832
rect 58066 656820 58072 656832
rect 58124 656820 58130 656872
rect 50982 656752 50988 656804
rect 51040 656792 51046 656804
rect 58434 656792 58440 656804
rect 51040 656764 58440 656792
rect 51040 656752 51046 656764
rect 58434 656752 58440 656764
rect 58492 656752 58498 656804
rect 42150 656140 42156 656192
rect 42208 656180 42214 656192
rect 43070 656180 43076 656192
rect 42208 656152 43076 656180
rect 42208 656140 42214 656152
rect 43070 656140 43076 656152
rect 43128 656140 43134 656192
rect 674650 649544 674656 649596
rect 674708 649584 674714 649596
rect 675386 649584 675392 649596
rect 674708 649556 675392 649584
rect 674708 649544 674714 649556
rect 675386 649544 675392 649556
rect 675444 649544 675450 649596
rect 654410 648592 654416 648644
rect 654468 648632 654474 648644
rect 674742 648632 674748 648644
rect 654468 648604 674748 648632
rect 654468 648592 654474 648604
rect 674742 648592 674748 648604
rect 674800 648592 674806 648644
rect 674282 647844 674288 647896
rect 674340 647884 674346 647896
rect 674926 647884 674932 647896
rect 674340 647856 674932 647884
rect 674340 647844 674346 647856
rect 674926 647844 674932 647856
rect 674984 647844 674990 647896
rect 674926 647708 674932 647760
rect 674984 647748 674990 647760
rect 675386 647748 675392 647760
rect 674984 647720 675392 647748
rect 674984 647708 674990 647720
rect 675386 647708 675392 647720
rect 675444 647708 675450 647760
rect 673454 646144 673460 646196
rect 673512 646184 673518 646196
rect 675202 646184 675208 646196
rect 673512 646156 675208 646184
rect 673512 646144 673518 646156
rect 675202 646144 675208 646156
rect 675260 646144 675266 646196
rect 656434 645872 656440 645924
rect 656492 645912 656498 645924
rect 675294 645912 675300 645924
rect 656492 645884 675300 645912
rect 656492 645872 656498 645884
rect 675294 645872 675300 645884
rect 675352 645872 675358 645924
rect 673730 645192 673736 645244
rect 673788 645232 673794 645244
rect 675386 645232 675392 645244
rect 673788 645204 675392 645232
rect 673788 645192 673794 645204
rect 675386 645192 675392 645204
rect 675444 645192 675450 645244
rect 41506 644648 41512 644700
rect 41564 644688 41570 644700
rect 50982 644688 50988 644700
rect 41564 644660 50988 644688
rect 41564 644648 41570 644660
rect 50982 644648 50988 644660
rect 51040 644648 51046 644700
rect 673638 644580 673644 644632
rect 673696 644620 673702 644632
rect 675386 644620 675392 644632
rect 673696 644592 675392 644620
rect 673696 644580 673702 644592
rect 675386 644580 675392 644592
rect 675444 644580 675450 644632
rect 41506 644240 41512 644292
rect 41564 644280 41570 644292
rect 48222 644280 48228 644292
rect 41564 644252 48228 644280
rect 41564 644240 41570 644252
rect 48222 644240 48228 644252
rect 48280 644240 48286 644292
rect 673178 644240 673184 644292
rect 673236 644280 673242 644292
rect 673546 644280 673552 644292
rect 673236 644252 673552 644280
rect 673236 644240 673242 644252
rect 673546 644240 673552 644252
rect 673604 644240 673610 644292
rect 673546 644104 673552 644156
rect 673604 644144 673610 644156
rect 675386 644144 675392 644156
rect 673604 644116 675392 644144
rect 673604 644104 673610 644116
rect 675386 644104 675392 644116
rect 675444 644104 675450 644156
rect 41782 644036 41788 644088
rect 41840 644076 41846 644088
rect 46014 644076 46020 644088
rect 41840 644048 46020 644076
rect 41840 644036 41846 644048
rect 46014 644036 46020 644048
rect 46072 644036 46078 644088
rect 41506 643968 41512 644020
rect 41564 644008 41570 644020
rect 43990 644008 43996 644020
rect 41564 643980 43996 644008
rect 41564 643968 41570 643980
rect 43990 643968 43996 643980
rect 44048 643968 44054 644020
rect 675202 643940 675208 643952
rect 674668 643912 675208 643940
rect 674668 643396 674696 643912
rect 675202 643900 675208 643912
rect 675260 643900 675266 643952
rect 675294 643832 675300 643884
rect 675352 643832 675358 643884
rect 674742 643492 674748 643544
rect 674800 643532 674806 643544
rect 674800 643504 674880 643532
rect 674800 643492 674806 643504
rect 674742 643396 674748 643408
rect 674668 643368 674748 643396
rect 674742 643356 674748 643368
rect 674800 643356 674806 643408
rect 674852 643396 674880 643504
rect 675312 643476 675340 643832
rect 675294 643424 675300 643476
rect 675352 643424 675358 643476
rect 675386 643396 675392 643408
rect 674852 643368 675392 643396
rect 675386 643356 675392 643368
rect 675444 643356 675450 643408
rect 41782 643220 41788 643272
rect 41840 643260 41846 643272
rect 43806 643260 43812 643272
rect 41840 643232 43812 643260
rect 41840 643220 41846 643232
rect 43806 643220 43812 643232
rect 43864 643220 43870 643272
rect 41506 643016 41512 643068
rect 41564 643056 41570 643068
rect 43530 643056 43536 643068
rect 41564 643028 43536 643056
rect 41564 643016 41570 643028
rect 43530 643016 43536 643028
rect 43588 643016 43594 643068
rect 41506 642812 41512 642864
rect 41564 642852 41570 642864
rect 43438 642852 43444 642864
rect 41564 642824 43444 642852
rect 41564 642812 41570 642824
rect 43438 642812 43444 642824
rect 43496 642812 43502 642864
rect 41782 642676 41788 642728
rect 41840 642716 41846 642728
rect 44082 642716 44088 642728
rect 41840 642688 44088 642716
rect 41840 642676 41846 642688
rect 44082 642676 44088 642688
rect 44140 642676 44146 642728
rect 673270 642200 673276 642252
rect 673328 642240 673334 642252
rect 674282 642240 674288 642252
rect 673328 642212 674288 642240
rect 673328 642200 673334 642212
rect 674282 642200 674288 642212
rect 674340 642200 674346 642252
rect 674282 642064 674288 642116
rect 674340 642104 674346 642116
rect 675386 642104 675392 642116
rect 674340 642076 675392 642104
rect 674340 642064 674346 642076
rect 675386 642064 675392 642076
rect 675444 642064 675450 642116
rect 41506 640568 41512 640620
rect 41564 640608 41570 640620
rect 43714 640608 43720 640620
rect 41564 640580 43720 640608
rect 41564 640568 41570 640580
rect 43714 640568 43720 640580
rect 43772 640568 43778 640620
rect 41782 640500 41788 640552
rect 41840 640540 41846 640552
rect 43254 640540 43260 640552
rect 41840 640512 43260 640540
rect 41840 640500 41846 640512
rect 43254 640500 43260 640512
rect 43312 640500 43318 640552
rect 41782 640364 41788 640416
rect 41840 640404 41846 640416
rect 42702 640404 42708 640416
rect 41840 640376 42708 640404
rect 41840 640364 41846 640376
rect 42702 640364 42708 640376
rect 42760 640364 42766 640416
rect 41598 640296 41604 640348
rect 41656 640336 41662 640348
rect 43346 640336 43352 640348
rect 41656 640308 43352 640336
rect 41656 640296 41662 640308
rect 43346 640296 43352 640308
rect 43404 640296 43410 640348
rect 674742 639248 674748 639260
rect 674668 639220 674748 639248
rect 41506 639072 41512 639124
rect 41564 639112 41570 639124
rect 43622 639112 43628 639124
rect 41564 639084 43628 639112
rect 41564 639072 41570 639084
rect 43622 639072 43628 639084
rect 43680 639072 43686 639124
rect 674668 639044 674696 639220
rect 674742 639208 674748 639220
rect 674800 639208 674806 639260
rect 674742 639072 674748 639124
rect 674800 639112 674806 639124
rect 675294 639112 675300 639124
rect 674800 639084 675300 639112
rect 674800 639072 674806 639084
rect 675294 639072 675300 639084
rect 675352 639072 675358 639124
rect 674668 639016 674788 639044
rect 41782 638460 41788 638512
rect 41840 638500 41846 638512
rect 43438 638500 43444 638512
rect 41840 638472 43444 638500
rect 41840 638460 41846 638472
rect 43438 638460 43444 638472
rect 43496 638460 43502 638512
rect 674760 638228 674788 639016
rect 675294 638664 675300 638716
rect 675352 638664 675358 638716
rect 675312 638444 675340 638664
rect 675294 638392 675300 638444
rect 675352 638392 675358 638444
rect 674834 638228 674840 638240
rect 674760 638200 674840 638228
rect 674834 638188 674840 638200
rect 674892 638188 674898 638240
rect 674926 638188 674932 638240
rect 674984 638228 674990 638240
rect 675570 638228 675576 638240
rect 674984 638200 675576 638228
rect 674984 638188 674990 638200
rect 675570 638188 675576 638200
rect 675628 638188 675634 638240
rect 674650 638120 674656 638172
rect 674708 638160 674714 638172
rect 675478 638160 675484 638172
rect 674708 638132 675484 638160
rect 674708 638120 674714 638132
rect 675478 638120 675484 638132
rect 675536 638120 675542 638172
rect 41506 637984 41512 638036
rect 41564 638024 41570 638036
rect 43162 638024 43168 638036
rect 41564 637996 43168 638024
rect 41564 637984 41570 637996
rect 43162 637984 43168 637996
rect 43220 637984 43226 638036
rect 673730 637984 673736 638036
rect 673788 638024 673794 638036
rect 674650 638024 674656 638036
rect 673788 637996 674656 638024
rect 673788 637984 673794 637996
rect 674650 637984 674656 637996
rect 674708 637984 674714 638036
rect 41506 637712 41512 637764
rect 41564 637752 41570 637764
rect 43070 637752 43076 637764
rect 41564 637724 43076 637752
rect 41564 637712 41570 637724
rect 43070 637712 43076 637724
rect 43128 637712 43134 637764
rect 674834 637508 674840 637560
rect 674892 637548 674898 637560
rect 679250 637548 679256 637560
rect 674892 637520 679256 637548
rect 674892 637508 674898 637520
rect 679250 637508 679256 637520
rect 679308 637508 679314 637560
rect 673362 637440 673368 637492
rect 673420 637480 673426 637492
rect 679342 637480 679348 637492
rect 673420 637452 679348 637480
rect 673420 637440 673426 637452
rect 679342 637440 679348 637452
rect 679400 637440 679406 637492
rect 673270 637372 673276 637424
rect 673328 637412 673334 637424
rect 679158 637412 679164 637424
rect 673328 637384 679164 637412
rect 673328 637372 673334 637384
rect 679158 637372 679164 637384
rect 679216 637372 679222 637424
rect 673178 637304 673184 637356
rect 673236 637344 673242 637356
rect 679066 637344 679072 637356
rect 673236 637316 679072 637344
rect 673236 637304 673242 637316
rect 679066 637304 679072 637316
rect 679124 637304 679130 637356
rect 41598 635400 41604 635452
rect 41656 635440 41662 635452
rect 43898 635440 43904 635452
rect 41656 635412 43904 635440
rect 41656 635400 41662 635412
rect 43898 635400 43904 635412
rect 43956 635400 43962 635452
rect 675110 635400 675116 635452
rect 675168 635400 675174 635452
rect 41598 635128 41604 635180
rect 41656 635168 41662 635180
rect 44082 635168 44088 635180
rect 41656 635140 44088 635168
rect 41656 635128 41662 635140
rect 44082 635128 44088 635140
rect 44140 635128 44146 635180
rect 675128 635112 675156 635400
rect 675110 635060 675116 635112
rect 675168 635060 675174 635112
rect 41506 634856 41512 634908
rect 41564 634896 41570 634908
rect 43530 634896 43536 634908
rect 41564 634868 43536 634896
rect 41564 634856 41570 634868
rect 43530 634856 43536 634868
rect 43588 634856 43594 634908
rect 41598 634788 41604 634840
rect 41656 634828 41662 634840
rect 43990 634828 43996 634840
rect 41656 634800 43996 634828
rect 41656 634788 41662 634800
rect 43990 634788 43996 634800
rect 44048 634788 44054 634840
rect 41506 633224 41512 633276
rect 41564 633264 41570 633276
rect 45922 633264 45928 633276
rect 41564 633236 45928 633264
rect 41564 633224 41570 633236
rect 45922 633224 45928 633236
rect 45980 633224 45986 633276
rect 43162 632000 43168 632052
rect 43220 632040 43226 632052
rect 43220 632012 44036 632040
rect 43220 632000 43226 632012
rect 43070 631932 43076 631984
rect 43128 631972 43134 631984
rect 43128 631944 43944 631972
rect 43128 631932 43134 631944
rect 38102 631864 38108 631916
rect 38160 631904 38166 631916
rect 43162 631904 43168 631916
rect 38160 631876 43168 631904
rect 38160 631864 38166 631876
rect 43162 631864 43168 631876
rect 43220 631864 43226 631916
rect 38194 631796 38200 631848
rect 38252 631836 38258 631848
rect 43070 631836 43076 631848
rect 38252 631808 43076 631836
rect 38252 631796 38258 631808
rect 43070 631796 43076 631808
rect 43128 631796 43134 631848
rect 43916 631768 43944 631944
rect 44008 631848 44036 632012
rect 43990 631796 43996 631848
rect 44048 631796 44054 631848
rect 44082 631768 44088 631780
rect 43916 631740 44088 631768
rect 44082 631728 44088 631740
rect 44140 631728 44146 631780
rect 42426 629688 42432 629740
rect 42484 629728 42490 629740
rect 43898 629728 43904 629740
rect 42484 629700 43904 629728
rect 42484 629688 42490 629700
rect 43898 629688 43904 629700
rect 43956 629688 43962 629740
rect 43438 629552 43444 629604
rect 43496 629592 43502 629604
rect 43898 629592 43904 629604
rect 43496 629564 43904 629592
rect 43496 629552 43502 629564
rect 43898 629552 43904 629564
rect 43956 629552 43962 629604
rect 41874 629416 41880 629468
rect 41932 629456 41938 629468
rect 43438 629456 43444 629468
rect 41932 629428 43444 629456
rect 41932 629416 41938 629428
rect 43438 629416 43444 629428
rect 43496 629416 43502 629468
rect 42242 626696 42248 626748
rect 42300 626736 42306 626748
rect 42702 626736 42708 626748
rect 42300 626708 42708 626736
rect 42300 626696 42306 626708
rect 42702 626696 42708 626708
rect 42760 626696 42766 626748
rect 42702 626560 42708 626612
rect 42760 626600 42766 626612
rect 58526 626600 58532 626612
rect 42760 626572 58532 626600
rect 42760 626560 42766 626572
rect 58526 626560 58532 626572
rect 58584 626560 58590 626612
rect 42150 625268 42156 625320
rect 42208 625308 42214 625320
rect 42334 625308 42340 625320
rect 42208 625280 42340 625308
rect 42208 625268 42214 625280
rect 42334 625268 42340 625280
rect 42392 625268 42398 625320
rect 42334 624452 42340 624504
rect 42392 624492 42398 624504
rect 42702 624492 42708 624504
rect 42392 624464 42708 624492
rect 42392 624452 42398 624464
rect 42702 624452 42708 624464
rect 42760 624452 42766 624504
rect 42242 624248 42248 624300
rect 42300 624288 42306 624300
rect 42702 624288 42708 624300
rect 42300 624260 42708 624288
rect 42300 624248 42306 624260
rect 42702 624248 42708 624260
rect 42760 624248 42766 624300
rect 655790 624112 655796 624164
rect 655848 624152 655854 624164
rect 676214 624152 676220 624164
rect 655848 624124 676220 624152
rect 655848 624112 655854 624124
rect 676214 624112 676220 624124
rect 676272 624112 676278 624164
rect 655606 623976 655612 624028
rect 655664 624016 655670 624028
rect 678974 624016 678980 624028
rect 655664 623988 678980 624016
rect 655664 623976 655670 623988
rect 678974 623976 678980 623988
rect 679032 623976 679038 624028
rect 673362 623908 673368 623960
rect 673420 623948 673426 623960
rect 676030 623948 676036 623960
rect 673420 623920 676036 623948
rect 673420 623908 673426 623920
rect 676030 623908 676036 623920
rect 676088 623908 676094 623960
rect 655422 623840 655428 623892
rect 655480 623880 655486 623892
rect 676122 623880 676128 623892
rect 655480 623852 676128 623880
rect 655480 623840 655486 623852
rect 676122 623840 676128 623852
rect 676180 623840 676186 623892
rect 675110 623704 675116 623756
rect 675168 623744 675174 623756
rect 676030 623744 676036 623756
rect 675168 623716 676036 623744
rect 675168 623704 675174 623716
rect 676030 623704 676036 623716
rect 676088 623704 676094 623756
rect 42150 623432 42156 623484
rect 42208 623472 42214 623484
rect 43530 623472 43536 623484
rect 42208 623444 43536 623472
rect 42208 623432 42214 623444
rect 43530 623432 43536 623444
rect 43588 623432 43594 623484
rect 43530 623296 43536 623348
rect 43588 623336 43594 623348
rect 44174 623336 44180 623348
rect 43588 623308 44180 623336
rect 43588 623296 43594 623308
rect 44174 623296 44180 623308
rect 44232 623296 44238 623348
rect 42150 622820 42156 622872
rect 42208 622860 42214 622872
rect 42334 622860 42340 622872
rect 42208 622832 42340 622860
rect 42208 622820 42214 622832
rect 42334 622820 42340 622832
rect 42392 622820 42398 622872
rect 673270 621936 673276 621988
rect 673328 621976 673334 621988
rect 676214 621976 676220 621988
rect 673328 621948 676220 621976
rect 673328 621936 673334 621948
rect 676214 621936 676220 621948
rect 676272 621936 676278 621988
rect 673454 621324 673460 621376
rect 673512 621364 673518 621376
rect 676030 621364 676036 621376
rect 673512 621336 676036 621364
rect 673512 621324 673518 621336
rect 676030 621324 676036 621336
rect 676088 621324 676094 621376
rect 674834 620916 674840 620968
rect 674892 620956 674898 620968
rect 676030 620956 676036 620968
rect 674892 620928 676036 620956
rect 674892 620916 674898 620928
rect 676030 620916 676036 620928
rect 676088 620916 676094 620968
rect 42058 620780 42064 620832
rect 42116 620820 42122 620832
rect 43530 620820 43536 620832
rect 42116 620792 43536 620820
rect 42116 620780 42122 620792
rect 43530 620780 43536 620792
rect 43588 620780 43594 620832
rect 42058 620304 42064 620356
rect 42116 620344 42122 620356
rect 43898 620344 43904 620356
rect 42116 620316 43904 620344
rect 42116 620304 42122 620316
rect 43898 620304 43904 620316
rect 43956 620304 43962 620356
rect 42426 619148 42432 619200
rect 42484 619188 42490 619200
rect 43070 619188 43076 619200
rect 42484 619160 43076 619188
rect 42484 619148 42490 619160
rect 43070 619148 43076 619160
rect 43128 619148 43134 619200
rect 42334 618196 42340 618248
rect 42392 618236 42398 618248
rect 58158 618236 58164 618248
rect 42392 618208 58164 618236
rect 42392 618196 42398 618208
rect 58158 618196 58164 618208
rect 58216 618196 58222 618248
rect 674466 618196 674472 618248
rect 674524 618236 674530 618248
rect 676030 618236 676036 618248
rect 674524 618208 676036 618236
rect 674524 618196 674530 618208
rect 676030 618196 676036 618208
rect 676088 618196 676094 618248
rect 673822 618128 673828 618180
rect 673880 618168 673886 618180
rect 676122 618168 676128 618180
rect 673880 618140 676128 618168
rect 673880 618128 673886 618140
rect 676122 618128 676128 618140
rect 676180 618128 676186 618180
rect 674558 618060 674564 618112
rect 674616 618100 674622 618112
rect 676030 618100 676036 618112
rect 674616 618072 676036 618100
rect 674616 618060 674622 618072
rect 676030 618060 676036 618072
rect 676088 618060 676094 618112
rect 42426 617312 42432 617364
rect 42484 617352 42490 617364
rect 43162 617352 43168 617364
rect 42484 617324 43168 617352
rect 42484 617312 42490 617324
rect 43162 617312 43168 617324
rect 43220 617312 43226 617364
rect 42426 616700 42432 616752
rect 42484 616740 42490 616752
rect 43438 616740 43444 616752
rect 42484 616712 43444 616740
rect 42484 616700 42490 616712
rect 43438 616700 43444 616712
rect 43496 616700 43502 616752
rect 42426 616020 42432 616072
rect 42484 616060 42490 616072
rect 43990 616060 43996 616072
rect 42484 616032 43996 616060
rect 42484 616020 42490 616032
rect 43990 616020 43996 616032
rect 44048 616020 44054 616072
rect 42334 615476 42340 615528
rect 42392 615516 42398 615528
rect 58526 615516 58532 615528
rect 42392 615488 58532 615516
rect 42392 615476 42398 615488
rect 58526 615476 58532 615488
rect 58584 615476 58590 615528
rect 46014 615408 46020 615460
rect 46072 615448 46078 615460
rect 58158 615448 58164 615460
rect 46072 615420 58164 615448
rect 46072 615408 46078 615420
rect 58158 615408 58164 615420
rect 58216 615408 58222 615460
rect 672258 614592 672264 614644
rect 672316 614632 672322 614644
rect 678974 614632 678980 614644
rect 672316 614604 678980 614632
rect 672316 614592 672322 614604
rect 678974 614592 678980 614604
rect 679032 614592 679038 614644
rect 42150 614184 42156 614236
rect 42208 614224 42214 614236
rect 42702 614224 42708 614236
rect 42208 614196 42708 614224
rect 42208 614184 42214 614196
rect 42702 614184 42708 614196
rect 42760 614184 42766 614236
rect 42242 614048 42248 614100
rect 42300 614088 42306 614100
rect 43622 614088 43628 614100
rect 42300 614060 43628 614088
rect 42300 614048 42306 614060
rect 43622 614048 43628 614060
rect 43680 614048 43686 614100
rect 42150 613436 42156 613488
rect 42208 613476 42214 613488
rect 44082 613476 44088 613488
rect 42208 613448 44088 613476
rect 42208 613436 42214 613448
rect 44082 613436 44088 613448
rect 44140 613436 44146 613488
rect 655422 612824 655428 612876
rect 655480 612864 655486 612876
rect 675662 612864 675668 612876
rect 655480 612836 675668 612864
rect 655480 612824 655486 612836
rect 675662 612824 675668 612836
rect 675720 612824 675726 612876
rect 48222 612688 48228 612740
rect 48280 612728 48286 612740
rect 58342 612728 58348 612740
rect 48280 612700 58348 612728
rect 48280 612688 48286 612700
rect 58342 612688 58348 612700
rect 58400 612688 58406 612740
rect 50982 612620 50988 612672
rect 51040 612660 51046 612672
rect 58526 612660 58532 612672
rect 51040 612632 58532 612660
rect 51040 612620 51046 612632
rect 58526 612620 58532 612632
rect 58584 612620 58590 612672
rect 674558 609084 674564 609136
rect 674616 609124 674622 609136
rect 675754 609124 675760 609136
rect 674616 609096 675760 609124
rect 674616 609084 674622 609096
rect 675754 609084 675760 609096
rect 675812 609084 675818 609136
rect 673730 609016 673736 609068
rect 673788 609056 673794 609068
rect 675478 609056 675484 609068
rect 673788 609028 675484 609056
rect 673788 609016 673794 609028
rect 675478 609016 675484 609028
rect 675536 609016 675542 609068
rect 674466 608948 674472 609000
rect 674524 608988 674530 609000
rect 675570 608988 675576 609000
rect 674524 608960 675576 608988
rect 674524 608948 674530 608960
rect 675570 608948 675576 608960
rect 675628 608948 675634 609000
rect 673822 606908 673828 606960
rect 673880 606948 673886 606960
rect 675294 606948 675300 606960
rect 673880 606920 675300 606948
rect 673880 606908 673886 606920
rect 675294 606908 675300 606920
rect 675352 606908 675358 606960
rect 655238 601740 655244 601792
rect 655296 601780 655302 601792
rect 675110 601780 675116 601792
rect 655296 601752 675116 601780
rect 655296 601740 655302 601752
rect 675110 601740 675116 601752
rect 675168 601740 675174 601792
rect 41782 601672 41788 601724
rect 41840 601712 41846 601724
rect 50982 601712 50988 601724
rect 41840 601684 50988 601712
rect 41840 601672 41846 601684
rect 50982 601672 50988 601684
rect 51040 601672 51046 601724
rect 655606 601672 655612 601724
rect 655664 601712 655670 601724
rect 675018 601712 675024 601724
rect 655664 601684 675024 601712
rect 655664 601672 655670 601684
rect 675018 601672 675024 601684
rect 675076 601672 675082 601724
rect 41782 601264 41788 601316
rect 41840 601304 41846 601316
rect 48222 601304 48228 601316
rect 41840 601276 48228 601304
rect 41840 601264 41846 601276
rect 48222 601264 48228 601276
rect 48280 601264 48286 601316
rect 41506 600992 41512 601044
rect 41564 601032 41570 601044
rect 43806 601032 43812 601044
rect 41564 601004 43812 601032
rect 41564 600992 41570 601004
rect 43806 600992 43812 601004
rect 43864 600992 43870 601044
rect 41782 600856 41788 600908
rect 41840 600896 41846 600908
rect 46106 600896 46112 600908
rect 41840 600868 46112 600896
rect 41840 600856 41846 600868
rect 46106 600856 46112 600868
rect 46164 600856 46170 600908
rect 41506 600312 41512 600364
rect 41564 600352 41570 600364
rect 43346 600352 43352 600364
rect 41564 600324 43352 600352
rect 41564 600312 41570 600324
rect 43346 600312 43352 600324
rect 43404 600312 43410 600364
rect 673546 599768 673552 599820
rect 673604 599808 673610 599820
rect 675478 599808 675484 599820
rect 673604 599780 675484 599808
rect 673604 599768 673610 599780
rect 675478 599768 675484 599780
rect 675536 599768 675542 599820
rect 41782 599020 41788 599072
rect 41840 599060 41846 599072
rect 43990 599060 43996 599072
rect 41840 599032 43996 599060
rect 41840 599020 41846 599032
rect 43990 599020 43996 599032
rect 44048 599020 44054 599072
rect 41506 598952 41512 599004
rect 41564 598992 41570 599004
rect 43346 598992 43352 599004
rect 41564 598964 43352 598992
rect 41564 598952 41570 598964
rect 43346 598952 43352 598964
rect 43404 598952 43410 599004
rect 41782 598884 41788 598936
rect 41840 598924 41846 598936
rect 43254 598924 43260 598936
rect 41840 598896 43260 598924
rect 41840 598884 41846 598896
rect 43254 598884 43260 598896
rect 43312 598884 43318 598936
rect 675110 598680 675116 598732
rect 675168 598720 675174 598732
rect 675386 598720 675392 598732
rect 675168 598692 675392 598720
rect 675168 598680 675174 598692
rect 675386 598680 675392 598692
rect 675444 598680 675450 598732
rect 673454 598544 673460 598596
rect 673512 598584 673518 598596
rect 675478 598584 675484 598596
rect 673512 598556 675484 598584
rect 673512 598544 673518 598556
rect 675478 598544 675484 598556
rect 675536 598544 675542 598596
rect 41506 598476 41512 598528
rect 41564 598516 41570 598528
rect 43714 598516 43720 598528
rect 41564 598488 43720 598516
rect 41564 598476 41570 598488
rect 43714 598476 43720 598488
rect 43772 598476 43778 598528
rect 674558 598476 674564 598528
rect 674616 598516 674622 598528
rect 675110 598516 675116 598528
rect 674616 598488 675116 598516
rect 674616 598476 674622 598488
rect 675110 598476 675116 598488
rect 675168 598476 675174 598528
rect 674558 598340 674564 598392
rect 674616 598380 674622 598392
rect 675294 598380 675300 598392
rect 674616 598352 675300 598380
rect 674616 598340 674622 598352
rect 675294 598340 675300 598352
rect 675352 598340 675358 598392
rect 675018 598068 675024 598120
rect 675076 598108 675082 598120
rect 675294 598108 675300 598120
rect 675076 598080 675300 598108
rect 675076 598068 675082 598080
rect 675294 598068 675300 598080
rect 675352 598068 675358 598120
rect 673178 597252 673184 597304
rect 673236 597292 673242 597304
rect 673822 597292 673828 597304
rect 673236 597264 673828 597292
rect 673236 597252 673242 597264
rect 673822 597252 673828 597264
rect 673880 597252 673886 597304
rect 673822 597116 673828 597168
rect 673880 597156 673886 597168
rect 675386 597156 675392 597168
rect 673880 597128 675392 597156
rect 673880 597116 673886 597128
rect 675386 597116 675392 597128
rect 675444 597116 675450 597168
rect 41506 597048 41512 597100
rect 41564 597088 41570 597100
rect 44082 597088 44088 597100
rect 41564 597060 44088 597088
rect 41564 597048 41570 597060
rect 44082 597048 44088 597060
rect 44140 597048 44146 597100
rect 675110 597048 675116 597100
rect 675168 597088 675174 597100
rect 675168 597060 675248 597088
rect 675168 597048 675174 597060
rect 675220 596896 675248 597060
rect 675202 596844 675208 596896
rect 675260 596844 675266 596896
rect 41506 596640 41512 596692
rect 41564 596680 41570 596692
rect 43806 596680 43812 596692
rect 41564 596652 43812 596680
rect 41564 596640 41570 596652
rect 43806 596640 43812 596652
rect 43864 596640 43870 596692
rect 41506 596368 41512 596420
rect 41564 596408 41570 596420
rect 43622 596408 43628 596420
rect 41564 596380 43628 596408
rect 41564 596368 41570 596380
rect 43622 596368 43628 596380
rect 43680 596368 43686 596420
rect 674466 596300 674472 596352
rect 674524 596340 674530 596352
rect 675294 596340 675300 596352
rect 674524 596312 675300 596340
rect 674524 596300 674530 596312
rect 675294 596300 675300 596312
rect 675352 596300 675358 596352
rect 41506 595416 41512 595468
rect 41564 595456 41570 595468
rect 43438 595456 43444 595468
rect 41564 595428 43444 595456
rect 41564 595416 41570 595428
rect 43438 595416 43444 595428
rect 43496 595416 43502 595468
rect 674466 595280 674472 595332
rect 674524 595320 674530 595332
rect 675386 595320 675392 595332
rect 674524 595292 675392 595320
rect 674524 595280 674530 595292
rect 675386 595280 675392 595292
rect 675444 595280 675450 595332
rect 41506 594600 41512 594652
rect 41564 594640 41570 594652
rect 43530 594640 43536 594652
rect 41564 594612 43536 594640
rect 41564 594600 41570 594612
rect 43530 594600 43536 594612
rect 43588 594600 43594 594652
rect 41506 594056 41512 594108
rect 41564 594096 41570 594108
rect 43162 594096 43168 594108
rect 41564 594068 43168 594096
rect 41564 594056 41570 594068
rect 43162 594056 43168 594068
rect 43220 594056 43226 594108
rect 41782 593512 41788 593564
rect 41840 593552 41846 593564
rect 43070 593552 43076 593564
rect 41840 593524 43076 593552
rect 41840 593512 41846 593524
rect 43070 593512 43076 593524
rect 43128 593512 43134 593564
rect 673546 593512 673552 593564
rect 673604 593552 673610 593564
rect 673604 593524 673776 593552
rect 673604 593512 673610 593524
rect 673748 593496 673776 593524
rect 673730 593444 673736 593496
rect 673788 593444 673794 593496
rect 673178 593376 673184 593428
rect 673236 593416 673242 593428
rect 673546 593416 673552 593428
rect 673236 593388 673552 593416
rect 673236 593376 673242 593388
rect 673546 593376 673552 593388
rect 673604 593376 673610 593428
rect 675662 593376 675668 593428
rect 675720 593376 675726 593428
rect 675202 593172 675208 593224
rect 675260 593212 675266 593224
rect 675680 593212 675708 593376
rect 675260 593184 675708 593212
rect 675260 593172 675266 593184
rect 41506 592152 41512 592204
rect 41564 592192 41570 592204
rect 43714 592192 43720 592204
rect 41564 592164 43720 592192
rect 41564 592152 41570 592164
rect 43714 592152 43720 592164
rect 43772 592152 43778 592204
rect 42334 591880 42340 591932
rect 42392 591920 42398 591932
rect 43530 591920 43536 591932
rect 42392 591892 43536 591920
rect 42392 591880 42398 591892
rect 43530 591880 43536 591892
rect 43588 591880 43594 591932
rect 41506 591744 41512 591796
rect 41564 591784 41570 591796
rect 43530 591784 43536 591796
rect 41564 591756 43536 591784
rect 41564 591744 41570 591756
rect 43530 591744 43536 591756
rect 43588 591744 43594 591796
rect 41506 591200 41512 591252
rect 41564 591240 41570 591252
rect 43254 591240 43260 591252
rect 41564 591212 43260 591240
rect 41564 591200 41570 591212
rect 43254 591200 43260 591212
rect 43312 591200 43318 591252
rect 41506 589976 41512 590028
rect 41564 590016 41570 590028
rect 46014 590016 46020 590028
rect 41564 589988 46020 590016
rect 41564 589976 41570 589988
rect 46014 589976 46020 589988
rect 46072 589976 46078 590028
rect 42150 588480 42156 588532
rect 42208 588520 42214 588532
rect 43898 588520 43904 588532
rect 42208 588492 43904 588520
rect 42208 588480 42214 588492
rect 43898 588480 43904 588492
rect 43956 588480 43962 588532
rect 673270 587936 673276 587988
rect 673328 587976 673334 587988
rect 679066 587976 679072 587988
rect 673328 587948 679072 587976
rect 673328 587936 673334 587948
rect 679066 587936 679072 587948
rect 679124 587936 679130 587988
rect 673362 587868 673368 587920
rect 673420 587908 673426 587920
rect 678974 587908 678980 587920
rect 673420 587880 678980 587908
rect 673420 587868 673426 587880
rect 678974 587868 678980 587880
rect 679032 587868 679038 587920
rect 38010 587800 38016 587852
rect 38068 587840 38074 587852
rect 42702 587840 42708 587852
rect 38068 587812 42708 587840
rect 38068 587800 38074 587812
rect 42702 587800 42708 587812
rect 42760 587800 42766 587852
rect 38102 587732 38108 587784
rect 38160 587772 38166 587784
rect 41414 587772 41420 587784
rect 38160 587744 41420 587772
rect 38160 587732 38166 587744
rect 41414 587732 41420 587744
rect 41472 587732 41478 587784
rect 41414 585216 41420 585268
rect 41472 585256 41478 585268
rect 44174 585256 44180 585268
rect 41472 585228 44180 585256
rect 41472 585216 41478 585228
rect 44174 585216 44180 585228
rect 44232 585216 44238 585268
rect 42334 585148 42340 585200
rect 42392 585188 42398 585200
rect 58526 585188 58532 585200
rect 42392 585160 58532 585188
rect 42392 585148 42398 585160
rect 58526 585148 58532 585160
rect 58584 585148 58590 585200
rect 42426 584196 42432 584248
rect 42484 584236 42490 584248
rect 42484 584208 42656 584236
rect 42484 584196 42490 584208
rect 42628 583692 42656 584208
rect 43898 583856 43904 583908
rect 43956 583896 43962 583908
rect 43956 583868 44128 583896
rect 43956 583856 43962 583868
rect 42702 583720 42708 583772
rect 42760 583760 42766 583772
rect 43162 583760 43168 583772
rect 42760 583732 43168 583760
rect 42760 583720 42766 583732
rect 43162 583720 43168 583732
rect 43220 583720 43226 583772
rect 44100 583704 44128 583868
rect 674466 583856 674472 583908
rect 674524 583896 674530 583908
rect 674524 583868 675432 583896
rect 674524 583856 674530 583868
rect 673454 583720 673460 583772
rect 673512 583760 673518 583772
rect 674466 583760 674472 583772
rect 673512 583732 674472 583760
rect 673512 583720 673518 583732
rect 674466 583720 674472 583732
rect 674524 583720 674530 583772
rect 675404 583704 675432 583868
rect 42628 583664 43208 583692
rect 43180 583636 43208 583664
rect 44082 583652 44088 583704
rect 44140 583652 44146 583704
rect 675386 583652 675392 583704
rect 675444 583652 675450 583704
rect 43162 583584 43168 583636
rect 43220 583584 43226 583636
rect 42242 582564 42248 582616
rect 42300 582604 42306 582616
rect 59262 582604 59268 582616
rect 42300 582576 59268 582604
rect 42300 582564 42306 582576
rect 59262 582564 59268 582576
rect 59320 582564 59326 582616
rect 673546 582292 673552 582344
rect 673604 582332 673610 582344
rect 676030 582332 676036 582344
rect 673604 582304 676036 582332
rect 673604 582292 673610 582304
rect 676030 582292 676036 582304
rect 676088 582292 676094 582344
rect 42150 582088 42156 582140
rect 42208 582128 42214 582140
rect 43622 582128 43628 582140
rect 42208 582100 43628 582128
rect 42208 582088 42214 582100
rect 43622 582088 43628 582100
rect 43680 582088 43686 582140
rect 43162 581952 43168 582004
rect 43220 581992 43226 582004
rect 43622 581992 43628 582004
rect 43220 581964 43628 581992
rect 43220 581952 43226 581964
rect 43622 581952 43628 581964
rect 43680 581952 43686 582004
rect 42242 581272 42248 581324
rect 42300 581272 42306 581324
rect 42260 581120 42288 581272
rect 42242 581068 42248 581120
rect 42300 581068 42306 581120
rect 42150 580252 42156 580304
rect 42208 580292 42214 580304
rect 43070 580292 43076 580304
rect 42208 580264 43076 580292
rect 42208 580252 42214 580264
rect 43070 580252 43076 580264
rect 43128 580252 43134 580304
rect 43070 580116 43076 580168
rect 43128 580156 43134 580168
rect 43806 580156 43812 580168
rect 43128 580128 43812 580156
rect 43128 580116 43134 580128
rect 43806 580116 43812 580128
rect 43864 580116 43870 580168
rect 656066 580048 656072 580100
rect 656124 580088 656130 580100
rect 676214 580088 676220 580100
rect 656124 580060 676220 580088
rect 656124 580048 656130 580060
rect 676214 580048 676220 580060
rect 676272 580048 676278 580100
rect 655882 579912 655888 579964
rect 655940 579952 655946 579964
rect 676122 579952 676128 579964
rect 655940 579924 676128 579952
rect 655940 579912 655946 579924
rect 676122 579912 676128 579924
rect 676180 579912 676186 579964
rect 655514 579776 655520 579828
rect 655572 579816 655578 579828
rect 676306 579816 676312 579828
rect 655572 579788 676312 579816
rect 655572 579776 655578 579788
rect 676306 579776 676312 579788
rect 676364 579776 676370 579828
rect 42242 578960 42248 579012
rect 42300 579000 42306 579012
rect 43530 579000 43536 579012
rect 42300 578972 43536 579000
rect 42300 578960 42306 578972
rect 43530 578960 43536 578972
rect 43588 578960 43594 579012
rect 43530 578824 43536 578876
rect 43588 578864 43594 578876
rect 44082 578864 44088 578876
rect 43588 578836 44088 578864
rect 43588 578824 43594 578836
rect 44082 578824 44088 578836
rect 44140 578824 44146 578876
rect 42150 578756 42156 578808
rect 42208 578796 42214 578808
rect 43254 578796 43260 578808
rect 42208 578768 43260 578796
rect 42208 578756 42214 578768
rect 43254 578756 43260 578768
rect 43312 578756 43318 578808
rect 42150 578416 42156 578468
rect 42208 578456 42214 578468
rect 43714 578456 43720 578468
rect 42208 578428 43720 578456
rect 42208 578416 42214 578428
rect 43714 578416 43720 578428
rect 43772 578416 43778 578468
rect 674834 576920 674840 576972
rect 674892 576960 674898 576972
rect 676030 576960 676036 576972
rect 674892 576932 676036 576960
rect 674892 576920 674898 576932
rect 676030 576920 676036 576932
rect 676088 576920 676094 576972
rect 675110 576784 675116 576836
rect 675168 576824 675174 576836
rect 676030 576824 676036 576836
rect 675168 576796 676036 576824
rect 675168 576784 675174 576796
rect 676030 576784 676036 576796
rect 676088 576784 676094 576836
rect 674742 576716 674748 576768
rect 674800 576756 674806 576768
rect 675938 576756 675944 576768
rect 674800 576728 675944 576756
rect 674800 576716 674806 576728
rect 675938 576716 675944 576728
rect 675996 576716 676002 576768
rect 673822 576648 673828 576700
rect 673880 576688 673886 576700
rect 675110 576688 675116 576700
rect 673880 576660 675116 576688
rect 673880 576648 673886 576660
rect 675110 576648 675116 576660
rect 675168 576648 675174 576700
rect 674650 575220 674656 575272
rect 674708 575260 674714 575272
rect 676030 575260 676036 575272
rect 674708 575232 676036 575260
rect 674708 575220 674714 575232
rect 676030 575220 676036 575232
rect 676088 575220 676094 575272
rect 674926 574812 674932 574864
rect 674984 574852 674990 574864
rect 676030 574852 676036 574864
rect 674984 574824 676036 574852
rect 674984 574812 674990 574824
rect 676030 574812 676036 574824
rect 676088 574812 676094 574864
rect 42334 574132 42340 574184
rect 42392 574172 42398 574184
rect 43162 574172 43168 574184
rect 42392 574144 43168 574172
rect 42392 574132 42398 574144
rect 43162 574132 43168 574144
rect 43220 574132 43226 574184
rect 42426 574064 42432 574116
rect 42484 574104 42490 574116
rect 60642 574104 60648 574116
rect 42484 574076 60648 574104
rect 42484 574064 42490 574076
rect 60642 574064 60648 574076
rect 60700 574064 60706 574116
rect 42150 573792 42156 573844
rect 42208 573832 42214 573844
rect 44082 573832 44088 573844
rect 42208 573804 44088 573832
rect 42208 573792 42214 573804
rect 44082 573792 44088 573804
rect 44140 573792 44146 573844
rect 674282 573588 674288 573640
rect 674340 573628 674346 573640
rect 676030 573628 676036 573640
rect 674340 573600 676036 573628
rect 674340 573588 674346 573600
rect 676030 573588 676036 573600
rect 676088 573588 676094 573640
rect 673638 572772 673644 572824
rect 673696 572812 673702 572824
rect 676030 572812 676036 572824
rect 673696 572784 676036 572812
rect 673696 572772 673702 572784
rect 676030 572772 676036 572784
rect 676088 572772 676094 572824
rect 42058 572636 42064 572688
rect 42116 572676 42122 572688
rect 43438 572676 43444 572688
rect 42116 572648 43444 572676
rect 42116 572636 42122 572648
rect 43438 572636 43444 572648
rect 43496 572636 43502 572688
rect 42242 571956 42248 572008
rect 42300 571996 42306 572008
rect 42702 571996 42708 572008
rect 42300 571968 42708 571996
rect 42300 571956 42306 571968
rect 42702 571956 42708 571968
rect 42760 571956 42766 572008
rect 46106 571276 46112 571328
rect 46164 571316 46170 571328
rect 58066 571316 58072 571328
rect 46164 571288 58072 571316
rect 46164 571276 46170 571288
rect 58066 571276 58072 571288
rect 58124 571276 58130 571328
rect 50982 571208 50988 571260
rect 51040 571248 51046 571260
rect 58342 571248 58348 571260
rect 51040 571220 58348 571248
rect 51040 571208 51046 571220
rect 58342 571208 58348 571220
rect 58400 571208 58406 571260
rect 42058 570936 42064 570988
rect 42116 570976 42122 570988
rect 43070 570976 43076 570988
rect 42116 570948 43076 570976
rect 42116 570936 42122 570948
rect 43070 570936 43076 570948
rect 43128 570936 43134 570988
rect 42058 569576 42064 569628
rect 42116 569616 42122 569628
rect 43530 569616 43536 569628
rect 42116 569588 43536 569616
rect 42116 569576 42122 569588
rect 43530 569576 43536 569588
rect 43588 569576 43594 569628
rect 674282 568760 674288 568812
rect 674340 568800 674346 568812
rect 675386 568800 675392 568812
rect 674340 568772 675392 568800
rect 674340 568760 674346 568772
rect 675386 568760 675392 568772
rect 675444 568760 675450 568812
rect 655882 568624 655888 568676
rect 655940 568664 655946 568676
rect 675386 568664 675392 568676
rect 655940 568636 675392 568664
rect 655940 568624 655946 568636
rect 675386 568624 675392 568636
rect 675444 568624 675450 568676
rect 672350 568556 672356 568608
rect 672408 568596 672414 568608
rect 678974 568596 678980 568608
rect 672408 568568 678980 568596
rect 672408 568556 672414 568568
rect 678974 568556 678980 568568
rect 679032 568556 679038 568608
rect 48222 568488 48228 568540
rect 48280 568528 48286 568540
rect 58250 568528 58256 568540
rect 48280 568500 58256 568528
rect 48280 568488 48286 568500
rect 58250 568488 58256 568500
rect 58308 568488 58314 568540
rect 673638 559512 673644 559564
rect 673696 559552 673702 559564
rect 675478 559552 675484 559564
rect 673696 559524 675484 559552
rect 673696 559512 673702 559524
rect 675478 559512 675484 559524
rect 675536 559512 675542 559564
rect 41506 558288 41512 558340
rect 41564 558328 41570 558340
rect 50982 558328 50988 558340
rect 41564 558300 50988 558328
rect 41564 558288 41570 558300
rect 50982 558288 50988 558300
rect 51040 558288 51046 558340
rect 673454 558220 673460 558272
rect 673512 558260 673518 558272
rect 675386 558260 675392 558272
rect 673512 558232 675392 558260
rect 673512 558220 673518 558232
rect 675386 558220 675392 558232
rect 675444 558220 675450 558272
rect 41506 557880 41512 557932
rect 41564 557920 41570 557932
rect 48314 557920 48320 557932
rect 41564 557892 48320 557920
rect 41564 557880 41570 557892
rect 48314 557880 48320 557892
rect 48372 557880 48378 557932
rect 41506 557540 41512 557592
rect 41564 557580 41570 557592
rect 46106 557580 46112 557592
rect 41564 557552 46112 557580
rect 41564 557540 41570 557552
rect 46106 557540 46112 557552
rect 46164 557540 46170 557592
rect 654226 557540 654232 557592
rect 654284 557580 654290 557592
rect 674742 557580 674748 557592
rect 654284 557552 674748 557580
rect 654284 557540 654290 557552
rect 674742 557540 674748 557552
rect 674800 557540 674806 557592
rect 673546 557472 673552 557524
rect 673604 557512 673610 557524
rect 675386 557512 675392 557524
rect 673604 557484 675392 557512
rect 673604 557472 673610 557484
rect 675386 557472 675392 557484
rect 675444 557472 675450 557524
rect 41782 557268 41788 557320
rect 41840 557308 41846 557320
rect 43990 557308 43996 557320
rect 41840 557280 43996 557308
rect 41840 557268 41846 557280
rect 43990 557268 43996 557280
rect 44048 557268 44054 557320
rect 41782 556792 41788 556844
rect 41840 556832 41846 556844
rect 43346 556832 43352 556844
rect 41840 556804 43352 556832
rect 41840 556792 41846 556804
rect 43346 556792 43352 556804
rect 43404 556792 43410 556844
rect 41506 556656 41512 556708
rect 41564 556696 41570 556708
rect 43622 556696 43628 556708
rect 41564 556668 43628 556696
rect 41564 556656 41570 556668
rect 43622 556656 43628 556668
rect 43680 556656 43686 556708
rect 674650 555024 674656 555076
rect 674708 555064 674714 555076
rect 675386 555064 675392 555076
rect 674708 555036 675392 555064
rect 674708 555024 674714 555036
rect 675386 555024 675392 555036
rect 675444 555024 675450 555076
rect 673822 554888 673828 554940
rect 673880 554928 673886 554940
rect 675294 554928 675300 554940
rect 673880 554900 675300 554928
rect 673880 554888 673886 554900
rect 675294 554888 675300 554900
rect 675352 554888 675358 554940
rect 38562 554752 38568 554804
rect 38620 554792 38626 554804
rect 43898 554792 43904 554804
rect 38620 554764 43904 554792
rect 38620 554752 38626 554764
rect 43898 554752 43904 554764
rect 43956 554752 43962 554804
rect 654134 554752 654140 554804
rect 654192 554792 654198 554804
rect 675294 554792 675300 554804
rect 654192 554764 675300 554792
rect 654192 554752 654198 554764
rect 675294 554752 675300 554764
rect 675352 554752 675358 554804
rect 674282 553732 674288 553784
rect 674340 553772 674346 553784
rect 675386 553772 675392 553784
rect 674340 553744 675392 553772
rect 674340 553732 674346 553744
rect 675386 553732 675392 553744
rect 675444 553732 675450 553784
rect 673362 553528 673368 553580
rect 673420 553568 673426 553580
rect 673638 553568 673644 553580
rect 673420 553540 673644 553568
rect 673420 553528 673426 553540
rect 673638 553528 673644 553540
rect 673696 553528 673702 553580
rect 674742 553460 674748 553512
rect 674800 553500 674806 553512
rect 675386 553500 675392 553512
rect 674800 553472 675392 553500
rect 674800 553460 674806 553472
rect 675386 553460 675392 553472
rect 675444 553460 675450 553512
rect 673638 553392 673644 553444
rect 673696 553432 673702 553444
rect 675478 553432 675484 553444
rect 673696 553404 675484 553432
rect 673696 553392 673702 553404
rect 675478 553392 675484 553404
rect 675536 553392 675542 553444
rect 41506 552304 41512 552356
rect 41564 552344 41570 552356
rect 43254 552344 43260 552356
rect 41564 552316 43260 552344
rect 41564 552304 41570 552316
rect 43254 552304 43260 552316
rect 43312 552304 43318 552356
rect 674742 551896 674748 551948
rect 674800 551936 674806 551948
rect 675386 551936 675392 551948
rect 674800 551908 675392 551936
rect 674800 551896 674806 551908
rect 675386 551896 675392 551908
rect 675444 551896 675450 551948
rect 41414 549720 41420 549772
rect 41472 549760 41478 549772
rect 43346 549760 43352 549772
rect 41472 549732 43352 549760
rect 41472 549720 41478 549732
rect 43346 549720 43352 549732
rect 43404 549720 43410 549772
rect 41506 549584 41512 549636
rect 41564 549624 41570 549636
rect 43070 549624 43076 549636
rect 41564 549596 43076 549624
rect 41564 549584 41570 549596
rect 43070 549584 43076 549596
rect 43128 549584 43134 549636
rect 41506 549312 41512 549364
rect 41564 549352 41570 549364
rect 43438 549352 43444 549364
rect 41564 549324 43444 549352
rect 41564 549312 41570 549324
rect 43438 549312 43444 549324
rect 43496 549312 43502 549364
rect 41506 548632 41512 548684
rect 41564 548672 41570 548684
rect 43898 548672 43904 548684
rect 41564 548644 43904 548672
rect 41564 548632 41570 548644
rect 43898 548632 43904 548644
rect 43956 548632 43962 548684
rect 675662 548224 675668 548276
rect 675720 548224 675726 548276
rect 674650 547952 674656 548004
rect 674708 547992 674714 548004
rect 674834 547992 674840 548004
rect 674708 547964 674840 547992
rect 674708 547952 674714 547964
rect 674834 547952 674840 547964
rect 674892 547952 674898 548004
rect 675294 547884 675300 547936
rect 675352 547924 675358 547936
rect 675680 547924 675708 548224
rect 675352 547896 675708 547924
rect 675352 547884 675358 547896
rect 674282 547816 674288 547868
rect 674340 547856 674346 547868
rect 674650 547856 674656 547868
rect 674340 547828 674656 547856
rect 674340 547816 674346 547828
rect 674650 547816 674656 547828
rect 674708 547816 674714 547868
rect 673730 547680 673736 547732
rect 673788 547680 673794 547732
rect 673822 547680 673828 547732
rect 673880 547720 673886 547732
rect 674282 547720 674288 547732
rect 673880 547692 674288 547720
rect 673880 547680 673886 547692
rect 674282 547680 674288 547692
rect 674340 547680 674346 547732
rect 673748 547528 673776 547680
rect 673730 547476 673736 547528
rect 673788 547476 673794 547528
rect 41506 547000 41512 547052
rect 41564 547040 41570 547052
rect 43162 547040 43168 547052
rect 41564 547012 43168 547040
rect 41564 547000 41570 547012
rect 43162 547000 43168 547012
rect 43220 547000 43226 547052
rect 41506 546864 41512 546916
rect 41564 546904 41570 546916
rect 48222 546904 48228 546916
rect 41564 546876 48228 546904
rect 41564 546864 41570 546876
rect 48222 546864 48228 546876
rect 48280 546864 48286 546916
rect 674926 543736 674932 543788
rect 674984 543776 674990 543788
rect 679342 543776 679348 543788
rect 674984 543748 679348 543776
rect 674984 543736 674990 543748
rect 679342 543736 679348 543748
rect 679400 543736 679406 543788
rect 43162 541288 43168 541340
rect 43220 541328 43226 541340
rect 43346 541328 43352 541340
rect 43220 541300 43352 541328
rect 43220 541288 43226 541300
rect 43346 541288 43352 541300
rect 43404 541288 43410 541340
rect 43070 541016 43076 541068
rect 43128 541056 43134 541068
rect 59262 541056 59268 541068
rect 43128 541028 59268 541056
rect 43128 541016 43134 541028
rect 59262 541016 59268 541028
rect 59320 541016 59326 541068
rect 42702 540948 42708 541000
rect 42760 540988 42766 541000
rect 59446 540988 59452 541000
rect 42760 540960 59452 540988
rect 42760 540948 42766 540960
rect 59446 540948 59452 540960
rect 59504 540948 59510 541000
rect 674282 539452 674288 539504
rect 674340 539492 674346 539504
rect 675570 539492 675576 539504
rect 674340 539464 675576 539492
rect 674340 539452 674346 539464
rect 675570 539452 675576 539464
rect 675628 539452 675634 539504
rect 42058 538908 42064 538960
rect 42116 538948 42122 538960
rect 43254 538948 43260 538960
rect 42116 538920 43260 538948
rect 42116 538908 42122 538920
rect 43254 538908 43260 538920
rect 43312 538908 43318 538960
rect 42242 538432 42248 538484
rect 42300 538472 42306 538484
rect 43070 538472 43076 538484
rect 42300 538444 43076 538472
rect 42300 538432 42306 538444
rect 43070 538432 43076 538444
rect 43128 538432 43134 538484
rect 42150 538228 42156 538280
rect 42208 538268 42214 538280
rect 42702 538268 42708 538280
rect 42208 538240 42708 538268
rect 42208 538228 42214 538240
rect 42702 538228 42708 538240
rect 42760 538228 42766 538280
rect 42058 537072 42064 537124
rect 42116 537112 42122 537124
rect 43162 537112 43168 537124
rect 42116 537084 43168 537112
rect 42116 537072 42122 537084
rect 43162 537072 43168 537084
rect 43220 537072 43226 537124
rect 673454 537072 673460 537124
rect 673512 537112 673518 537124
rect 674282 537112 674288 537124
rect 673512 537084 674288 537112
rect 673512 537072 673518 537084
rect 674282 537072 674288 537084
rect 674340 537072 674346 537124
rect 673454 536732 673460 536784
rect 673512 536772 673518 536784
rect 673638 536772 673644 536784
rect 673512 536744 673644 536772
rect 673512 536732 673518 536744
rect 673638 536732 673644 536744
rect 673696 536732 673702 536784
rect 674834 536732 674840 536784
rect 674892 536772 674898 536784
rect 675294 536772 675300 536784
rect 674892 536744 675300 536772
rect 674892 536732 674898 536744
rect 675294 536732 675300 536744
rect 675352 536732 675358 536784
rect 673454 536596 673460 536648
rect 673512 536636 673518 536648
rect 675386 536636 675392 536648
rect 673512 536608 675392 536636
rect 673512 536596 673518 536608
rect 675386 536596 675392 536608
rect 675444 536596 675450 536648
rect 655974 535712 655980 535764
rect 656032 535752 656038 535764
rect 676030 535752 676036 535764
rect 656032 535724 676036 535752
rect 656032 535712 656038 535724
rect 676030 535712 676036 535724
rect 676088 535712 676094 535764
rect 42150 535576 42156 535628
rect 42208 535616 42214 535628
rect 43346 535616 43352 535628
rect 42208 535588 43352 535616
rect 42208 535576 42214 535588
rect 43346 535576 43352 535588
rect 43404 535576 43410 535628
rect 655698 535576 655704 535628
rect 655756 535616 655762 535628
rect 676214 535616 676220 535628
rect 655756 535588 676220 535616
rect 655756 535576 655762 535588
rect 676214 535576 676220 535588
rect 676272 535576 676278 535628
rect 42058 535032 42064 535084
rect 42116 535072 42122 535084
rect 43438 535072 43444 535084
rect 42116 535044 43444 535072
rect 42116 535032 42122 535044
rect 43438 535032 43444 535044
rect 43496 535032 43502 535084
rect 42150 534420 42156 534472
rect 42208 534460 42214 534472
rect 43898 534460 43904 534472
rect 42208 534432 43904 534460
rect 42208 534420 42214 534432
rect 43898 534420 43904 534432
rect 43956 534420 43962 534472
rect 42150 533944 42156 533996
rect 42208 533984 42214 533996
rect 43070 533984 43076 533996
rect 42208 533956 43076 533984
rect 42208 533944 42214 533956
rect 43070 533944 43076 533956
rect 43128 533944 43134 533996
rect 655790 532856 655796 532908
rect 655848 532896 655854 532908
rect 679158 532896 679164 532908
rect 655848 532868 679164 532896
rect 655848 532856 655854 532868
rect 679158 532856 679164 532868
rect 679216 532856 679222 532908
rect 675018 532652 675024 532704
rect 675076 532692 675082 532704
rect 676030 532692 676036 532704
rect 675076 532664 676036 532692
rect 675076 532652 675082 532664
rect 676030 532652 676036 532664
rect 676088 532652 676094 532704
rect 42150 531428 42156 531480
rect 42208 531468 42214 531480
rect 43530 531468 43536 531480
rect 42208 531440 43536 531468
rect 42208 531428 42214 531440
rect 43530 531428 43536 531440
rect 43588 531428 43594 531480
rect 42150 530884 42156 530936
rect 42208 530924 42214 530936
rect 42702 530924 42708 530936
rect 42208 530896 42708 530924
rect 42208 530884 42214 530896
rect 42702 530884 42708 530896
rect 42760 530884 42766 530936
rect 42426 530068 42432 530120
rect 42484 530068 42490 530120
rect 42444 530040 42472 530068
rect 42352 530012 42472 530040
rect 42242 529592 42248 529644
rect 42300 529632 42306 529644
rect 42352 529632 42380 530012
rect 42426 529932 42432 529984
rect 42484 529972 42490 529984
rect 58526 529972 58532 529984
rect 42484 529944 58532 529972
rect 42484 529932 42490 529944
rect 58526 529932 58532 529944
rect 58584 529932 58590 529984
rect 46106 529864 46112 529916
rect 46164 529904 46170 529916
rect 58342 529904 58348 529916
rect 46164 529876 58348 529904
rect 46164 529864 46170 529876
rect 58342 529864 58348 529876
rect 58400 529864 58406 529916
rect 675202 529864 675208 529916
rect 675260 529904 675266 529916
rect 676030 529904 676036 529916
rect 675260 529876 676036 529904
rect 675260 529864 675266 529876
rect 676030 529864 676036 529876
rect 676088 529864 676094 529916
rect 42300 529604 42380 529632
rect 42300 529592 42306 529604
rect 675110 529456 675116 529508
rect 675168 529496 675174 529508
rect 676030 529496 676036 529508
rect 675168 529468 676036 529496
rect 675168 529456 675174 529468
rect 676030 529456 676036 529468
rect 676088 529456 676094 529508
rect 674558 527824 674564 527876
rect 674616 527864 674622 527876
rect 676030 527864 676036 527876
rect 674616 527836 676036 527864
rect 674616 527824 674622 527836
rect 676030 527824 676036 527836
rect 676088 527824 676094 527876
rect 42150 527756 42156 527808
rect 42208 527796 42214 527808
rect 43162 527796 43168 527808
rect 42208 527768 43168 527796
rect 42208 527756 42214 527768
rect 43162 527756 43168 527768
rect 43220 527756 43226 527808
rect 48314 527076 48320 527128
rect 48372 527116 48378 527128
rect 58066 527116 58072 527128
rect 48372 527088 58072 527116
rect 48372 527076 48378 527088
rect 58066 527076 58072 527088
rect 58124 527076 58130 527128
rect 674466 527076 674472 527128
rect 674524 527116 674530 527128
rect 676030 527116 676036 527128
rect 674524 527088 676036 527116
rect 674524 527076 674530 527088
rect 676030 527076 676036 527088
rect 676088 527076 676094 527128
rect 50982 527008 50988 527060
rect 51040 527048 51046 527060
rect 57974 527048 57980 527060
rect 51040 527020 57980 527048
rect 51040 527008 51046 527020
rect 57974 527008 57980 527020
rect 58032 527008 58038 527060
rect 673730 527008 673736 527060
rect 673788 527048 673794 527060
rect 675938 527048 675944 527060
rect 673788 527020 675944 527048
rect 673788 527008 673794 527020
rect 675938 527008 675944 527020
rect 675996 527008 676002 527060
rect 42334 526600 42340 526652
rect 42392 526640 42398 526652
rect 43070 526640 43076 526652
rect 42392 526612 43076 526640
rect 42392 526600 42398 526612
rect 43070 526600 43076 526612
rect 43128 526600 43134 526652
rect 672442 524424 672448 524476
rect 672500 524464 672506 524476
rect 679066 524464 679072 524476
rect 672500 524436 679072 524464
rect 672500 524424 672506 524436
rect 679066 524424 679072 524436
rect 679124 524424 679130 524476
rect 676122 521568 676128 521620
rect 676180 521608 676186 521620
rect 678974 521608 678980 521620
rect 676180 521580 678980 521608
rect 676180 521568 676186 521580
rect 678974 521568 678980 521580
rect 679032 521568 679038 521620
rect 677390 521500 677396 521552
rect 677448 521540 677454 521552
rect 679158 521540 679164 521552
rect 677448 521512 679164 521540
rect 677448 521500 677454 521512
rect 679158 521500 679164 521512
rect 679216 521500 679222 521552
rect 677298 521432 677304 521484
rect 677356 521472 677362 521484
rect 679342 521472 679348 521484
rect 677356 521444 679348 521472
rect 677356 521432 677362 521444
rect 679342 521432 679348 521444
rect 679400 521432 679406 521484
rect 677482 521364 677488 521416
rect 677540 521404 677546 521416
rect 679250 521404 679256 521416
rect 677540 521376 679256 521404
rect 677540 521364 677546 521376
rect 679250 521364 679256 521376
rect 679308 521364 679314 521416
rect 655606 491648 655612 491700
rect 655664 491688 655670 491700
rect 676030 491688 676036 491700
rect 655664 491660 676036 491688
rect 655664 491648 655670 491660
rect 676030 491648 676036 491660
rect 676088 491648 676094 491700
rect 655514 491512 655520 491564
rect 655572 491552 655578 491564
rect 676030 491552 676036 491564
rect 655572 491524 676036 491552
rect 655572 491512 655578 491524
rect 676030 491512 676036 491524
rect 676088 491512 676094 491564
rect 655422 491376 655428 491428
rect 655480 491416 655486 491428
rect 675938 491416 675944 491428
rect 655480 491388 675944 491416
rect 655480 491376 655486 491388
rect 675938 491376 675944 491388
rect 675996 491376 676002 491428
rect 676214 491240 676220 491292
rect 676272 491280 676278 491292
rect 677298 491280 677304 491292
rect 676272 491252 677304 491280
rect 676272 491240 676278 491252
rect 677298 491240 677304 491252
rect 677356 491240 677362 491292
rect 676214 490764 676220 490816
rect 676272 490804 676278 490816
rect 677482 490804 677488 490816
rect 676272 490776 677488 490804
rect 676272 490764 676278 490776
rect 677482 490764 677488 490776
rect 677540 490764 677546 490816
rect 676214 489948 676220 490000
rect 676272 489988 676278 490000
rect 677390 489988 677396 490000
rect 676272 489960 677396 489988
rect 676272 489948 676278 489960
rect 677390 489948 677396 489960
rect 677448 489948 677454 490000
rect 676030 489336 676036 489388
rect 676088 489376 676094 489388
rect 676088 489348 676168 489376
rect 676088 489336 676094 489348
rect 676140 489184 676168 489348
rect 676122 489132 676128 489184
rect 676180 489132 676186 489184
rect 674926 488452 674932 488504
rect 674984 488492 674990 488504
rect 676030 488492 676036 488504
rect 674984 488464 676036 488492
rect 674984 488452 674990 488464
rect 676030 488452 676036 488464
rect 676088 488452 676094 488504
rect 674282 488384 674288 488436
rect 674340 488424 674346 488436
rect 675846 488424 675852 488436
rect 674340 488396 675852 488424
rect 674340 488384 674346 488396
rect 675846 488384 675852 488396
rect 675904 488384 675910 488436
rect 673454 488316 673460 488368
rect 673512 488356 673518 488368
rect 675478 488356 675484 488368
rect 673512 488328 675484 488356
rect 673512 488316 673518 488328
rect 675478 488316 675484 488328
rect 675536 488316 675542 488368
rect 674834 485732 674840 485784
rect 674892 485772 674898 485784
rect 676030 485772 676036 485784
rect 674892 485744 676036 485772
rect 674892 485732 674898 485744
rect 676030 485732 676036 485744
rect 676088 485732 676094 485784
rect 673638 485664 673644 485716
rect 673696 485704 673702 485716
rect 675846 485704 675852 485716
rect 673696 485676 675852 485704
rect 673696 485664 673702 485676
rect 675846 485664 675852 485676
rect 675904 485664 675910 485716
rect 674742 485460 674748 485512
rect 674800 485500 674806 485512
rect 676030 485500 676036 485512
rect 674800 485472 676036 485500
rect 674800 485460 674806 485472
rect 676030 485460 676036 485472
rect 676088 485460 676094 485512
rect 674650 483828 674656 483880
rect 674708 483868 674714 483880
rect 676030 483868 676036 483880
rect 674708 483840 676036 483868
rect 674708 483828 674714 483840
rect 676030 483828 676036 483840
rect 676088 483828 676094 483880
rect 673546 483420 673552 483472
rect 673604 483460 673610 483472
rect 676030 483460 676036 483472
rect 673604 483432 676036 483460
rect 673604 483420 673610 483432
rect 676030 483420 676036 483432
rect 676088 483420 676094 483472
rect 673822 482944 673828 482996
rect 673880 482984 673886 482996
rect 676030 482984 676036 482996
rect 673880 482956 676036 482984
rect 673880 482944 673886 482956
rect 676030 482944 676036 482956
rect 676088 482944 676094 482996
rect 672534 480700 672540 480752
rect 672592 480740 672598 480752
rect 676030 480740 676036 480752
rect 672592 480712 676036 480740
rect 672592 480700 672598 480712
rect 676030 480700 676036 480712
rect 676088 480700 676094 480752
rect 41782 430856 41788 430908
rect 41840 430896 41846 430908
rect 50982 430896 50988 430908
rect 41840 430868 50988 430896
rect 41840 430856 41846 430868
rect 50982 430856 50988 430868
rect 51040 430856 51046 430908
rect 41782 430448 41788 430500
rect 41840 430488 41846 430500
rect 48406 430488 48412 430500
rect 41840 430460 48412 430488
rect 41840 430448 41846 430460
rect 48406 430448 48412 430460
rect 48464 430448 48470 430500
rect 41782 430040 41788 430092
rect 41840 430080 41846 430092
rect 46106 430080 46112 430092
rect 41840 430052 46112 430080
rect 41840 430040 41846 430052
rect 46106 430040 46112 430052
rect 46164 430040 46170 430092
rect 41782 429904 41788 429956
rect 41840 429944 41846 429956
rect 43346 429944 43352 429956
rect 41840 429916 43352 429944
rect 41840 429904 41846 429916
rect 43346 429904 43352 429916
rect 43404 429904 43410 429956
rect 41782 429020 41788 429072
rect 41840 429060 41846 429072
rect 43898 429060 43904 429072
rect 41840 429032 43904 429060
rect 41840 429020 41846 429032
rect 43898 429020 43904 429032
rect 43956 429020 43962 429072
rect 41782 428884 41788 428936
rect 41840 428924 41846 428936
rect 43714 428924 43720 428936
rect 41840 428896 43720 428924
rect 41840 428884 41846 428896
rect 43714 428884 43720 428896
rect 43772 428884 43778 428936
rect 41782 426504 41788 426556
rect 41840 426544 41846 426556
rect 43714 426544 43720 426556
rect 41840 426516 43720 426544
rect 41840 426504 41846 426516
rect 43714 426504 43720 426516
rect 43772 426504 43778 426556
rect 41782 426368 41788 426420
rect 41840 426408 41846 426420
rect 43806 426408 43812 426420
rect 41840 426380 43812 426408
rect 41840 426368 41846 426380
rect 43806 426368 43812 426380
rect 43864 426368 43870 426420
rect 41782 425416 41788 425468
rect 41840 425456 41846 425468
rect 42702 425456 42708 425468
rect 41840 425428 42708 425456
rect 41840 425416 41846 425428
rect 42702 425416 42708 425428
rect 42760 425416 42766 425468
rect 41782 425144 41788 425196
rect 41840 425184 41846 425196
rect 43254 425184 43260 425196
rect 41840 425156 43260 425184
rect 41840 425144 41846 425156
rect 43254 425144 43260 425156
rect 43312 425144 43318 425196
rect 41874 423648 41880 423700
rect 41932 423688 41938 423700
rect 43530 423688 43536 423700
rect 41932 423660 43536 423688
rect 41932 423648 41938 423660
rect 43530 423648 43536 423660
rect 43588 423648 43594 423700
rect 41874 423512 41880 423564
rect 41932 423552 41938 423564
rect 43070 423552 43076 423564
rect 41932 423524 43076 423552
rect 41932 423512 41938 423524
rect 43070 423512 43076 423524
rect 43128 423512 43134 423564
rect 41874 422900 41880 422952
rect 41932 422940 41938 422952
rect 43622 422940 43628 422952
rect 41932 422912 43628 422940
rect 41932 422900 41938 422912
rect 43622 422900 43628 422912
rect 43680 422900 43686 422952
rect 41874 422628 41880 422680
rect 41932 422668 41938 422680
rect 43438 422668 43444 422680
rect 41932 422640 43444 422668
rect 41932 422628 41938 422640
rect 43438 422628 43444 422640
rect 43496 422628 43502 422680
rect 41782 422424 41788 422476
rect 41840 422464 41846 422476
rect 43990 422464 43996 422476
rect 41840 422436 43996 422464
rect 41840 422424 41846 422436
rect 43990 422424 43996 422436
rect 44048 422424 44054 422476
rect 41782 422288 41788 422340
rect 41840 422328 41846 422340
rect 44082 422328 44088 422340
rect 41840 422300 44088 422328
rect 41840 422288 41846 422300
rect 44082 422288 44088 422300
rect 44140 422288 44146 422340
rect 41782 421540 41788 421592
rect 41840 421580 41846 421592
rect 43346 421580 43352 421592
rect 41840 421552 43352 421580
rect 41840 421540 41846 421552
rect 43346 421540 43352 421552
rect 43404 421540 43410 421592
rect 41782 419432 41788 419484
rect 41840 419472 41846 419484
rect 48314 419472 48320 419484
rect 41840 419444 48320 419472
rect 41840 419432 41846 419444
rect 48314 419432 48320 419444
rect 48372 419432 48378 419484
rect 41874 416304 41880 416356
rect 41932 416344 41938 416356
rect 43162 416344 43168 416356
rect 41932 416316 43168 416344
rect 41932 416304 41938 416316
rect 43162 416304 43168 416316
rect 43220 416304 43226 416356
rect 43990 413924 43996 413976
rect 44048 413964 44054 413976
rect 44266 413964 44272 413976
rect 44048 413936 44272 413964
rect 44048 413924 44054 413936
rect 44266 413924 44272 413936
rect 44324 413924 44330 413976
rect 44082 413856 44088 413908
rect 44140 413896 44146 413908
rect 44174 413896 44180 413908
rect 44140 413868 44180 413896
rect 44140 413856 44146 413868
rect 44174 413856 44180 413868
rect 44232 413856 44238 413908
rect 42058 413788 42064 413840
rect 42116 413828 42122 413840
rect 43990 413828 43996 413840
rect 42116 413800 43996 413828
rect 42116 413788 42122 413800
rect 43990 413788 43996 413800
rect 44048 413788 44054 413840
rect 42426 413720 42432 413772
rect 42484 413760 42490 413772
rect 44082 413760 44088 413772
rect 42484 413732 44088 413760
rect 42484 413720 42490 413732
rect 44082 413720 44088 413732
rect 44140 413720 44146 413772
rect 41966 413380 41972 413432
rect 42024 413380 42030 413432
rect 41984 413216 42012 413380
rect 41984 413188 42288 413216
rect 42260 413024 42288 413188
rect 42242 412972 42248 413024
rect 42300 412972 42306 413024
rect 43254 411272 43260 411324
rect 43312 411312 43318 411324
rect 43898 411312 43904 411324
rect 43312 411284 43904 411312
rect 43312 411272 43318 411284
rect 43898 411272 43904 411284
rect 43956 411272 43962 411324
rect 43898 411136 43904 411188
rect 43956 411176 43962 411188
rect 44174 411176 44180 411188
rect 43956 411148 44180 411176
rect 43956 411136 43962 411148
rect 44174 411136 44180 411148
rect 44232 411136 44238 411188
rect 42150 409708 42156 409760
rect 42208 409748 42214 409760
rect 42334 409748 42340 409760
rect 42208 409720 42340 409748
rect 42208 409708 42214 409720
rect 42334 409708 42340 409720
rect 42392 409708 42398 409760
rect 42150 409436 42156 409488
rect 42208 409476 42214 409488
rect 43438 409476 43444 409488
rect 42208 409448 43444 409476
rect 42208 409436 42214 409448
rect 43438 409436 43444 409448
rect 43496 409436 43502 409488
rect 43070 409300 43076 409352
rect 43128 409340 43134 409352
rect 43438 409340 43444 409352
rect 43128 409312 43444 409340
rect 43128 409300 43134 409312
rect 43438 409300 43444 409312
rect 43496 409300 43502 409352
rect 42150 407872 42156 407924
rect 42208 407912 42214 407924
rect 43070 407912 43076 407924
rect 42208 407884 43076 407912
rect 42208 407872 42214 407884
rect 43070 407872 43076 407884
rect 43128 407872 43134 407924
rect 42242 407532 42248 407584
rect 42300 407572 42306 407584
rect 43898 407572 43904 407584
rect 42300 407544 43904 407572
rect 42300 407532 42306 407544
rect 43898 407532 43904 407544
rect 43956 407532 43962 407584
rect 42058 406988 42064 407040
rect 42116 407028 42122 407040
rect 43162 407028 43168 407040
rect 42116 407000 43168 407028
rect 42116 406988 42122 407000
rect 43162 406988 43168 407000
rect 43220 406988 43226 407040
rect 42242 406920 42248 406972
rect 42300 406960 42306 406972
rect 44266 406960 44272 406972
rect 42300 406932 44272 406960
rect 42300 406920 42306 406932
rect 44266 406920 44272 406932
rect 44324 406920 44330 406972
rect 42334 405628 42340 405680
rect 42392 405668 42398 405680
rect 58434 405668 58440 405680
rect 42392 405640 58440 405668
rect 42392 405628 42398 405640
rect 58434 405628 58440 405640
rect 58492 405628 58498 405680
rect 42334 405492 42340 405544
rect 42392 405532 42398 405544
rect 43346 405532 43352 405544
rect 42392 405504 43352 405532
rect 42392 405492 42398 405504
rect 43346 405492 43352 405504
rect 43404 405492 43410 405544
rect 42426 405152 42432 405204
rect 42484 405192 42490 405204
rect 42702 405192 42708 405204
rect 42484 405164 42708 405192
rect 42484 405152 42490 405164
rect 42702 405152 42708 405164
rect 42760 405152 42766 405204
rect 42334 403316 42340 403368
rect 42392 403356 42398 403368
rect 43622 403356 43628 403368
rect 42392 403328 43628 403356
rect 42392 403316 42398 403328
rect 43622 403316 43628 403328
rect 43680 403316 43686 403368
rect 655698 403112 655704 403164
rect 655756 403152 655762 403164
rect 676122 403152 676128 403164
rect 655756 403124 676128 403152
rect 655756 403112 655762 403124
rect 676122 403112 676128 403124
rect 676180 403112 676186 403164
rect 655514 403044 655520 403096
rect 655572 403084 655578 403096
rect 676214 403084 676220 403096
rect 655572 403056 676220 403084
rect 655572 403044 655578 403056
rect 676214 403044 676220 403056
rect 676272 403044 676278 403096
rect 655422 402976 655428 403028
rect 655480 403016 655486 403028
rect 676122 403016 676128 403028
rect 655480 402988 676128 403016
rect 655480 402976 655486 402988
rect 676122 402976 676128 402988
rect 676180 402976 676186 403028
rect 43070 402908 43076 402960
rect 43128 402948 43134 402960
rect 58526 402948 58532 402960
rect 43128 402920 58532 402948
rect 43128 402908 43134 402920
rect 58526 402908 58532 402920
rect 58584 402908 58590 402960
rect 42242 402568 42248 402620
rect 42300 402608 42306 402620
rect 43530 402608 43536 402620
rect 42300 402580 43536 402608
rect 42300 402568 42306 402580
rect 43530 402568 43536 402580
rect 43588 402568 43594 402620
rect 42150 402500 42156 402552
rect 42208 402540 42214 402552
rect 43438 402540 43444 402552
rect 42208 402512 43444 402540
rect 42208 402500 42214 402512
rect 43438 402500 43444 402512
rect 43496 402500 43502 402552
rect 42150 401820 42156 401872
rect 42208 401860 42214 401872
rect 43162 401860 43168 401872
rect 42208 401832 43168 401860
rect 42208 401820 42214 401832
rect 43162 401820 43168 401832
rect 43220 401820 43226 401872
rect 42150 400188 42156 400240
rect 42208 400228 42214 400240
rect 43806 400228 43812 400240
rect 42208 400200 43812 400228
rect 42208 400188 42214 400200
rect 43806 400188 43812 400200
rect 43864 400188 43870 400240
rect 46106 400120 46112 400172
rect 46164 400160 46170 400172
rect 58434 400160 58440 400172
rect 46164 400132 58440 400160
rect 46164 400120 46170 400132
rect 58434 400120 58440 400132
rect 58492 400120 58498 400172
rect 48406 400052 48412 400104
rect 48464 400092 48470 400104
rect 58342 400092 58348 400104
rect 48464 400064 58348 400092
rect 48464 400052 48470 400064
rect 58342 400052 58348 400064
rect 58400 400052 58406 400104
rect 50982 399984 50988 400036
rect 51040 400024 51046 400036
rect 58526 400024 58532 400036
rect 51040 399996 58532 400024
rect 51040 399984 51046 399996
rect 58526 399984 58532 399996
rect 58584 399984 58590 400036
rect 674282 399440 674288 399492
rect 674340 399480 674346 399492
rect 676030 399480 676036 399492
rect 674340 399452 676036 399480
rect 674340 399440 674346 399452
rect 676030 399440 676036 399452
rect 676088 399440 676094 399492
rect 674558 398216 674564 398268
rect 674616 398256 674622 398268
rect 676030 398256 676036 398268
rect 674616 398228 676036 398256
rect 674616 398216 674622 398228
rect 676030 398216 676036 398228
rect 676088 398216 676094 398268
rect 675018 397604 675024 397656
rect 675076 397644 675082 397656
rect 675938 397644 675944 397656
rect 675076 397616 675944 397644
rect 675076 397604 675082 397616
rect 675938 397604 675944 397616
rect 675996 397604 676002 397656
rect 673638 397536 673644 397588
rect 673696 397576 673702 397588
rect 676122 397576 676128 397588
rect 673696 397548 676128 397576
rect 673696 397536 673702 397548
rect 676122 397536 676128 397548
rect 676180 397536 676186 397588
rect 674650 397468 674656 397520
rect 674708 397508 674714 397520
rect 676030 397508 676036 397520
rect 674708 397480 676036 397508
rect 674708 397468 674714 397480
rect 676030 397468 676036 397480
rect 676088 397468 676094 397520
rect 674466 396992 674472 397044
rect 674524 397032 674530 397044
rect 676030 397032 676036 397044
rect 674524 397004 676036 397032
rect 674524 396992 674530 397004
rect 676030 396992 676036 397004
rect 676088 396992 676094 397044
rect 673454 395360 673460 395412
rect 673512 395400 673518 395412
rect 675662 395400 675668 395412
rect 673512 395372 675668 395400
rect 673512 395360 673518 395372
rect 675662 395360 675668 395372
rect 675720 395360 675726 395412
rect 674742 394952 674748 395004
rect 674800 394992 674806 395004
rect 675938 394992 675944 395004
rect 674800 394964 675944 394992
rect 674800 394952 674806 394964
rect 675938 394952 675944 394964
rect 675996 394952 676002 395004
rect 673546 394884 673552 394936
rect 673604 394924 673610 394936
rect 675662 394924 675668 394936
rect 673604 394896 675668 394924
rect 673604 394884 673610 394896
rect 675662 394884 675668 394896
rect 675720 394884 675726 394936
rect 674834 394816 674840 394868
rect 674892 394856 674898 394868
rect 676122 394856 676128 394868
rect 674892 394828 676128 394856
rect 674892 394816 674898 394828
rect 676122 394816 676128 394828
rect 676180 394816 676186 394868
rect 675110 394748 675116 394800
rect 675168 394788 675174 394800
rect 675938 394788 675944 394800
rect 675168 394760 675944 394788
rect 675168 394748 675174 394760
rect 675938 394748 675944 394760
rect 675996 394748 676002 394800
rect 675202 394680 675208 394732
rect 675260 394720 675266 394732
rect 676030 394720 676036 394732
rect 675260 394692 676036 394720
rect 675260 394680 675266 394692
rect 676030 394680 676036 394692
rect 676088 394680 676094 394732
rect 42150 394612 42156 394664
rect 42208 394652 42214 394664
rect 60366 394652 60372 394664
rect 42208 394624 60372 394652
rect 42208 394612 42214 394624
rect 60366 394612 60372 394624
rect 60424 394612 60430 394664
rect 673730 394136 673736 394188
rect 673788 394176 673794 394188
rect 676030 394176 676036 394188
rect 673788 394148 676036 394176
rect 673788 394136 673794 394148
rect 676030 394136 676036 394148
rect 676088 394136 676094 394188
rect 672626 392028 672632 392080
rect 672684 392068 672690 392080
rect 678974 392068 678980 392080
rect 672684 392040 678980 392068
rect 672684 392028 672690 392040
rect 678974 392028 678980 392040
rect 679032 392028 679038 392080
rect 673822 391960 673828 392012
rect 673880 392000 673886 392012
rect 676030 392000 676036 392012
rect 673880 391972 676036 392000
rect 673880 391960 673886 391972
rect 676030 391960 676036 391972
rect 676088 391960 676094 392012
rect 674926 390532 674932 390584
rect 674984 390572 674990 390584
rect 675754 390572 675760 390584
rect 674984 390544 675760 390572
rect 674984 390532 674990 390544
rect 675754 390532 675760 390544
rect 675812 390532 675818 390584
rect 41506 388016 41512 388068
rect 41564 388056 41570 388068
rect 43254 388056 43260 388068
rect 41564 388028 43260 388056
rect 41564 388016 41570 388028
rect 43254 388016 43260 388028
rect 43312 388016 43318 388068
rect 41414 387472 41420 387524
rect 41472 387512 41478 387524
rect 50982 387512 50988 387524
rect 41472 387484 50988 387512
rect 41472 387472 41478 387484
rect 50982 387472 50988 387484
rect 51040 387472 51046 387524
rect 41414 387064 41420 387116
rect 41472 387104 41478 387116
rect 48498 387104 48504 387116
rect 41472 387076 48504 387104
rect 41472 387064 41478 387076
rect 48498 387064 48504 387076
rect 48556 387064 48562 387116
rect 41782 386792 41788 386844
rect 41840 386832 41846 386844
rect 46106 386832 46112 386844
rect 41840 386804 46112 386832
rect 41840 386792 41846 386804
rect 46106 386792 46112 386804
rect 46164 386792 46170 386844
rect 675754 386588 675760 386640
rect 675812 386588 675818 386640
rect 41782 386316 41788 386368
rect 41840 386356 41846 386368
rect 43714 386356 43720 386368
rect 41840 386328 43720 386356
rect 41840 386316 41846 386328
rect 43714 386316 43720 386328
rect 43772 386316 43778 386368
rect 675018 386112 675024 386164
rect 675076 386112 675082 386164
rect 41506 386044 41512 386096
rect 41564 386084 41570 386096
rect 44082 386084 44088 386096
rect 41564 386056 44088 386084
rect 41564 386044 41570 386056
rect 44082 386044 44088 386056
rect 44140 386044 44146 386096
rect 675036 386084 675064 386112
rect 674944 386056 675064 386084
rect 41506 385772 41512 385824
rect 41564 385812 41570 385824
rect 43990 385812 43996 385824
rect 41564 385784 43996 385812
rect 41564 385772 41570 385784
rect 43990 385772 43996 385784
rect 44048 385772 44054 385824
rect 674944 385064 674972 386056
rect 675772 386028 675800 386588
rect 675018 385976 675024 386028
rect 675076 386016 675082 386028
rect 675386 386016 675392 386028
rect 675076 385988 675392 386016
rect 675076 385976 675082 385988
rect 675386 385976 675392 385988
rect 675444 385976 675450 386028
rect 675754 385976 675760 386028
rect 675812 385976 675818 386028
rect 675202 385568 675208 385620
rect 675260 385608 675266 385620
rect 675386 385608 675392 385620
rect 675260 385580 675392 385608
rect 675260 385568 675266 385580
rect 675386 385568 675392 385580
rect 675444 385568 675450 385620
rect 674208 385036 674972 385064
rect 674208 384860 674236 385036
rect 674282 384956 674288 385008
rect 674340 384996 674346 385008
rect 675202 384996 675208 385008
rect 674340 384968 675208 384996
rect 674340 384956 674346 384968
rect 675202 384956 675208 384968
rect 675260 384956 675266 385008
rect 674282 384860 674288 384872
rect 674208 384832 674288 384860
rect 674282 384820 674288 384832
rect 674340 384820 674346 384872
rect 674558 384752 674564 384804
rect 674616 384792 674622 384804
rect 675386 384792 675392 384804
rect 674616 384764 675392 384792
rect 674616 384752 674622 384764
rect 675386 384752 675392 384764
rect 675444 384752 675450 384804
rect 41874 383732 41880 383784
rect 41932 383772 41938 383784
rect 44082 383772 44088 383784
rect 41932 383744 44088 383772
rect 41932 383732 41938 383744
rect 44082 383732 44088 383744
rect 44140 383732 44146 383784
rect 41506 383664 41512 383716
rect 41564 383704 41570 383716
rect 43806 383704 43812 383716
rect 41564 383676 43812 383704
rect 41564 383664 41570 383676
rect 43806 383664 43812 383676
rect 43864 383664 43870 383716
rect 674650 383120 674656 383172
rect 674708 383160 674714 383172
rect 675386 383160 675392 383172
rect 674708 383132 675392 383160
rect 674708 383120 674714 383132
rect 675386 383120 675392 383132
rect 675444 383120 675450 383172
rect 41506 382712 41512 382764
rect 41564 382752 41570 382764
rect 43714 382752 43720 382764
rect 41564 382724 43720 382752
rect 41564 382712 41570 382724
rect 43714 382712 43720 382724
rect 43772 382712 43778 382764
rect 674834 382440 674840 382492
rect 674892 382480 674898 382492
rect 675386 382480 675392 382492
rect 674892 382452 675392 382480
rect 674892 382440 674898 382452
rect 675386 382440 675392 382452
rect 675444 382440 675450 382492
rect 41506 381896 41512 381948
rect 41564 381936 41570 381948
rect 42702 381936 42708 381948
rect 41564 381908 42708 381936
rect 41564 381896 41570 381908
rect 42702 381896 42708 381908
rect 42760 381896 42766 381948
rect 674742 381896 674748 381948
rect 674800 381936 674806 381948
rect 675386 381936 675392 381948
rect 674800 381908 675392 381936
rect 674800 381896 674806 381908
rect 675386 381896 675392 381908
rect 675444 381896 675450 381948
rect 41506 381760 41512 381812
rect 41564 381800 41570 381812
rect 43070 381800 43076 381812
rect 41564 381772 43076 381800
rect 41564 381760 41570 381772
rect 43070 381760 43076 381772
rect 43128 381760 43134 381812
rect 41506 381216 41512 381268
rect 41564 381256 41570 381268
rect 43622 381256 43628 381268
rect 41564 381228 43628 381256
rect 41564 381216 41570 381228
rect 43622 381216 43628 381228
rect 43680 381216 43686 381268
rect 675110 381216 675116 381268
rect 675168 381256 675174 381268
rect 675168 381228 675432 381256
rect 675168 381216 675174 381228
rect 675404 381132 675432 381228
rect 674926 381080 674932 381132
rect 674984 381120 674990 381132
rect 675110 381120 675116 381132
rect 674984 381092 675116 381120
rect 674984 381080 674990 381092
rect 675110 381080 675116 381092
rect 675168 381080 675174 381132
rect 675386 381080 675392 381132
rect 675444 381080 675450 381132
rect 673638 381012 673644 381064
rect 673696 381052 673702 381064
rect 673696 381024 674512 381052
rect 673696 381012 673702 381024
rect 674484 380928 674512 381024
rect 673638 380876 673644 380928
rect 673696 380916 673702 380928
rect 674282 380916 674288 380928
rect 673696 380888 674288 380916
rect 673696 380876 673702 380888
rect 674282 380876 674288 380888
rect 674340 380876 674346 380928
rect 674466 380876 674472 380928
rect 674524 380876 674530 380928
rect 41506 380128 41512 380180
rect 41564 380168 41570 380180
rect 43622 380168 43628 380180
rect 41564 380140 43628 380168
rect 41564 380128 41570 380140
rect 43622 380128 43628 380140
rect 43680 380128 43686 380180
rect 41506 379448 41512 379500
rect 41564 379488 41570 379500
rect 43990 379488 43996 379500
rect 41564 379460 43996 379488
rect 41564 379448 41570 379460
rect 43990 379448 43996 379460
rect 44048 379448 44054 379500
rect 41414 378904 41420 378956
rect 41472 378944 41478 378956
rect 43346 378944 43352 378956
rect 41472 378916 43352 378944
rect 41472 378904 41478 378916
rect 43346 378904 43352 378916
rect 43404 378904 43410 378956
rect 673638 378768 673644 378820
rect 673696 378808 673702 378820
rect 675386 378808 675392 378820
rect 673696 378780 675392 378808
rect 673696 378768 673702 378780
rect 675386 378768 675392 378780
rect 675444 378768 675450 378820
rect 41506 378496 41512 378548
rect 41564 378536 41570 378548
rect 43162 378536 43168 378548
rect 41564 378508 43168 378536
rect 41564 378496 41570 378508
rect 43162 378496 43168 378508
rect 43220 378496 43226 378548
rect 41598 378224 41604 378276
rect 41656 378264 41662 378276
rect 43438 378264 43444 378276
rect 41656 378236 43444 378264
rect 41656 378224 41662 378236
rect 43438 378224 43444 378236
rect 43496 378224 43502 378276
rect 673730 377952 673736 378004
rect 673788 377992 673794 378004
rect 675478 377992 675484 378004
rect 673788 377964 675484 377992
rect 673788 377952 673794 377964
rect 675478 377952 675484 377964
rect 675536 377952 675542 378004
rect 673546 377408 673552 377460
rect 673604 377448 673610 377460
rect 675386 377448 675392 377460
rect 673604 377420 675392 377448
rect 673604 377408 673610 377420
rect 675386 377408 675392 377420
rect 675444 377408 675450 377460
rect 673822 376932 673828 376984
rect 673880 376972 673886 376984
rect 675478 376972 675484 376984
rect 673880 376944 675484 376972
rect 673880 376932 673886 376944
rect 675478 376932 675484 376944
rect 675536 376932 675542 376984
rect 41414 376048 41420 376100
rect 41472 376088 41478 376100
rect 48406 376088 48412 376100
rect 41472 376060 48412 376088
rect 41472 376048 41478 376060
rect 48406 376048 48412 376060
rect 48464 376048 48470 376100
rect 673454 375708 673460 375760
rect 673512 375748 673518 375760
rect 675386 375748 675392 375760
rect 673512 375720 675392 375748
rect 673512 375708 673518 375720
rect 675386 375708 675392 375720
rect 675444 375708 675450 375760
rect 42426 374892 42432 374944
rect 42484 374932 42490 374944
rect 44082 374932 44088 374944
rect 42484 374904 44088 374932
rect 42484 374892 42490 374904
rect 44082 374892 44088 374904
rect 44140 374892 44146 374944
rect 674466 373872 674472 373924
rect 674524 373912 674530 373924
rect 675386 373912 675392 373924
rect 674524 373884 675392 373912
rect 674524 373872 674530 373884
rect 675386 373872 675392 373884
rect 675444 373872 675450 373924
rect 654502 372512 654508 372564
rect 654560 372552 654566 372564
rect 675018 372552 675024 372564
rect 654560 372524 675024 372552
rect 654560 372512 654566 372524
rect 675018 372512 675024 372524
rect 675076 372512 675082 372564
rect 674650 372036 674656 372088
rect 674708 372076 674714 372088
rect 675386 372076 675392 372088
rect 674708 372048 675392 372076
rect 674708 372036 674714 372048
rect 675386 372036 675392 372048
rect 675444 372036 675450 372088
rect 41506 371968 41512 372020
rect 41564 372008 41570 372020
rect 43254 372008 43260 372020
rect 41564 371980 43260 372008
rect 41564 371968 41570 371980
rect 43254 371968 43260 371980
rect 43312 371968 43318 372020
rect 43622 371356 43628 371408
rect 43680 371396 43686 371408
rect 43680 371368 43944 371396
rect 43680 371356 43686 371368
rect 43622 371220 43628 371272
rect 43680 371260 43686 371272
rect 43806 371260 43812 371272
rect 43680 371232 43812 371260
rect 43680 371220 43686 371232
rect 43806 371220 43812 371232
rect 43864 371220 43870 371272
rect 43916 371000 43944 371368
rect 43898 370948 43904 371000
rect 43956 370948 43962 371000
rect 675202 370744 675208 370796
rect 675260 370784 675266 370796
rect 675662 370784 675668 370796
rect 675260 370756 675668 370784
rect 675260 370744 675266 370756
rect 675662 370744 675668 370756
rect 675720 370744 675726 370796
rect 675110 370676 675116 370728
rect 675168 370716 675174 370728
rect 675754 370716 675760 370728
rect 675168 370688 675760 370716
rect 675168 370676 675174 370688
rect 675754 370676 675760 370688
rect 675812 370676 675818 370728
rect 41322 370540 41328 370592
rect 41380 370580 41386 370592
rect 41380 370552 42656 370580
rect 41380 370540 41386 370552
rect 41966 370200 41972 370252
rect 42024 370200 42030 370252
rect 41984 370036 42012 370200
rect 41984 370008 42288 370036
rect 42260 369288 42288 370008
rect 42334 369860 42340 369912
rect 42392 369900 42398 369912
rect 42628 369900 42656 370552
rect 42392 369872 42656 369900
rect 42392 369860 42398 369872
rect 42334 369316 42340 369368
rect 42392 369356 42398 369368
rect 42702 369356 42708 369368
rect 42392 369328 42708 369356
rect 42392 369316 42398 369328
rect 42702 369316 42708 369328
rect 42760 369316 42766 369368
rect 42260 369260 42748 369288
rect 42720 369232 42748 369260
rect 42702 369180 42708 369232
rect 42760 369180 42766 369232
rect 42150 368092 42156 368144
rect 42208 368132 42214 368144
rect 42334 368132 42340 368144
rect 42208 368104 42340 368132
rect 42208 368092 42214 368104
rect 42334 368092 42340 368104
rect 42392 368092 42398 368144
rect 42702 366664 42708 366716
rect 42760 366704 42766 366716
rect 42760 366676 43300 366704
rect 42760 366664 42766 366676
rect 42150 366528 42156 366580
rect 42208 366568 42214 366580
rect 42702 366568 42708 366580
rect 42208 366540 42708 366568
rect 42208 366528 42214 366540
rect 42702 366528 42708 366540
rect 42760 366528 42766 366580
rect 42150 366256 42156 366308
rect 42208 366296 42214 366308
rect 43162 366296 43168 366308
rect 42208 366268 43168 366296
rect 42208 366256 42214 366268
rect 43162 366256 43168 366268
rect 43220 366256 43226 366308
rect 43272 366228 43300 366676
rect 43180 366200 43300 366228
rect 43180 366172 43208 366200
rect 43162 366120 43168 366172
rect 43220 366120 43226 366172
rect 42334 365072 42340 365084
rect 42260 365044 42340 365072
rect 42260 364880 42288 365044
rect 42334 365032 42340 365044
rect 42392 365032 42398 365084
rect 42242 364828 42248 364880
rect 42300 364828 42306 364880
rect 42242 364692 42248 364744
rect 42300 364732 42306 364744
rect 43346 364732 43352 364744
rect 42300 364704 43352 364732
rect 42300 364692 42306 364704
rect 43346 364692 43352 364704
rect 43404 364692 43410 364744
rect 43346 364556 43352 364608
rect 43404 364596 43410 364608
rect 43990 364596 43996 364608
rect 43404 364568 43996 364596
rect 43404 364556 43410 364568
rect 43990 364556 43996 364568
rect 44048 364556 44054 364608
rect 43162 364284 43168 364336
rect 43220 364324 43226 364336
rect 43898 364324 43904 364336
rect 43220 364296 43904 364324
rect 43220 364284 43226 364296
rect 43898 364284 43904 364296
rect 43956 364284 43962 364336
rect 42150 363808 42156 363860
rect 42208 363848 42214 363860
rect 43254 363848 43260 363860
rect 42208 363820 43260 363848
rect 42208 363808 42214 363820
rect 43254 363808 43260 363820
rect 43312 363808 43318 363860
rect 42150 363128 42156 363180
rect 42208 363168 42214 363180
rect 43530 363168 43536 363180
rect 42208 363140 43536 363168
rect 42208 363128 42214 363140
rect 43530 363128 43536 363140
rect 43588 363128 43594 363180
rect 42426 361904 42432 361956
rect 42484 361944 42490 361956
rect 43070 361944 43076 361956
rect 42484 361916 43076 361944
rect 42484 361904 42490 361916
rect 43070 361904 43076 361916
rect 43128 361904 43134 361956
rect 42702 361496 42708 361548
rect 42760 361536 42766 361548
rect 58158 361536 58164 361548
rect 42760 361508 58164 361536
rect 42760 361496 42766 361508
rect 58158 361496 58164 361508
rect 58216 361496 58222 361548
rect 42334 361292 42340 361344
rect 42392 361332 42398 361344
rect 58526 361332 58532 361344
rect 42392 361304 58532 361332
rect 42392 361292 42398 361304
rect 58526 361292 58532 361304
rect 58584 361292 58590 361344
rect 42334 360884 42340 360936
rect 42392 360924 42398 360936
rect 43530 360924 43536 360936
rect 42392 360896 43536 360924
rect 42392 360884 42398 360896
rect 43530 360884 43536 360896
rect 43588 360884 43594 360936
rect 42334 360136 42340 360188
rect 42392 360176 42398 360188
rect 43990 360176 43996 360188
rect 42392 360148 43996 360176
rect 42392 360136 42398 360148
rect 43990 360136 43996 360148
rect 44048 360136 44054 360188
rect 42150 359932 42156 359984
rect 42208 359972 42214 359984
rect 43346 359972 43352 359984
rect 42208 359944 43352 359972
rect 42208 359932 42214 359944
rect 43346 359932 43352 359944
rect 43404 359932 43410 359984
rect 46106 358708 46112 358760
rect 46164 358748 46170 358760
rect 58526 358748 58532 358760
rect 46164 358720 58532 358748
rect 46164 358708 46170 358720
rect 58526 358708 58532 358720
rect 58584 358708 58590 358760
rect 42426 358300 42432 358352
rect 42484 358340 42490 358352
rect 43898 358340 43904 358352
rect 42484 358312 43904 358340
rect 42484 358300 42490 358312
rect 43898 358300 43904 358312
rect 43956 358300 43962 358352
rect 655514 356396 655520 356448
rect 655572 356436 655578 356448
rect 676030 356436 676036 356448
rect 655572 356408 676036 356436
rect 655572 356396 655578 356408
rect 676030 356396 676036 356408
rect 676088 356396 676094 356448
rect 655422 356260 655428 356312
rect 655480 356300 655486 356312
rect 675846 356300 675852 356312
rect 655480 356272 675852 356300
rect 655480 356260 655486 356272
rect 675846 356260 675852 356272
rect 675904 356260 675910 356312
rect 655606 356192 655612 356244
rect 655664 356232 655670 356244
rect 675938 356232 675944 356244
rect 655664 356204 675944 356232
rect 655664 356192 655670 356204
rect 675938 356192 675944 356204
rect 675996 356192 676002 356244
rect 673362 356124 673368 356176
rect 673420 356164 673426 356176
rect 676030 356164 676036 356176
rect 673420 356136 676036 356164
rect 673420 356124 673426 356136
rect 676030 356124 676036 356136
rect 676088 356124 676094 356176
rect 48498 355988 48504 356040
rect 48556 356028 48562 356040
rect 58434 356028 58440 356040
rect 48556 356000 58440 356028
rect 48556 355988 48562 356000
rect 58434 355988 58440 356000
rect 58492 355988 58498 356040
rect 50982 355920 50988 355972
rect 51040 355960 51046 355972
rect 58526 355960 58532 355972
rect 51040 355932 58532 355960
rect 51040 355920 51046 355932
rect 58526 355920 58532 355932
rect 58584 355920 58590 355972
rect 674650 353472 674656 353524
rect 674708 353512 674714 353524
rect 676030 353512 676036 353524
rect 674708 353484 676036 353512
rect 674708 353472 674714 353484
rect 676030 353472 676036 353484
rect 676088 353472 676094 353524
rect 674926 353268 674932 353320
rect 674984 353308 674990 353320
rect 676030 353308 676036 353320
rect 674984 353280 676036 353308
rect 674984 353268 674990 353280
rect 676030 353268 676036 353280
rect 676088 353268 676094 353320
rect 674558 352248 674564 352300
rect 674616 352288 674622 352300
rect 675938 352288 675944 352300
rect 674616 352260 675944 352288
rect 674616 352248 674622 352260
rect 675938 352248 675944 352260
rect 675996 352248 676002 352300
rect 674834 351840 674840 351892
rect 674892 351880 674898 351892
rect 676030 351880 676036 351892
rect 674892 351852 676036 351880
rect 674892 351840 674898 351852
rect 676030 351840 676036 351852
rect 676088 351840 676094 351892
rect 673638 351432 673644 351484
rect 673696 351472 673702 351484
rect 675938 351472 675944 351484
rect 673696 351444 675944 351472
rect 673696 351432 673702 351444
rect 675938 351432 675944 351444
rect 675996 351432 676002 351484
rect 673546 350752 673552 350804
rect 673604 350792 673610 350804
rect 675662 350792 675668 350804
rect 673604 350764 675668 350792
rect 673604 350752 673610 350764
rect 675662 350752 675668 350764
rect 675720 350752 675726 350804
rect 674282 350684 674288 350736
rect 674340 350724 674346 350736
rect 675846 350724 675852 350736
rect 674340 350696 675852 350724
rect 674340 350684 674346 350696
rect 675846 350684 675852 350696
rect 675904 350684 675910 350736
rect 674742 350616 674748 350668
rect 674800 350656 674806 350668
rect 675938 350656 675944 350668
rect 674800 350628 675944 350656
rect 674800 350616 674806 350628
rect 675938 350616 675944 350628
rect 675996 350616 676002 350668
rect 675018 350548 675024 350600
rect 675076 350588 675082 350600
rect 676030 350588 676036 350600
rect 675076 350560 676036 350588
rect 675076 350548 675082 350560
rect 676030 350548 676036 350560
rect 676088 350548 676094 350600
rect 42150 350480 42156 350532
rect 42208 350520 42214 350532
rect 57974 350520 57980 350532
rect 42208 350492 57980 350520
rect 42208 350480 42214 350492
rect 57974 350480 57980 350492
rect 58032 350480 58038 350532
rect 673822 349800 673828 349852
rect 673880 349840 673886 349852
rect 676030 349840 676036 349852
rect 673880 349812 676036 349840
rect 673880 349800 673886 349812
rect 676030 349800 676036 349812
rect 676088 349800 676094 349852
rect 673454 347896 673460 347948
rect 673512 347936 673518 347948
rect 675846 347936 675852 347948
rect 673512 347908 675852 347936
rect 673512 347896 673518 347908
rect 675846 347896 675852 347908
rect 675904 347896 675910 347948
rect 673730 347828 673736 347880
rect 673788 347868 673794 347880
rect 675938 347868 675944 347880
rect 673788 347840 675944 347868
rect 673788 347828 673794 347840
rect 675938 347828 675944 347840
rect 675996 347828 676002 347880
rect 674466 347760 674472 347812
rect 674524 347800 674530 347812
rect 676030 347800 676036 347812
rect 674524 347772 676036 347800
rect 674524 347760 674530 347772
rect 676030 347760 676036 347772
rect 676088 347760 676094 347812
rect 672718 347216 672724 347268
rect 672776 347256 672782 347268
rect 676030 347256 676036 347268
rect 672776 347228 676036 347256
rect 672776 347216 672782 347228
rect 676030 347216 676036 347228
rect 676088 347216 676094 347268
rect 41874 344972 41880 345024
rect 41932 345012 41938 345024
rect 44082 345012 44088 345024
rect 41932 344984 44088 345012
rect 41932 344972 41938 344984
rect 44082 344972 44088 344984
rect 44140 344972 44146 345024
rect 41506 344224 41512 344276
rect 41564 344264 41570 344276
rect 50982 344264 50988 344276
rect 41564 344236 50988 344264
rect 41564 344224 41570 344236
rect 50982 344224 50988 344236
rect 51040 344224 51046 344276
rect 41782 344088 41788 344140
rect 41840 344128 41846 344140
rect 43806 344128 43812 344140
rect 41840 344100 43812 344128
rect 41840 344088 41846 344100
rect 43806 344088 43812 344100
rect 43864 344088 43870 344140
rect 41506 343816 41512 343868
rect 41564 343856 41570 343868
rect 48498 343856 48504 343868
rect 41564 343828 48504 343856
rect 41564 343816 41570 343828
rect 48498 343816 48504 343828
rect 48556 343816 48562 343868
rect 41506 343408 41512 343460
rect 41564 343448 41570 343460
rect 46106 343448 46112 343460
rect 41564 343420 46112 343448
rect 41564 343408 41570 343420
rect 46106 343408 46112 343420
rect 46164 343408 46170 343460
rect 41506 342592 41512 342644
rect 41564 342632 41570 342644
rect 43898 342632 43904 342644
rect 41564 342604 43904 342632
rect 41564 342592 41570 342604
rect 43898 342592 43904 342604
rect 43956 342592 43962 342644
rect 673270 342524 673276 342576
rect 673328 342564 673334 342576
rect 673546 342564 673552 342576
rect 673328 342536 673552 342564
rect 673328 342524 673334 342536
rect 673546 342524 673552 342536
rect 673604 342524 673610 342576
rect 673454 342456 673460 342508
rect 673512 342456 673518 342508
rect 673472 342304 673500 342456
rect 673454 342252 673460 342304
rect 673512 342252 673518 342304
rect 673638 342252 673644 342304
rect 673696 342292 673702 342304
rect 674558 342292 674564 342304
rect 673696 342264 674564 342292
rect 673696 342252 673702 342264
rect 674558 342252 674564 342264
rect 674616 342252 674622 342304
rect 41506 341844 41512 341896
rect 41564 341884 41570 341896
rect 43622 341884 43628 341896
rect 41564 341856 43628 341884
rect 41564 341844 41570 341856
rect 43622 341844 43628 341856
rect 43680 341844 43686 341896
rect 41506 341436 41512 341488
rect 41564 341476 41570 341488
rect 43714 341476 43720 341488
rect 41564 341448 43720 341476
rect 41564 341436 41570 341448
rect 43714 341436 43720 341448
rect 43772 341436 43778 341488
rect 674558 341436 674564 341488
rect 674616 341476 674622 341488
rect 675754 341476 675760 341488
rect 674616 341448 675760 341476
rect 674616 341436 674622 341448
rect 675754 341436 675760 341448
rect 675812 341436 675818 341488
rect 41782 341368 41788 341420
rect 41840 341408 41846 341420
rect 43530 341408 43536 341420
rect 41840 341380 43536 341408
rect 41840 341368 41846 341380
rect 43530 341368 43536 341380
rect 43588 341368 43594 341420
rect 675110 341368 675116 341420
rect 675168 341408 675174 341420
rect 675386 341408 675392 341420
rect 675168 341380 675392 341408
rect 675168 341368 675174 341380
rect 675386 341368 675392 341380
rect 675444 341368 675450 341420
rect 674926 340960 674932 341012
rect 674984 341000 674990 341012
rect 675478 341000 675484 341012
rect 674984 340972 675484 341000
rect 674984 340960 674990 340972
rect 675478 340960 675484 340972
rect 675536 340960 675542 341012
rect 675018 340892 675024 340944
rect 675076 340892 675082 340944
rect 675036 340672 675064 340892
rect 675018 340620 675024 340672
rect 675076 340620 675082 340672
rect 675110 340620 675116 340672
rect 675168 340660 675174 340672
rect 675386 340660 675392 340672
rect 675168 340632 675392 340660
rect 675168 340620 675174 340632
rect 675386 340620 675392 340632
rect 675444 340620 675450 340672
rect 675018 340212 675024 340264
rect 675076 340252 675082 340264
rect 675386 340252 675392 340264
rect 675076 340224 675392 340252
rect 675076 340212 675082 340224
rect 675386 340212 675392 340224
rect 675444 340212 675450 340264
rect 673270 340076 673276 340128
rect 673328 340116 673334 340128
rect 675018 340116 675024 340128
rect 673328 340088 675024 340116
rect 673328 340076 673334 340088
rect 675018 340076 675024 340088
rect 675076 340076 675082 340128
rect 674650 339532 674656 339584
rect 674708 339572 674714 339584
rect 675478 339572 675484 339584
rect 674708 339544 675484 339572
rect 674708 339532 674714 339544
rect 675478 339532 675484 339544
rect 675536 339532 675542 339584
rect 41782 339464 41788 339516
rect 41840 339504 41846 339516
rect 43346 339504 43352 339516
rect 41840 339476 43352 339504
rect 41840 339464 41846 339476
rect 43346 339464 43352 339476
rect 43404 339464 43410 339516
rect 674834 337900 674840 337952
rect 674892 337940 674898 337952
rect 675478 337940 675484 337952
rect 674892 337912 675484 337940
rect 674892 337900 674898 337912
rect 675478 337900 675484 337912
rect 675536 337900 675542 337952
rect 674742 337084 674748 337136
rect 674800 337124 674806 337136
rect 675386 337124 675392 337136
rect 674800 337096 675392 337124
rect 674800 337084 674806 337096
rect 675386 337084 675392 337096
rect 675444 337084 675450 337136
rect 674282 336540 674288 336592
rect 674340 336580 674346 336592
rect 675386 336580 675392 336592
rect 674340 336552 675392 336580
rect 674340 336540 674346 336552
rect 675386 336540 675392 336552
rect 675444 336540 675450 336592
rect 674466 336064 674472 336116
rect 674524 336104 674530 336116
rect 675478 336104 675484 336116
rect 674524 336076 675484 336104
rect 674524 336064 674530 336076
rect 675478 336064 675484 336076
rect 675536 336064 675542 336116
rect 655974 335316 655980 335368
rect 656032 335356 656038 335368
rect 675110 335356 675116 335368
rect 656032 335328 675116 335356
rect 656032 335316 656038 335328
rect 675110 335316 675116 335328
rect 675168 335316 675174 335368
rect 673638 333548 673644 333600
rect 673696 333588 673702 333600
rect 675386 333588 675392 333600
rect 673696 333560 675392 333588
rect 673696 333548 673702 333560
rect 675386 333548 675392 333560
rect 675444 333548 675450 333600
rect 41874 333072 41880 333124
rect 41932 333112 41938 333124
rect 48590 333112 48596 333124
rect 41932 333084 48596 333112
rect 41932 333072 41938 333084
rect 48590 333072 48596 333084
rect 48648 333072 48654 333124
rect 673730 332732 673736 332784
rect 673788 332772 673794 332784
rect 675386 332772 675392 332784
rect 673788 332744 675392 332772
rect 673788 332732 673794 332744
rect 675386 332732 675392 332744
rect 675444 332732 675450 332784
rect 675110 332528 675116 332580
rect 675168 332568 675174 332580
rect 675294 332568 675300 332580
rect 675168 332540 675300 332568
rect 675168 332528 675174 332540
rect 675294 332528 675300 332540
rect 675352 332528 675358 332580
rect 674558 332392 674564 332444
rect 674616 332432 674622 332444
rect 675294 332432 675300 332444
rect 674616 332404 675300 332432
rect 674616 332392 674622 332404
rect 675294 332392 675300 332404
rect 675352 332392 675358 332444
rect 673822 332188 673828 332240
rect 673880 332228 673886 332240
rect 675386 332228 675392 332240
rect 673880 332200 675392 332228
rect 673880 332188 673886 332200
rect 675386 332188 675392 332200
rect 675444 332188 675450 332240
rect 673454 331576 673460 331628
rect 673512 331616 673518 331628
rect 675386 331616 675392 331628
rect 673512 331588 675392 331616
rect 673512 331576 673518 331588
rect 675386 331576 675392 331588
rect 675444 331576 675450 331628
rect 41506 331168 41512 331220
rect 41564 331208 41570 331220
rect 42702 331208 42708 331220
rect 41564 331180 42708 331208
rect 41564 331168 41570 331180
rect 42702 331168 42708 331180
rect 42760 331168 42766 331220
rect 41414 331100 41420 331152
rect 41472 331140 41478 331152
rect 43162 331140 43168 331152
rect 41472 331112 43168 331140
rect 41472 331100 41478 331112
rect 43162 331100 43168 331112
rect 43220 331100 43226 331152
rect 41690 330896 41696 330948
rect 41748 330936 41754 330948
rect 43438 330936 43444 330948
rect 41748 330908 43444 330936
rect 41748 330896 41754 330908
rect 43438 330896 43444 330908
rect 43496 330896 43502 330948
rect 675018 330556 675024 330608
rect 675076 330596 675082 330608
rect 675386 330596 675392 330608
rect 675076 330568 675392 330596
rect 675076 330556 675082 330568
rect 675386 330556 675392 330568
rect 675444 330556 675450 330608
rect 30282 330284 30288 330336
rect 30340 330324 30346 330336
rect 42242 330324 42248 330336
rect 30340 330296 42248 330324
rect 30340 330284 30346 330296
rect 42242 330284 42248 330296
rect 42300 330284 42306 330336
rect 33042 330216 33048 330268
rect 33100 330256 33106 330268
rect 42334 330256 42340 330268
rect 33100 330228 42340 330256
rect 33100 330216 33106 330228
rect 42334 330216 42340 330228
rect 42392 330216 42398 330268
rect 30190 330012 30196 330064
rect 30248 330052 30254 330064
rect 43622 330052 43628 330064
rect 30248 330024 43628 330052
rect 30248 330012 30254 330024
rect 43622 330012 43628 330024
rect 43680 330012 43686 330064
rect 41782 329400 41788 329452
rect 41840 329440 41846 329452
rect 43254 329440 43260 329452
rect 41840 329412 43260 329440
rect 41840 329400 41846 329412
rect 43254 329400 43260 329412
rect 43312 329400 43318 329452
rect 41598 329332 41604 329384
rect 41656 329372 41662 329384
rect 43070 329372 43076 329384
rect 41656 329344 43076 329372
rect 41656 329332 41662 329344
rect 43070 329332 43076 329344
rect 43128 329332 43134 329384
rect 674926 328720 674932 328772
rect 674984 328760 674990 328772
rect 675386 328760 675392 328772
rect 674984 328732 675392 328760
rect 674984 328720 674990 328732
rect 675386 328720 675392 328732
rect 675444 328720 675450 328772
rect 673546 326884 673552 326936
rect 673604 326924 673610 326936
rect 675386 326924 675392 326936
rect 673604 326896 675392 326924
rect 673604 326884 673610 326896
rect 675386 326884 675392 326896
rect 675444 326884 675450 326936
rect 43070 323184 43076 323196
rect 42996 323156 43076 323184
rect 42058 323076 42064 323128
rect 42116 323116 42122 323128
rect 42702 323116 42708 323128
rect 42116 323088 42708 323116
rect 42116 323076 42122 323088
rect 42702 323076 42708 323088
rect 42760 323076 42766 323128
rect 42702 322940 42708 322992
rect 42760 322980 42766 322992
rect 42996 322980 43024 323156
rect 43070 323144 43076 323156
rect 43128 323144 43134 323196
rect 42760 322952 43024 322980
rect 42760 322940 42766 322952
rect 42242 321988 42248 322040
rect 42300 322028 42306 322040
rect 43254 322028 43260 322040
rect 42300 322000 43260 322028
rect 42300 321988 42306 322000
rect 43254 321988 43260 322000
rect 43312 321988 43318 322040
rect 42242 321784 42248 321836
rect 42300 321824 42306 321836
rect 43162 321824 43168 321836
rect 42300 321796 43168 321824
rect 42300 321784 42306 321796
rect 43162 321784 43168 321796
rect 43220 321784 43226 321836
rect 42150 321580 42156 321632
rect 42208 321620 42214 321632
rect 43438 321620 43444 321632
rect 42208 321592 43444 321620
rect 42208 321580 42214 321592
rect 43438 321580 43444 321592
rect 43496 321580 43502 321632
rect 42242 320560 42248 320612
rect 42300 320600 42306 320612
rect 43070 320600 43076 320612
rect 42300 320572 43076 320600
rect 42300 320560 42306 320572
rect 43070 320560 43076 320572
rect 43128 320560 43134 320612
rect 42242 319948 42248 320000
rect 42300 319988 42306 320000
rect 43622 319988 43628 320000
rect 42300 319960 43628 319988
rect 42300 319948 42306 319960
rect 43622 319948 43628 319960
rect 43680 319948 43686 320000
rect 42426 318724 42432 318776
rect 42484 318764 42490 318776
rect 42702 318764 42708 318776
rect 42484 318736 42708 318764
rect 42484 318724 42490 318736
rect 42702 318724 42708 318736
rect 42760 318724 42766 318776
rect 43254 318724 43260 318776
rect 43312 318764 43318 318776
rect 58526 318764 58532 318776
rect 43312 318736 58532 318764
rect 43312 318724 43318 318736
rect 58526 318724 58532 318736
rect 58584 318724 58590 318776
rect 42334 317364 42340 317416
rect 42392 317404 42398 317416
rect 58066 317404 58072 317416
rect 42392 317376 58072 317404
rect 42392 317364 42398 317376
rect 58066 317364 58072 317376
rect 58124 317364 58130 317416
rect 46106 314576 46112 314628
rect 46164 314616 46170 314628
rect 58526 314616 58532 314628
rect 46164 314588 58532 314616
rect 46164 314576 46170 314588
rect 58526 314576 58532 314588
rect 58584 314576 58590 314628
rect 675202 314576 675208 314628
rect 675260 314616 675266 314628
rect 676030 314616 676036 314628
rect 675260 314588 676036 314616
rect 675260 314576 675266 314588
rect 676030 314576 676036 314588
rect 676088 314576 676094 314628
rect 50982 314508 50988 314560
rect 51040 314548 51046 314560
rect 58158 314548 58164 314560
rect 51040 314520 58164 314548
rect 51040 314508 51046 314520
rect 58158 314508 58164 314520
rect 58216 314508 58222 314560
rect 655422 312060 655428 312112
rect 655480 312100 655486 312112
rect 676214 312100 676220 312112
rect 655480 312072 676220 312100
rect 655480 312060 655486 312072
rect 676214 312060 676220 312072
rect 676272 312060 676278 312112
rect 655698 311992 655704 312044
rect 655756 312032 655762 312044
rect 676306 312032 676312 312044
rect 655756 312004 676312 312032
rect 655756 311992 655762 312004
rect 676306 311992 676312 312004
rect 676364 311992 676370 312044
rect 655514 311924 655520 311976
rect 655572 311964 655578 311976
rect 676122 311964 676128 311976
rect 655572 311936 676128 311964
rect 655572 311924 655578 311936
rect 676122 311924 676128 311936
rect 676180 311924 676186 311976
rect 672994 311856 673000 311908
rect 673052 311896 673058 311908
rect 676214 311896 676220 311908
rect 673052 311868 676220 311896
rect 673052 311856 673058 311868
rect 676214 311856 676220 311868
rect 676272 311856 676278 311908
rect 48498 311788 48504 311840
rect 48556 311828 48562 311840
rect 58526 311828 58532 311840
rect 48556 311800 58532 311828
rect 48556 311788 48562 311800
rect 58526 311788 58532 311800
rect 58584 311788 58590 311840
rect 673362 311652 673368 311704
rect 673420 311692 673426 311704
rect 676030 311692 676036 311704
rect 673420 311664 676036 311692
rect 673420 311652 673426 311664
rect 676030 311652 676036 311664
rect 676088 311652 676094 311704
rect 675110 311516 675116 311568
rect 675168 311556 675174 311568
rect 676030 311556 676036 311568
rect 675168 311528 676036 311556
rect 675168 311516 675174 311528
rect 676030 311516 676036 311528
rect 676088 311516 676094 311568
rect 673270 311040 673276 311092
rect 673328 311080 673334 311092
rect 676214 311080 676220 311092
rect 673328 311052 676220 311080
rect 673328 311040 673334 311052
rect 676214 311040 676220 311052
rect 676272 311040 676278 311092
rect 673178 310224 673184 310276
rect 673236 310264 673242 310276
rect 676214 310264 676220 310276
rect 673236 310236 676220 310264
rect 673236 310224 673242 310236
rect 676214 310224 676220 310236
rect 676272 310224 676278 310276
rect 673086 309408 673092 309460
rect 673144 309448 673150 309460
rect 676214 309448 676220 309460
rect 673144 309420 676220 309448
rect 673144 309408 673150 309420
rect 676214 309408 676220 309420
rect 676272 309408 676278 309460
rect 674650 309136 674656 309188
rect 674708 309176 674714 309188
rect 676030 309176 676036 309188
rect 674708 309148 676036 309176
rect 674708 309136 674714 309148
rect 676030 309136 676036 309148
rect 676088 309136 676094 309188
rect 673546 308048 673552 308100
rect 673604 308088 673610 308100
rect 676030 308088 676036 308100
rect 673604 308060 676036 308088
rect 673604 308048 673610 308060
rect 676030 308048 676036 308060
rect 676088 308048 676094 308100
rect 674926 307232 674932 307284
rect 674984 307272 674990 307284
rect 676030 307272 676036 307284
rect 674984 307244 676036 307272
rect 674984 307232 674990 307244
rect 676030 307232 676036 307244
rect 676088 307232 676094 307284
rect 674834 306824 674840 306876
rect 674892 306864 674898 306876
rect 676030 306864 676036 306876
rect 674892 306836 676036 306864
rect 674892 306824 674898 306836
rect 676030 306824 676036 306836
rect 676088 306824 676094 306876
rect 674282 306416 674288 306468
rect 674340 306456 674346 306468
rect 676122 306456 676128 306468
rect 674340 306428 676128 306456
rect 674340 306416 674346 306428
rect 676122 306416 676128 306428
rect 676180 306416 676186 306468
rect 675018 306348 675024 306400
rect 675076 306388 675082 306400
rect 676030 306388 676036 306400
rect 675076 306360 676036 306388
rect 675076 306348 675082 306360
rect 676030 306348 676036 306360
rect 676088 306348 676094 306400
rect 42058 306280 42064 306332
rect 42116 306320 42122 306332
rect 58342 306320 58348 306332
rect 42116 306292 58348 306320
rect 42116 306280 42122 306292
rect 58342 306280 58348 306292
rect 58400 306280 58406 306332
rect 673822 305056 673828 305108
rect 673880 305096 673886 305108
rect 676122 305096 676128 305108
rect 673880 305068 676128 305096
rect 673880 305056 673886 305068
rect 676122 305056 676128 305068
rect 676180 305056 676186 305108
rect 675110 304784 675116 304836
rect 675168 304824 675174 304836
rect 676030 304824 676036 304836
rect 675168 304796 676036 304824
rect 675168 304784 675174 304796
rect 676030 304784 676036 304796
rect 676088 304784 676094 304836
rect 673730 304308 673736 304360
rect 673788 304348 673794 304360
rect 676122 304348 676128 304360
rect 673788 304320 676128 304348
rect 673788 304308 673794 304320
rect 676122 304308 676128 304320
rect 676180 304308 676186 304360
rect 675202 304172 675208 304224
rect 675260 304212 675266 304224
rect 676030 304212 676036 304224
rect 675260 304184 676036 304212
rect 675260 304172 675266 304184
rect 676030 304172 676036 304184
rect 676088 304172 676094 304224
rect 674466 303900 674472 303952
rect 674524 303940 674530 303952
rect 676122 303940 676128 303952
rect 674524 303912 676128 303940
rect 674524 303900 674530 303912
rect 676122 303900 676128 303912
rect 676180 303900 676186 303952
rect 673638 303696 673644 303748
rect 673696 303736 673702 303748
rect 676030 303736 676036 303748
rect 673696 303708 676036 303736
rect 673696 303696 673702 303708
rect 676030 303696 676036 303708
rect 676088 303696 676094 303748
rect 672810 300840 672816 300892
rect 672868 300880 672874 300892
rect 678974 300880 678980 300892
rect 672868 300852 678980 300880
rect 672868 300840 672874 300852
rect 678974 300840 678980 300852
rect 679032 300840 679038 300892
rect 674834 300160 674840 300212
rect 674892 300160 674898 300212
rect 41782 300092 41788 300144
rect 41840 300132 41846 300144
rect 43898 300132 43904 300144
rect 41840 300104 43904 300132
rect 41840 300092 41846 300104
rect 43898 300092 43904 300104
rect 43956 300092 43962 300144
rect 674852 300008 674880 300160
rect 675018 300024 675024 300076
rect 675076 300024 675082 300076
rect 41782 299956 41788 300008
rect 41840 299996 41846 300008
rect 43530 299996 43536 300008
rect 41840 299968 43536 299996
rect 41840 299956 41846 299968
rect 43530 299956 43536 299968
rect 43588 299956 43594 300008
rect 674834 299956 674840 300008
rect 674892 299956 674898 300008
rect 675036 299872 675064 300024
rect 675018 299820 675024 299872
rect 675076 299820 675082 299872
rect 42058 299344 42064 299396
rect 42116 299384 42122 299396
rect 43254 299384 43260 299396
rect 42116 299356 43260 299384
rect 42116 299344 42122 299356
rect 43254 299344 43260 299356
rect 43312 299344 43318 299396
rect 41782 299072 41788 299124
rect 41840 299112 41846 299124
rect 43346 299112 43352 299124
rect 41840 299084 43352 299112
rect 41840 299072 41846 299084
rect 43346 299072 43352 299084
rect 43404 299072 43410 299124
rect 655054 298120 655060 298172
rect 655112 298160 655118 298172
rect 675386 298160 675392 298172
rect 655112 298132 675392 298160
rect 655112 298120 655118 298132
rect 675386 298120 675392 298132
rect 675444 298120 675450 298172
rect 41782 297304 41788 297356
rect 41840 297344 41846 297356
rect 43622 297344 43628 297356
rect 41840 297316 43628 297344
rect 41840 297304 41846 297316
rect 43622 297304 43628 297316
rect 43680 297304 43686 297356
rect 41782 296216 41788 296268
rect 41840 296256 41846 296268
rect 43806 296256 43812 296268
rect 41840 296228 43812 296256
rect 41840 296216 41846 296228
rect 43806 296216 43812 296228
rect 43864 296216 43870 296268
rect 675018 295400 675024 295452
rect 675076 295440 675082 295452
rect 675294 295440 675300 295452
rect 675076 295412 675300 295440
rect 675076 295400 675082 295412
rect 675294 295400 675300 295412
rect 675352 295400 675358 295452
rect 42334 295332 42340 295384
rect 42392 295372 42398 295384
rect 58526 295372 58532 295384
rect 42392 295344 58532 295372
rect 42392 295332 42398 295344
rect 58526 295332 58532 295344
rect 58584 295332 58590 295384
rect 674742 294720 674748 294772
rect 674800 294760 674806 294772
rect 675294 294760 675300 294772
rect 674800 294732 675300 294760
rect 674800 294720 674806 294732
rect 675294 294720 675300 294732
rect 675352 294720 675358 294772
rect 674650 294516 674656 294568
rect 674708 294556 674714 294568
rect 675386 294556 675392 294568
rect 674708 294528 675392 294556
rect 674708 294516 674714 294528
rect 675386 294516 675392 294528
rect 675444 294516 675450 294568
rect 42058 293632 42064 293684
rect 42116 293672 42122 293684
rect 43990 293672 43996 293684
rect 42116 293644 43996 293672
rect 42116 293632 42122 293644
rect 43990 293632 43996 293644
rect 44048 293632 44054 293684
rect 42058 293428 42064 293480
rect 42116 293468 42122 293480
rect 44082 293468 44088 293480
rect 42116 293440 44088 293468
rect 42116 293428 42122 293440
rect 44082 293428 44088 293440
rect 44140 293428 44146 293480
rect 43530 292612 43536 292664
rect 43588 292652 43594 292664
rect 58434 292652 58440 292664
rect 43588 292624 58440 292652
rect 43588 292612 43594 292624
rect 58434 292612 58440 292624
rect 58492 292612 58498 292664
rect 41966 292476 41972 292528
rect 42024 292516 42030 292528
rect 57974 292516 57980 292528
rect 42024 292488 57980 292516
rect 42024 292476 42030 292488
rect 57974 292476 57980 292488
rect 58032 292476 58038 292528
rect 41874 292408 41880 292460
rect 41932 292448 41938 292460
rect 58526 292448 58532 292460
rect 41932 292420 58532 292448
rect 41932 292408 41938 292420
rect 58526 292408 58532 292420
rect 58584 292408 58590 292460
rect 41874 292272 41880 292324
rect 41932 292312 41938 292324
rect 43070 292312 43076 292324
rect 41932 292284 43076 292312
rect 41932 292272 41938 292284
rect 43070 292272 43076 292284
rect 43128 292272 43134 292324
rect 674926 291524 674932 291576
rect 674984 291564 674990 291576
rect 675386 291564 675392 291576
rect 674984 291536 675392 291564
rect 674984 291524 674990 291536
rect 675386 291524 675392 291536
rect 675444 291524 675450 291576
rect 41782 291048 41788 291100
rect 41840 291088 41846 291100
rect 51074 291088 51080 291100
rect 41840 291060 51080 291088
rect 41840 291048 41846 291060
rect 51074 291048 51080 291060
rect 51132 291048 51138 291100
rect 41782 290640 41788 290692
rect 41840 290680 41846 290692
rect 51166 290680 51172 290692
rect 41840 290652 51172 290680
rect 41840 290640 41846 290652
rect 51166 290640 51172 290652
rect 51224 290640 51230 290692
rect 674466 290436 674472 290488
rect 674524 290476 674530 290488
rect 675110 290476 675116 290488
rect 674524 290448 675116 290476
rect 674524 290436 674530 290448
rect 675110 290436 675116 290448
rect 675168 290436 675174 290488
rect 41782 289824 41788 289876
rect 41840 289864 41846 289876
rect 48774 289864 48780 289876
rect 41840 289836 48780 289864
rect 41840 289824 41846 289836
rect 48774 289824 48780 289836
rect 48832 289824 48838 289876
rect 27522 289756 27528 289808
rect 27580 289796 27586 289808
rect 57974 289796 57980 289808
rect 27580 289768 57980 289796
rect 27580 289756 27586 289768
rect 57974 289756 57980 289768
rect 58032 289756 58038 289808
rect 674282 288600 674288 288652
rect 674340 288640 674346 288652
rect 675386 288640 675392 288652
rect 674340 288612 675392 288640
rect 674340 288600 674346 288612
rect 675386 288600 675392 288612
rect 675444 288600 675450 288652
rect 654502 288532 654508 288584
rect 654560 288572 654566 288584
rect 666830 288572 666836 288584
rect 654560 288544 666836 288572
rect 654560 288532 654566 288544
rect 666830 288532 666836 288544
rect 666888 288532 666894 288584
rect 673730 287376 673736 287428
rect 673788 287416 673794 287428
rect 675110 287416 675116 287428
rect 673788 287388 675116 287416
rect 673788 287376 673794 287388
rect 675110 287376 675116 287388
rect 675168 287376 675174 287428
rect 48682 287104 48688 287156
rect 48740 287144 48746 287156
rect 58158 287144 58164 287156
rect 48740 287116 58164 287144
rect 48740 287104 48746 287116
rect 58158 287104 58164 287116
rect 58216 287104 58222 287156
rect 656802 287104 656808 287156
rect 656860 287144 656866 287156
rect 669406 287144 669412 287156
rect 656860 287116 669412 287144
rect 656860 287104 656866 287116
rect 669406 287104 669412 287116
rect 669464 287104 669470 287156
rect 46290 287036 46296 287088
rect 46348 287076 46354 287088
rect 58526 287076 58532 287088
rect 46348 287048 58532 287076
rect 46348 287036 46354 287048
rect 58526 287036 58532 287048
rect 58584 287036 58590 287088
rect 654870 287036 654876 287088
rect 654928 287076 654934 287088
rect 669498 287076 669504 287088
rect 654928 287048 669504 287076
rect 654928 287036 654934 287048
rect 669498 287036 669504 287048
rect 669556 287036 669562 287088
rect 35802 286968 35808 287020
rect 35860 287008 35866 287020
rect 42242 287008 42248 287020
rect 35860 286980 42248 287008
rect 35860 286968 35866 286980
rect 42242 286968 42248 286980
rect 42300 286968 42306 287020
rect 42150 286900 42156 286952
rect 42208 286940 42214 286952
rect 43438 286940 43444 286952
rect 42208 286912 43444 286940
rect 42208 286900 42214 286912
rect 43438 286900 43444 286912
rect 43496 286900 43502 286952
rect 41966 286832 41972 286884
rect 42024 286872 42030 286884
rect 43346 286872 43352 286884
rect 42024 286844 43352 286872
rect 42024 286832 42030 286844
rect 43346 286832 43352 286844
rect 43404 286832 43410 286884
rect 673822 286764 673828 286816
rect 673880 286804 673886 286816
rect 675110 286804 675116 286816
rect 673880 286776 675116 286804
rect 673880 286764 673886 286776
rect 675110 286764 675116 286776
rect 675168 286764 675174 286816
rect 673638 286560 673644 286612
rect 673696 286600 673702 286612
rect 675386 286600 675392 286612
rect 673696 286572 675392 286600
rect 673696 286560 673702 286572
rect 675386 286560 675392 286572
rect 675444 286560 675450 286612
rect 42058 286152 42064 286204
rect 42116 286192 42122 286204
rect 43162 286192 43168 286204
rect 42116 286164 43168 286192
rect 42116 286152 42122 286164
rect 43162 286152 43168 286164
rect 43220 286152 43226 286204
rect 41690 285744 41696 285796
rect 41748 285784 41754 285796
rect 43806 285784 43812 285796
rect 41748 285756 43812 285784
rect 41748 285744 41754 285756
rect 43806 285744 43812 285756
rect 43864 285744 43870 285796
rect 42426 285608 42432 285660
rect 42484 285648 42490 285660
rect 43714 285648 43720 285660
rect 42484 285620 43720 285648
rect 42484 285608 42490 285620
rect 43714 285608 43720 285620
rect 43772 285608 43778 285660
rect 655422 284928 655428 284980
rect 655480 284968 655486 284980
rect 669590 284968 669596 284980
rect 655480 284940 669596 284968
rect 655480 284928 655486 284940
rect 669590 284928 669596 284940
rect 669648 284928 669654 284980
rect 56502 284792 56508 284844
rect 56560 284832 56566 284844
rect 57974 284832 57980 284844
rect 56560 284804 57980 284832
rect 56560 284792 56566 284804
rect 57974 284792 57980 284804
rect 58032 284792 58038 284844
rect 654870 284656 654876 284708
rect 654928 284696 654934 284708
rect 666738 284696 666744 284708
rect 654928 284668 666744 284696
rect 654928 284656 654934 284668
rect 666738 284656 666744 284668
rect 666796 284656 666802 284708
rect 51258 284316 51264 284368
rect 51316 284356 51322 284368
rect 58526 284356 58532 284368
rect 51316 284328 58532 284356
rect 51316 284316 51322 284328
rect 58526 284316 58532 284328
rect 58584 284316 58590 284368
rect 43990 284248 43996 284300
rect 44048 284288 44054 284300
rect 44266 284288 44272 284300
rect 44048 284260 44272 284288
rect 44048 284248 44054 284260
rect 44266 284248 44272 284260
rect 44324 284248 44330 284300
rect 43070 284112 43076 284164
rect 43128 284152 43134 284164
rect 43990 284152 43996 284164
rect 43128 284124 43996 284152
rect 43128 284112 43134 284124
rect 43990 284112 43996 284124
rect 44048 284112 44054 284164
rect 41874 283772 41880 283824
rect 41932 283772 41938 283824
rect 41892 283620 41920 283772
rect 673546 283704 673552 283756
rect 673604 283744 673610 283756
rect 675478 283744 675484 283756
rect 673604 283716 675484 283744
rect 673604 283704 673610 283716
rect 675478 283704 675484 283716
rect 675536 283704 675542 283756
rect 41874 283568 41880 283620
rect 41932 283568 41938 283620
rect 43070 281596 43076 281648
rect 43128 281636 43134 281648
rect 44266 281636 44272 281648
rect 43128 281608 44272 281636
rect 43128 281596 43134 281608
rect 44266 281596 44272 281608
rect 44324 281596 44330 281648
rect 50982 281596 50988 281648
rect 51040 281636 51046 281648
rect 58250 281636 58256 281648
rect 51040 281608 58256 281636
rect 51040 281596 51046 281608
rect 58250 281596 58256 281608
rect 58308 281596 58314 281648
rect 656802 281596 656808 281648
rect 656860 281636 656866 281648
rect 669222 281636 669228 281648
rect 656860 281608 669228 281636
rect 656860 281596 656866 281608
rect 669222 281596 669228 281608
rect 669280 281596 669286 281648
rect 48498 281528 48504 281580
rect 48556 281568 48562 281580
rect 58526 281568 58532 281580
rect 48556 281540 58532 281568
rect 48556 281528 48562 281540
rect 58526 281528 58532 281540
rect 58584 281528 58590 281580
rect 42334 280440 42340 280492
rect 42392 280480 42398 280492
rect 43346 280480 43352 280492
rect 42392 280452 43352 280480
rect 42392 280440 42398 280452
rect 43346 280440 43352 280452
rect 43404 280440 43410 280492
rect 42242 280372 42248 280424
rect 42300 280412 42306 280424
rect 43530 280412 43536 280424
rect 42300 280384 43536 280412
rect 42300 280372 42306 280384
rect 43530 280372 43536 280384
rect 43588 280372 43594 280424
rect 654686 280168 654692 280220
rect 654744 280208 654750 280220
rect 669314 280208 669320 280220
rect 654744 280180 669320 280208
rect 654744 280168 654750 280180
rect 669314 280168 669320 280180
rect 669372 280168 669378 280220
rect 42150 279828 42156 279880
rect 42208 279868 42214 279880
rect 43162 279868 43168 279880
rect 42208 279840 43168 279868
rect 42208 279828 42214 279840
rect 43162 279828 43168 279840
rect 43220 279828 43226 279880
rect 654870 278944 654876 278996
rect 654928 278984 654934 278996
rect 666646 278984 666652 278996
rect 654928 278956 666652 278984
rect 654928 278944 654934 278956
rect 666646 278944 666652 278956
rect 666704 278944 666710 278996
rect 46198 278808 46204 278860
rect 46256 278848 46262 278860
rect 58158 278848 58164 278860
rect 46256 278820 58164 278848
rect 46256 278808 46262 278820
rect 58158 278808 58164 278820
rect 58216 278808 58222 278860
rect 46106 278740 46112 278792
rect 46164 278780 46170 278792
rect 58250 278780 58256 278792
rect 46164 278752 58256 278780
rect 46164 278740 46170 278752
rect 58250 278740 58256 278752
rect 58308 278740 58314 278792
rect 42058 278400 42064 278452
rect 42116 278440 42122 278452
rect 42702 278440 42708 278452
rect 42116 278412 42708 278440
rect 42116 278400 42122 278412
rect 42702 278400 42708 278412
rect 42760 278400 42766 278452
rect 42150 277856 42156 277908
rect 42208 277896 42214 277908
rect 43438 277896 43444 277908
rect 42208 277868 43444 277896
rect 42208 277856 42214 277868
rect 43438 277856 43444 277868
rect 43496 277856 43502 277908
rect 45646 277312 45652 277364
rect 45704 277352 45710 277364
rect 666554 277352 666560 277364
rect 45704 277324 666560 277352
rect 45704 277312 45710 277324
rect 666554 277312 666560 277324
rect 666612 277312 666618 277364
rect 42334 276768 42340 276820
rect 42392 276808 42398 276820
rect 43806 276808 43812 276820
rect 42392 276780 43812 276808
rect 42392 276768 42398 276780
rect 43806 276768 43812 276780
rect 43864 276768 43870 276820
rect 342530 275952 342536 276004
rect 342588 275992 342594 276004
rect 464154 275992 464160 276004
rect 342588 275964 464160 275992
rect 342588 275952 342594 275964
rect 464154 275952 464160 275964
rect 464212 275952 464218 276004
rect 345106 275884 345112 275936
rect 345164 275924 345170 275936
rect 471238 275924 471244 275936
rect 345164 275896 471244 275924
rect 345164 275884 345170 275896
rect 471238 275884 471244 275896
rect 471296 275884 471302 275936
rect 347774 275816 347780 275868
rect 347832 275856 347838 275868
rect 478322 275856 478328 275868
rect 347832 275828 478328 275856
rect 347832 275816 347838 275828
rect 478322 275816 478328 275828
rect 478380 275816 478386 275868
rect 346394 275748 346400 275800
rect 346452 275788 346458 275800
rect 474826 275788 474832 275800
rect 346452 275760 474832 275788
rect 346452 275748 346458 275760
rect 474826 275748 474832 275760
rect 474884 275748 474890 275800
rect 351638 275680 351644 275732
rect 351696 275720 351702 275732
rect 488994 275720 489000 275732
rect 351696 275692 489000 275720
rect 351696 275680 351702 275692
rect 488994 275680 489000 275692
rect 489052 275680 489058 275732
rect 353202 275612 353208 275664
rect 353260 275652 353266 275664
rect 492582 275652 492588 275664
rect 353260 275624 492588 275652
rect 353260 275612 353266 275624
rect 492582 275612 492588 275624
rect 492640 275612 492646 275664
rect 42426 275544 42432 275596
rect 42484 275584 42490 275596
rect 43990 275584 43996 275596
rect 42484 275556 43996 275584
rect 42484 275544 42490 275556
rect 43990 275544 43996 275556
rect 44048 275544 44054 275596
rect 357066 275544 357072 275596
rect 357124 275584 357130 275596
rect 503162 275584 503168 275596
rect 357124 275556 503168 275584
rect 357124 275544 357130 275556
rect 503162 275544 503168 275556
rect 503220 275544 503226 275596
rect 358446 275476 358452 275528
rect 358504 275516 358510 275528
rect 506750 275516 506756 275528
rect 358504 275488 506756 275516
rect 358504 275476 358510 275488
rect 506750 275476 506756 275488
rect 506808 275476 506814 275528
rect 361114 275408 361120 275460
rect 361172 275448 361178 275460
rect 513834 275448 513840 275460
rect 361172 275420 513840 275448
rect 361172 275408 361178 275420
rect 513834 275408 513840 275420
rect 513892 275408 513898 275460
rect 363782 275340 363788 275392
rect 363840 275380 363846 275392
rect 520918 275380 520924 275392
rect 363840 275352 520924 275380
rect 363840 275340 363846 275352
rect 520918 275340 520924 275352
rect 520976 275340 520982 275392
rect 366450 275272 366456 275324
rect 366508 275312 366514 275324
rect 528002 275312 528008 275324
rect 366508 275284 528008 275312
rect 366508 275272 366514 275284
rect 528002 275272 528008 275284
rect 528060 275272 528066 275324
rect 371786 275204 371792 275256
rect 371844 275244 371850 275256
rect 371844 275216 390600 275244
rect 371844 275204 371850 275216
rect 375282 275136 375288 275188
rect 375340 275176 375346 275188
rect 390572 275176 390600 275216
rect 390646 275204 390652 275256
rect 390704 275244 390710 275256
rect 535086 275244 535092 275256
rect 390704 275216 535092 275244
rect 390704 275204 390710 275216
rect 535086 275204 535092 275216
rect 535144 275204 535150 275256
rect 542170 275176 542176 275188
rect 375340 275148 390508 275176
rect 390572 275148 542176 275176
rect 375340 275136 375346 275148
rect 377766 275068 377772 275120
rect 377824 275108 377830 275120
rect 390480 275108 390508 275148
rect 542170 275136 542176 275148
rect 542228 275136 542234 275188
rect 550450 275108 550456 275120
rect 377824 275080 390416 275108
rect 390480 275080 550456 275108
rect 377824 275068 377830 275080
rect 390388 275040 390416 275080
rect 550450 275068 550456 275080
rect 550508 275068 550514 275120
rect 557534 275040 557540 275052
rect 390388 275012 557540 275040
rect 557534 275000 557540 275012
rect 557592 275000 557598 275052
rect 380342 274932 380348 274984
rect 380400 274972 380406 274984
rect 564618 274972 564624 274984
rect 380400 274944 564624 274972
rect 380400 274932 380406 274944
rect 564618 274932 564624 274944
rect 564676 274932 564682 274984
rect 383286 274864 383292 274916
rect 383344 274904 383350 274916
rect 571702 274904 571708 274916
rect 383344 274876 571708 274904
rect 383344 274864 383350 274876
rect 571702 274864 571708 274876
rect 571760 274864 571766 274916
rect 317506 274796 317512 274848
rect 317564 274836 317570 274848
rect 398006 274836 398012 274848
rect 317564 274808 398012 274836
rect 317564 274796 317570 274808
rect 398006 274796 398012 274808
rect 398064 274796 398070 274848
rect 610710 274836 610716 274848
rect 400186 274808 610716 274836
rect 320174 274728 320180 274780
rect 320232 274768 320238 274780
rect 390462 274768 390468 274780
rect 320232 274740 390468 274768
rect 320232 274728 320238 274740
rect 390462 274728 390468 274740
rect 390520 274728 390526 274780
rect 397638 274728 397644 274780
rect 397696 274768 397702 274780
rect 400186 274768 400214 274808
rect 610710 274796 610716 274808
rect 610768 274796 610774 274848
rect 397696 274740 400214 274768
rect 397696 274728 397702 274740
rect 402974 274728 402980 274780
rect 403032 274768 403038 274780
rect 624970 274768 624976 274780
rect 403032 274740 624976 274768
rect 403032 274728 403038 274740
rect 624970 274728 624976 274740
rect 625028 274728 625034 274780
rect 321002 274660 321008 274712
rect 321060 274700 321066 274712
rect 407482 274700 407488 274712
rect 321060 274672 407488 274700
rect 321060 274660 321066 274672
rect 407482 274660 407488 274672
rect 407540 274660 407546 274712
rect 409230 274660 409236 274712
rect 409288 274700 409294 274712
rect 409288 274672 419534 274700
rect 409288 274660 409294 274672
rect 322566 274592 322572 274644
rect 322624 274632 322630 274644
rect 410978 274632 410984 274644
rect 322624 274604 410984 274632
rect 322624 274592 322630 274604
rect 410978 274592 410984 274604
rect 411036 274592 411042 274644
rect 419506 274632 419534 274672
rect 429102 274660 429108 274712
rect 429160 274700 429166 274712
rect 634354 274700 634360 274712
rect 429160 274672 634360 274700
rect 429160 274660 429166 274672
rect 634354 274660 634360 274672
rect 634412 274660 634418 274712
rect 641438 274632 641444 274644
rect 419506 274604 641444 274632
rect 641438 274592 641444 274604
rect 641496 274592 641502 274644
rect 341058 274524 341064 274576
rect 341116 274564 341122 274576
rect 460658 274564 460664 274576
rect 341116 274536 460664 274564
rect 341116 274524 341122 274536
rect 460658 274524 460664 274536
rect 460716 274524 460722 274576
rect 338390 274456 338396 274508
rect 338448 274496 338454 274508
rect 453574 274496 453580 274508
rect 338448 274468 453580 274496
rect 338448 274456 338454 274468
rect 453574 274456 453580 274468
rect 453632 274456 453638 274508
rect 337102 274388 337108 274440
rect 337160 274428 337166 274440
rect 449986 274428 449992 274440
rect 337160 274400 449992 274428
rect 337160 274388 337166 274400
rect 449986 274388 449992 274400
rect 450044 274388 450050 274440
rect 336090 274320 336096 274372
rect 336148 274360 336154 274372
rect 446490 274360 446496 274372
rect 336148 274332 446496 274360
rect 336148 274320 336154 274332
rect 446490 274320 446496 274332
rect 446548 274320 446554 274372
rect 334342 274252 334348 274304
rect 334400 274292 334406 274304
rect 334400 274264 351868 274292
rect 334400 274252 334406 274264
rect 351840 274224 351868 274264
rect 351914 274252 351920 274304
rect 351972 274292 351978 274304
rect 439314 274292 439320 274304
rect 351972 274264 439320 274292
rect 351972 274252 351978 274264
rect 439314 274252 439320 274264
rect 439372 274252 439378 274304
rect 351840 274196 429148 274224
rect 333054 274116 333060 274168
rect 333112 274156 333118 274168
rect 351730 274156 351736 274168
rect 333112 274128 351736 274156
rect 333112 274116 333118 274128
rect 351730 274116 351736 274128
rect 351788 274116 351794 274168
rect 351822 274116 351828 274168
rect 351880 274156 351886 274168
rect 429120 274156 429148 274196
rect 442902 274156 442908 274168
rect 351880 274128 426480 274156
rect 429120 274128 442908 274156
rect 351880 274116 351886 274128
rect 330386 274048 330392 274100
rect 330444 274088 330450 274100
rect 426452 274088 426480 274128
rect 442902 274116 442908 274128
rect 442960 274116 442966 274168
rect 433426 274088 433432 274100
rect 330444 274060 425928 274088
rect 426452 274060 433432 274088
rect 330444 274048 330450 274060
rect 331674 273980 331680 274032
rect 331732 274020 331738 274032
rect 425900 274020 425928 274060
rect 433426 274048 433432 274060
rect 433484 274048 433490 274100
rect 432230 274020 432236 274032
rect 331732 273992 425836 274020
rect 425900 273992 432236 274020
rect 331732 273980 331738 273992
rect 327718 273912 327724 273964
rect 327776 273952 327782 273964
rect 425146 273952 425152 273964
rect 327776 273924 425152 273952
rect 327776 273912 327782 273924
rect 425146 273912 425152 273924
rect 425204 273912 425210 273964
rect 425808 273952 425836 273992
rect 432230 273980 432236 273992
rect 432288 273980 432294 274032
rect 435818 273952 435824 273964
rect 425808 273924 435824 273952
rect 435818 273912 435824 273924
rect 435876 273912 435882 273964
rect 329006 273844 329012 273896
rect 329064 273884 329070 273896
rect 428734 273884 428740 273896
rect 329064 273856 428740 273884
rect 329064 273844 329070 273856
rect 428734 273844 428740 273856
rect 428792 273844 428798 273896
rect 325050 273776 325056 273828
rect 325108 273816 325114 273828
rect 418062 273816 418068 273828
rect 325108 273788 418068 273816
rect 325108 273776 325114 273788
rect 418062 273776 418068 273788
rect 418120 273776 418126 273828
rect 42426 273708 42432 273760
rect 42484 273748 42490 273760
rect 44082 273748 44088 273760
rect 42484 273720 44088 273748
rect 42484 273708 42490 273720
rect 44082 273708 44088 273720
rect 44140 273708 44146 273760
rect 325510 273708 325516 273760
rect 325568 273748 325574 273760
rect 419258 273748 419264 273760
rect 325568 273720 419264 273748
rect 325568 273708 325574 273720
rect 419258 273708 419264 273720
rect 419316 273708 419322 273760
rect 326338 273640 326344 273692
rect 326396 273680 326402 273692
rect 421650 273680 421656 273692
rect 326396 273652 421656 273680
rect 326396 273640 326402 273652
rect 421650 273640 421656 273652
rect 421708 273640 421714 273692
rect 323670 273572 323676 273624
rect 323728 273612 323734 273624
rect 414566 273612 414572 273624
rect 323728 273584 414572 273612
rect 323728 273572 323734 273584
rect 414566 273572 414572 273584
rect 414624 273572 414630 273624
rect 330846 273504 330852 273556
rect 330904 273544 330910 273556
rect 351822 273544 351828 273556
rect 330904 273516 351828 273544
rect 330904 273504 330910 273516
rect 351822 273504 351828 273516
rect 351880 273504 351886 273556
rect 390462 273504 390468 273556
rect 390520 273544 390526 273556
rect 405090 273544 405096 273556
rect 390520 273516 405096 273544
rect 390520 273504 390526 273516
rect 405090 273504 405096 273516
rect 405148 273504 405154 273556
rect 406562 273504 406568 273556
rect 406620 273544 406626 273556
rect 429102 273544 429108 273556
rect 406620 273516 429108 273544
rect 406620 273504 406626 273516
rect 429102 273504 429108 273516
rect 429160 273504 429166 273556
rect 369118 273436 369124 273488
rect 369176 273476 369182 273488
rect 390646 273476 390652 273488
rect 369176 273448 390652 273476
rect 369176 273436 369182 273448
rect 390646 273436 390652 273448
rect 390704 273436 390710 273488
rect 154482 273164 154488 273216
rect 154540 273204 154546 273216
rect 211062 273204 211068 273216
rect 154540 273176 211068 273204
rect 154540 273164 154546 273176
rect 211062 273164 211068 273176
rect 211120 273164 211126 273216
rect 224494 273204 224500 273216
rect 211172 273176 224500 273204
rect 42426 273096 42432 273148
rect 42484 273136 42490 273148
rect 43070 273136 43076 273148
rect 42484 273108 43076 273136
rect 42484 273096 42490 273108
rect 43070 273096 43076 273108
rect 43128 273096 43134 273148
rect 176838 273096 176844 273148
rect 176896 273136 176902 273148
rect 210970 273136 210976 273148
rect 176896 273108 210976 273136
rect 176896 273096 176902 273108
rect 210970 273096 210976 273108
rect 211028 273096 211034 273148
rect 152182 273028 152188 273080
rect 152240 273068 152246 273080
rect 211172 273068 211200 273176
rect 224494 273164 224500 273176
rect 224552 273164 224558 273216
rect 263226 273164 263232 273216
rect 263284 273204 263290 273216
rect 266722 273204 266728 273216
rect 263284 273176 266728 273204
rect 263284 273164 263290 273176
rect 266722 273164 266728 273176
rect 266780 273164 266786 273216
rect 292114 273164 292120 273216
rect 292172 273204 292178 273216
rect 330570 273204 330576 273216
rect 292172 273176 330576 273204
rect 292172 273164 292178 273176
rect 330570 273164 330576 273176
rect 330628 273164 330634 273216
rect 352650 273164 352656 273216
rect 352708 273204 352714 273216
rect 491386 273204 491392 273216
rect 352708 273176 491392 273204
rect 352708 273164 352714 273176
rect 491386 273164 491392 273176
rect 491444 273164 491450 273216
rect 491478 273164 491484 273216
rect 491536 273204 491542 273216
rect 507946 273204 507952 273216
rect 491536 273176 507952 273204
rect 491536 273164 491542 273176
rect 507946 273164 507952 273176
rect 508004 273164 508010 273216
rect 260926 273096 260932 273148
rect 260984 273136 260990 273148
rect 265802 273136 265808 273148
rect 260984 273108 265808 273136
rect 260984 273096 260990 273108
rect 265802 273096 265808 273108
rect 265860 273096 265866 273148
rect 293862 273096 293868 273148
rect 293920 273136 293926 273148
rect 335354 273136 335360 273148
rect 293920 273108 335360 273136
rect 293920 273096 293926 273108
rect 335354 273096 335360 273108
rect 335412 273096 335418 273148
rect 344922 273096 344928 273148
rect 344980 273136 344986 273148
rect 470134 273136 470140 273148
rect 344980 273108 470140 273136
rect 344980 273096 344986 273108
rect 470134 273096 470140 273108
rect 470192 273096 470198 273148
rect 471974 273096 471980 273148
rect 472032 273136 472038 273148
rect 614298 273136 614304 273148
rect 472032 273108 614304 273136
rect 472032 273096 472038 273108
rect 614298 273096 614304 273108
rect 614356 273096 614362 273148
rect 152240 273040 211200 273068
rect 152240 273028 152246 273040
rect 211246 273028 211252 273080
rect 211304 273068 211310 273080
rect 217962 273068 217968 273080
rect 211304 273040 217968 273068
rect 211304 273028 211310 273040
rect 217962 273028 217968 273040
rect 218020 273028 218026 273080
rect 243170 273028 243176 273080
rect 243228 273068 243234 273080
rect 259178 273068 259184 273080
rect 243228 273040 259184 273068
rect 243228 273028 243234 273040
rect 259178 273028 259184 273040
rect 259236 273028 259242 273080
rect 259730 273028 259736 273080
rect 259788 273068 259794 273080
rect 265434 273068 265440 273080
rect 259788 273040 265440 273068
rect 259788 273028 259794 273040
rect 265434 273028 265440 273040
rect 265492 273028 265498 273080
rect 296070 273028 296076 273080
rect 296128 273068 296134 273080
rect 341242 273068 341248 273080
rect 296128 273040 341248 273068
rect 296128 273028 296134 273040
rect 341242 273028 341248 273040
rect 341300 273028 341306 273080
rect 356054 273028 356060 273080
rect 356112 273068 356118 273080
rect 358814 273068 358820 273080
rect 356112 273040 358820 273068
rect 356112 273028 356118 273040
rect 358814 273028 358820 273040
rect 358872 273028 358878 273080
rect 358906 273028 358912 273080
rect 358964 273068 358970 273080
rect 497274 273068 497280 273080
rect 358964 273040 497280 273068
rect 358964 273028 358970 273040
rect 497274 273028 497280 273040
rect 497332 273028 497338 273080
rect 497918 273028 497924 273080
rect 497976 273068 497982 273080
rect 600130 273068 600136 273080
rect 497976 273040 600136 273068
rect 497976 273028 497982 273040
rect 600130 273028 600136 273040
rect 600188 273028 600194 273080
rect 147398 272960 147404 273012
rect 147456 273000 147462 273012
rect 222654 273000 222660 273012
rect 147456 272972 222660 273000
rect 147456 272960 147462 272972
rect 222654 272960 222660 272972
rect 222712 272960 222718 273012
rect 240778 272960 240784 273012
rect 240836 273000 240842 273012
rect 258258 273000 258264 273012
rect 240836 272972 258264 273000
rect 240836 272960 240842 272972
rect 258258 272960 258264 272972
rect 258316 272960 258322 273012
rect 301866 272960 301872 273012
rect 301924 273000 301930 273012
rect 356606 273000 356612 273012
rect 301924 272972 356612 273000
rect 301924 272960 301930 272972
rect 356606 272960 356612 272972
rect 356664 272960 356670 273012
rect 360562 272960 360568 273012
rect 360620 273000 360626 273012
rect 511442 273000 511448 273012
rect 360620 272972 511448 273000
rect 360620 272960 360626 272972
rect 511442 272960 511448 272972
rect 511500 272960 511506 273012
rect 149790 272892 149796 272944
rect 149848 272932 149854 272944
rect 214742 272932 214748 272944
rect 149848 272904 214748 272932
rect 149848 272892 149854 272904
rect 214742 272892 214748 272904
rect 214800 272892 214806 272944
rect 214834 272892 214840 272944
rect 214892 272932 214898 272944
rect 220446 272932 220452 272944
rect 214892 272904 220452 272932
rect 214892 272892 214898 272904
rect 220446 272892 220452 272904
rect 220504 272892 220510 272944
rect 234890 272892 234896 272944
rect 234948 272932 234954 272944
rect 256050 272932 256056 272944
rect 234948 272904 256056 272932
rect 234948 272892 234954 272904
rect 256050 272892 256056 272904
rect 256108 272892 256114 272944
rect 303522 272892 303528 272944
rect 303580 272932 303586 272944
rect 360194 272932 360200 272944
rect 303580 272904 360200 272932
rect 303580 272892 303586 272904
rect 360194 272892 360200 272904
rect 360252 272892 360258 272944
rect 363138 272892 363144 272944
rect 363196 272932 363202 272944
rect 518526 272932 518532 272944
rect 363196 272904 518532 272932
rect 363196 272892 363202 272904
rect 518526 272892 518532 272904
rect 518584 272892 518590 272944
rect 146202 272824 146208 272876
rect 146260 272864 146266 272876
rect 223022 272864 223028 272876
rect 146260 272836 223028 272864
rect 146260 272824 146266 272836
rect 223022 272824 223028 272836
rect 223080 272824 223086 272876
rect 233694 272824 233700 272876
rect 233752 272864 233758 272876
rect 255590 272864 255596 272876
rect 233752 272836 255596 272864
rect 233752 272824 233758 272836
rect 255590 272824 255596 272836
rect 255648 272824 255654 272876
rect 294874 272824 294880 272876
rect 294932 272864 294938 272876
rect 337746 272864 337752 272876
rect 294932 272836 337752 272864
rect 294932 272824 294938 272836
rect 337746 272824 337752 272836
rect 337804 272824 337810 272876
rect 347498 272824 347504 272876
rect 347556 272864 347562 272876
rect 477218 272864 477224 272876
rect 347556 272836 477224 272864
rect 347556 272824 347562 272836
rect 477218 272824 477224 272836
rect 477276 272824 477282 272876
rect 477310 272824 477316 272876
rect 477368 272864 477374 272876
rect 632054 272864 632060 272876
rect 477368 272836 632060 272864
rect 477368 272824 477374 272836
rect 632054 272824 632060 272836
rect 632112 272824 632118 272876
rect 139118 272756 139124 272808
rect 139176 272796 139182 272808
rect 220354 272796 220360 272808
rect 139176 272768 220360 272796
rect 139176 272756 139182 272768
rect 220354 272756 220360 272768
rect 220412 272756 220418 272808
rect 236086 272756 236092 272808
rect 236144 272796 236150 272808
rect 256418 272796 256424 272808
rect 236144 272768 256424 272796
rect 236144 272756 236150 272768
rect 256418 272756 256424 272768
rect 256476 272756 256482 272808
rect 295058 272756 295064 272808
rect 295116 272796 295122 272808
rect 338850 272796 338856 272808
rect 295116 272768 338856 272796
rect 295116 272756 295122 272768
rect 338850 272756 338856 272768
rect 338908 272756 338914 272808
rect 342162 272756 342168 272808
rect 342220 272796 342226 272808
rect 462958 272796 462964 272808
rect 342220 272768 462964 272796
rect 342220 272756 342226 272768
rect 462958 272756 462964 272768
rect 463016 272756 463022 272808
rect 463326 272756 463332 272808
rect 463384 272796 463390 272808
rect 621382 272796 621388 272808
rect 463384 272768 621388 272796
rect 463384 272756 463390 272768
rect 621382 272756 621388 272768
rect 621440 272756 621446 272808
rect 141510 272688 141516 272740
rect 141568 272728 141574 272740
rect 221182 272728 221188 272740
rect 141568 272700 221188 272728
rect 141568 272688 141574 272700
rect 221182 272688 221188 272700
rect 221240 272688 221246 272740
rect 232498 272688 232504 272740
rect 232556 272728 232562 272740
rect 255130 272728 255136 272740
rect 232556 272700 255136 272728
rect 232556 272688 232562 272700
rect 255130 272688 255136 272700
rect 255188 272688 255194 272740
rect 324222 272688 324228 272740
rect 324280 272728 324286 272740
rect 362494 272728 362500 272740
rect 324280 272700 362500 272728
rect 324280 272688 324286 272700
rect 362494 272688 362500 272700
rect 362552 272688 362558 272740
rect 362586 272688 362592 272740
rect 362644 272728 362650 272740
rect 370774 272728 370780 272740
rect 362644 272700 370780 272728
rect 362644 272688 362650 272700
rect 370774 272688 370780 272700
rect 370832 272688 370838 272740
rect 375650 272688 375656 272740
rect 375708 272728 375714 272740
rect 381446 272728 381452 272740
rect 375708 272700 381452 272728
rect 375708 272688 375714 272700
rect 381446 272688 381452 272700
rect 381504 272688 381510 272740
rect 391934 272688 391940 272740
rect 391992 272728 391998 272740
rect 555234 272728 555240 272740
rect 391992 272700 555240 272728
rect 391992 272688 391998 272700
rect 555234 272688 555240 272700
rect 555292 272688 555298 272740
rect 119062 272620 119068 272672
rect 119120 272660 119126 272672
rect 119120 272632 137600 272660
rect 119120 272620 119126 272632
rect 126146 272552 126152 272604
rect 126204 272592 126210 272604
rect 137572 272592 137600 272632
rect 140314 272620 140320 272672
rect 140372 272660 140378 272672
rect 219986 272660 219992 272672
rect 140372 272632 219992 272660
rect 140372 272620 140378 272632
rect 219986 272620 219992 272632
rect 220044 272620 220050 272672
rect 306742 272620 306748 272672
rect 306800 272660 306806 272672
rect 369578 272660 369584 272672
rect 306800 272632 369584 272660
rect 306800 272620 306806 272632
rect 369578 272620 369584 272632
rect 369636 272620 369642 272672
rect 369670 272620 369676 272672
rect 369728 272660 369734 272672
rect 532694 272660 532700 272672
rect 369728 272632 532700 272660
rect 369728 272620 369734 272632
rect 532694 272620 532700 272632
rect 532752 272620 532758 272672
rect 126204 272564 129734 272592
rect 137572 272564 193352 272592
rect 126204 272552 126210 272564
rect 129706 272524 129734 272564
rect 187694 272524 187700 272536
rect 129706 272496 187700 272524
rect 187694 272484 187700 272496
rect 187752 272484 187758 272536
rect 89530 272416 89536 272468
rect 89588 272456 89594 272468
rect 177114 272456 177120 272468
rect 89588 272428 177120 272456
rect 89588 272416 89594 272428
rect 177114 272416 177120 272428
rect 177172 272416 177178 272468
rect 193324 272456 193352 272564
rect 193490 272552 193496 272604
rect 193548 272592 193554 272604
rect 203610 272592 203616 272604
rect 193548 272564 203616 272592
rect 193548 272552 193554 272564
rect 203610 272552 203616 272564
rect 203668 272552 203674 272604
rect 214742 272552 214748 272604
rect 214800 272592 214806 272604
rect 224402 272592 224408 272604
rect 214800 272564 224408 272592
rect 214800 272552 214806 272564
rect 224402 272552 224408 272564
rect 224460 272552 224466 272604
rect 293402 272552 293408 272604
rect 293460 272592 293466 272604
rect 334158 272592 334164 272604
rect 293460 272564 334164 272592
rect 293460 272552 293466 272564
rect 334158 272552 334164 272564
rect 334216 272552 334222 272604
rect 336642 272552 336648 272604
rect 336700 272592 336706 272604
rect 448790 272592 448796 272604
rect 336700 272564 448796 272592
rect 336700 272552 336706 272564
rect 448790 272552 448796 272564
rect 448848 272552 448854 272604
rect 448882 272552 448888 272604
rect 448940 272592 448946 272604
rect 628466 272592 628472 272604
rect 448940 272564 628472 272592
rect 448940 272552 448946 272564
rect 628466 272552 628472 272564
rect 628524 272552 628530 272604
rect 197262 272484 197268 272536
rect 197320 272524 197326 272536
rect 197320 272496 207014 272524
rect 197320 272484 197326 272496
rect 206830 272456 206836 272468
rect 193324 272428 206836 272456
rect 206830 272416 206836 272428
rect 206888 272416 206894 272468
rect 206986 272456 207014 272496
rect 211062 272484 211068 272536
rect 211120 272524 211126 272536
rect 225322 272524 225328 272536
rect 211120 272496 225328 272524
rect 211120 272484 211126 272496
rect 225322 272484 225328 272496
rect 225380 272484 225386 272536
rect 229002 272484 229008 272536
rect 229060 272524 229066 272536
rect 253750 272524 253756 272536
rect 229060 272496 253756 272524
rect 229060 272484 229066 272496
rect 253750 272484 253756 272496
rect 253808 272484 253814 272536
rect 307202 272484 307208 272536
rect 307260 272524 307266 272536
rect 307260 272496 322244 272524
rect 307260 272484 307266 272496
rect 232038 272456 232044 272468
rect 206986 272428 232044 272456
rect 232038 272416 232044 272428
rect 232096 272416 232102 272468
rect 237282 272416 237288 272468
rect 237340 272456 237346 272468
rect 256878 272456 256884 272468
rect 237340 272428 256884 272456
rect 237340 272416 237346 272428
rect 256878 272416 256884 272428
rect 256936 272416 256942 272468
rect 306282 272416 306288 272468
rect 306340 272456 306346 272468
rect 322216 272456 322244 272496
rect 322290 272484 322296 272536
rect 322348 272524 322354 272536
rect 367278 272524 367284 272536
rect 322348 272496 367284 272524
rect 322348 272484 322354 272496
rect 367278 272484 367284 272496
rect 367336 272484 367342 272536
rect 379330 272484 379336 272536
rect 379388 272524 379394 272536
rect 562318 272524 562324 272536
rect 379388 272496 562324 272524
rect 379388 272484 379394 272496
rect 562318 272484 562324 272496
rect 562376 272484 562382 272536
rect 362586 272456 362592 272468
rect 306340 272428 320128 272456
rect 322216 272428 362592 272456
rect 306340 272416 306346 272428
rect 111978 272348 111984 272400
rect 112036 272388 112042 272400
rect 201586 272388 201592 272400
rect 112036 272360 201592 272388
rect 112036 272348 112042 272360
rect 201586 272348 201592 272360
rect 201644 272348 201650 272400
rect 288158 272348 288164 272400
rect 288216 272388 288222 272400
rect 319990 272388 319996 272400
rect 288216 272360 319996 272388
rect 288216 272348 288222 272360
rect 319990 272348 319996 272360
rect 320048 272348 320054 272400
rect 320100 272388 320128 272428
rect 362586 272416 362592 272428
rect 362644 272416 362650 272468
rect 362862 272416 362868 272468
rect 362920 272456 362926 272468
rect 384942 272456 384948 272468
rect 362920 272428 384948 272456
rect 362920 272416 362926 272428
rect 384942 272416 384948 272428
rect 385000 272416 385006 272468
rect 386414 272416 386420 272468
rect 386472 272456 386478 272468
rect 569402 272456 569408 272468
rect 386472 272428 569408 272456
rect 386472 272416 386478 272428
rect 569402 272416 569408 272428
rect 569460 272416 569466 272468
rect 322290 272388 322296 272400
rect 320100 272360 322296 272388
rect 322290 272348 322296 272360
rect 322348 272348 322354 272400
rect 322842 272348 322848 272400
rect 322900 272388 322906 272400
rect 383838 272388 383844 272400
rect 322900 272360 383844 272388
rect 322900 272348 322906 272360
rect 383838 272348 383844 272360
rect 383896 272348 383902 272400
rect 384666 272348 384672 272400
rect 384724 272388 384730 272400
rect 576486 272388 576492 272400
rect 384724 272360 576492 272388
rect 384724 272348 384730 272360
rect 576486 272348 576492 272360
rect 576544 272348 576550 272400
rect 117866 272280 117872 272332
rect 117924 272320 117930 272332
rect 117924 272292 201632 272320
rect 117924 272280 117930 272292
rect 88334 272212 88340 272264
rect 88392 272252 88398 272264
rect 184934 272252 184940 272264
rect 88392 272224 184940 272252
rect 88392 272212 88398 272224
rect 184934 272212 184940 272224
rect 184992 272212 184998 272264
rect 185210 272212 185216 272264
rect 185268 272252 185274 272264
rect 197262 272252 197268 272264
rect 185268 272224 197268 272252
rect 185268 272212 185274 272224
rect 197262 272212 197268 272224
rect 197320 272212 197326 272264
rect 102502 272144 102508 272196
rect 102560 272184 102566 272196
rect 201494 272184 201500 272196
rect 102560 272156 201500 272184
rect 102560 272144 102566 272156
rect 201494 272144 201500 272156
rect 201552 272144 201558 272196
rect 201604 272184 201632 272292
rect 210970 272280 210976 272332
rect 211028 272320 211034 272332
rect 227070 272320 227076 272332
rect 211028 272292 227076 272320
rect 211028 272280 211034 272292
rect 227070 272280 227076 272292
rect 227128 272280 227134 272332
rect 230198 272280 230204 272332
rect 230256 272320 230262 272332
rect 254210 272320 254216 272332
rect 230256 272292 254216 272320
rect 230256 272280 230262 272292
rect 254210 272280 254216 272292
rect 254268 272280 254274 272332
rect 309318 272320 309324 272332
rect 284266 272292 309324 272320
rect 284266 272264 284294 272292
rect 309318 272280 309324 272292
rect 309376 272280 309382 272332
rect 309870 272280 309876 272332
rect 309928 272320 309934 272332
rect 377858 272320 377864 272332
rect 309928 272292 377864 272320
rect 309928 272280 309934 272292
rect 377858 272280 377864 272292
rect 377916 272280 377922 272332
rect 390002 272280 390008 272332
rect 390060 272320 390066 272332
rect 590654 272320 590660 272332
rect 390060 272292 590660 272320
rect 390060 272280 390066 272292
rect 590654 272280 590660 272292
rect 590712 272280 590718 272332
rect 209682 272252 209688 272264
rect 201788 272224 209688 272252
rect 201788 272184 201816 272224
rect 209682 272212 209688 272224
rect 209740 272212 209746 272264
rect 238478 272212 238484 272264
rect 238536 272252 238542 272264
rect 257246 272252 257252 272264
rect 238536 272224 257252 272252
rect 238536 272212 238542 272224
rect 257246 272212 257252 272224
rect 257304 272212 257310 272264
rect 284202 272212 284208 272264
rect 284260 272224 284294 272264
rect 284260 272212 284266 272224
rect 292574 272212 292580 272264
rect 292632 272252 292638 272264
rect 331766 272252 331772 272264
rect 292632 272224 331772 272252
rect 292632 272212 292638 272224
rect 331766 272212 331772 272224
rect 331824 272212 331830 272264
rect 434622 272252 434628 272264
rect 331876 272224 434628 272252
rect 201604 272156 201816 272184
rect 205358 272144 205364 272196
rect 205416 272184 205422 272196
rect 244918 272184 244924 272196
rect 205416 272156 244924 272184
rect 205416 272144 205422 272156
rect 244918 272144 244924 272156
rect 244976 272144 244982 272196
rect 285858 272144 285864 272196
rect 285916 272184 285922 272196
rect 314102 272184 314108 272196
rect 285916 272156 314108 272184
rect 285916 272144 285922 272156
rect 314102 272144 314108 272156
rect 314160 272144 314166 272196
rect 331306 272144 331312 272196
rect 331364 272184 331370 272196
rect 331876 272184 331904 272224
rect 434622 272212 434628 272224
rect 434680 272212 434686 272264
rect 436094 272212 436100 272264
rect 436152 272252 436158 272264
rect 639138 272252 639144 272264
rect 436152 272224 639144 272252
rect 436152 272212 436158 272224
rect 639138 272212 639144 272224
rect 639196 272212 639202 272264
rect 362862 272184 362868 272196
rect 331364 272156 331904 272184
rect 331968 272156 362868 272184
rect 331364 272144 331370 272156
rect 97810 272076 97816 272128
rect 97868 272116 97874 272128
rect 198826 272116 198832 272128
rect 97868 272088 198832 272116
rect 97868 272076 97874 272088
rect 198826 272076 198832 272088
rect 198884 272076 198890 272128
rect 204162 272076 204168 272128
rect 204220 272116 204226 272128
rect 240134 272116 240140 272128
rect 204220 272088 240140 272116
rect 204220 272076 204226 272088
rect 240134 272076 240140 272088
rect 240192 272076 240198 272128
rect 288526 272076 288532 272128
rect 288584 272116 288590 272128
rect 321186 272116 321192 272128
rect 288584 272088 321192 272116
rect 288584 272076 288590 272088
rect 321186 272076 321192 272088
rect 321244 272076 321250 272128
rect 331968 272116 331996 272156
rect 362862 272144 362868 272156
rect 362920 272144 362926 272196
rect 367094 272144 367100 272196
rect 367152 272184 367158 272196
rect 387334 272184 387340 272196
rect 367152 272156 387340 272184
rect 367152 272144 367158 272156
rect 387334 272144 387340 272156
rect 387392 272144 387398 272196
rect 392762 272144 392768 272196
rect 392820 272184 392826 272196
rect 597738 272184 597744 272196
rect 392820 272156 597744 272184
rect 392820 272144 392826 272156
rect 597738 272144 597744 272156
rect 597796 272144 597802 272196
rect 324332 272088 331996 272116
rect 96614 272008 96620 272060
rect 96672 272048 96678 272060
rect 198734 272048 198740 272060
rect 96672 272020 198740 272048
rect 96672 272008 96678 272020
rect 198734 272008 198740 272020
rect 198792 272008 198798 272060
rect 202966 272008 202972 272060
rect 203024 272048 203030 272060
rect 243998 272048 244004 272060
rect 203024 272020 244004 272048
rect 203024 272008 203030 272020
rect 243998 272008 244004 272020
rect 244056 272008 244062 272060
rect 286686 272008 286692 272060
rect 286744 272048 286750 272060
rect 316402 272048 316408 272060
rect 286744 272020 316408 272048
rect 286744 272008 286750 272020
rect 316402 272008 316408 272020
rect 316460 272008 316466 272060
rect 317322 272008 317328 272060
rect 317380 272048 317386 272060
rect 324332 272048 324360 272088
rect 332318 272076 332324 272128
rect 332376 272116 332382 272128
rect 390922 272116 390928 272128
rect 332376 272088 390928 272116
rect 332376 272076 332382 272088
rect 390922 272076 390928 272088
rect 390980 272076 390986 272128
rect 398098 272076 398104 272128
rect 398156 272116 398162 272128
rect 611906 272116 611912 272128
rect 398156 272088 611912 272116
rect 398156 272076 398162 272088
rect 611906 272076 611912 272088
rect 611964 272076 611970 272128
rect 317380 272020 324360 272048
rect 317380 272008 317386 272020
rect 332226 272008 332232 272060
rect 332284 272048 332290 272060
rect 392118 272048 392124 272060
rect 332284 272020 392124 272048
rect 332284 272008 332290 272020
rect 392118 272008 392124 272020
rect 392176 272008 392182 272060
rect 406102 272008 406108 272060
rect 406160 272048 406166 272060
rect 406160 272020 413784 272048
rect 406160 272008 406166 272020
rect 77662 271940 77668 271992
rect 77720 271980 77726 271992
rect 193214 271980 193220 271992
rect 77720 271952 193220 271980
rect 77720 271940 77726 271952
rect 193214 271940 193220 271952
rect 193272 271940 193278 271992
rect 198274 271940 198280 271992
rect 198332 271980 198338 271992
rect 242250 271980 242256 271992
rect 198332 271952 242256 271980
rect 198332 271940 198338 271952
rect 242250 271940 242256 271952
rect 242308 271940 242314 271992
rect 244366 271940 244372 271992
rect 244424 271980 244430 271992
rect 259546 271980 259552 271992
rect 244424 271952 259552 271980
rect 244424 271940 244430 271952
rect 259546 271940 259552 271952
rect 259604 271940 259610 271992
rect 262122 271940 262128 271992
rect 262180 271980 262186 271992
rect 266262 271980 266268 271992
rect 262180 271952 266268 271980
rect 262180 271940 262186 271952
rect 266262 271940 266268 271952
rect 266320 271940 266326 271992
rect 286594 271940 286600 271992
rect 286652 271980 286658 271992
rect 315206 271980 315212 271992
rect 286652 271952 315212 271980
rect 286652 271940 286658 271952
rect 315206 271940 315212 271952
rect 315264 271940 315270 271992
rect 320542 271940 320548 271992
rect 320600 271980 320606 271992
rect 320600 271952 322612 271980
rect 320600 271940 320606 271952
rect 156874 271872 156880 271924
rect 156932 271912 156938 271924
rect 176838 271912 176844 271924
rect 156932 271884 176844 271912
rect 156932 271872 156938 271884
rect 176838 271872 176844 271884
rect 176896 271872 176902 271924
rect 176930 271872 176936 271924
rect 176988 271912 176994 271924
rect 193122 271912 193128 271924
rect 176988 271884 193128 271912
rect 176988 271872 176994 271884
rect 193122 271872 193128 271884
rect 193180 271872 193186 271924
rect 194686 271872 194692 271924
rect 194744 271912 194750 271924
rect 240870 271912 240876 271924
rect 194744 271884 240876 271912
rect 194744 271872 194750 271884
rect 240870 271872 240876 271884
rect 240928 271872 240934 271924
rect 289170 271872 289176 271924
rect 289228 271912 289234 271924
rect 322382 271912 322388 271924
rect 289228 271884 322388 271912
rect 289228 271872 289234 271884
rect 322382 271872 322388 271884
rect 322440 271872 322446 271924
rect 322584 271912 322612 271952
rect 332134 271940 332140 271992
rect 332192 271980 332198 271992
rect 399202 271980 399208 271992
rect 332192 271952 399208 271980
rect 332192 271940 332198 271952
rect 399202 271940 399208 271952
rect 399260 271940 399266 271992
rect 409598 271940 409604 271992
rect 409656 271980 409662 271992
rect 413756 271980 413784 272020
rect 413830 272008 413836 272060
rect 413888 272048 413894 272060
rect 618990 272048 618996 272060
rect 413888 272020 618996 272048
rect 413888 272008 413894 272020
rect 618990 272008 618996 272020
rect 619048 272008 619054 272060
rect 633250 271980 633256 271992
rect 409656 271952 413692 271980
rect 413756 271952 633256 271980
rect 409656 271940 409662 271952
rect 406286 271912 406292 271924
rect 322584 271884 406292 271912
rect 406286 271872 406292 271884
rect 406344 271872 406350 271924
rect 411438 271872 411444 271924
rect 411496 271912 411502 271924
rect 413664 271912 413692 271952
rect 633250 271940 633256 271952
rect 633308 271940 633314 271992
rect 642634 271912 642640 271924
rect 411496 271884 413508 271912
rect 413664 271884 642640 271912
rect 411496 271872 411502 271884
rect 42426 271804 42432 271856
rect 42484 271844 42490 271856
rect 59262 271844 59268 271856
rect 42484 271816 59268 271844
rect 42484 271804 42490 271816
rect 59262 271804 59268 271816
rect 59320 271804 59326 271856
rect 67082 271804 67088 271856
rect 67140 271844 67146 271856
rect 67140 271816 190132 271844
rect 67140 271804 67146 271816
rect 127342 271736 127348 271788
rect 127400 271776 127406 271788
rect 189902 271776 189908 271788
rect 127400 271748 189908 271776
rect 127400 271736 127406 271748
rect 189902 271736 189908 271748
rect 189960 271736 189966 271788
rect 190104 271776 190132 271816
rect 191190 271804 191196 271856
rect 191248 271844 191254 271856
rect 239490 271844 239496 271856
rect 191248 271816 239496 271844
rect 191248 271804 191254 271816
rect 239490 271804 239496 271816
rect 239548 271804 239554 271856
rect 247862 271804 247868 271856
rect 247920 271844 247926 271856
rect 260926 271844 260932 271856
rect 247920 271816 260932 271844
rect 247920 271804 247926 271816
rect 260926 271804 260932 271816
rect 260984 271804 260990 271856
rect 264422 271804 264428 271856
rect 264480 271844 264486 271856
rect 267182 271844 267188 271856
rect 264480 271816 267188 271844
rect 264480 271804 264486 271816
rect 267182 271804 267188 271816
rect 267240 271804 267246 271856
rect 289630 271804 289636 271856
rect 289688 271844 289694 271856
rect 323486 271844 323492 271856
rect 289688 271816 323492 271844
rect 289688 271804 289694 271816
rect 323486 271804 323492 271816
rect 323544 271804 323550 271856
rect 323578 271804 323584 271856
rect 323636 271844 323642 271856
rect 413370 271844 413376 271856
rect 323636 271816 413376 271844
rect 323636 271804 323642 271816
rect 413370 271804 413376 271816
rect 413428 271804 413434 271856
rect 413480 271844 413508 271884
rect 642634 271872 642640 271884
rect 642692 271872 642698 271924
rect 647418 271844 647424 271856
rect 413480 271816 647424 271844
rect 647418 271804 647424 271816
rect 647476 271804 647482 271856
rect 192478 271776 192484 271788
rect 190104 271748 192484 271776
rect 192478 271736 192484 271748
rect 192536 271736 192542 271788
rect 200574 271736 200580 271788
rect 200632 271776 200638 271788
rect 243262 271776 243268 271788
rect 200632 271748 243268 271776
rect 200632 271736 200638 271748
rect 243262 271736 243268 271748
rect 243320 271736 243326 271788
rect 249058 271736 249064 271788
rect 249116 271776 249122 271788
rect 261386 271776 261392 271788
rect 249116 271748 261392 271776
rect 249116 271736 249122 271748
rect 261386 271736 261392 271748
rect 261444 271736 261450 271788
rect 292022 271736 292028 271788
rect 292080 271776 292086 271788
rect 329466 271776 329472 271788
rect 292080 271748 329472 271776
rect 292080 271736 292086 271748
rect 329466 271736 329472 271748
rect 329524 271736 329530 271788
rect 352190 271736 352196 271788
rect 352248 271776 352254 271788
rect 490190 271776 490196 271788
rect 352248 271748 490196 271776
rect 352248 271736 352254 271748
rect 490190 271736 490196 271748
rect 490248 271736 490254 271788
rect 159266 271668 159272 271720
rect 159324 271708 159330 271720
rect 227530 271708 227536 271720
rect 159324 271680 227536 271708
rect 159324 271668 159330 271680
rect 227530 271668 227536 271680
rect 227588 271668 227594 271720
rect 239582 271668 239588 271720
rect 239640 271708 239646 271720
rect 239640 271680 251404 271708
rect 239640 271668 239646 271680
rect 163958 271600 163964 271652
rect 164016 271640 164022 271652
rect 229738 271640 229744 271652
rect 164016 271612 229744 271640
rect 164016 271600 164022 271612
rect 229738 271600 229744 271612
rect 229796 271600 229802 271652
rect 245562 271600 245568 271652
rect 245620 271640 245626 271652
rect 251174 271640 251180 271652
rect 245620 271612 251180 271640
rect 245620 271600 245626 271612
rect 251174 271600 251180 271612
rect 251232 271600 251238 271652
rect 161566 271532 161572 271584
rect 161624 271572 161630 271584
rect 227990 271572 227996 271584
rect 161624 271544 227996 271572
rect 161624 271532 161630 271544
rect 227990 271532 227996 271544
rect 228048 271532 228054 271584
rect 171042 271464 171048 271516
rect 171100 271504 171106 271516
rect 229278 271504 229284 271516
rect 171100 271476 229284 271504
rect 171100 271464 171106 271476
rect 229278 271464 229284 271476
rect 229336 271464 229342 271516
rect 241974 271464 241980 271516
rect 242032 271504 242038 271516
rect 251266 271504 251272 271516
rect 242032 271476 251272 271504
rect 242032 271464 242038 271476
rect 251266 271464 251272 271476
rect 251324 271464 251330 271516
rect 251376 271504 251404 271680
rect 251450 271668 251456 271720
rect 251508 271708 251514 271720
rect 262214 271708 262220 271720
rect 251508 271680 262220 271708
rect 251508 271668 251514 271680
rect 262214 271668 262220 271680
rect 262272 271668 262278 271720
rect 291194 271668 291200 271720
rect 291252 271708 291258 271720
rect 328270 271708 328276 271720
rect 291252 271680 328276 271708
rect 291252 271668 291258 271680
rect 328270 271668 328276 271680
rect 328328 271668 328334 271720
rect 350166 271668 350172 271720
rect 350224 271708 350230 271720
rect 484302 271708 484308 271720
rect 350224 271680 484308 271708
rect 350224 271668 350230 271680
rect 484302 271668 484308 271680
rect 484360 271668 484366 271720
rect 485682 271668 485688 271720
rect 485740 271708 485746 271720
rect 607214 271708 607220 271720
rect 485740 271680 607220 271708
rect 485740 271668 485746 271680
rect 607214 271668 607220 271680
rect 607272 271668 607278 271720
rect 253842 271600 253848 271652
rect 253900 271640 253906 271652
rect 263134 271640 263140 271652
rect 253900 271612 263140 271640
rect 253900 271600 253906 271612
rect 263134 271600 263140 271612
rect 263192 271600 263198 271652
rect 290274 271600 290280 271652
rect 290332 271640 290338 271652
rect 325878 271640 325884 271652
rect 290332 271612 325884 271640
rect 290332 271600 290338 271612
rect 325878 271600 325884 271612
rect 325936 271600 325942 271652
rect 349614 271600 349620 271652
rect 349672 271640 349678 271652
rect 483106 271640 483112 271652
rect 349672 271612 483112 271640
rect 349672 271600 349678 271612
rect 483106 271600 483112 271612
rect 483164 271600 483170 271652
rect 257338 271532 257344 271584
rect 257396 271572 257402 271584
rect 264514 271572 264520 271584
rect 257396 271544 264520 271572
rect 257396 271532 257402 271544
rect 264514 271532 264520 271544
rect 264572 271532 264578 271584
rect 290734 271532 290740 271584
rect 290792 271572 290798 271584
rect 327074 271572 327080 271584
rect 290792 271544 327080 271572
rect 290792 271532 290798 271544
rect 327074 271532 327080 271544
rect 327132 271532 327138 271584
rect 346854 271532 346860 271584
rect 346912 271572 346918 271584
rect 476022 271572 476028 271584
rect 346912 271544 476028 271572
rect 346912 271532 346918 271544
rect 476022 271532 476028 271544
rect 476080 271532 476086 271584
rect 257798 271504 257804 271516
rect 251376 271476 257804 271504
rect 257798 271464 257804 271476
rect 257856 271464 257862 271516
rect 258534 271464 258540 271516
rect 258592 271504 258598 271516
rect 264882 271504 264888 271516
rect 258592 271476 264888 271504
rect 258592 271464 258598 271476
rect 264882 271464 264888 271476
rect 264940 271464 264946 271516
rect 266814 271464 266820 271516
rect 266872 271504 266878 271516
rect 268010 271504 268016 271516
rect 266872 271476 268016 271504
rect 266872 271464 266878 271476
rect 268010 271464 268016 271476
rect 268068 271464 268074 271516
rect 289814 271464 289820 271516
rect 289872 271504 289878 271516
rect 324682 271504 324688 271516
rect 289872 271476 324688 271504
rect 289872 271464 289878 271476
rect 324682 271464 324688 271476
rect 324740 271464 324746 271516
rect 344186 271464 344192 271516
rect 344244 271504 344250 271516
rect 468938 271504 468944 271516
rect 344244 271476 468944 271504
rect 344244 271464 344250 271476
rect 468938 271464 468944 271476
rect 468996 271464 469002 271516
rect 168742 271396 168748 271448
rect 168800 271436 168806 271448
rect 230382 271436 230388 271448
rect 168800 271408 230388 271436
rect 168800 271396 168806 271408
rect 230382 271396 230388 271408
rect 230440 271396 230446 271448
rect 253382 271436 253388 271448
rect 245626 271408 253388 271436
rect 166350 271328 166356 271380
rect 166408 271368 166414 271380
rect 224034 271368 224040 271380
rect 166408 271340 224040 271368
rect 166408 271328 166414 271340
rect 224034 271328 224040 271340
rect 224092 271328 224098 271380
rect 227806 271328 227812 271380
rect 227864 271368 227870 271380
rect 245626 271368 245654 271408
rect 253382 271396 253388 271408
rect 253440 271396 253446 271448
rect 254946 271396 254952 271448
rect 255004 271436 255010 271448
rect 263594 271436 263600 271448
rect 255004 271408 263600 271436
rect 255004 271396 255010 271408
rect 263594 271396 263600 271408
rect 263652 271396 263658 271448
rect 287606 271396 287612 271448
rect 287664 271436 287670 271448
rect 318794 271436 318800 271448
rect 287664 271408 318800 271436
rect 287664 271396 287670 271408
rect 318794 271396 318800 271408
rect 318852 271396 318858 271448
rect 322658 271396 322664 271448
rect 322716 271436 322722 271448
rect 332318 271436 332324 271448
rect 322716 271408 332324 271436
rect 322716 271396 322722 271408
rect 332318 271396 332324 271408
rect 332376 271396 332382 271448
rect 342070 271396 342076 271448
rect 342128 271436 342134 271448
rect 342128 271408 448468 271436
rect 342128 271396 342134 271408
rect 227864 271340 245654 271368
rect 227864 271328 227870 271340
rect 252646 271328 252652 271380
rect 252704 271368 252710 271380
rect 262858 271368 262864 271380
rect 252704 271340 262864 271368
rect 252704 271328 252710 271340
rect 262858 271328 262864 271340
rect 262916 271328 262922 271380
rect 285398 271328 285404 271380
rect 285456 271368 285462 271380
rect 312906 271368 312912 271380
rect 285456 271340 312912 271368
rect 285456 271328 285462 271340
rect 312906 271328 312912 271340
rect 312964 271328 312970 271380
rect 315206 271328 315212 271380
rect 315264 271368 315270 271380
rect 332226 271368 332232 271380
rect 315264 271340 332232 271368
rect 315264 271328 315270 271340
rect 332226 271328 332232 271340
rect 332284 271328 332290 271380
rect 339218 271328 339224 271380
rect 339276 271368 339282 271380
rect 448440 271368 448468 271408
rect 452654 271396 452660 271448
rect 452712 271436 452718 271448
rect 458266 271436 458272 271448
rect 452712 271408 458272 271436
rect 452712 271396 452718 271408
rect 458266 271396 458272 271408
rect 458324 271396 458330 271448
rect 339276 271340 447364 271368
rect 448440 271340 458174 271368
rect 339276 271328 339282 271340
rect 173434 271260 173440 271312
rect 173492 271300 173498 271312
rect 227622 271300 227628 271312
rect 173492 271272 227628 271300
rect 173492 271260 173498 271272
rect 227622 271260 227628 271272
rect 227680 271260 227686 271312
rect 231302 271260 231308 271312
rect 231360 271300 231366 271312
rect 231360 271272 245654 271300
rect 231360 271260 231366 271272
rect 178126 271192 178132 271244
rect 178184 271232 178190 271244
rect 231854 271232 231860 271244
rect 178184 271204 231860 271232
rect 178184 271192 178190 271204
rect 231854 271192 231860 271204
rect 231912 271192 231918 271244
rect 245626 271232 245654 271272
rect 250254 271260 250260 271312
rect 250312 271300 250318 271312
rect 261846 271300 261852 271312
rect 250312 271272 261852 271300
rect 250312 271260 250318 271272
rect 261846 271260 261852 271272
rect 261904 271260 261910 271312
rect 287146 271260 287152 271312
rect 287204 271300 287210 271312
rect 317598 271300 317604 271312
rect 287204 271272 317604 271300
rect 287204 271260 287210 271272
rect 317598 271260 317604 271272
rect 317656 271260 317662 271312
rect 317874 271260 317880 271312
rect 317932 271300 317938 271312
rect 332134 271300 332140 271312
rect 317932 271272 332140 271300
rect 317932 271260 317938 271272
rect 332134 271260 332140 271272
rect 332192 271260 332198 271312
rect 337470 271260 337476 271312
rect 337528 271300 337534 271312
rect 337528 271272 445064 271300
rect 337528 271260 337534 271272
rect 254670 271232 254676 271244
rect 245626 271204 254676 271232
rect 254670 271192 254676 271204
rect 254728 271192 254734 271244
rect 304074 271192 304080 271244
rect 304132 271232 304138 271244
rect 324222 271232 324228 271244
rect 304132 271204 324228 271232
rect 304132 271192 304138 271204
rect 324222 271192 324228 271204
rect 324280 271192 324286 271244
rect 333974 271192 333980 271244
rect 334032 271232 334038 271244
rect 441706 271232 441712 271244
rect 334032 271204 441712 271232
rect 334032 271192 334038 271204
rect 441706 271192 441712 271204
rect 441764 271192 441770 271244
rect 175826 271124 175832 271176
rect 175884 271164 175890 271176
rect 229094 271164 229100 271176
rect 175884 271136 229100 271164
rect 175884 271124 175890 271136
rect 229094 271124 229100 271136
rect 229152 271124 229158 271176
rect 246758 271124 246764 271176
rect 246816 271164 246822 271176
rect 260466 271164 260472 271176
rect 246816 271136 260472 271164
rect 246816 271124 246822 271136
rect 260466 271124 260472 271136
rect 260524 271124 260530 271176
rect 334802 271124 334808 271176
rect 334860 271164 334866 271176
rect 444098 271164 444104 271176
rect 334860 271136 444104 271164
rect 334860 271124 334866 271136
rect 444098 271124 444104 271136
rect 444156 271124 444162 271176
rect 445036 271164 445064 271272
rect 447336 271232 447364 271340
rect 458146 271300 458174 271340
rect 461854 271300 461860 271312
rect 458146 271272 461860 271300
rect 461854 271260 461860 271272
rect 461912 271260 461918 271312
rect 455874 271232 455880 271244
rect 447336 271204 455880 271232
rect 455874 271192 455880 271204
rect 455932 271192 455938 271244
rect 451182 271164 451188 271176
rect 445036 271136 451188 271164
rect 451182 271124 451188 271136
rect 451240 271124 451246 271176
rect 186406 271056 186412 271108
rect 186464 271096 186470 271108
rect 231946 271096 231952 271108
rect 186464 271068 231952 271096
rect 186464 271056 186470 271068
rect 231946 271056 231952 271068
rect 232004 271056 232010 271108
rect 251266 271056 251272 271108
rect 251324 271096 251330 271108
rect 258718 271096 258724 271108
rect 251324 271068 258724 271096
rect 251324 271056 251330 271068
rect 258718 271056 258724 271068
rect 258776 271056 258782 271108
rect 329466 271056 329472 271108
rect 329524 271096 329530 271108
rect 429930 271096 429936 271108
rect 329524 271068 429936 271096
rect 329524 271056 329530 271068
rect 429930 271056 429936 271068
rect 429988 271056 429994 271108
rect 442534 271056 442540 271108
rect 442592 271096 442598 271108
rect 454678 271096 454684 271108
rect 442592 271068 454684 271096
rect 442592 271056 442598 271068
rect 454678 271056 454684 271068
rect 454736 271056 454742 271108
rect 180518 270988 180524 271040
rect 180576 271028 180582 271040
rect 227806 271028 227812 271040
rect 180576 271000 227812 271028
rect 180576 270988 180582 271000
rect 227806 270988 227812 271000
rect 227864 270988 227870 271040
rect 251174 270988 251180 271040
rect 251232 271028 251238 271040
rect 260006 271028 260012 271040
rect 251232 271000 260012 271028
rect 251232 270988 251238 271000
rect 260006 270988 260012 271000
rect 260064 270988 260070 271040
rect 328638 270988 328644 271040
rect 328696 271028 328702 271040
rect 427538 271028 427544 271040
rect 328696 271000 427544 271028
rect 328696 270988 328702 271000
rect 427538 270988 427544 271000
rect 427596 270988 427602 271040
rect 187602 270920 187608 270972
rect 187660 270960 187666 270972
rect 230750 270960 230756 270972
rect 187660 270932 230756 270960
rect 187660 270920 187666 270932
rect 230750 270920 230756 270932
rect 230808 270920 230814 270972
rect 325970 270920 325976 270972
rect 326028 270960 326034 270972
rect 420454 270960 420460 270972
rect 326028 270932 420460 270960
rect 326028 270920 326034 270932
rect 420454 270920 420460 270932
rect 420512 270920 420518 270972
rect 420822 270920 420828 270972
rect 420880 270960 420886 270972
rect 447594 270960 447600 270972
rect 420880 270932 447600 270960
rect 420880 270920 420886 270932
rect 447594 270920 447600 270932
rect 447652 270920 447658 270972
rect 184106 270852 184112 270904
rect 184164 270892 184170 270904
rect 227438 270892 227444 270904
rect 184164 270864 227444 270892
rect 184164 270852 184170 270864
rect 227438 270852 227444 270864
rect 227496 270852 227502 270904
rect 325786 270852 325792 270904
rect 325844 270892 325850 270904
rect 376754 270892 376760 270904
rect 325844 270864 376760 270892
rect 325844 270852 325850 270864
rect 376754 270852 376760 270864
rect 376812 270852 376818 270904
rect 385678 270852 385684 270904
rect 385736 270892 385742 270904
rect 437014 270892 437020 270904
rect 385736 270864 437020 270892
rect 385736 270852 385742 270864
rect 437014 270852 437020 270864
rect 437072 270852 437078 270904
rect 189994 270784 190000 270836
rect 190052 270824 190058 270836
rect 229830 270824 229836 270836
rect 190052 270796 229836 270824
rect 190052 270784 190058 270796
rect 229830 270784 229836 270796
rect 229888 270784 229894 270836
rect 325694 270784 325700 270836
rect 325752 270824 325758 270836
rect 325752 270796 351868 270824
rect 325752 270784 325758 270796
rect 179322 270716 179328 270768
rect 179380 270756 179386 270768
rect 184106 270756 184112 270768
rect 179380 270728 184112 270756
rect 179380 270716 179386 270728
rect 184106 270716 184112 270728
rect 184164 270716 184170 270768
rect 187694 270716 187700 270768
rect 187752 270756 187758 270768
rect 187752 270728 197400 270756
rect 187752 270716 187758 270728
rect 71774 270648 71780 270700
rect 71832 270688 71838 270700
rect 194594 270688 194600 270700
rect 71832 270660 194600 270688
rect 71832 270648 71838 270660
rect 194594 270648 194600 270660
rect 194652 270648 194658 270700
rect 189902 270580 189908 270632
rect 189960 270620 189966 270632
rect 197170 270620 197176 270632
rect 189960 270592 197176 270620
rect 189960 270580 189966 270592
rect 197170 270580 197176 270592
rect 197228 270580 197234 270632
rect 197372 270620 197400 270728
rect 199470 270716 199476 270768
rect 199528 270756 199534 270768
rect 242618 270756 242624 270768
rect 199528 270728 242624 270756
rect 199528 270716 199534 270728
rect 242618 270716 242624 270728
rect 242676 270716 242682 270768
rect 317230 270716 317236 270768
rect 317288 270756 317294 270768
rect 345934 270756 345940 270768
rect 317288 270728 345940 270756
rect 317288 270716 317294 270728
rect 345934 270716 345940 270728
rect 345992 270716 345998 270768
rect 201770 270648 201776 270700
rect 201828 270688 201834 270700
rect 243538 270688 243544 270700
rect 201828 270660 243544 270688
rect 201828 270648 201834 270660
rect 243538 270648 243544 270660
rect 243596 270648 243602 270700
rect 256142 270648 256148 270700
rect 256200 270688 256206 270700
rect 264054 270688 264060 270700
rect 256200 270660 264060 270688
rect 256200 270648 256206 270660
rect 264054 270648 264060 270660
rect 264112 270648 264118 270700
rect 319898 270648 319904 270700
rect 319956 270688 319962 270700
rect 349522 270688 349528 270700
rect 319956 270660 349528 270688
rect 319956 270648 319962 270660
rect 349522 270648 349528 270660
rect 349580 270648 349586 270700
rect 351840 270688 351868 270796
rect 354858 270784 354864 270836
rect 354916 270824 354922 270836
rect 358906 270824 358912 270836
rect 354916 270796 358912 270824
rect 354916 270784 354922 270796
rect 358906 270784 358912 270796
rect 358964 270784 358970 270836
rect 381354 270784 381360 270836
rect 381412 270824 381418 270836
rect 422846 270824 422852 270836
rect 381412 270796 422852 270824
rect 381412 270784 381418 270796
rect 422846 270784 422852 270796
rect 422904 270784 422910 270836
rect 360838 270716 360844 270768
rect 360896 270756 360902 270768
rect 373166 270756 373172 270768
rect 360896 270728 373172 270756
rect 360896 270716 360902 270728
rect 373166 270716 373172 270728
rect 373224 270716 373230 270768
rect 375558 270716 375564 270768
rect 375616 270756 375622 270768
rect 408586 270756 408592 270768
rect 375616 270728 408592 270756
rect 375616 270716 375622 270728
rect 408586 270716 408592 270728
rect 408644 270716 408650 270768
rect 366082 270688 366088 270700
rect 351840 270660 366088 270688
rect 366082 270648 366088 270660
rect 366140 270648 366146 270700
rect 369854 270648 369860 270700
rect 369912 270688 369918 270700
rect 401502 270688 401508 270700
rect 369912 270660 401508 270688
rect 369912 270648 369918 270660
rect 401502 270648 401508 270660
rect 401560 270648 401566 270700
rect 207658 270620 207664 270632
rect 197372 270592 207664 270620
rect 207658 270580 207664 270592
rect 207716 270580 207722 270632
rect 207750 270580 207756 270632
rect 207808 270620 207814 270632
rect 215202 270620 215208 270632
rect 207808 270592 215208 270620
rect 207808 270580 207814 270592
rect 215202 270580 215208 270592
rect 215260 270580 215266 270632
rect 218330 270580 218336 270632
rect 218388 270620 218394 270632
rect 223390 270620 223396 270632
rect 218388 270592 223396 270620
rect 218388 270580 218394 270592
rect 223390 270580 223396 270592
rect 223448 270580 223454 270632
rect 226610 270580 226616 270632
rect 226668 270620 226674 270632
rect 252922 270620 252928 270632
rect 226668 270592 252928 270620
rect 226668 270580 226674 270592
rect 252922 270580 252928 270592
rect 252980 270580 252986 270632
rect 313182 270580 313188 270632
rect 313240 270620 313246 270632
rect 342438 270620 342444 270632
rect 313240 270592 342444 270620
rect 313240 270580 313246 270592
rect 342438 270580 342444 270592
rect 342496 270580 342502 270632
rect 375374 270580 375380 270632
rect 375432 270620 375438 270632
rect 394418 270620 394424 270632
rect 375432 270592 394424 270620
rect 375432 270580 375438 270592
rect 394418 270580 394424 270592
rect 394476 270580 394482 270632
rect 400766 270580 400772 270632
rect 400824 270620 400830 270632
rect 413830 270620 413836 270632
rect 400824 270592 413836 270620
rect 400824 270580 400830 270592
rect 413830 270580 413836 270592
rect 413888 270580 413894 270632
rect 150986 270512 150992 270564
rect 151044 270552 151050 270564
rect 151044 270524 154528 270552
rect 151044 270512 151050 270524
rect 154500 270484 154528 270524
rect 192386 270512 192392 270564
rect 192444 270552 192450 270564
rect 239950 270552 239956 270564
rect 192444 270524 239956 270552
rect 192444 270512 192450 270524
rect 239950 270512 239956 270524
rect 240008 270512 240014 270564
rect 364334 270512 364340 270564
rect 364392 270552 364398 270564
rect 380250 270552 380256 270564
rect 364392 270524 380256 270552
rect 364392 270512 364398 270524
rect 380250 270512 380256 270524
rect 380308 270512 380314 270564
rect 207566 270484 207572 270496
rect 154500 270456 207572 270484
rect 207566 270444 207572 270456
rect 207624 270444 207630 270496
rect 207658 270444 207664 270496
rect 207716 270484 207722 270496
rect 214650 270484 214656 270496
rect 207716 270456 214656 270484
rect 207716 270444 207722 270456
rect 214650 270444 214656 270456
rect 214708 270444 214714 270496
rect 227622 270444 227628 270496
rect 227680 270484 227686 270496
rect 232866 270484 232872 270496
rect 227680 270456 232872 270484
rect 227680 270444 227686 270456
rect 232866 270444 232872 270456
rect 232924 270444 232930 270496
rect 265618 270444 265624 270496
rect 265676 270484 265682 270496
rect 267550 270484 267556 270496
rect 265676 270456 267556 270484
rect 265676 270444 265682 270456
rect 267550 270444 267556 270456
rect 267608 270444 267614 270496
rect 269390 270444 269396 270496
rect 269448 270484 269454 270496
rect 270310 270484 270316 270496
rect 269448 270456 270316 270484
rect 269448 270444 269454 270456
rect 270310 270444 270316 270456
rect 270368 270444 270374 270496
rect 270678 270444 270684 270496
rect 270736 270484 270742 270496
rect 273898 270484 273904 270496
rect 270736 270456 273904 270484
rect 270736 270444 270742 270456
rect 273898 270444 273904 270456
rect 273956 270444 273962 270496
rect 274266 270444 274272 270496
rect 274324 270484 274330 270496
rect 283374 270484 283380 270496
rect 274324 270456 283380 270484
rect 274324 270444 274330 270456
rect 283374 270444 283380 270456
rect 283432 270444 283438 270496
rect 294322 270444 294328 270496
rect 294380 270484 294386 270496
rect 336550 270484 336556 270496
rect 294380 270456 336556 270484
rect 294380 270444 294386 270456
rect 336550 270444 336556 270456
rect 336608 270444 336614 270496
rect 351270 270444 351276 270496
rect 351328 270484 351334 270496
rect 351328 270456 357204 270484
rect 351328 270444 351334 270456
rect 148594 270376 148600 270428
rect 148652 270416 148658 270428
rect 223206 270416 223212 270428
rect 148652 270388 223212 270416
rect 148652 270376 148658 270388
rect 223206 270376 223212 270388
rect 223264 270376 223270 270428
rect 229278 270376 229284 270428
rect 229336 270416 229342 270428
rect 232406 270416 232412 270428
rect 229336 270388 232412 270416
rect 229336 270376 229342 270388
rect 232406 270376 232412 270388
rect 232464 270376 232470 270428
rect 271138 270376 271144 270428
rect 271196 270416 271202 270428
rect 275094 270416 275100 270428
rect 271196 270388 275100 270416
rect 271196 270376 271202 270388
rect 275094 270376 275100 270388
rect 275152 270376 275158 270428
rect 277486 270376 277492 270428
rect 277544 270416 277550 270428
rect 291562 270416 291568 270428
rect 277544 270388 291568 270416
rect 277544 270376 277550 270388
rect 291562 270376 291568 270388
rect 291620 270376 291626 270428
rect 295610 270376 295616 270428
rect 295668 270416 295674 270428
rect 340046 270416 340052 270428
rect 295668 270388 340052 270416
rect 295668 270376 295674 270388
rect 340046 270376 340052 270388
rect 340104 270376 340110 270428
rect 349062 270376 349068 270428
rect 349120 270416 349126 270428
rect 356054 270416 356060 270428
rect 349120 270388 356060 270416
rect 349120 270376 349126 270388
rect 356054 270376 356060 270388
rect 356112 270376 356118 270428
rect 145098 270308 145104 270360
rect 145156 270348 145162 270360
rect 222194 270348 222200 270360
rect 145156 270320 222200 270348
rect 145156 270308 145162 270320
rect 222194 270308 222200 270320
rect 222252 270308 222258 270360
rect 224218 270308 224224 270360
rect 224276 270348 224282 270360
rect 252002 270348 252008 270360
rect 224276 270320 252008 270348
rect 224276 270308 224282 270320
rect 252002 270308 252008 270320
rect 252060 270308 252066 270360
rect 271598 270308 271604 270360
rect 271656 270348 271662 270360
rect 276198 270348 276204 270360
rect 271656 270320 276204 270348
rect 271656 270308 271662 270320
rect 276198 270308 276204 270320
rect 276256 270308 276262 270360
rect 277854 270308 277860 270360
rect 277912 270348 277918 270360
rect 277912 270320 282500 270348
rect 277912 270308 277918 270320
rect 143902 270240 143908 270292
rect 143960 270280 143966 270292
rect 221274 270280 221280 270292
rect 143960 270252 221280 270280
rect 143960 270240 143966 270252
rect 221274 270240 221280 270252
rect 221332 270240 221338 270292
rect 225414 270240 225420 270292
rect 225472 270280 225478 270292
rect 252462 270280 252468 270292
rect 225472 270252 252468 270280
rect 225472 270240 225478 270252
rect 252462 270240 252468 270252
rect 252520 270240 252526 270292
rect 272058 270240 272064 270292
rect 272116 270280 272122 270292
rect 277394 270280 277400 270292
rect 272116 270252 277400 270280
rect 272116 270240 272122 270252
rect 277394 270240 277400 270252
rect 277452 270240 277458 270292
rect 278682 270240 278688 270292
rect 278740 270280 278746 270292
rect 278740 270252 282408 270280
rect 278740 270240 278746 270252
rect 135622 270172 135628 270224
rect 135680 270212 135686 270224
rect 219066 270212 219072 270224
rect 135680 270184 219072 270212
rect 135680 270172 135686 270184
rect 219066 270172 219072 270184
rect 219124 270172 219130 270224
rect 219526 270172 219532 270224
rect 219584 270212 219590 270224
rect 250254 270212 250260 270224
rect 219584 270184 250260 270212
rect 219584 270172 219590 270184
rect 250254 270172 250260 270184
rect 250312 270172 250318 270224
rect 272518 270172 272524 270224
rect 272576 270212 272582 270224
rect 278590 270212 278596 270224
rect 272576 270184 278596 270212
rect 272576 270172 272582 270184
rect 278590 270172 278596 270184
rect 278648 270172 278654 270224
rect 279142 270172 279148 270224
rect 279200 270212 279206 270224
rect 279200 270184 282316 270212
rect 279200 270172 279206 270184
rect 142706 270104 142712 270156
rect 142764 270144 142770 270156
rect 221734 270144 221740 270156
rect 142764 270116 221740 270144
rect 142764 270104 142770 270116
rect 221734 270104 221740 270116
rect 221792 270104 221798 270156
rect 221918 270104 221924 270156
rect 221976 270144 221982 270156
rect 251082 270144 251088 270156
rect 221976 270116 251088 270144
rect 221976 270104 221982 270116
rect 251082 270104 251088 270116
rect 251140 270104 251146 270156
rect 272978 270104 272984 270156
rect 273036 270144 273042 270156
rect 279786 270144 279792 270156
rect 273036 270116 279792 270144
rect 273036 270104 273042 270116
rect 279786 270104 279792 270116
rect 279844 270104 279850 270156
rect 136818 270036 136824 270088
rect 136876 270076 136882 270088
rect 218606 270076 218612 270088
rect 136876 270048 218612 270076
rect 136876 270036 136882 270048
rect 218606 270036 218612 270048
rect 218664 270036 218670 270088
rect 223390 270036 223396 270088
rect 223448 270076 223454 270088
rect 249794 270076 249800 270088
rect 223448 270048 249800 270076
rect 223448 270036 223454 270048
rect 249794 270036 249800 270048
rect 249852 270036 249858 270088
rect 273714 270036 273720 270088
rect 273772 270076 273778 270088
rect 280982 270076 280988 270088
rect 273772 270048 280988 270076
rect 273772 270036 273778 270048
rect 280982 270036 280988 270048
rect 281040 270036 281046 270088
rect 137922 269968 137928 270020
rect 137980 270008 137986 270020
rect 219526 270008 219532 270020
rect 137980 269980 219532 270008
rect 137980 269968 137986 269980
rect 219526 269968 219532 269980
rect 219584 269968 219590 270020
rect 220722 269968 220728 270020
rect 220780 270008 220786 270020
rect 250714 270008 250720 270020
rect 220780 269980 250720 270008
rect 220780 269968 220786 269980
rect 250714 269968 250720 269980
rect 250772 269968 250778 270020
rect 273806 269968 273812 270020
rect 273864 270008 273870 270020
rect 282178 270008 282184 270020
rect 273864 269980 282184 270008
rect 273864 269968 273870 269980
rect 282178 269968 282184 269980
rect 282236 269968 282242 270020
rect 282288 270008 282316 270184
rect 282380 270144 282408 270252
rect 282472 270212 282500 270320
rect 297450 270308 297456 270360
rect 297508 270348 297514 270360
rect 344830 270348 344836 270360
rect 297508 270320 344836 270348
rect 297508 270308 297514 270320
rect 344830 270308 344836 270320
rect 344888 270308 344894 270360
rect 350902 270308 350908 270360
rect 350960 270348 350966 270360
rect 357176 270348 357204 270456
rect 362862 270444 362868 270496
rect 362920 270484 362926 270496
rect 480714 270484 480720 270496
rect 362920 270456 480720 270484
rect 362920 270444 362926 270456
rect 480714 270444 480720 270456
rect 480772 270444 480778 270496
rect 358906 270376 358912 270428
rect 358964 270416 358970 270428
rect 491478 270416 491484 270428
rect 358964 270388 491484 270416
rect 358964 270376 358970 270388
rect 491478 270376 491484 270388
rect 491536 270376 491542 270428
rect 487798 270348 487804 270360
rect 350960 270320 353294 270348
rect 357176 270320 487804 270348
rect 350960 270308 350966 270320
rect 282546 270240 282552 270292
rect 282604 270280 282610 270292
rect 290458 270280 290464 270292
rect 282604 270252 290464 270280
rect 282604 270240 282610 270252
rect 290458 270240 290464 270252
rect 290516 270240 290522 270292
rect 296990 270240 296996 270292
rect 297048 270280 297054 270292
rect 343634 270280 343640 270292
rect 297048 270252 343640 270280
rect 297048 270240 297054 270252
rect 343634 270240 343640 270252
rect 343692 270240 343698 270292
rect 353266 270280 353294 270320
rect 487798 270308 487804 270320
rect 487856 270308 487862 270360
rect 486602 270280 486608 270292
rect 353266 270252 486608 270280
rect 486602 270240 486608 270252
rect 486660 270240 486666 270292
rect 292758 270212 292764 270224
rect 282472 270184 292764 270212
rect 292758 270172 292764 270184
rect 292816 270172 292822 270224
rect 298278 270172 298284 270224
rect 298336 270212 298342 270224
rect 347130 270212 347136 270224
rect 298336 270184 347136 270212
rect 298336 270172 298342 270184
rect 347130 270172 347136 270184
rect 347188 270172 347194 270224
rect 348602 270172 348608 270224
rect 348660 270212 348666 270224
rect 351914 270212 351920 270224
rect 348660 270184 351920 270212
rect 348660 270172 348666 270184
rect 351914 270172 351920 270184
rect 351972 270172 351978 270224
rect 353570 270172 353576 270224
rect 353628 270212 353634 270224
rect 493686 270212 493692 270224
rect 353628 270184 493692 270212
rect 353628 270172 353634 270184
rect 493686 270172 493692 270184
rect 493744 270172 493750 270224
rect 295150 270144 295156 270156
rect 282380 270116 295156 270144
rect 295150 270104 295156 270116
rect 295208 270104 295214 270156
rect 298830 270104 298836 270156
rect 298888 270144 298894 270156
rect 348326 270144 348332 270156
rect 298888 270116 348332 270144
rect 298888 270104 298894 270116
rect 348326 270104 348332 270116
rect 348384 270104 348390 270156
rect 348786 270104 348792 270156
rect 348844 270144 348850 270156
rect 355410 270144 355416 270156
rect 348844 270116 355416 270144
rect 348844 270104 348850 270116
rect 355410 270104 355416 270116
rect 355468 270104 355474 270156
rect 494882 270144 494888 270156
rect 355520 270116 494888 270144
rect 282362 270036 282368 270088
rect 282420 270076 282426 270088
rect 293954 270076 293960 270088
rect 282420 270048 293960 270076
rect 282420 270036 282426 270048
rect 293954 270036 293960 270048
rect 294012 270036 294018 270088
rect 300578 270036 300584 270088
rect 300636 270076 300642 270088
rect 353110 270076 353116 270088
rect 300636 270048 353116 270076
rect 300636 270036 300642 270048
rect 353110 270036 353116 270048
rect 353168 270036 353174 270088
rect 353938 270036 353944 270088
rect 353996 270076 354002 270088
rect 355520 270076 355548 270116
rect 494882 270104 494888 270116
rect 494940 270104 494946 270156
rect 353996 270048 355548 270076
rect 353996 270036 354002 270048
rect 356238 270036 356244 270088
rect 356296 270076 356302 270088
rect 500862 270076 500868 270088
rect 356296 270048 500868 270076
rect 356296 270036 356302 270048
rect 500862 270036 500868 270048
rect 500920 270036 500926 270088
rect 296346 270008 296352 270020
rect 282288 269980 296352 270008
rect 296346 269968 296352 269980
rect 296404 269968 296410 270020
rect 300118 269968 300124 270020
rect 300176 270008 300182 270020
rect 351546 270008 351552 270020
rect 300176 269980 351552 270008
rect 300176 269968 300182 269980
rect 351546 269968 351552 269980
rect 351604 269968 351610 270020
rect 360838 270008 360844 270020
rect 351656 269980 360844 270008
rect 130838 269900 130844 269952
rect 130896 269940 130902 269952
rect 216858 269940 216864 269952
rect 130896 269912 216864 269940
rect 130896 269900 130902 269912
rect 216858 269900 216864 269912
rect 216916 269900 216922 269952
rect 223114 269900 223120 269952
rect 223172 269940 223178 269952
rect 251542 269940 251548 269952
rect 223172 269912 251548 269940
rect 223172 269900 223178 269912
rect 251542 269900 251548 269912
rect 251600 269900 251606 269952
rect 279602 269900 279608 269952
rect 279660 269940 279666 269952
rect 297542 269940 297548 269952
rect 279660 269912 297548 269940
rect 279660 269900 279666 269912
rect 297542 269900 297548 269912
rect 297600 269900 297606 269952
rect 301406 269900 301412 269952
rect 301464 269940 301470 269952
rect 348786 269940 348792 269952
rect 301464 269912 348792 269940
rect 301464 269900 301470 269912
rect 348786 269900 348792 269912
rect 348844 269900 348850 269952
rect 129642 269832 129648 269884
rect 129700 269872 129706 269884
rect 215846 269872 215852 269884
rect 129700 269844 215852 269872
rect 129700 269832 129706 269844
rect 215846 269832 215852 269844
rect 215904 269832 215910 269884
rect 220446 269832 220452 269884
rect 220504 269872 220510 269884
rect 248414 269872 248420 269884
rect 220504 269844 248420 269872
rect 220504 269832 220510 269844
rect 248414 269832 248420 269844
rect 248472 269832 248478 269884
rect 278314 269832 278320 269884
rect 278372 269872 278378 269884
rect 282362 269872 282368 269884
rect 278372 269844 282368 269872
rect 278372 269832 278378 269844
rect 282362 269832 282368 269844
rect 282420 269832 282426 269884
rect 282454 269832 282460 269884
rect 282512 269872 282518 269884
rect 286870 269872 286876 269884
rect 282512 269844 286876 269872
rect 282512 269832 282518 269844
rect 286870 269832 286876 269844
rect 286928 269832 286934 269884
rect 308214 269832 308220 269884
rect 308272 269872 308278 269884
rect 351656 269872 351684 269980
rect 360838 269968 360844 269980
rect 360896 269968 360902 270020
rect 361574 269968 361580 270020
rect 361632 270008 361638 270020
rect 515030 270008 515036 270020
rect 361632 269980 515036 270008
rect 361632 269968 361638 269980
rect 515030 269968 515036 269980
rect 515088 269968 515094 270020
rect 364334 269940 364340 269952
rect 308272 269844 351684 269872
rect 351840 269912 364340 269940
rect 308272 269832 308278 269844
rect 128538 269764 128544 269816
rect 128596 269804 128602 269816
rect 216398 269804 216404 269816
rect 128596 269776 216404 269804
rect 128596 269764 128602 269776
rect 216398 269764 216404 269776
rect 216456 269764 216462 269816
rect 217962 269764 217968 269816
rect 218020 269804 218026 269816
rect 247126 269804 247132 269816
rect 218020 269776 247132 269804
rect 218020 269764 218026 269776
rect 247126 269764 247132 269776
rect 247184 269764 247190 269816
rect 280522 269764 280528 269816
rect 280580 269804 280586 269816
rect 299842 269804 299848 269816
rect 280580 269776 299848 269804
rect 280580 269764 280586 269776
rect 299842 269764 299848 269776
rect 299900 269764 299906 269816
rect 302786 269764 302792 269816
rect 302844 269804 302850 269816
rect 349062 269804 349068 269816
rect 302844 269776 349068 269804
rect 302844 269764 302850 269776
rect 349062 269764 349068 269776
rect 349120 269764 349126 269816
rect 122558 269696 122564 269748
rect 122616 269736 122622 269748
rect 213270 269736 213276 269748
rect 122616 269708 213276 269736
rect 122616 269696 122622 269708
rect 213270 269696 213276 269708
rect 213328 269696 213334 269748
rect 215938 269696 215944 269748
rect 215996 269736 216002 269748
rect 248874 269736 248880 269748
rect 215996 269708 248880 269736
rect 215996 269696 216002 269708
rect 248874 269696 248880 269708
rect 248932 269696 248938 269748
rect 280062 269696 280068 269748
rect 280120 269736 280126 269748
rect 298738 269736 298744 269748
rect 280120 269708 298744 269736
rect 280120 269696 280126 269708
rect 298738 269696 298744 269708
rect 298796 269696 298802 269748
rect 310790 269696 310796 269748
rect 310848 269736 310854 269748
rect 351840 269736 351868 269912
rect 364334 269900 364340 269912
rect 364392 269900 364398 269952
rect 364702 269900 364708 269952
rect 364760 269940 364766 269952
rect 523310 269940 523316 269952
rect 364760 269912 523316 269940
rect 364760 269900 364766 269912
rect 523310 269900 523316 269912
rect 523368 269900 523374 269952
rect 351914 269832 351920 269884
rect 351972 269872 351978 269884
rect 362862 269872 362868 269884
rect 351972 269844 362868 269872
rect 351972 269832 351978 269844
rect 362862 269832 362868 269844
rect 362920 269832 362926 269884
rect 367370 269832 367376 269884
rect 367428 269872 367434 269884
rect 530394 269872 530400 269884
rect 367428 269844 530400 269872
rect 367428 269832 367434 269844
rect 530394 269832 530400 269844
rect 530452 269832 530458 269884
rect 370038 269764 370044 269816
rect 370096 269804 370102 269816
rect 537478 269804 537484 269816
rect 370096 269776 537484 269804
rect 370096 269764 370102 269776
rect 537478 269764 537484 269776
rect 537536 269764 537542 269816
rect 363690 269736 363696 269748
rect 310848 269708 351868 269736
rect 351932 269708 363696 269736
rect 310848 269696 310854 269708
rect 101306 269628 101312 269680
rect 101364 269668 101370 269680
rect 205266 269668 205272 269680
rect 101364 269640 205272 269668
rect 101364 269628 101370 269640
rect 205266 269628 205272 269640
rect 205324 269628 205330 269680
rect 215202 269628 215208 269680
rect 215260 269668 215266 269680
rect 245746 269668 245752 269680
rect 215260 269640 245752 269668
rect 215260 269628 215266 269640
rect 245746 269628 245752 269640
rect 245804 269628 245810 269680
rect 281810 269628 281816 269680
rect 281868 269668 281874 269680
rect 303430 269668 303436 269680
rect 281868 269640 303436 269668
rect 281868 269628 281874 269640
rect 303430 269628 303436 269640
rect 303488 269628 303494 269680
rect 313458 269628 313464 269680
rect 313516 269668 313522 269680
rect 351822 269668 351828 269680
rect 313516 269640 351828 269668
rect 313516 269628 313522 269640
rect 351822 269628 351828 269640
rect 351880 269628 351886 269680
rect 115474 269560 115480 269612
rect 115532 269600 115538 269612
rect 210602 269600 210608 269612
rect 115532 269572 210608 269600
rect 115532 269560 115538 269572
rect 210602 269560 210608 269572
rect 210660 269560 210666 269612
rect 217134 269560 217140 269612
rect 217192 269600 217198 269612
rect 249334 269600 249340 269612
rect 217192 269572 249340 269600
rect 217192 269560 217198 269572
rect 249334 269560 249340 269572
rect 249392 269560 249398 269612
rect 281442 269560 281448 269612
rect 281500 269600 281506 269612
rect 302234 269600 302240 269612
rect 281500 269572 302240 269600
rect 281500 269560 281506 269572
rect 302234 269560 302240 269572
rect 302292 269560 302298 269612
rect 304534 269560 304540 269612
rect 304592 269600 304598 269612
rect 351932 269600 351960 269708
rect 363690 269696 363696 269708
rect 363748 269696 363754 269748
rect 372706 269696 372712 269748
rect 372764 269736 372770 269748
rect 544562 269736 544568 269748
rect 372764 269708 544568 269736
rect 372764 269696 372770 269708
rect 544562 269696 544568 269708
rect 544620 269696 544626 269748
rect 352006 269628 352012 269680
rect 352064 269668 352070 269680
rect 367094 269668 367100 269680
rect 352064 269640 367100 269668
rect 352064 269628 352070 269640
rect 367094 269628 367100 269640
rect 367152 269628 367158 269680
rect 375466 269628 375472 269680
rect 375524 269668 375530 269680
rect 551646 269668 551652 269680
rect 375524 269640 551652 269668
rect 375524 269628 375530 269640
rect 551646 269628 551652 269640
rect 551704 269628 551710 269680
rect 304592 269572 351960 269600
rect 304592 269560 304598 269572
rect 352466 269560 352472 269612
rect 352524 269600 352530 269612
rect 361666 269600 361672 269612
rect 352524 269572 361672 269600
rect 352524 269560 352530 269572
rect 361666 269560 361672 269572
rect 361724 269560 361730 269612
rect 362862 269560 362868 269612
rect 362920 269600 362926 269612
rect 385678 269600 385684 269612
rect 362920 269572 385684 269600
rect 362920 269560 362926 269572
rect 385678 269560 385684 269572
rect 385736 269560 385742 269612
rect 558730 269600 558736 269612
rect 390480 269572 558736 269600
rect 100110 269492 100116 269544
rect 100168 269532 100174 269544
rect 205726 269532 205732 269544
rect 100168 269504 205732 269532
rect 100168 269492 100174 269504
rect 205726 269492 205732 269504
rect 205784 269492 205790 269544
rect 212442 269492 212448 269544
rect 212500 269532 212506 269544
rect 247586 269532 247592 269544
rect 212500 269504 247592 269532
rect 212500 269492 212506 269504
rect 247586 269492 247592 269504
rect 247644 269492 247650 269544
rect 280982 269492 280988 269544
rect 281040 269532 281046 269544
rect 301038 269532 301044 269544
rect 281040 269504 301044 269532
rect 281040 269492 281046 269504
rect 301038 269492 301044 269504
rect 301096 269492 301102 269544
rect 316126 269492 316132 269544
rect 316184 269532 316190 269544
rect 375374 269532 375380 269544
rect 316184 269504 375380 269532
rect 316184 269492 316190 269504
rect 375374 269492 375380 269504
rect 375432 269492 375438 269544
rect 377858 269492 377864 269544
rect 377916 269532 377922 269544
rect 390480 269532 390508 269572
rect 558730 269560 558736 269572
rect 558788 269560 558794 269612
rect 579982 269532 579988 269544
rect 377916 269504 390508 269532
rect 390664 269504 579988 269532
rect 377916 269492 377922 269504
rect 94222 269424 94228 269476
rect 94280 269464 94286 269476
rect 202598 269464 202604 269476
rect 94280 269436 202604 269464
rect 94280 269424 94286 269436
rect 202598 269424 202604 269436
rect 202656 269424 202662 269476
rect 210050 269424 210056 269476
rect 210108 269464 210114 269476
rect 246666 269464 246672 269476
rect 210108 269436 246672 269464
rect 210108 269424 210114 269436
rect 246666 269424 246672 269436
rect 246724 269424 246730 269476
rect 275646 269424 275652 269476
rect 275704 269464 275710 269476
rect 282454 269464 282460 269476
rect 275704 269436 282460 269464
rect 275704 269424 275710 269436
rect 282454 269424 282460 269436
rect 282512 269424 282518 269476
rect 282730 269424 282736 269476
rect 282788 269464 282794 269476
rect 305822 269464 305828 269476
rect 282788 269436 305828 269464
rect 282788 269424 282794 269436
rect 305822 269424 305828 269436
rect 305880 269424 305886 269476
rect 308582 269424 308588 269476
rect 308640 269464 308646 269476
rect 374362 269464 374368 269476
rect 308640 269436 374368 269464
rect 308640 269424 308646 269436
rect 374362 269424 374368 269436
rect 374420 269424 374426 269476
rect 91830 269356 91836 269408
rect 91888 269396 91894 269408
rect 202138 269396 202144 269408
rect 91888 269368 202144 269396
rect 91888 269356 91894 269368
rect 202138 269356 202144 269368
rect 202196 269356 202202 269408
rect 208854 269356 208860 269408
rect 208912 269396 208918 269408
rect 246206 269396 246212 269408
rect 208912 269368 246212 269396
rect 208912 269356 208918 269368
rect 246206 269356 246212 269368
rect 246264 269356 246270 269408
rect 282270 269356 282276 269408
rect 282328 269396 282334 269408
rect 304626 269396 304632 269408
rect 282328 269368 304632 269396
rect 282328 269356 282334 269368
rect 304626 269356 304632 269368
rect 304684 269356 304690 269408
rect 311250 269356 311256 269408
rect 311308 269396 311314 269408
rect 375650 269396 375656 269408
rect 311308 269368 375656 269396
rect 311308 269356 311314 269368
rect 375650 269356 375656 269368
rect 375708 269356 375714 269408
rect 386046 269356 386052 269408
rect 386104 269396 386110 269408
rect 390664 269396 390692 269504
rect 579982 269492 579988 269504
rect 580040 269492 580046 269544
rect 587066 269464 587072 269476
rect 386104 269368 390692 269396
rect 390756 269436 587072 269464
rect 386104 269356 386110 269368
rect 82446 269288 82452 269340
rect 82504 269328 82510 269340
rect 198550 269328 198556 269340
rect 82504 269300 198556 269328
rect 82504 269288 82510 269300
rect 198550 269288 198556 269300
rect 198608 269288 198614 269340
rect 206554 269288 206560 269340
rect 206612 269328 206618 269340
rect 229002 269328 229008 269340
rect 206612 269300 229008 269328
rect 206612 269288 206618 269300
rect 229002 269288 229008 269300
rect 229060 269288 229066 269340
rect 229094 269288 229100 269340
rect 229152 269328 229158 269340
rect 233326 269328 233332 269340
rect 229152 269300 233332 269328
rect 229152 269288 229158 269300
rect 233326 269288 233332 269300
rect 233384 269288 233390 269340
rect 276934 269288 276940 269340
rect 276992 269328 276998 269340
rect 282546 269328 282552 269340
rect 276992 269300 282552 269328
rect 276992 269288 276998 269300
rect 282546 269288 282552 269300
rect 282604 269288 282610 269340
rect 283650 269288 283656 269340
rect 283708 269328 283714 269340
rect 308122 269328 308128 269340
rect 283708 269300 308128 269328
rect 283708 269288 283714 269300
rect 308122 269288 308128 269300
rect 308180 269288 308186 269340
rect 313918 269288 313924 269340
rect 313976 269328 313982 269340
rect 388530 269328 388536 269340
rect 313976 269300 388536 269328
rect 313976 269288 313982 269300
rect 388530 269288 388536 269300
rect 388588 269288 388594 269340
rect 388714 269288 388720 269340
rect 388772 269328 388778 269340
rect 390756 269328 390784 269436
rect 587066 269424 587072 269436
rect 587124 269424 587130 269476
rect 391382 269356 391388 269408
rect 391440 269396 391446 269408
rect 594242 269396 594248 269408
rect 391440 269368 594248 269396
rect 391440 269356 391446 269368
rect 594242 269356 594248 269368
rect 594300 269356 594306 269408
rect 388772 269300 390784 269328
rect 388772 269288 388778 269300
rect 394050 269288 394056 269340
rect 394108 269328 394114 269340
rect 601326 269328 601332 269340
rect 394108 269300 601332 269328
rect 394108 269288 394114 269300
rect 601326 269288 601332 269300
rect 601384 269288 601390 269340
rect 75362 269220 75368 269272
rect 75420 269260 75426 269272
rect 195422 269260 195428 269272
rect 75420 269232 195428 269260
rect 75420 269220 75426 269232
rect 195422 269220 195428 269232
rect 195480 269220 195486 269272
rect 203610 269220 203616 269272
rect 203668 269260 203674 269272
rect 240410 269260 240416 269272
rect 203668 269232 240416 269260
rect 203668 269220 203674 269232
rect 240410 269220 240416 269232
rect 240468 269220 240474 269272
rect 283190 269220 283196 269272
rect 283248 269260 283254 269272
rect 307018 269260 307024 269272
rect 283248 269232 307024 269260
rect 283248 269220 283254 269232
rect 307018 269220 307024 269232
rect 307076 269220 307082 269272
rect 319254 269220 319260 269272
rect 319312 269260 319318 269272
rect 319312 269232 333100 269260
rect 319312 269220 319318 269232
rect 197078 269152 197084 269204
rect 197136 269192 197142 269204
rect 241790 269192 241796 269204
rect 197136 269164 241796 269192
rect 197136 269152 197142 269164
rect 241790 269152 241796 269164
rect 241848 269152 241854 269204
rect 284938 269152 284944 269204
rect 284996 269192 285002 269204
rect 311710 269192 311716 269204
rect 284996 269164 311716 269192
rect 284996 269152 285002 269164
rect 311710 269152 311716 269164
rect 311768 269152 311774 269204
rect 332962 269192 332968 269204
rect 314626 269164 332968 269192
rect 65886 269084 65892 269136
rect 65944 269124 65950 269136
rect 192386 269124 192392 269136
rect 65944 269096 192392 269124
rect 65944 269084 65950 269096
rect 192386 269084 192392 269096
rect 192444 269084 192450 269136
rect 195882 269084 195888 269136
rect 195940 269124 195946 269136
rect 241330 269124 241336 269136
rect 195940 269096 241336 269124
rect 195940 269084 195946 269096
rect 241330 269084 241336 269096
rect 241388 269084 241394 269136
rect 284570 269084 284576 269136
rect 284628 269124 284634 269136
rect 310514 269124 310520 269136
rect 284628 269096 310520 269124
rect 284628 269084 284634 269096
rect 310514 269084 310520 269096
rect 310572 269084 310578 269136
rect 153378 269016 153384 269068
rect 153436 269056 153442 269068
rect 225782 269056 225788 269068
rect 153436 269028 225788 269056
rect 153436 269016 153442 269028
rect 225782 269016 225788 269028
rect 225840 269016 225846 269068
rect 229002 269016 229008 269068
rect 229060 269056 229066 269068
rect 245286 269056 245292 269068
rect 229060 269028 245292 269056
rect 229060 269016 229066 269028
rect 245286 269016 245292 269028
rect 245344 269016 245350 269068
rect 292942 269016 292948 269068
rect 293000 269056 293006 269068
rect 314626 269056 314654 269164
rect 332962 269152 332968 269164
rect 333020 269152 333026 269204
rect 333072 269192 333100 269232
rect 333146 269220 333152 269272
rect 333204 269260 333210 269272
rect 395614 269260 395620 269272
rect 333204 269232 395620 269260
rect 333204 269220 333210 269232
rect 395614 269220 395620 269232
rect 395672 269220 395678 269272
rect 396718 269220 396724 269272
rect 396776 269260 396782 269272
rect 608410 269260 608416 269272
rect 396776 269232 608416 269260
rect 396776 269220 396782 269232
rect 608410 269220 608416 269232
rect 608468 269220 608474 269272
rect 333072 269164 401456 269192
rect 321922 269084 321928 269136
rect 321980 269124 321986 269136
rect 401318 269124 401324 269136
rect 321980 269096 401324 269124
rect 321980 269084 321986 269096
rect 401318 269084 401324 269096
rect 401376 269084 401382 269136
rect 401428 269124 401456 269164
rect 402054 269152 402060 269204
rect 402112 269192 402118 269204
rect 622578 269192 622584 269204
rect 402112 269164 622584 269192
rect 402112 269152 402118 269164
rect 622578 269152 622584 269164
rect 622636 269152 622642 269204
rect 402698 269124 402704 269136
rect 401428 269096 402704 269124
rect 402698 269084 402704 269096
rect 402756 269084 402762 269136
rect 410058 269084 410064 269136
rect 410116 269124 410122 269136
rect 643830 269124 643836 269136
rect 410116 269096 643836 269124
rect 410116 269084 410122 269096
rect 643830 269084 643836 269096
rect 643888 269084 643894 269136
rect 293000 269028 314654 269056
rect 293000 269016 293006 269028
rect 332594 269016 332600 269068
rect 332652 269056 332658 269068
rect 351730 269056 351736 269068
rect 332652 269028 351736 269056
rect 332652 269016 332658 269028
rect 351730 269016 351736 269028
rect 351788 269016 351794 269068
rect 361666 269016 361672 269068
rect 361724 269056 361730 269068
rect 479518 269056 479524 269068
rect 361724 269028 479524 269056
rect 361724 269016 361730 269028
rect 479518 269016 479524 269028
rect 479576 269016 479582 269068
rect 158070 268948 158076 269000
rect 158128 268988 158134 269000
rect 226610 268988 226616 269000
rect 158128 268960 226616 268988
rect 158128 268948 158134 268960
rect 226610 268948 226616 268960
rect 226668 268948 226674 269000
rect 232038 268948 232044 269000
rect 232096 268988 232102 269000
rect 237742 268988 237748 269000
rect 232096 268960 237748 268988
rect 232096 268948 232102 268960
rect 237742 268948 237748 268960
rect 237800 268948 237806 269000
rect 305454 268948 305460 269000
rect 305512 268988 305518 269000
rect 325694 268988 325700 269000
rect 305512 268960 325700 268988
rect 305512 268948 305518 268960
rect 325694 268948 325700 268960
rect 325752 268948 325758 269000
rect 345474 268948 345480 269000
rect 345532 268988 345538 269000
rect 472434 268988 472440 269000
rect 345532 268960 472440 268988
rect 345532 268948 345538 268960
rect 472434 268948 472440 268960
rect 472492 268948 472498 269000
rect 155678 268880 155684 268932
rect 155736 268920 155742 268932
rect 226150 268920 226156 268932
rect 155736 268892 226156 268920
rect 155736 268880 155742 268892
rect 226150 268880 226156 268892
rect 226208 268880 226214 268932
rect 299198 268880 299204 268932
rect 299256 268920 299262 268932
rect 319898 268920 319904 268932
rect 299256 268892 319904 268920
rect 299256 268880 299262 268892
rect 319898 268880 319904 268892
rect 319956 268880 319962 268932
rect 329926 268880 329932 268932
rect 329984 268920 329990 268932
rect 351914 268920 351920 268932
rect 329984 268892 351920 268920
rect 329984 268880 329990 268892
rect 351914 268880 351920 268892
rect 351972 268880 351978 268932
rect 473630 268920 473636 268932
rect 352024 268892 473636 268920
rect 160462 268812 160468 268864
rect 160520 268852 160526 268864
rect 228450 268852 228456 268864
rect 160520 268824 228456 268852
rect 160520 268812 160526 268824
rect 228450 268812 228456 268824
rect 228508 268812 228514 268864
rect 297910 268812 297916 268864
rect 297968 268852 297974 268864
rect 317230 268852 317236 268864
rect 297968 268824 317236 268852
rect 297968 268812 297974 268824
rect 317230 268812 317236 268824
rect 317288 268812 317294 268864
rect 345934 268812 345940 268864
rect 345992 268852 345998 268864
rect 352024 268852 352052 268892
rect 473630 268880 473636 268892
rect 473688 268880 473694 268932
rect 345992 268824 352052 268852
rect 345992 268812 345998 268824
rect 352098 268812 352104 268864
rect 352156 268852 352162 268864
rect 466546 268852 466552 268864
rect 352156 268824 466552 268852
rect 352156 268812 352162 268824
rect 466546 268812 466552 268824
rect 466604 268812 466610 268864
rect 165154 268744 165160 268796
rect 165212 268784 165218 268796
rect 229278 268784 229284 268796
rect 165212 268756 229284 268784
rect 165212 268744 165218 268756
rect 229278 268744 229284 268756
rect 229336 268744 229342 268796
rect 316586 268744 316592 268796
rect 316644 268784 316650 268796
rect 333146 268784 333152 268796
rect 316644 268756 333152 268784
rect 316644 268744 316650 268756
rect 333146 268744 333152 268756
rect 333204 268744 333210 268796
rect 348234 268744 348240 268796
rect 348292 268784 348298 268796
rect 352466 268784 352472 268796
rect 348292 268756 352472 268784
rect 348292 268744 348298 268756
rect 352466 268744 352472 268756
rect 352524 268744 352530 268796
rect 352558 268744 352564 268796
rect 352616 268784 352622 268796
rect 465350 268784 465356 268796
rect 352616 268756 465356 268784
rect 352616 268744 352622 268756
rect 465350 268744 465356 268756
rect 465408 268744 465414 268796
rect 162762 268676 162768 268728
rect 162820 268716 162826 268728
rect 228818 268716 228824 268728
rect 162820 268688 228824 268716
rect 162820 268676 162826 268688
rect 228818 268676 228824 268688
rect 228876 268676 228882 268728
rect 229830 268676 229836 268728
rect 229888 268716 229894 268728
rect 238662 268716 238668 268728
rect 229888 268688 238668 268716
rect 229888 268676 229894 268688
rect 238662 268676 238668 268688
rect 238720 268676 238726 268728
rect 296530 268676 296536 268728
rect 296588 268716 296594 268728
rect 313182 268716 313188 268728
rect 296588 268688 313188 268716
rect 296588 268676 296594 268688
rect 313182 268676 313188 268688
rect 313240 268676 313246 268728
rect 340598 268676 340604 268728
rect 340656 268716 340662 268728
rect 459462 268716 459468 268728
rect 340656 268688 459468 268716
rect 340656 268676 340662 268688
rect 459462 268676 459468 268688
rect 459520 268676 459526 268728
rect 167546 268608 167552 268660
rect 167604 268648 167610 268660
rect 231118 268648 231124 268660
rect 167604 268620 231124 268648
rect 167604 268608 167610 268620
rect 231118 268608 231124 268620
rect 231176 268608 231182 268660
rect 231946 268608 231952 268660
rect 232004 268648 232010 268660
rect 237282 268648 237288 268660
rect 232004 268620 237288 268648
rect 232004 268608 232010 268620
rect 237282 268608 237288 268620
rect 237340 268608 237346 268660
rect 312078 268608 312084 268660
rect 312136 268648 312142 268660
rect 322842 268648 322848 268660
rect 312136 268620 322848 268648
rect 312136 268608 312142 268620
rect 322842 268608 322848 268620
rect 322900 268608 322906 268660
rect 340138 268608 340144 268660
rect 340196 268648 340202 268660
rect 452654 268648 452660 268660
rect 340196 268620 452660 268648
rect 340196 268608 340202 268620
rect 452654 268608 452660 268620
rect 452712 268608 452718 268660
rect 169846 268540 169852 268592
rect 169904 268580 169910 268592
rect 231486 268580 231492 268592
rect 169904 268552 231492 268580
rect 169904 268540 169910 268552
rect 231486 268540 231492 268552
rect 231544 268540 231550 268592
rect 240134 268540 240140 268592
rect 240192 268580 240198 268592
rect 244458 268580 244464 268592
rect 240192 268552 244464 268580
rect 240192 268540 240198 268552
rect 244458 268540 244464 268552
rect 244516 268540 244522 268592
rect 337930 268540 337936 268592
rect 337988 268580 337994 268592
rect 452378 268580 452384 268592
rect 337988 268552 452384 268580
rect 337988 268540 337994 268552
rect 452378 268540 452384 268552
rect 452436 268540 452442 268592
rect 172238 268472 172244 268524
rect 172296 268512 172302 268524
rect 231946 268512 231952 268524
rect 172296 268484 231952 268512
rect 172296 268472 172302 268484
rect 231946 268472 231952 268484
rect 232004 268472 232010 268524
rect 269850 268472 269856 268524
rect 269908 268512 269914 268524
rect 271506 268512 271512 268524
rect 269908 268484 271512 268512
rect 269908 268472 269914 268484
rect 271506 268472 271512 268484
rect 271564 268472 271570 268524
rect 312538 268472 312544 268524
rect 312596 268512 312602 268524
rect 317322 268512 317328 268524
rect 312596 268484 317328 268512
rect 312596 268472 312602 268484
rect 317322 268472 317328 268484
rect 317380 268472 317386 268524
rect 335262 268472 335268 268524
rect 335320 268512 335326 268524
rect 445294 268512 445300 268524
rect 335320 268484 445300 268512
rect 335320 268472 335326 268484
rect 445294 268472 445300 268484
rect 445352 268472 445358 268524
rect 174630 268404 174636 268456
rect 174688 268444 174694 268456
rect 233786 268444 233792 268456
rect 174688 268416 233792 268444
rect 174688 268404 174694 268416
rect 233786 268404 233792 268416
rect 233844 268404 233850 268456
rect 338850 268404 338856 268456
rect 338908 268444 338914 268456
rect 442534 268444 442540 268456
rect 338908 268416 442540 268444
rect 338908 268404 338914 268416
rect 442534 268404 442540 268416
rect 442592 268404 442598 268456
rect 181714 268336 181720 268388
rect 181772 268376 181778 268388
rect 236454 268376 236460 268388
rect 181772 268348 236460 268376
rect 181772 268336 181778 268348
rect 236454 268336 236460 268348
rect 236512 268336 236518 268388
rect 276474 268336 276480 268388
rect 276532 268376 276538 268388
rect 289262 268376 289268 268388
rect 276532 268348 289268 268376
rect 276532 268336 276538 268348
rect 289262 268336 289268 268348
rect 289320 268336 289326 268388
rect 332134 268336 332140 268388
rect 332192 268376 332198 268388
rect 348142 268376 348148 268388
rect 332192 268348 348148 268376
rect 332192 268336 332198 268348
rect 348142 268336 348148 268348
rect 348200 268336 348206 268388
rect 351730 268336 351736 268388
rect 351788 268376 351794 268388
rect 438210 268376 438216 268388
rect 351788 268348 438216 268376
rect 351788 268336 351794 268348
rect 438210 268336 438216 268348
rect 438268 268336 438274 268388
rect 184106 268268 184112 268320
rect 184164 268308 184170 268320
rect 234614 268308 234620 268320
rect 184164 268280 234620 268308
rect 184164 268268 184170 268280
rect 234614 268268 234620 268280
rect 234672 268268 234678 268320
rect 274726 268268 274732 268320
rect 274784 268308 274790 268320
rect 284478 268308 284484 268320
rect 274784 268280 284484 268308
rect 274784 268268 274790 268280
rect 284478 268268 284484 268280
rect 284536 268268 284542 268320
rect 336458 268268 336464 268320
rect 336516 268308 336522 268320
rect 351822 268308 351828 268320
rect 336516 268280 351828 268308
rect 336516 268268 336522 268280
rect 351822 268268 351828 268280
rect 351880 268268 351886 268320
rect 351914 268268 351920 268320
rect 351972 268308 351978 268320
rect 431126 268308 431132 268320
rect 351972 268280 431132 268308
rect 351972 268268 351978 268280
rect 431126 268268 431132 268280
rect 431184 268268 431190 268320
rect 193214 268200 193220 268252
rect 193272 268240 193278 268252
rect 196342 268240 196348 268252
rect 193272 268212 196348 268240
rect 193272 268200 193278 268212
rect 196342 268200 196348 268212
rect 196400 268200 196406 268252
rect 239122 268240 239128 268252
rect 197924 268212 239128 268240
rect 182910 268132 182916 268184
rect 182968 268172 182974 268184
rect 197262 268172 197268 268184
rect 182968 268144 197268 268172
rect 182968 268132 182974 268144
rect 197262 268132 197268 268144
rect 197320 268132 197326 268184
rect 188798 268064 188804 268116
rect 188856 268104 188862 268116
rect 197924 268104 197952 268212
rect 239122 268200 239128 268212
rect 239180 268200 239186 268252
rect 275186 268200 275192 268252
rect 275244 268240 275250 268252
rect 285674 268240 285680 268252
rect 275244 268212 285680 268240
rect 275244 268200 275250 268212
rect 285674 268200 285680 268212
rect 285732 268200 285738 268252
rect 309410 268200 309416 268252
rect 309468 268240 309474 268252
rect 325786 268240 325792 268252
rect 309468 268212 325792 268240
rect 309468 268200 309474 268212
rect 325786 268200 325792 268212
rect 325844 268200 325850 268252
rect 327258 268200 327264 268252
rect 327316 268240 327322 268252
rect 423950 268240 423956 268252
rect 327316 268212 423956 268240
rect 327316 268200 327322 268212
rect 423950 268200 423956 268212
rect 424008 268200 424014 268252
rect 235994 268172 236000 268184
rect 206296 268144 236000 268172
rect 188856 268076 197952 268104
rect 188856 268064 188862 268076
rect 198826 268064 198832 268116
rect 198884 268104 198890 268116
rect 203886 268104 203892 268116
rect 198884 268076 203892 268104
rect 198884 268064 198890 268076
rect 203886 268064 203892 268076
rect 203944 268064 203950 268116
rect 177114 267996 177120 268048
rect 177172 268036 177178 268048
rect 200758 268036 200764 268048
rect 177172 268008 200764 268036
rect 177172 267996 177178 268008
rect 200758 267996 200764 268008
rect 200816 267996 200822 268048
rect 201494 267996 201500 268048
rect 201552 268036 201558 268048
rect 206186 268036 206192 268048
rect 201552 268008 206192 268036
rect 201552 267996 201558 268008
rect 206186 267996 206192 268008
rect 206244 267996 206250 268048
rect 74166 267928 74172 267980
rect 74224 267968 74230 267980
rect 195882 267968 195888 267980
rect 74224 267940 195888 267968
rect 74224 267928 74230 267940
rect 195882 267928 195888 267940
rect 195940 267928 195946 267980
rect 197262 267928 197268 267980
rect 197320 267968 197326 267980
rect 206296 267968 206324 268144
rect 235994 268132 236000 268144
rect 236052 268132 236058 268184
rect 270310 268132 270316 268184
rect 270368 268172 270374 268184
rect 272702 268172 272708 268184
rect 270368 268144 272708 268172
rect 270368 268132 270374 268144
rect 272702 268132 272708 268144
rect 272760 268132 272766 268184
rect 324590 268132 324596 268184
rect 324648 268172 324654 268184
rect 324648 268144 401180 268172
rect 324648 268132 324654 268144
rect 234154 268104 234160 268116
rect 206480 268076 234160 268104
rect 206480 267968 206508 268076
rect 234154 268064 234160 268076
rect 234212 268064 234218 268116
rect 321462 268064 321468 268116
rect 321520 268104 321526 268116
rect 321520 268076 342254 268104
rect 321520 268064 321526 268076
rect 206554 267996 206560 268048
rect 206612 268036 206618 268048
rect 215478 268036 215484 268048
rect 206612 268008 215484 268036
rect 206612 267996 206618 268008
rect 215478 267996 215484 268008
rect 215536 267996 215542 268048
rect 248046 268036 248052 268048
rect 226306 268008 248052 268036
rect 209222 267968 209228 267980
rect 197320 267940 206324 267968
rect 206388 267940 206508 267968
rect 206664 267940 209228 267968
rect 197320 267928 197326 267940
rect 193122 267860 193128 267912
rect 193180 267900 193186 267912
rect 206388 267900 206416 267940
rect 206664 267900 206692 267940
rect 209222 267928 209228 267940
rect 209280 267928 209286 267980
rect 209682 267928 209688 267980
rect 209740 267968 209746 267980
rect 212350 267968 212356 267980
rect 209740 267940 212356 267968
rect 209740 267928 209746 267940
rect 212350 267928 212356 267940
rect 212408 267928 212414 267980
rect 213638 267928 213644 267980
rect 213696 267968 213702 267980
rect 226306 267968 226334 268008
rect 248046 267996 248052 268008
rect 248104 267996 248110 268048
rect 342226 268036 342254 268076
rect 343266 268064 343272 268116
rect 343324 268104 343330 268116
rect 351730 268104 351736 268116
rect 343324 268076 351736 268104
rect 343324 268064 343330 268076
rect 351730 268064 351736 268076
rect 351788 268064 351794 268116
rect 351822 268064 351828 268116
rect 351880 268104 351886 268116
rect 351880 268076 400214 268104
rect 351880 268064 351886 268076
rect 375558 268036 375564 268048
rect 342226 268008 375564 268036
rect 375558 267996 375564 268008
rect 375616 267996 375622 268048
rect 381998 267996 382004 268048
rect 382056 268036 382062 268048
rect 386414 268036 386420 268048
rect 382056 268008 386420 268036
rect 382056 267996 382062 268008
rect 386414 267996 386420 268008
rect 386472 267996 386478 268048
rect 213696 267940 226334 267968
rect 213696 267928 213702 267940
rect 227806 267928 227812 267980
rect 227864 267968 227870 267980
rect 235534 267968 235540 267980
rect 227864 267940 235540 267968
rect 227864 267928 227870 267940
rect 235534 267928 235540 267940
rect 235592 267928 235598 267980
rect 326798 267928 326804 267980
rect 326856 267968 326862 267980
rect 381354 267968 381360 267980
rect 326856 267940 381360 267968
rect 326856 267928 326862 267940
rect 381354 267928 381360 267940
rect 381412 267928 381418 267980
rect 400186 267968 400214 268076
rect 401152 268036 401180 268144
rect 401318 268132 401324 268184
rect 401376 268172 401382 268184
rect 409782 268172 409788 268184
rect 401376 268144 409788 268172
rect 401376 268132 401382 268144
rect 409782 268132 409788 268144
rect 409840 268132 409846 268184
rect 420822 268104 420828 268116
rect 419506 268076 420828 268104
rect 416866 268036 416872 268048
rect 401152 268008 416872 268036
rect 416866 267996 416872 268008
rect 416924 267996 416930 268048
rect 419506 267968 419534 268076
rect 420822 268064 420828 268076
rect 420880 268064 420886 268116
rect 656250 268064 656256 268116
rect 656308 268104 656314 268116
rect 676214 268104 676220 268116
rect 656308 268076 676220 268104
rect 656308 268064 656314 268076
rect 676214 268064 676220 268076
rect 676272 268064 676278 268116
rect 400186 267940 419534 267968
rect 656066 267928 656072 267980
rect 656124 267968 656130 267980
rect 676030 267968 676036 267980
rect 656124 267940 676036 267968
rect 656124 267928 656130 267940
rect 676030 267928 676036 267940
rect 676088 267928 676094 267980
rect 193180 267872 206416 267900
rect 206480 267872 206692 267900
rect 193180 267860 193186 267872
rect 201586 267792 201592 267844
rect 201644 267832 201650 267844
rect 206480 267832 206508 267872
rect 206830 267860 206836 267912
rect 206888 267900 206894 267912
rect 211890 267900 211896 267912
rect 206888 267872 211896 267900
rect 206888 267860 206894 267872
rect 211890 267860 211896 267872
rect 211948 267860 211954 267912
rect 227438 267860 227444 267912
rect 227496 267900 227502 267912
rect 236914 267900 236920 267912
rect 227496 267872 236920 267900
rect 227496 267860 227502 267872
rect 236914 267860 236920 267872
rect 236972 267860 236978 267912
rect 276290 267860 276296 267912
rect 276348 267900 276354 267912
rect 288066 267900 288072 267912
rect 276348 267872 288072 267900
rect 276348 267860 276354 267872
rect 288066 267860 288072 267872
rect 288124 267860 288130 267912
rect 348142 267860 348148 267912
rect 348200 267900 348206 267912
rect 362862 267900 362868 267912
rect 348200 267872 362868 267900
rect 348200 267860 348206 267872
rect 362862 267860 362868 267872
rect 362920 267860 362926 267912
rect 368198 267860 368204 267912
rect 368256 267900 368262 267912
rect 369670 267900 369676 267912
rect 368256 267872 369676 267900
rect 368256 267860 368262 267872
rect 369670 267860 369676 267872
rect 369728 267860 369734 267912
rect 201644 267804 206508 267832
rect 201644 267792 201650 267804
rect 206738 267792 206744 267844
rect 206796 267832 206802 267844
rect 208854 267832 208860 267844
rect 206796 267804 208860 267832
rect 206796 267792 206802 267804
rect 208854 267792 208860 267804
rect 208912 267792 208918 267844
rect 231854 267792 231860 267844
rect 231912 267832 231918 267844
rect 235074 267832 235080 267844
rect 231912 267804 235080 267832
rect 231912 267792 231918 267804
rect 235074 267792 235080 267804
rect 235132 267792 235138 267844
rect 318794 267792 318800 267844
rect 318852 267832 318858 267844
rect 369854 267832 369860 267844
rect 318852 267804 369860 267832
rect 318852 267792 318858 267804
rect 369854 267792 369860 267804
rect 369912 267792 369918 267844
rect 376662 267792 376668 267844
rect 376720 267832 376726 267844
rect 391934 267832 391940 267844
rect 376720 267804 391940 267832
rect 376720 267792 376726 267804
rect 391934 267792 391940 267804
rect 391992 267792 391998 267844
rect 197170 267724 197176 267776
rect 197228 267764 197234 267776
rect 206554 267764 206560 267776
rect 197228 267736 206560 267764
rect 197228 267724 197234 267736
rect 206554 267724 206560 267736
rect 206612 267724 206618 267776
rect 207566 267724 207572 267776
rect 207624 267764 207630 267776
rect 223942 267764 223948 267776
rect 207624 267736 223948 267764
rect 207624 267724 207630 267736
rect 223942 267724 223948 267736
rect 224000 267724 224006 267776
rect 224034 267724 224040 267776
rect 224092 267764 224098 267776
rect 230198 267764 230204 267776
rect 224092 267736 230204 267764
rect 224092 267724 224098 267736
rect 230198 267724 230204 267736
rect 230256 267724 230262 267776
rect 230750 267724 230756 267776
rect 230808 267764 230814 267776
rect 238202 267764 238208 267776
rect 230808 267736 238208 267764
rect 230808 267724 230814 267736
rect 238202 267724 238208 267736
rect 238260 267724 238266 267776
rect 314838 267724 314844 267776
rect 314896 267764 314902 267776
rect 322658 267764 322664 267776
rect 314896 267736 322664 267764
rect 314896 267724 314902 267736
rect 322658 267724 322664 267736
rect 322716 267724 322722 267776
rect 342806 267724 342812 267776
rect 342864 267764 342870 267776
rect 352558 267764 352564 267776
rect 342864 267736 352564 267764
rect 342864 267724 342870 267736
rect 352558 267724 352564 267736
rect 352616 267724 352622 267776
rect 655882 267724 655888 267776
rect 655940 267764 655946 267776
rect 676122 267764 676128 267776
rect 655940 267736 676128 267764
rect 655940 267724 655946 267736
rect 676122 267724 676128 267736
rect 676180 267724 676186 267776
rect 367738 267656 367744 267708
rect 367796 267696 367802 267708
rect 531590 267696 531596 267708
rect 367796 267668 531596 267696
rect 367796 267656 367802 267668
rect 531590 267656 531596 267668
rect 531648 267656 531654 267708
rect 370498 267588 370504 267640
rect 370556 267628 370562 267640
rect 538674 267628 538680 267640
rect 370556 267600 538680 267628
rect 370556 267588 370562 267600
rect 538674 267588 538680 267600
rect 538732 267588 538738 267640
rect 373166 267520 373172 267572
rect 373224 267560 373230 267572
rect 545758 267560 545764 267572
rect 373224 267532 545764 267560
rect 373224 267520 373230 267532
rect 545758 267520 545764 267532
rect 545816 267520 545822 267572
rect 373534 267452 373540 267504
rect 373592 267492 373598 267504
rect 546954 267492 546960 267504
rect 373592 267464 546960 267492
rect 373592 267452 373598 267464
rect 546954 267452 546960 267464
rect 547012 267452 547018 267504
rect 672994 267452 673000 267504
rect 673052 267492 673058 267504
rect 676030 267492 676036 267504
rect 673052 267464 676036 267492
rect 673052 267452 673058 267464
rect 676030 267452 676036 267464
rect 676088 267452 676094 267504
rect 374454 267384 374460 267436
rect 374512 267424 374518 267436
rect 549254 267424 549260 267436
rect 374512 267396 549260 267424
rect 374512 267384 374518 267396
rect 549254 267384 549260 267396
rect 549312 267384 549318 267436
rect 376202 267316 376208 267368
rect 376260 267356 376266 267368
rect 554038 267356 554044 267368
rect 376260 267328 554044 267356
rect 376260 267316 376266 267328
rect 554038 267316 554044 267328
rect 554096 267316 554102 267368
rect 375834 267248 375840 267300
rect 375892 267288 375898 267300
rect 552842 267288 552848 267300
rect 375892 267260 552848 267288
rect 375892 267248 375898 267260
rect 552842 267248 552848 267260
rect 552900 267248 552906 267300
rect 299658 267180 299664 267232
rect 299716 267220 299722 267232
rect 350718 267220 350724 267232
rect 299716 267192 350724 267220
rect 299716 267180 299722 267192
rect 350718 267180 350724 267192
rect 350776 267180 350782 267232
rect 377122 267180 377128 267232
rect 377180 267220 377186 267232
rect 556338 267220 556344 267232
rect 377180 267192 556344 267220
rect 377180 267180 377186 267192
rect 556338 267180 556344 267192
rect 556396 267180 556402 267232
rect 300946 267112 300952 267164
rect 301004 267152 301010 267164
rect 354214 267152 354220 267164
rect 301004 267124 354220 267152
rect 301004 267112 301010 267124
rect 354214 267112 354220 267124
rect 354272 267112 354278 267164
rect 378502 267112 378508 267164
rect 378560 267152 378566 267164
rect 559926 267152 559932 267164
rect 378560 267124 559932 267152
rect 378560 267112 378566 267124
rect 559926 267112 559932 267124
rect 559984 267112 559990 267164
rect 302326 267044 302332 267096
rect 302384 267084 302390 267096
rect 357802 267084 357808 267096
rect 302384 267056 357808 267084
rect 302384 267044 302390 267056
rect 357802 267044 357808 267056
rect 357860 267044 357866 267096
rect 378870 267044 378876 267096
rect 378928 267084 378934 267096
rect 561122 267084 561128 267096
rect 378928 267056 561128 267084
rect 378928 267044 378934 267056
rect 561122 267044 561128 267056
rect 561180 267044 561186 267096
rect 303706 266976 303712 267028
rect 303764 267016 303770 267028
rect 361390 267016 361396 267028
rect 303764 266988 361396 267016
rect 303764 266976 303770 266988
rect 361390 266976 361396 266988
rect 361448 266976 361454 267028
rect 379790 266976 379796 267028
rect 379848 267016 379854 267028
rect 563422 267016 563428 267028
rect 379848 266988 563428 267016
rect 379848 266976 379854 266988
rect 563422 266976 563428 266988
rect 563480 266976 563486 267028
rect 304994 266908 305000 266960
rect 305052 266948 305058 266960
rect 364886 266948 364892 266960
rect 305052 266920 364892 266948
rect 305052 266908 305058 266920
rect 364886 266908 364892 266920
rect 364944 266908 364950 266960
rect 381630 266908 381636 266960
rect 381688 266948 381694 266960
rect 568206 266948 568212 266960
rect 381688 266920 568212 266948
rect 381688 266908 381694 266920
rect 568206 266908 568212 266920
rect 568264 266908 568270 266960
rect 306374 266840 306380 266892
rect 306432 266880 306438 266892
rect 368474 266880 368480 266892
rect 306432 266852 368480 266880
rect 306432 266840 306438 266852
rect 368474 266840 368480 266852
rect 368532 266840 368538 266892
rect 381170 266840 381176 266892
rect 381228 266880 381234 266892
rect 567010 266880 567016 266892
rect 381228 266852 567016 266880
rect 381228 266840 381234 266852
rect 567010 266840 567016 266852
rect 567068 266840 567074 266892
rect 307662 266772 307668 266824
rect 307720 266812 307726 266824
rect 371970 266812 371976 266824
rect 307720 266784 371976 266812
rect 307720 266772 307726 266784
rect 371970 266772 371976 266784
rect 372028 266772 372034 266824
rect 382458 266772 382464 266824
rect 382516 266812 382522 266824
rect 570598 266812 570604 266824
rect 382516 266784 570604 266812
rect 382516 266772 382522 266784
rect 570598 266772 570604 266784
rect 570656 266772 570662 266824
rect 309042 266704 309048 266756
rect 309100 266744 309106 266756
rect 375742 266744 375748 266756
rect 309100 266716 375748 266744
rect 309100 266704 309106 266716
rect 375742 266704 375748 266716
rect 375800 266704 375806 266756
rect 384298 266704 384304 266756
rect 384356 266744 384362 266756
rect 575290 266744 575296 266756
rect 384356 266716 575296 266744
rect 384356 266704 384362 266716
rect 575290 266704 575296 266716
rect 575348 266704 575354 266756
rect 310330 266636 310336 266688
rect 310388 266676 310394 266688
rect 379054 266676 379060 266688
rect 310388 266648 379060 266676
rect 310388 266636 310394 266648
rect 379054 266636 379060 266648
rect 379112 266636 379118 266688
rect 383838 266636 383844 266688
rect 383896 266676 383902 266688
rect 574094 266676 574100 266688
rect 383896 266648 574100 266676
rect 383896 266636 383902 266648
rect 574094 266636 574100 266648
rect 574152 266636 574158 266688
rect 673270 266636 673276 266688
rect 673328 266676 673334 266688
rect 676030 266676 676036 266688
rect 673328 266648 676036 266676
rect 673328 266636 673334 266648
rect 676030 266636 676036 266648
rect 676088 266636 676094 266688
rect 123754 266568 123760 266620
rect 123812 266608 123818 266620
rect 214190 266608 214196 266620
rect 123812 266580 214196 266608
rect 123812 266568 123818 266580
rect 214190 266568 214196 266580
rect 214248 266568 214254 266620
rect 311710 266568 311716 266620
rect 311768 266608 311774 266620
rect 382642 266608 382648 266620
rect 311768 266580 382648 266608
rect 311768 266568 311774 266580
rect 382642 266568 382648 266580
rect 382700 266568 382706 266620
rect 385126 266568 385132 266620
rect 385184 266608 385190 266620
rect 577682 266608 577688 266620
rect 385184 266580 577688 266608
rect 385184 266568 385190 266580
rect 577682 266568 577688 266580
rect 577740 266568 577746 266620
rect 116670 266500 116676 266552
rect 116728 266540 116734 266552
rect 211522 266540 211528 266552
rect 116728 266512 211528 266540
rect 116728 266500 116734 266512
rect 211522 266500 211528 266512
rect 211580 266500 211586 266552
rect 312998 266500 313004 266552
rect 313056 266540 313062 266552
rect 386138 266540 386144 266552
rect 313056 266512 386144 266540
rect 313056 266500 313062 266512
rect 386138 266500 386144 266512
rect 386196 266500 386202 266552
rect 386506 266500 386512 266552
rect 386564 266540 386570 266552
rect 581178 266540 581184 266552
rect 386564 266512 581184 266540
rect 386564 266500 386570 266512
rect 581178 266500 581184 266512
rect 581236 266500 581242 266552
rect 72970 266432 72976 266484
rect 73028 266472 73034 266484
rect 195054 266472 195060 266484
rect 73028 266444 195060 266472
rect 73028 266432 73034 266444
rect 195054 266432 195060 266444
rect 195112 266432 195118 266484
rect 389174 266432 389180 266484
rect 389232 266472 389238 266484
rect 588262 266472 588268 266484
rect 389232 266444 588268 266472
rect 389232 266432 389238 266444
rect 588262 266432 588268 266444
rect 588320 266432 588326 266484
rect 113174 266364 113180 266416
rect 113232 266404 113238 266416
rect 210142 266404 210148 266416
rect 113232 266376 210148 266404
rect 113232 266364 113238 266376
rect 210142 266364 210148 266376
rect 210200 266364 210206 266416
rect 315666 266364 315672 266416
rect 315724 266404 315730 266416
rect 315724 266376 387104 266404
rect 315724 266364 315730 266376
rect 68186 266296 68192 266348
rect 68244 266336 68250 266348
rect 193214 266336 193220 266348
rect 68244 266308 193220 266336
rect 68244 266296 68250 266308
rect 193214 266296 193220 266308
rect 193272 266296 193278 266348
rect 317046 266296 317052 266348
rect 317104 266336 317110 266348
rect 386874 266336 386880 266348
rect 317104 266308 386880 266336
rect 317104 266296 317110 266308
rect 386874 266296 386880 266308
rect 386932 266296 386938 266348
rect 387076 266336 387104 266376
rect 392302 266364 392308 266416
rect 392360 266404 392366 266416
rect 596542 266404 596548 266416
rect 392360 266376 596548 266404
rect 392360 266364 392366 266376
rect 596542 266364 596548 266376
rect 596600 266364 596606 266416
rect 393222 266336 393228 266348
rect 387076 266308 393228 266336
rect 393222 266296 393228 266308
rect 393280 266296 393286 266348
rect 395798 266296 395804 266348
rect 395856 266336 395862 266348
rect 606018 266336 606024 266348
rect 395856 266308 606024 266336
rect 395856 266296 395862 266308
rect 606018 266296 606024 266308
rect 606076 266296 606082 266348
rect 365070 266228 365076 266280
rect 365128 266268 365134 266280
rect 524506 266268 524512 266280
rect 365128 266240 524512 266268
rect 365128 266228 365134 266240
rect 524506 266228 524512 266240
rect 524564 266228 524570 266280
rect 362402 266160 362408 266212
rect 362460 266200 362466 266212
rect 517330 266200 517336 266212
rect 362460 266172 517336 266200
rect 362460 266160 362466 266172
rect 517330 266160 517336 266172
rect 517388 266160 517394 266212
rect 359734 266092 359740 266144
rect 359792 266132 359798 266144
rect 510246 266132 510252 266144
rect 359792 266104 510252 266132
rect 359792 266092 359798 266104
rect 510246 266092 510252 266104
rect 510304 266092 510310 266144
rect 355778 266024 355784 266076
rect 355836 266064 355842 266076
rect 499666 266064 499672 266076
rect 355836 266036 499672 266064
rect 355836 266024 355842 266036
rect 499666 266024 499672 266036
rect 499724 266024 499730 266076
rect 354398 265956 354404 266008
rect 354456 265996 354462 266008
rect 496078 265996 496084 266008
rect 354456 265968 496084 265996
rect 354456 265956 354462 265968
rect 496078 265956 496084 265968
rect 496136 265956 496142 266008
rect 350258 265888 350264 265940
rect 350316 265928 350322 265940
rect 485498 265928 485504 265940
rect 350316 265900 485504 265928
rect 350316 265888 350322 265900
rect 485498 265888 485504 265900
rect 485556 265888 485562 265940
rect 349062 265820 349068 265872
rect 349120 265860 349126 265872
rect 481910 265860 481916 265872
rect 349120 265832 481916 265860
rect 349120 265820 349126 265832
rect 481910 265820 481916 265832
rect 481968 265820 481974 265872
rect 673178 265820 673184 265872
rect 673236 265860 673242 265872
rect 676030 265860 676036 265872
rect 673236 265832 676036 265860
rect 673236 265820 673242 265832
rect 676030 265820 676036 265832
rect 676088 265820 676094 265872
rect 343726 265752 343732 265804
rect 343784 265792 343790 265804
rect 467742 265792 467748 265804
rect 343784 265764 467748 265792
rect 343784 265752 343790 265764
rect 467742 265752 467748 265764
rect 467800 265752 467806 265804
rect 339770 265684 339776 265736
rect 339828 265724 339834 265736
rect 457070 265724 457076 265736
rect 339828 265696 457076 265724
rect 339828 265684 339834 265696
rect 457070 265684 457076 265696
rect 457128 265684 457134 265736
rect 333514 265616 333520 265668
rect 333572 265656 333578 265668
rect 440510 265656 440516 265668
rect 333572 265628 440516 265656
rect 333572 265616 333578 265628
rect 440510 265616 440516 265628
rect 440568 265616 440574 265668
rect 328178 265548 328184 265600
rect 328236 265588 328242 265600
rect 426342 265588 426348 265600
rect 328236 265560 426348 265588
rect 328236 265548 328242 265560
rect 426342 265548 426348 265560
rect 426400 265548 426406 265600
rect 324130 265480 324136 265532
rect 324188 265520 324194 265532
rect 415762 265520 415768 265532
rect 324188 265492 415768 265520
rect 324188 265480 324194 265492
rect 415762 265480 415768 265492
rect 415820 265480 415826 265532
rect 322842 265412 322848 265464
rect 322900 265452 322906 265464
rect 412174 265452 412180 265464
rect 322900 265424 412180 265452
rect 322900 265412 322906 265424
rect 412174 265412 412180 265424
rect 412232 265412 412238 265464
rect 319714 265344 319720 265396
rect 319772 265384 319778 265396
rect 403894 265384 403900 265396
rect 319772 265356 403900 265384
rect 319772 265344 319778 265356
rect 403894 265344 403900 265356
rect 403952 265344 403958 265396
rect 404262 265344 404268 265396
rect 404320 265384 404326 265396
rect 448882 265384 448888 265396
rect 404320 265356 448888 265384
rect 404320 265344 404326 265356
rect 448882 265344 448888 265356
rect 448940 265344 448946 265396
rect 318334 265276 318340 265328
rect 318392 265316 318398 265328
rect 400306 265316 400312 265328
rect 318392 265288 400312 265316
rect 318392 265276 318398 265288
rect 400306 265276 400312 265288
rect 400364 265276 400370 265328
rect 401594 265276 401600 265328
rect 401652 265316 401658 265328
rect 463326 265316 463332 265328
rect 401652 265288 463332 265316
rect 401652 265276 401658 265288
rect 463326 265276 463332 265288
rect 463384 265276 463390 265328
rect 314378 265208 314384 265260
rect 314436 265248 314442 265260
rect 314436 265220 353294 265248
rect 314436 265208 314442 265220
rect 353266 265180 353294 265220
rect 386874 265208 386880 265260
rect 386932 265248 386938 265260
rect 396810 265248 396816 265260
rect 386932 265220 396816 265248
rect 386932 265208 386938 265220
rect 396810 265208 396816 265220
rect 396868 265208 396874 265260
rect 389726 265180 389732 265192
rect 353266 265152 389732 265180
rect 389726 265140 389732 265152
rect 389784 265140 389790 265192
rect 673086 264936 673092 264988
rect 673144 264976 673150 264988
rect 676214 264976 676220 264988
rect 673144 264948 676220 264976
rect 673144 264936 673150 264948
rect 676214 264936 676220 264948
rect 676272 264936 676278 264988
rect 674282 264256 674288 264308
rect 674340 264296 674346 264308
rect 676030 264296 676036 264308
rect 674340 264268 676036 264296
rect 674340 264256 674346 264268
rect 676030 264256 676036 264268
rect 676088 264256 676094 264308
rect 674466 263032 674472 263084
rect 674524 263072 674530 263084
rect 676030 263072 676036 263084
rect 674524 263044 676036 263072
rect 674524 263032 674530 263044
rect 676030 263032 676036 263044
rect 676088 263032 676094 263084
rect 674926 262352 674932 262404
rect 674984 262392 674990 262404
rect 675938 262392 675944 262404
rect 674984 262364 675944 262392
rect 674984 262352 674990 262364
rect 675938 262352 675944 262364
rect 675996 262352 676002 262404
rect 673638 262284 673644 262336
rect 673696 262324 673702 262336
rect 676122 262324 676128 262336
rect 673696 262296 676128 262324
rect 673696 262284 673702 262296
rect 676122 262284 676128 262296
rect 676180 262284 676186 262336
rect 674558 262216 674564 262268
rect 674616 262256 674622 262268
rect 676030 262256 676036 262268
rect 674616 262228 676036 262256
rect 674616 262216 674622 262228
rect 676030 262216 676036 262228
rect 676088 262216 676094 262268
rect 673822 261400 673828 261452
rect 673880 261440 673886 261452
rect 676030 261440 676036 261452
rect 673880 261412 676036 261440
rect 673880 261400 673886 261412
rect 676030 261400 676036 261412
rect 676088 261400 676094 261452
rect 673454 260176 673460 260228
rect 673512 260216 673518 260228
rect 675938 260216 675944 260228
rect 673512 260188 675944 260216
rect 673512 260176 673518 260188
rect 675938 260176 675944 260188
rect 675996 260176 676002 260228
rect 675018 259768 675024 259820
rect 675076 259808 675082 259820
rect 676030 259808 676036 259820
rect 675076 259780 676036 259808
rect 675076 259768 675082 259780
rect 676030 259768 676036 259780
rect 676088 259768 676094 259820
rect 673546 259564 673552 259616
rect 673604 259604 673610 259616
rect 675938 259604 675944 259616
rect 673604 259576 675944 259604
rect 673604 259564 673610 259576
rect 675938 259564 675944 259576
rect 675996 259564 676002 259616
rect 674742 259496 674748 259548
rect 674800 259536 674806 259548
rect 676122 259536 676128 259548
rect 674800 259508 676128 259536
rect 674800 259496 674806 259508
rect 676122 259496 676128 259508
rect 676180 259496 676186 259548
rect 674834 259428 674840 259480
rect 674892 259468 674898 259480
rect 676030 259468 676036 259480
rect 674892 259440 676036 259468
rect 674892 259428 674898 259440
rect 676030 259428 676036 259440
rect 676088 259428 676094 259480
rect 41782 258816 41788 258868
rect 41840 258856 41846 258868
rect 43254 258856 43260 258868
rect 41840 258828 43260 258856
rect 41840 258816 41846 258828
rect 43254 258816 43260 258828
rect 43312 258816 43318 258868
rect 41874 257660 41880 257712
rect 41932 257700 41938 257712
rect 51258 257700 51264 257712
rect 41932 257672 51264 257700
rect 41932 257660 41938 257672
rect 51258 257660 51264 257672
rect 51316 257660 51322 257712
rect 41598 257524 41604 257576
rect 41656 257564 41662 257576
rect 46290 257564 46296 257576
rect 41656 257536 46296 257564
rect 41656 257524 41662 257536
rect 46290 257524 46296 257536
rect 46348 257524 46354 257576
rect 672902 256844 672908 256896
rect 672960 256884 672966 256896
rect 678974 256884 678980 256896
rect 672960 256856 678980 256884
rect 672960 256844 672966 256856
rect 678974 256844 678980 256856
rect 679032 256844 679038 256896
rect 673730 256776 673736 256828
rect 673788 256816 673794 256828
rect 676122 256816 676128 256828
rect 673788 256788 676128 256816
rect 673788 256776 673794 256788
rect 676122 256776 676128 256788
rect 676180 256776 676186 256828
rect 41506 256708 41512 256760
rect 41564 256748 41570 256760
rect 56502 256748 56508 256760
rect 41564 256720 56508 256748
rect 41564 256708 41570 256720
rect 56502 256708 56508 256720
rect 56560 256708 56566 256760
rect 674650 256708 674656 256760
rect 674708 256748 674714 256760
rect 676030 256748 676036 256760
rect 674708 256720 676036 256748
rect 674708 256708 674714 256720
rect 676030 256708 676036 256720
rect 676088 256708 676094 256760
rect 41506 256300 41512 256352
rect 41564 256340 41570 256352
rect 43714 256340 43720 256352
rect 41564 256312 43720 256340
rect 41564 256300 41570 256312
rect 43714 256300 43720 256312
rect 43772 256300 43778 256352
rect 41506 255688 41512 255740
rect 41564 255728 41570 255740
rect 43622 255728 43628 255740
rect 41564 255700 43628 255728
rect 41564 255688 41570 255700
rect 43622 255688 43628 255700
rect 43680 255688 43686 255740
rect 675110 255280 675116 255332
rect 675168 255320 675174 255332
rect 675754 255320 675760 255332
rect 675168 255292 675760 255320
rect 675168 255280 675174 255292
rect 675754 255280 675760 255292
rect 675812 255280 675818 255332
rect 41506 254872 41512 254924
rect 41564 254912 41570 254924
rect 43898 254912 43904 254924
rect 41564 254884 43904 254912
rect 41564 254872 41570 254884
rect 43898 254872 43904 254884
rect 43956 254872 43962 254924
rect 41874 254124 41880 254176
rect 41932 254164 41938 254176
rect 43898 254164 43904 254176
rect 41932 254136 43904 254164
rect 41932 254124 41938 254136
rect 43898 254124 43904 254136
rect 43956 254124 43962 254176
rect 41874 253988 41880 254040
rect 41932 254028 41938 254040
rect 43622 254028 43628 254040
rect 41932 254000 43628 254028
rect 41932 253988 41938 254000
rect 43622 253988 43628 254000
rect 43680 253988 43686 254040
rect 41782 253920 41788 253972
rect 41840 253960 41846 253972
rect 43162 253960 43168 253972
rect 41840 253932 43168 253960
rect 41840 253920 41846 253932
rect 43162 253920 43168 253932
rect 43220 253920 43226 253972
rect 675478 251336 675484 251388
rect 675536 251336 675542 251388
rect 675754 251336 675760 251388
rect 675812 251336 675818 251388
rect 416774 251200 416780 251252
rect 416832 251240 416838 251252
rect 567102 251240 567108 251252
rect 416832 251212 567108 251240
rect 416832 251200 416838 251212
rect 567102 251200 567108 251212
rect 567160 251200 567166 251252
rect 673362 250928 673368 250980
rect 673420 250968 673426 250980
rect 674926 250968 674932 250980
rect 673420 250940 674932 250968
rect 673420 250928 673426 250940
rect 674926 250928 674932 250940
rect 674984 250928 674990 250980
rect 675386 250928 675392 250980
rect 675444 250968 675450 250980
rect 675496 250968 675524 251336
rect 675444 250940 675524 250968
rect 675444 250928 675450 250940
rect 674926 250792 674932 250844
rect 674984 250832 674990 250844
rect 675478 250832 675484 250844
rect 674984 250804 675484 250832
rect 674984 250792 674990 250804
rect 675478 250792 675484 250804
rect 675536 250792 675542 250844
rect 675772 250232 675800 251336
rect 675754 250180 675760 250232
rect 675812 250180 675818 250232
rect 674466 249568 674472 249620
rect 674524 249608 674530 249620
rect 675386 249608 675392 249620
rect 674524 249580 675392 249608
rect 674524 249568 674530 249580
rect 675386 249568 675392 249580
rect 675444 249568 675450 249620
rect 673822 249432 673828 249484
rect 673880 249472 673886 249484
rect 674466 249472 674472 249484
rect 673880 249444 674472 249472
rect 673880 249432 673886 249444
rect 674466 249432 674472 249444
rect 674524 249432 674530 249484
rect 673362 249296 673368 249348
rect 673420 249336 673426 249348
rect 673822 249336 673828 249348
rect 673420 249308 673828 249336
rect 673420 249296 673426 249308
rect 673822 249296 673828 249308
rect 673880 249296 673886 249348
rect 416774 248412 416780 248464
rect 416832 248452 416838 248464
rect 567286 248452 567292 248464
rect 416832 248424 567292 248452
rect 416832 248412 416838 248424
rect 567286 248412 567292 248424
rect 567344 248412 567350 248464
rect 674558 247868 674564 247920
rect 674616 247908 674622 247920
rect 675386 247908 675392 247920
rect 674616 247880 675392 247908
rect 674616 247868 674622 247880
rect 675386 247868 675392 247880
rect 675444 247868 675450 247920
rect 41506 247664 41512 247716
rect 41564 247704 41570 247716
rect 46290 247704 46296 247716
rect 41564 247676 46296 247704
rect 41564 247664 41570 247676
rect 46290 247664 46296 247676
rect 46348 247664 46354 247716
rect 41506 247256 41512 247308
rect 41564 247296 41570 247308
rect 45646 247296 45652 247308
rect 41564 247268 45652 247296
rect 41564 247256 41570 247268
rect 45646 247256 45652 247268
rect 45704 247256 45710 247308
rect 675018 247256 675024 247308
rect 675076 247296 675082 247308
rect 675076 247268 675432 247296
rect 675076 247256 675082 247268
rect 674650 247120 674656 247172
rect 674708 247160 674714 247172
rect 675018 247160 675024 247172
rect 674708 247132 675024 247160
rect 674708 247120 674714 247132
rect 675018 247120 675024 247132
rect 675076 247120 675082 247172
rect 675404 247104 675432 247268
rect 675386 247052 675392 247104
rect 675444 247052 675450 247104
rect 674742 246508 674748 246560
rect 674800 246548 674806 246560
rect 675386 246548 675392 246560
rect 674800 246520 675392 246548
rect 674800 246508 674806 246520
rect 675386 246508 675392 246520
rect 675444 246508 675450 246560
rect 41506 246440 41512 246492
rect 41564 246480 41570 246492
rect 48866 246480 48872 246492
rect 41564 246452 48872 246480
rect 41564 246440 41570 246452
rect 48866 246440 48872 246452
rect 48924 246440 48930 246492
rect 180702 246440 180708 246492
rect 180760 246480 180766 246492
rect 184842 246480 184848 246492
rect 180760 246452 184848 246480
rect 180760 246440 180766 246452
rect 184842 246440 184848 246452
rect 184900 246440 184906 246492
rect 673638 246372 673644 246424
rect 673696 246412 673702 246424
rect 674742 246412 674748 246424
rect 673696 246384 674748 246412
rect 673696 246372 673702 246384
rect 674742 246372 674748 246384
rect 674800 246372 674806 246424
rect 673638 246236 673644 246288
rect 673696 246276 673702 246288
rect 673822 246276 673828 246288
rect 673696 246248 673828 246276
rect 673696 246236 673702 246248
rect 673822 246236 673828 246248
rect 673880 246236 673886 246288
rect 674282 246100 674288 246152
rect 674340 246140 674346 246152
rect 675202 246140 675208 246152
rect 674340 246112 675208 246140
rect 674340 246100 674346 246112
rect 675202 246100 675208 246112
rect 675260 246100 675266 246152
rect 674834 246032 674840 246084
rect 674892 246072 674898 246084
rect 675386 246072 675392 246084
rect 674892 246044 675392 246072
rect 674892 246032 674898 246044
rect 675386 246032 675392 246044
rect 675444 246032 675450 246084
rect 416774 245624 416780 245676
rect 416832 245664 416838 245676
rect 564342 245664 564348 245676
rect 416832 245636 564348 245664
rect 416832 245624 416838 245636
rect 564342 245624 564348 245636
rect 564400 245624 564406 245676
rect 41690 245556 41696 245608
rect 41748 245596 41754 245608
rect 42702 245596 42708 245608
rect 41748 245568 42708 245596
rect 41748 245556 41754 245568
rect 42702 245556 42708 245568
rect 42760 245556 42766 245608
rect 655698 245556 655704 245608
rect 655756 245596 655762 245608
rect 674926 245596 674932 245608
rect 655756 245568 674932 245596
rect 655756 245556 655762 245568
rect 674926 245556 674932 245568
rect 674984 245556 674990 245608
rect 41874 245080 41880 245132
rect 41932 245120 41938 245132
rect 43530 245120 43536 245132
rect 41932 245092 43536 245120
rect 41932 245080 41938 245092
rect 43530 245080 43536 245092
rect 43588 245080 43594 245132
rect 41782 244604 41788 244656
rect 41840 244644 41846 244656
rect 43346 244644 43352 244656
rect 41840 244616 43352 244644
rect 41840 244604 41846 244616
rect 43346 244604 43352 244616
rect 43404 244604 43410 244656
rect 673638 243584 673644 243636
rect 673696 243624 673702 243636
rect 675386 243624 675392 243636
rect 673696 243596 675392 243624
rect 673696 243584 673702 243596
rect 675386 243584 675392 243596
rect 675444 243584 675450 243636
rect 41322 242836 41328 242888
rect 41380 242876 41386 242888
rect 43254 242876 43260 242888
rect 41380 242848 43260 242876
rect 41380 242836 41386 242848
rect 43254 242836 43260 242848
rect 43312 242836 43318 242888
rect 41414 242768 41420 242820
rect 41472 242808 41478 242820
rect 43070 242808 43076 242820
rect 41472 242780 43076 242808
rect 41472 242768 41478 242780
rect 43070 242768 43076 242780
rect 43128 242768 43134 242820
rect 675018 242768 675024 242820
rect 675076 242808 675082 242820
rect 675386 242808 675392 242820
rect 675076 242780 675392 242808
rect 675076 242768 675082 242780
rect 675386 242768 675392 242780
rect 675444 242768 675450 242820
rect 41230 242700 41236 242752
rect 41288 242740 41294 242752
rect 42242 242740 42248 242752
rect 41288 242712 42248 242740
rect 41288 242700 41294 242712
rect 42242 242700 42248 242712
rect 42300 242700 42306 242752
rect 41598 242632 41604 242684
rect 41656 242672 41662 242684
rect 43438 242672 43444 242684
rect 41656 242644 43444 242672
rect 41656 242632 41662 242644
rect 43438 242632 43444 242644
rect 43496 242632 43502 242684
rect 38562 242564 38568 242616
rect 38620 242604 38626 242616
rect 43714 242604 43720 242616
rect 38620 242576 43720 242604
rect 38620 242564 38626 242576
rect 43714 242564 43720 242576
rect 43772 242564 43778 242616
rect 38470 242496 38476 242548
rect 38528 242536 38534 242548
rect 43806 242536 43812 242548
rect 38528 242508 43812 242536
rect 38528 242496 38534 242508
rect 43806 242496 43812 242508
rect 43864 242496 43870 242548
rect 35802 242428 35808 242480
rect 35860 242468 35866 242480
rect 43990 242468 43996 242480
rect 35860 242440 43996 242468
rect 35860 242428 35866 242440
rect 43990 242428 43996 242440
rect 44048 242428 44054 242480
rect 673546 242156 673552 242208
rect 673604 242196 673610 242208
rect 675386 242196 675392 242208
rect 673604 242168 675392 242196
rect 673604 242156 673610 242168
rect 675386 242156 675392 242168
rect 675444 242156 675450 242208
rect 673730 241748 673736 241800
rect 673788 241788 673794 241800
rect 675386 241788 675392 241800
rect 673788 241760 675392 241788
rect 673788 241748 673794 241760
rect 675386 241748 675392 241760
rect 675444 241748 675450 241800
rect 41138 240932 41144 240984
rect 41196 240972 41202 240984
rect 41196 240944 41828 240972
rect 41196 240932 41202 240944
rect 41800 240372 41828 240944
rect 673454 240524 673460 240576
rect 673512 240564 673518 240576
rect 675386 240564 675392 240576
rect 673512 240536 675392 240564
rect 673512 240524 673518 240536
rect 675386 240524 675392 240536
rect 675444 240524 675450 240576
rect 41782 240320 41788 240372
rect 41840 240320 41846 240372
rect 674742 238688 674748 238740
rect 674800 238728 674806 238740
rect 675386 238728 675392 238740
rect 674800 238700 675392 238728
rect 674800 238688 674806 238700
rect 675386 238688 675392 238700
rect 675444 238688 675450 238740
rect 42150 238484 42156 238536
rect 42208 238524 42214 238536
rect 42702 238524 42708 238536
rect 42208 238496 42708 238524
rect 42208 238484 42214 238496
rect 42702 238484 42708 238496
rect 42760 238484 42766 238536
rect 43530 237940 43536 237992
rect 43588 237980 43594 237992
rect 43898 237980 43904 237992
rect 43588 237952 43904 237980
rect 43588 237940 43594 237952
rect 43898 237940 43904 237952
rect 43956 237940 43962 237992
rect 184934 237436 184940 237448
rect 179432 237408 184940 237436
rect 177942 237328 177948 237380
rect 178000 237368 178006 237380
rect 179432 237368 179460 237408
rect 184934 237396 184940 237408
rect 184992 237396 184998 237448
rect 178000 237340 179460 237368
rect 178000 237328 178006 237340
rect 674466 236852 674472 236904
rect 674524 236892 674530 236904
rect 675386 236892 675392 236904
rect 674524 236864 675392 236892
rect 674524 236852 674530 236864
rect 675386 236852 675392 236864
rect 675444 236852 675450 236904
rect 42242 236036 42248 236088
rect 42300 236076 42306 236088
rect 43254 236076 43260 236088
rect 42300 236048 43260 236076
rect 42300 236036 42306 236048
rect 43254 236036 43260 236048
rect 43312 236036 43318 236088
rect 675018 235560 675024 235612
rect 675076 235600 675082 235612
rect 675754 235600 675760 235612
rect 675076 235572 675760 235600
rect 675076 235560 675082 235572
rect 675754 235560 675760 235572
rect 675812 235560 675818 235612
rect 42334 234200 42340 234252
rect 42392 234240 42398 234252
rect 43070 234240 43076 234252
rect 42392 234212 43076 234240
rect 42392 234200 42398 234212
rect 43070 234200 43076 234212
rect 43128 234200 43134 234252
rect 42150 233316 42156 233368
rect 42208 233356 42214 233368
rect 43346 233356 43352 233368
rect 42208 233328 43352 233356
rect 42208 233316 42214 233328
rect 43346 233316 43352 233328
rect 43404 233316 43410 233368
rect 74442 232500 74448 232552
rect 74500 232540 74506 232552
rect 177942 232540 177948 232552
rect 74500 232512 177948 232540
rect 74500 232500 74506 232512
rect 177942 232500 177948 232512
rect 178000 232500 178006 232552
rect 42426 232296 42432 232348
rect 42484 232336 42490 232348
rect 43438 232336 43444 232348
rect 42484 232308 43444 232336
rect 42484 232296 42490 232308
rect 43438 232296 43444 232308
rect 43496 232296 43502 232348
rect 46014 230936 46020 230988
rect 46072 230976 46078 230988
rect 654134 230976 654140 230988
rect 46072 230948 654140 230976
rect 46072 230936 46078 230948
rect 654134 230936 654140 230948
rect 654192 230936 654198 230988
rect 48314 230868 48320 230920
rect 48372 230908 48378 230920
rect 656986 230908 656992 230920
rect 48372 230880 656992 230908
rect 48372 230868 48378 230880
rect 656986 230868 656992 230880
rect 657044 230868 657050 230920
rect 48222 230800 48228 230852
rect 48280 230840 48286 230852
rect 656894 230840 656900 230852
rect 48280 230812 656900 230840
rect 48280 230800 48286 230812
rect 656894 230800 656900 230812
rect 656952 230800 656958 230852
rect 48590 230732 48596 230784
rect 48648 230772 48654 230784
rect 659654 230772 659660 230784
rect 48648 230744 659660 230772
rect 48648 230732 48654 230744
rect 659654 230732 659660 230744
rect 659712 230732 659718 230784
rect 51166 230664 51172 230716
rect 51224 230704 51230 230716
rect 662782 230704 662788 230716
rect 51224 230676 662788 230704
rect 51224 230664 51230 230676
rect 662782 230664 662788 230676
rect 662840 230664 662846 230716
rect 51074 230596 51080 230648
rect 51132 230636 51138 230648
rect 662874 230636 662880 230648
rect 51132 230608 662880 230636
rect 51132 230596 51138 230608
rect 662874 230596 662880 230608
rect 662932 230596 662938 230648
rect 42426 230528 42432 230580
rect 42484 230568 42490 230580
rect 43806 230568 43812 230580
rect 42484 230540 43812 230568
rect 42484 230528 42490 230540
rect 43806 230528 43812 230540
rect 43864 230528 43870 230580
rect 48406 230528 48412 230580
rect 48464 230568 48470 230580
rect 659746 230568 659752 230580
rect 48464 230540 659752 230568
rect 48464 230528 48470 230540
rect 659746 230528 659752 230540
rect 659804 230528 659810 230580
rect 48774 230460 48780 230512
rect 48832 230500 48838 230512
rect 662598 230500 662604 230512
rect 48832 230472 662604 230500
rect 48832 230460 48838 230472
rect 662598 230460 662604 230472
rect 662656 230460 662662 230512
rect 48866 230392 48872 230444
rect 48924 230432 48930 230444
rect 662690 230432 662696 230444
rect 48924 230404 662696 230432
rect 48924 230392 48930 230404
rect 662690 230392 662696 230404
rect 662748 230392 662754 230444
rect 42150 230324 42156 230376
rect 42208 230364 42214 230376
rect 43714 230364 43720 230376
rect 42208 230336 43720 230364
rect 42208 230324 42214 230336
rect 43714 230324 43720 230336
rect 43772 230324 43778 230376
rect 350166 230188 350172 230240
rect 350224 230228 350230 230240
rect 423858 230228 423864 230240
rect 350224 230200 423864 230228
rect 350224 230188 350230 230200
rect 423858 230188 423864 230200
rect 423916 230188 423922 230240
rect 348786 230120 348792 230172
rect 348844 230160 348850 230172
rect 420454 230160 420460 230172
rect 348844 230132 420460 230160
rect 348844 230120 348850 230132
rect 420454 230120 420460 230132
rect 420512 230120 420518 230172
rect 345934 230052 345940 230104
rect 345992 230092 345998 230104
rect 414014 230092 414020 230104
rect 345992 230064 414020 230092
rect 345992 230052 345998 230064
rect 414014 230052 414020 230064
rect 414072 230052 414078 230104
rect 351638 229984 351644 230036
rect 351696 230024 351702 230036
rect 427170 230024 427176 230036
rect 351696 229996 427176 230024
rect 351696 229984 351702 229996
rect 427170 229984 427176 229996
rect 427228 229984 427234 230036
rect 354490 229916 354496 229968
rect 354548 229956 354554 229968
rect 433886 229956 433892 229968
rect 354548 229928 433892 229956
rect 354548 229916 354554 229928
rect 433886 229916 433892 229928
rect 433944 229916 433950 229968
rect 353018 229848 353024 229900
rect 353076 229888 353082 229900
rect 430574 229888 430580 229900
rect 353076 229860 430580 229888
rect 353076 229848 353082 229860
rect 430574 229848 430580 229860
rect 430632 229848 430638 229900
rect 357342 229780 357348 229832
rect 357400 229820 357406 229832
rect 440694 229820 440700 229832
rect 357400 229792 440700 229820
rect 357400 229780 357406 229792
rect 440694 229780 440700 229792
rect 440752 229780 440758 229832
rect 359826 229712 359832 229764
rect 359884 229752 359890 229764
rect 445662 229752 445668 229764
rect 359884 229724 445668 229752
rect 359884 229712 359890 229724
rect 445662 229712 445668 229724
rect 445720 229712 445726 229764
rect 360194 229644 360200 229696
rect 360252 229684 360258 229696
rect 447410 229684 447416 229696
rect 360252 229656 447416 229684
rect 360252 229644 360258 229656
rect 447410 229644 447416 229656
rect 447468 229644 447474 229696
rect 364426 229576 364432 229628
rect 364484 229616 364490 229628
rect 457438 229616 457444 229628
rect 364484 229588 457444 229616
rect 364484 229576 364490 229588
rect 457438 229576 457444 229588
rect 457496 229576 457502 229628
rect 365530 229508 365536 229560
rect 365588 229548 365594 229560
rect 459186 229548 459192 229560
rect 365588 229520 459192 229548
rect 365588 229508 365594 229520
rect 459186 229508 459192 229520
rect 459244 229508 459250 229560
rect 364058 229440 364064 229492
rect 364116 229480 364122 229492
rect 455782 229480 455788 229492
rect 364116 229452 455788 229480
rect 364116 229440 364122 229452
rect 455782 229440 455788 229452
rect 455840 229440 455846 229492
rect 370130 229372 370136 229424
rect 370188 229412 370194 229424
rect 470962 229412 470968 229424
rect 370188 229384 470968 229412
rect 370188 229372 370194 229384
rect 470962 229372 470968 229384
rect 471020 229372 471026 229424
rect 371234 229304 371240 229356
rect 371292 229344 371298 229356
rect 472618 229344 472624 229356
rect 371292 229316 472624 229344
rect 371292 229304 371298 229316
rect 472618 229304 472624 229316
rect 472676 229304 472682 229356
rect 374822 229236 374828 229288
rect 374880 229276 374886 229288
rect 483014 229276 483020 229288
rect 374880 229248 483020 229276
rect 374880 229236 374886 229248
rect 483014 229236 483020 229248
rect 483072 229236 483078 229288
rect 388346 229168 388352 229220
rect 388404 229208 388410 229220
rect 515490 229208 515496 229220
rect 388404 229180 515496 229208
rect 388404 229168 388410 229180
rect 515490 229168 515496 229180
rect 515548 229168 515554 229220
rect 74442 229140 74448 229152
rect 66272 229112 74448 229140
rect 63494 229032 63500 229084
rect 63552 229072 63558 229084
rect 66272 229072 66300 229112
rect 74442 229100 74448 229112
rect 74500 229100 74506 229152
rect 396902 229100 396908 229152
rect 396960 229140 396966 229152
rect 535454 229140 535460 229152
rect 396960 229112 535460 229140
rect 396960 229100 396966 229112
rect 535454 229100 535460 229112
rect 535512 229100 535518 229152
rect 63552 229044 66300 229072
rect 63552 229032 63558 229044
rect 156966 229032 156972 229084
rect 157024 229072 157030 229084
rect 237190 229072 237196 229084
rect 157024 229044 237196 229072
rect 157024 229032 157030 229044
rect 237190 229032 237196 229044
rect 237248 229032 237254 229084
rect 256970 229032 256976 229084
rect 257028 229072 257034 229084
rect 264606 229072 264612 229084
rect 257028 229044 264612 229072
rect 257028 229032 257034 229044
rect 264606 229032 264612 229044
rect 264664 229032 264670 229084
rect 264698 229032 264704 229084
rect 264756 229072 264762 229084
rect 273898 229072 273904 229084
rect 264756 229044 273904 229072
rect 264756 229032 264762 229044
rect 273898 229032 273904 229044
rect 273956 229032 273962 229084
rect 296346 229032 296352 229084
rect 296404 229072 296410 229084
rect 298462 229072 298468 229084
rect 296404 229044 298468 229072
rect 296404 229032 296410 229044
rect 298462 229032 298468 229044
rect 298520 229032 298526 229084
rect 306650 229032 306656 229084
rect 306708 229072 306714 229084
rect 323854 229072 323860 229084
rect 306708 229044 323860 229072
rect 306708 229032 306714 229044
rect 323854 229032 323860 229044
rect 323912 229032 323918 229084
rect 338022 229032 338028 229084
rect 338080 229072 338086 229084
rect 373902 229072 373908 229084
rect 338080 229044 373908 229072
rect 338080 229032 338086 229044
rect 373902 229032 373908 229044
rect 373960 229032 373966 229084
rect 389726 229032 389732 229084
rect 389784 229072 389790 229084
rect 469122 229072 469128 229084
rect 389784 229044 469128 229072
rect 389784 229032 389790 229044
rect 469122 229032 469128 229044
rect 469180 229032 469186 229084
rect 152826 228964 152832 229016
rect 152884 229004 152890 229016
rect 233970 229004 233976 229016
rect 152884 228976 233976 229004
rect 152884 228964 152890 228976
rect 233970 228964 233976 228976
rect 234028 228964 234034 229016
rect 239858 228964 239864 229016
rect 239916 229004 239922 229016
rect 265342 229004 265348 229016
rect 239916 228976 265348 229004
rect 239916 228964 239922 228976
rect 265342 228964 265348 228976
rect 265400 228964 265406 229016
rect 290734 228964 290740 229016
rect 290792 229004 290798 229016
rect 292390 229004 292396 229016
rect 290792 228976 292396 229004
rect 290792 228964 290798 228976
rect 292390 228964 292396 228976
rect 292448 228964 292454 229016
rect 293218 228964 293224 229016
rect 293276 229004 293282 229016
rect 294598 229004 294604 229016
rect 293276 228976 294604 229004
rect 293276 228964 293282 228976
rect 294598 228964 294604 228976
rect 294656 228964 294662 229016
rect 297450 228964 297456 229016
rect 297508 229004 297514 229016
rect 299382 229004 299388 229016
rect 297508 228976 299388 229004
rect 297508 228964 297514 228976
rect 299382 228964 299388 228976
rect 299440 228964 299446 229016
rect 304166 228964 304172 229016
rect 304224 229004 304230 229016
rect 314654 229004 314660 229016
rect 304224 228976 314660 229004
rect 304224 228964 304230 228976
rect 314654 228964 314660 228976
rect 314712 228964 314718 229016
rect 321646 228964 321652 229016
rect 321704 229004 321710 229016
rect 340690 229004 340696 229016
rect 321704 228976 340696 229004
rect 321704 228964 321710 228976
rect 340690 228964 340696 228976
rect 340748 228964 340754 229016
rect 342346 228964 342352 229016
rect 342404 229004 342410 229016
rect 362954 229004 362960 229016
rect 342404 228976 362960 229004
rect 342404 228964 342410 228976
rect 362954 228964 362960 228976
rect 363012 228964 363018 229016
rect 363046 228964 363052 229016
rect 363104 229004 363110 229016
rect 365898 229004 365904 229016
rect 363104 228976 365904 229004
rect 363104 228964 363110 228976
rect 365898 228964 365904 228976
rect 365956 228964 365962 229016
rect 391934 228964 391940 229016
rect 391992 229004 391998 229016
rect 472066 229004 472072 229016
rect 391992 228976 472072 229004
rect 391992 228964 391998 228976
rect 472066 228964 472072 228976
rect 472124 228964 472130 229016
rect 156138 228896 156144 228948
rect 156196 228936 156202 228948
rect 235350 228936 235356 228948
rect 156196 228908 235356 228936
rect 156196 228896 156202 228908
rect 235350 228896 235356 228908
rect 235408 228896 235414 228948
rect 240318 228896 240324 228948
rect 240376 228936 240382 228948
rect 269574 228936 269580 228948
rect 240376 228908 269580 228936
rect 240376 228896 240382 228908
rect 269574 228896 269580 228908
rect 269632 228896 269638 228948
rect 304534 228896 304540 228948
rect 304592 228936 304598 228948
rect 316126 228936 316132 228948
rect 304592 228908 316132 228936
rect 304592 228896 304598 228908
rect 316126 228896 316132 228908
rect 316184 228896 316190 228948
rect 342714 228896 342720 228948
rect 342772 228936 342778 228948
rect 380986 228936 380992 228948
rect 342772 228908 380992 228936
rect 342772 228896 342778 228908
rect 380986 228896 380992 228908
rect 381044 228896 381050 228948
rect 398282 228896 398288 228948
rect 398340 228936 398346 228948
rect 477494 228936 477500 228948
rect 398340 228908 477500 228936
rect 398340 228896 398346 228908
rect 477494 228896 477500 228908
rect 477552 228896 477558 228948
rect 150250 228828 150256 228880
rect 150308 228868 150314 228880
rect 234338 228868 234344 228880
rect 150308 228840 234344 228868
rect 150308 228828 150314 228840
rect 234338 228828 234344 228840
rect 234396 228828 234402 228880
rect 239950 228828 239956 228880
rect 240008 228868 240014 228880
rect 266722 228868 266728 228880
rect 240008 228840 266728 228868
rect 240008 228828 240014 228840
rect 266722 228828 266728 228840
rect 266780 228828 266786 228880
rect 305638 228828 305644 228880
rect 305696 228868 305702 228880
rect 317874 228868 317880 228880
rect 305696 228840 317880 228868
rect 305696 228828 305702 228840
rect 317874 228828 317880 228840
rect 317932 228828 317938 228880
rect 340874 228828 340880 228880
rect 340932 228868 340938 228880
rect 380894 228868 380900 228880
rect 340932 228840 380900 228868
rect 340932 228828 340938 228840
rect 380894 228828 380900 228840
rect 380952 228828 380958 228880
rect 396166 228828 396172 228880
rect 396224 228868 396230 228880
rect 474826 228868 474832 228880
rect 396224 228840 474832 228868
rect 396224 228828 396230 228840
rect 474826 228828 474832 228840
rect 474884 228828 474890 228880
rect 121178 228760 121184 228812
rect 121236 228800 121242 228812
rect 203334 228800 203340 228812
rect 121236 228772 203340 228800
rect 121236 228760 121242 228772
rect 203334 228760 203340 228772
rect 203392 228760 203398 228812
rect 209590 228760 209596 228812
rect 209648 228800 209654 228812
rect 258166 228800 258172 228812
rect 209648 228772 258172 228800
rect 209648 228760 209654 228772
rect 258166 228760 258172 228772
rect 258224 228760 258230 228812
rect 258258 228760 258264 228812
rect 258316 228800 258322 228812
rect 277486 228800 277492 228812
rect 258316 228772 277492 228800
rect 258316 228760 258322 228772
rect 277486 228760 277492 228772
rect 277544 228760 277550 228812
rect 306006 228760 306012 228812
rect 306064 228800 306070 228812
rect 319530 228800 319536 228812
rect 306064 228772 319536 228800
rect 306064 228760 306070 228772
rect 319530 228760 319536 228772
rect 319588 228760 319594 228812
rect 337746 228760 337752 228812
rect 337804 228800 337810 228812
rect 383746 228800 383752 228812
rect 337804 228772 383752 228800
rect 337804 228760 337810 228772
rect 383746 228760 383752 228772
rect 383804 228760 383810 228812
rect 394050 228760 394056 228812
rect 394108 228800 394114 228812
rect 474734 228800 474740 228812
rect 394108 228772 474740 228800
rect 394108 228760 394114 228772
rect 474734 228760 474740 228772
rect 474792 228760 474798 228812
rect 151722 228692 151728 228744
rect 151780 228732 151786 228744
rect 234706 228732 234712 228744
rect 151780 228704 234712 228732
rect 151780 228692 151786 228704
rect 234706 228692 234712 228704
rect 234764 228692 234770 228744
rect 241974 228692 241980 228744
rect 242032 228732 242038 228744
rect 272150 228732 272156 228744
rect 242032 228704 272156 228732
rect 242032 228692 242038 228704
rect 272150 228692 272156 228704
rect 272208 228692 272214 228744
rect 298830 228692 298836 228744
rect 298888 228732 298894 228744
rect 302694 228732 302700 228744
rect 298888 228704 302700 228732
rect 298888 228692 298894 228704
rect 302694 228692 302700 228704
rect 302752 228692 302758 228744
rect 305270 228692 305276 228744
rect 305328 228732 305334 228744
rect 320358 228732 320364 228744
rect 305328 228704 320364 228732
rect 305328 228692 305334 228704
rect 320358 228692 320364 228704
rect 320416 228692 320422 228744
rect 322014 228692 322020 228744
rect 322072 228732 322078 228744
rect 359090 228732 359096 228744
rect 322072 228704 359096 228732
rect 322072 228692 322078 228704
rect 359090 228692 359096 228704
rect 359148 228692 359154 228744
rect 376570 228692 376576 228744
rect 376628 228732 376634 228744
rect 466362 228732 466368 228744
rect 376628 228704 466368 228732
rect 376628 228692 376634 228704
rect 466362 228692 466368 228704
rect 466420 228692 466426 228744
rect 146018 228624 146024 228676
rect 146076 228664 146082 228676
rect 231118 228664 231124 228676
rect 146076 228636 231124 228664
rect 146076 228624 146082 228636
rect 231118 228624 231124 228636
rect 231176 228624 231182 228676
rect 245286 228624 245292 228676
rect 245344 228664 245350 228676
rect 273530 228664 273536 228676
rect 245344 228636 273536 228664
rect 245344 228624 245350 228636
rect 273530 228624 273536 228636
rect 273588 228624 273594 228676
rect 308858 228624 308864 228676
rect 308916 228664 308922 228676
rect 316218 228664 316224 228676
rect 308916 228636 316224 228664
rect 308916 228624 308922 228636
rect 316218 228624 316224 228636
rect 316276 228624 316282 228676
rect 328822 228624 328828 228676
rect 328880 228664 328886 228676
rect 345934 228664 345940 228676
rect 328880 228636 345940 228664
rect 328880 228624 328886 228636
rect 345934 228624 345940 228636
rect 345992 228624 345998 228676
rect 375466 228624 375472 228676
rect 375524 228664 375530 228676
rect 484394 228664 484400 228676
rect 375524 228636 484400 228664
rect 375524 228624 375530 228636
rect 484394 228624 484400 228636
rect 484452 228624 484458 228676
rect 145190 228556 145196 228608
rect 145248 228596 145254 228608
rect 231854 228596 231860 228608
rect 145248 228568 231860 228596
rect 145248 228556 145254 228568
rect 231854 228556 231860 228568
rect 231912 228556 231918 228608
rect 238478 228556 238484 228608
rect 238536 228596 238542 228608
rect 268194 228596 268200 228608
rect 238536 228568 268200 228596
rect 238536 228556 238542 228568
rect 268194 228556 268200 228568
rect 268252 228556 268258 228608
rect 307386 228556 307392 228608
rect 307444 228596 307450 228608
rect 322934 228596 322940 228608
rect 307444 228568 322940 228596
rect 307444 228556 307450 228568
rect 322934 228556 322940 228568
rect 322992 228556 322998 228608
rect 336642 228556 336648 228608
rect 336700 228596 336706 228608
rect 376662 228596 376668 228608
rect 336700 228568 376668 228596
rect 336700 228556 336706 228568
rect 376662 228556 376668 228568
rect 376720 228556 376726 228608
rect 379422 228556 379428 228608
rect 379480 228596 379486 228608
rect 494514 228596 494520 228608
rect 379480 228568 494520 228596
rect 379480 228556 379486 228568
rect 494514 228556 494520 228568
rect 494572 228556 494578 228608
rect 138474 228488 138480 228540
rect 138532 228528 138538 228540
rect 229002 228528 229008 228540
rect 138532 228500 229008 228528
rect 138532 228488 138538 228500
rect 229002 228488 229008 228500
rect 229060 228488 229066 228540
rect 240134 228488 240140 228540
rect 240192 228528 240198 228540
rect 271046 228528 271052 228540
rect 240192 228500 271052 228528
rect 240192 228488 240198 228500
rect 271046 228488 271052 228500
rect 271104 228488 271110 228540
rect 307754 228488 307760 228540
rect 307812 228528 307818 228540
rect 325694 228528 325700 228540
rect 307812 228500 325700 228528
rect 307812 228488 307818 228500
rect 325694 228488 325700 228500
rect 325752 228488 325758 228540
rect 329190 228488 329196 228540
rect 329248 228528 329254 228540
rect 375926 228528 375932 228540
rect 329248 228500 375932 228528
rect 329248 228488 329254 228500
rect 375926 228488 375932 228500
rect 375984 228488 375990 228540
rect 384390 228488 384396 228540
rect 384448 228528 384454 228540
rect 506290 228528 506296 228540
rect 384448 228500 506296 228528
rect 384448 228488 384454 228500
rect 506290 228488 506296 228500
rect 506348 228488 506354 228540
rect 143442 228420 143448 228472
rect 143500 228460 143506 228472
rect 231486 228460 231492 228472
rect 143500 228432 231492 228460
rect 143500 228420 143506 228432
rect 231486 228420 231492 228432
rect 231544 228420 231550 228472
rect 235258 228420 235264 228472
rect 235316 228460 235322 228472
rect 269298 228460 269304 228472
rect 235316 228432 269304 228460
rect 235316 228420 235322 228432
rect 269298 228420 269304 228432
rect 269356 228420 269362 228472
rect 310238 228420 310244 228472
rect 310296 228460 310302 228472
rect 329650 228460 329656 228472
rect 310296 228432 329656 228460
rect 310296 228420 310302 228432
rect 329650 228420 329656 228432
rect 329708 228420 329714 228472
rect 362954 228420 362960 228472
rect 363012 228460 363018 228472
rect 378226 228460 378232 228472
rect 363012 228432 378232 228460
rect 363012 228420 363018 228432
rect 378226 228420 378232 228432
rect 378284 228420 378290 228472
rect 386506 228420 386512 228472
rect 386564 228460 386570 228472
rect 511350 228460 511356 228472
rect 386564 228432 511356 228460
rect 386564 228420 386570 228432
rect 511350 228420 511356 228432
rect 511408 228420 511414 228472
rect 136818 228352 136824 228404
rect 136876 228392 136882 228404
rect 228634 228392 228640 228404
rect 136876 228364 228640 228392
rect 136876 228352 136882 228364
rect 228634 228352 228640 228364
rect 228692 228352 228698 228404
rect 229278 228352 229284 228404
rect 229336 228392 229342 228404
rect 267458 228392 267464 228404
rect 229336 228364 267464 228392
rect 229336 228352 229342 228364
rect 267458 228352 267464 228364
rect 267516 228352 267522 228404
rect 298738 228352 298744 228404
rect 298796 228392 298802 228404
rect 301038 228392 301044 228404
rect 298796 228364 301044 228392
rect 298796 228352 298802 228364
rect 301038 228352 301044 228364
rect 301096 228352 301102 228404
rect 308122 228352 308128 228404
rect 308180 228392 308186 228404
rect 327074 228392 327080 228404
rect 308180 228364 327080 228392
rect 308180 228352 308186 228364
rect 327074 228352 327080 228364
rect 327132 228352 327138 228404
rect 333422 228352 333428 228404
rect 333480 228392 333486 228404
rect 385954 228392 385960 228404
rect 333480 228364 385960 228392
rect 333480 228352 333486 228364
rect 385954 228352 385960 228364
rect 386012 228352 386018 228404
rect 400490 228352 400496 228404
rect 400548 228392 400554 228404
rect 544102 228392 544108 228404
rect 400548 228364 544108 228392
rect 400548 228352 400554 228364
rect 544102 228352 544108 228364
rect 544160 228352 544166 228404
rect 130102 228284 130108 228336
rect 130160 228324 130166 228336
rect 225782 228324 225788 228336
rect 130160 228296 225788 228324
rect 130160 228284 130166 228296
rect 225782 228284 225788 228296
rect 225840 228284 225846 228336
rect 238570 228284 238576 228336
rect 238628 228324 238634 228336
rect 270678 228324 270684 228336
rect 238628 228296 270684 228324
rect 238628 228284 238634 228296
rect 270678 228284 270684 228296
rect 270736 228284 270742 228336
rect 309502 228284 309508 228336
rect 309560 228324 309566 228336
rect 330478 228324 330484 228336
rect 309560 228296 330484 228324
rect 309560 228284 309566 228296
rect 330478 228284 330484 228296
rect 330536 228284 330542 228336
rect 334894 228284 334900 228336
rect 334952 228324 334958 228336
rect 389082 228324 389088 228336
rect 334952 228296 389088 228324
rect 334952 228284 334958 228296
rect 389082 228284 389088 228296
rect 389140 228284 389146 228336
rect 401870 228284 401876 228336
rect 401928 228324 401934 228336
rect 547782 228324 547788 228336
rect 401928 228296 547788 228324
rect 401928 228284 401934 228296
rect 547782 228284 547788 228296
rect 547840 228284 547846 228336
rect 125042 228216 125048 228268
rect 125100 228256 125106 228268
rect 223298 228256 223304 228268
rect 125100 228228 223304 228256
rect 125100 228216 125106 228228
rect 223298 228216 223304 228228
rect 223356 228216 223362 228268
rect 227714 228216 227720 228268
rect 227772 228256 227778 228268
rect 267090 228256 267096 228268
rect 227772 228228 267096 228256
rect 227772 228216 227778 228228
rect 267090 228216 267096 228228
rect 267148 228216 267154 228268
rect 296714 228216 296720 228268
rect 296772 228256 296778 228268
rect 300210 228256 300216 228268
rect 296772 228228 300216 228256
rect 296772 228216 296778 228228
rect 300210 228216 300216 228228
rect 300268 228216 300274 228268
rect 302786 228216 302792 228268
rect 302844 228256 302850 228268
rect 311158 228256 311164 228268
rect 302844 228228 311164 228256
rect 302844 228216 302850 228228
rect 311158 228216 311164 228228
rect 311216 228216 311222 228268
rect 328822 228256 328828 228268
rect 316052 228228 328828 228256
rect 131758 228148 131764 228200
rect 131816 228188 131822 228200
rect 226150 228188 226156 228200
rect 131816 228160 226156 228188
rect 131816 228148 131822 228160
rect 226150 228148 226156 228160
rect 226208 228148 226214 228200
rect 231670 228148 231676 228200
rect 231728 228188 231734 228200
rect 267826 228188 267832 228200
rect 231728 228160 267832 228188
rect 231728 228148 231734 228160
rect 267826 228148 267832 228160
rect 267884 228148 267890 228200
rect 309226 228148 309232 228200
rect 309284 228188 309290 228200
rect 316052 228188 316080 228228
rect 328822 228216 328828 228228
rect 328880 228216 328886 228268
rect 337010 228216 337016 228268
rect 337068 228256 337074 228268
rect 391934 228256 391940 228268
rect 337068 228228 391940 228256
rect 337068 228216 337074 228228
rect 391934 228216 391940 228228
rect 391992 228216 391998 228268
rect 402606 228216 402612 228268
rect 402664 228256 402670 228268
rect 549254 228256 549260 228268
rect 402664 228228 549260 228256
rect 402664 228216 402670 228228
rect 549254 228216 549260 228228
rect 549312 228216 549318 228268
rect 309284 228160 316080 228188
rect 309284 228148 309290 228160
rect 316218 228148 316224 228200
rect 316276 228188 316282 228200
rect 326246 228188 326252 228200
rect 316276 228160 326252 228188
rect 316276 228148 316282 228160
rect 326246 228148 326252 228160
rect 326304 228148 326310 228200
rect 339126 228148 339132 228200
rect 339184 228188 339190 228200
rect 393774 228188 393780 228200
rect 339184 228160 393780 228188
rect 339184 228148 339190 228160
rect 393774 228148 393780 228160
rect 393832 228148 393838 228200
rect 403618 228148 403624 228200
rect 403676 228188 403682 228200
rect 552014 228188 552020 228200
rect 403676 228160 552020 228188
rect 403676 228148 403682 228160
rect 552014 228148 552020 228160
rect 552072 228148 552078 228200
rect 123386 228080 123392 228132
rect 123444 228120 123450 228132
rect 222930 228120 222936 228132
rect 123444 228092 222936 228120
rect 123444 228080 123450 228092
rect 222930 228080 222936 228092
rect 222988 228080 222994 228132
rect 223482 228080 223488 228132
rect 223540 228120 223546 228132
rect 263870 228120 263876 228132
rect 223540 228092 263876 228120
rect 223540 228080 223546 228092
rect 263870 228080 263876 228092
rect 263928 228080 263934 228132
rect 311710 228080 311716 228132
rect 311768 228120 311774 228132
rect 332962 228120 332968 228132
rect 311768 228092 332968 228120
rect 311768 228080 311774 228092
rect 332962 228080 332968 228092
rect 333020 228080 333026 228132
rect 336274 228080 336280 228132
rect 336332 228120 336338 228132
rect 389910 228120 389916 228132
rect 336332 228092 389916 228120
rect 336332 228080 336338 228092
rect 389910 228080 389916 228092
rect 389968 228080 389974 228132
rect 406838 228080 406844 228132
rect 406896 228120 406902 228132
rect 559282 228120 559288 228132
rect 406896 228092 559288 228120
rect 406896 228080 406902 228092
rect 559282 228080 559288 228092
rect 559340 228080 559346 228132
rect 108206 228012 108212 228064
rect 108264 228052 108270 228064
rect 216122 228052 216128 228064
rect 108264 228024 216128 228052
rect 108264 228012 108270 228024
rect 216122 228012 216128 228024
rect 216180 228012 216186 228064
rect 216674 228012 216680 228064
rect 216732 228052 216738 228064
rect 261018 228052 261024 228064
rect 216732 228024 261024 228052
rect 216732 228012 216738 228024
rect 261018 228012 261024 228024
rect 261076 228012 261082 228064
rect 311342 228012 311348 228064
rect 311400 228052 311406 228064
rect 331306 228052 331312 228064
rect 311400 228024 331312 228052
rect 311400 228012 311406 228024
rect 331306 228012 331312 228024
rect 331364 228012 331370 228064
rect 341242 228012 341248 228064
rect 341300 228052 341306 228064
rect 396166 228052 396172 228064
rect 341300 228024 396172 228052
rect 341300 228012 341306 228024
rect 396166 228012 396172 228024
rect 396224 228012 396230 228064
rect 406194 228012 406200 228064
rect 406252 228052 406258 228064
rect 557626 228052 557632 228064
rect 406252 228024 557632 228052
rect 406252 228012 406258 228024
rect 557626 228012 557632 228024
rect 557684 228012 557690 228064
rect 78766 227944 78772 227996
rect 78824 227984 78830 227996
rect 193398 227984 193404 227996
rect 78824 227956 193404 227984
rect 78824 227944 78830 227956
rect 193398 227944 193404 227956
rect 193456 227944 193462 227996
rect 199746 227984 199752 227996
rect 193508 227956 199752 227984
rect 72050 227876 72056 227928
rect 72108 227916 72114 227928
rect 193508 227916 193536 227956
rect 199746 227944 199752 227956
rect 199804 227944 199810 227996
rect 203242 227944 203248 227996
rect 203300 227984 203306 227996
rect 255314 227984 255320 227996
rect 203300 227956 255320 227984
rect 203300 227944 203306 227956
rect 255314 227944 255320 227956
rect 255372 227944 255378 227996
rect 257706 227944 257712 227996
rect 257764 227984 257770 227996
rect 276014 227984 276020 227996
rect 257764 227956 276020 227984
rect 257764 227944 257770 227956
rect 276014 227944 276020 227956
rect 276072 227944 276078 227996
rect 303154 227944 303160 227996
rect 303212 227984 303218 227996
rect 312814 227984 312820 227996
rect 303212 227956 312820 227984
rect 303212 227944 303218 227956
rect 312814 227944 312820 227956
rect 312872 227944 312878 227996
rect 332134 227984 332140 227996
rect 315684 227956 332140 227984
rect 72108 227888 193536 227916
rect 72108 227876 72114 227888
rect 193582 227876 193588 227928
rect 193640 227916 193646 227928
rect 193640 227888 197768 227916
rect 193640 227876 193646 227888
rect 64506 227808 64512 227860
rect 64564 227848 64570 227860
rect 197630 227848 197636 227860
rect 64564 227820 197636 227848
rect 64564 227808 64570 227820
rect 197630 227808 197636 227820
rect 197688 227808 197694 227860
rect 197740 227848 197768 227888
rect 199010 227876 199016 227928
rect 199068 227916 199074 227928
rect 254670 227916 254676 227928
rect 199068 227888 254676 227916
rect 199068 227876 199074 227888
rect 254670 227876 254676 227888
rect 254728 227876 254734 227928
rect 256602 227876 256608 227928
rect 256660 227916 256666 227928
rect 277118 227916 277124 227928
rect 256660 227888 277124 227916
rect 256660 227876 256666 227888
rect 277118 227876 277124 227888
rect 277176 227876 277182 227928
rect 301682 227876 301688 227928
rect 301740 227916 301746 227928
rect 309410 227916 309416 227928
rect 301740 227888 309416 227916
rect 301740 227876 301746 227888
rect 309410 227876 309416 227888
rect 309468 227876 309474 227928
rect 310606 227876 310612 227928
rect 310664 227916 310670 227928
rect 315684 227916 315712 227956
rect 332134 227944 332140 227956
rect 332192 227944 332198 227996
rect 338390 227944 338396 227996
rect 338448 227984 338454 227996
rect 395246 227984 395252 227996
rect 338448 227956 395252 227984
rect 338448 227944 338454 227956
rect 395246 227944 395252 227956
rect 395304 227944 395310 227996
rect 409046 227944 409052 227996
rect 409104 227984 409110 227996
rect 564434 227984 564440 227996
rect 409104 227956 564440 227984
rect 409104 227944 409110 227956
rect 564434 227944 564440 227956
rect 564492 227944 564498 227996
rect 334710 227916 334716 227928
rect 310664 227888 315712 227916
rect 315868 227888 334716 227916
rect 310664 227876 310670 227888
rect 202598 227848 202604 227860
rect 197740 227820 202604 227848
rect 202598 227808 202604 227820
rect 202656 227808 202662 227860
rect 204070 227808 204076 227860
rect 204128 227848 204134 227860
rect 257154 227848 257160 227860
rect 204128 227820 257160 227848
rect 204128 227808 204134 227820
rect 257154 227808 257160 227820
rect 257212 227808 257218 227860
rect 259638 227808 259644 227860
rect 259696 227848 259702 227860
rect 278866 227848 278872 227860
rect 259696 227820 278872 227848
rect 259696 227808 259702 227820
rect 278866 227808 278872 227820
rect 278924 227808 278930 227860
rect 65334 227740 65340 227792
rect 65392 227780 65398 227792
rect 196894 227780 196900 227792
rect 65392 227752 196900 227780
rect 65392 227740 65398 227752
rect 196894 227740 196900 227752
rect 196952 227740 196958 227792
rect 197354 227740 197360 227792
rect 197412 227780 197418 227792
rect 254302 227780 254308 227792
rect 197412 227752 254308 227780
rect 197412 227740 197418 227752
rect 254302 227740 254308 227752
rect 254360 227740 254366 227792
rect 256142 227740 256148 227792
rect 256200 227780 256206 227792
rect 274266 227780 274272 227792
rect 256200 227752 274272 227780
rect 256200 227740 256206 227752
rect 274266 227740 274272 227752
rect 274324 227740 274330 227792
rect 302050 227740 302056 227792
rect 302108 227780 302114 227792
rect 311986 227780 311992 227792
rect 302108 227752 311992 227780
rect 302108 227740 302114 227752
rect 311986 227740 311992 227752
rect 312044 227740 312050 227792
rect 312722 227740 312728 227792
rect 312780 227780 312786 227792
rect 315868 227780 315896 227888
rect 334710 227876 334716 227888
rect 334768 227876 334774 227928
rect 341610 227876 341616 227928
rect 341668 227916 341674 227928
rect 400030 227916 400036 227928
rect 341668 227888 400036 227916
rect 341668 227876 341674 227888
rect 400030 227876 400036 227888
rect 400088 227876 400094 227928
rect 407206 227876 407212 227928
rect 407264 227916 407270 227928
rect 560386 227916 560392 227928
rect 407264 227888 560392 227916
rect 407264 227876 407270 227888
rect 560386 227876 560392 227888
rect 560444 227876 560450 227928
rect 315942 227808 315948 227860
rect 316000 227848 316006 227860
rect 338114 227848 338120 227860
rect 316000 227820 338120 227848
rect 316000 227808 316006 227820
rect 338114 227808 338120 227820
rect 338172 227808 338178 227860
rect 340598 227808 340604 227860
rect 340656 227848 340662 227860
rect 402790 227848 402796 227860
rect 340656 227820 402796 227848
rect 340656 227808 340662 227820
rect 402790 227808 402796 227820
rect 402848 227808 402854 227860
rect 408310 227808 408316 227860
rect 408368 227848 408374 227860
rect 562870 227848 562876 227860
rect 408368 227820 562876 227848
rect 408368 227808 408374 227820
rect 562870 227808 562876 227820
rect 562928 227808 562934 227860
rect 312780 227752 315896 227780
rect 312780 227740 312786 227752
rect 318794 227740 318800 227792
rect 318852 227780 318858 227792
rect 339586 227780 339592 227792
rect 318852 227752 339592 227780
rect 318852 227740 318858 227752
rect 339586 227740 339592 227752
rect 339644 227740 339650 227792
rect 341978 227740 341984 227792
rect 342036 227780 342042 227792
rect 403710 227780 403716 227792
rect 342036 227752 403716 227780
rect 342036 227740 342042 227752
rect 403710 227740 403716 227752
rect 403768 227740 403774 227792
rect 410426 227740 410432 227792
rect 410484 227780 410490 227792
rect 567930 227780 567936 227792
rect 410484 227752 567936 227780
rect 410484 227740 410490 227752
rect 567930 227740 567936 227752
rect 567988 227740 567994 227792
rect 52730 227672 52736 227724
rect 52788 227712 52794 227724
rect 192938 227712 192944 227724
rect 52788 227684 192944 227712
rect 52788 227672 52794 227684
rect 192938 227672 192944 227684
rect 192996 227672 193002 227724
rect 193030 227672 193036 227724
rect 193088 227712 193094 227724
rect 251818 227712 251824 227724
rect 193088 227684 251824 227712
rect 193088 227672 193094 227684
rect 251818 227672 251824 227684
rect 251876 227672 251882 227724
rect 253658 227672 253664 227724
rect 253716 227712 253722 227724
rect 276750 227712 276756 227724
rect 253716 227684 276756 227712
rect 253716 227672 253722 227684
rect 276750 227672 276756 227684
rect 276808 227672 276814 227724
rect 320266 227672 320272 227724
rect 320324 227712 320330 227724
rect 341518 227712 341524 227724
rect 320324 227684 341524 227712
rect 320324 227672 320330 227684
rect 341518 227672 341524 227684
rect 341576 227672 341582 227724
rect 344462 227672 344468 227724
rect 344520 227712 344526 227724
rect 410334 227712 410340 227724
rect 344520 227684 410340 227712
rect 344520 227672 344526 227684
rect 410334 227672 410340 227684
rect 410392 227672 410398 227724
rect 411530 227672 411536 227724
rect 411588 227712 411594 227724
rect 570230 227712 570236 227724
rect 411588 227684 570236 227712
rect 411588 227672 411594 227684
rect 570230 227672 570236 227684
rect 570288 227672 570294 227724
rect 158714 227604 158720 227656
rect 158772 227644 158778 227656
rect 237558 227644 237564 227656
rect 158772 227616 237564 227644
rect 158772 227604 158778 227616
rect 237558 227604 237564 227616
rect 237616 227604 237622 227656
rect 243630 227604 243636 227656
rect 243688 227644 243694 227656
rect 272426 227644 272432 227656
rect 243688 227616 272432 227644
rect 243688 227604 243694 227616
rect 272426 227604 272432 227616
rect 272484 227604 272490 227656
rect 308490 227604 308496 227656
rect 308548 227644 308554 227656
rect 324590 227644 324596 227656
rect 308548 227616 324596 227644
rect 308548 227604 308554 227616
rect 324590 227604 324596 227616
rect 324648 227604 324654 227656
rect 339494 227604 339500 227656
rect 339552 227644 339558 227656
rect 376846 227644 376852 227656
rect 339552 227616 376852 227644
rect 339552 227604 339558 227616
rect 376846 227604 376852 227616
rect 376904 227604 376910 227656
rect 387242 227604 387248 227656
rect 387300 227644 387306 227656
rect 460934 227644 460940 227656
rect 387300 227616 460940 227644
rect 387300 227604 387306 227616
rect 460934 227604 460940 227616
rect 460992 227604 460998 227656
rect 165430 227536 165436 227588
rect 165488 227576 165494 227588
rect 240410 227576 240416 227588
rect 165488 227548 240416 227576
rect 165488 227536 165494 227548
rect 240410 227536 240416 227548
rect 240468 227536 240474 227588
rect 250346 227536 250352 227588
rect 250404 227576 250410 227588
rect 275278 227576 275284 227588
rect 250404 227548 275284 227576
rect 250404 227536 250410 227548
rect 275278 227536 275284 227548
rect 275336 227536 275342 227588
rect 307018 227536 307024 227588
rect 307076 227576 307082 227588
rect 321186 227576 321192 227588
rect 307076 227548 321192 227576
rect 307076 227536 307082 227548
rect 321186 227536 321192 227548
rect 321244 227536 321250 227588
rect 343726 227536 343732 227588
rect 343784 227576 343790 227588
rect 378134 227576 378140 227588
rect 343784 227548 378140 227576
rect 343784 227536 343790 227548
rect 378134 227536 378140 227548
rect 378192 227536 378198 227588
rect 385126 227536 385132 227588
rect 385184 227576 385190 227588
rect 458174 227576 458180 227588
rect 385184 227548 458180 227576
rect 385184 227536 385190 227548
rect 458174 227536 458180 227548
rect 458232 227536 458238 227588
rect 162762 227468 162768 227520
rect 162820 227508 162826 227520
rect 238202 227508 238208 227520
rect 162820 227480 238208 227508
rect 162820 227468 162826 227480
rect 238202 227468 238208 227480
rect 238260 227468 238266 227520
rect 248690 227468 248696 227520
rect 248748 227508 248754 227520
rect 275002 227508 275008 227520
rect 248748 227480 275008 227508
rect 248748 227468 248754 227480
rect 275002 227468 275008 227480
rect 275060 227468 275066 227520
rect 320634 227468 320640 227520
rect 320692 227508 320698 227520
rect 356054 227508 356060 227520
rect 320692 227480 356060 227508
rect 320692 227468 320698 227480
rect 356054 227468 356060 227480
rect 356112 227468 356118 227520
rect 383010 227468 383016 227520
rect 383068 227508 383074 227520
rect 453850 227508 453856 227520
rect 383068 227480 453856 227508
rect 383068 227468 383074 227480
rect 453850 227468 453856 227480
rect 453908 227468 453914 227520
rect 163682 227400 163688 227452
rect 163740 227440 163746 227452
rect 240042 227440 240048 227452
rect 163740 227412 240048 227440
rect 163740 227400 163746 227412
rect 240042 227400 240048 227412
rect 240100 227400 240106 227452
rect 252002 227400 252008 227452
rect 252060 227440 252066 227452
rect 276382 227440 276388 227452
rect 252060 227412 276388 227440
rect 252060 227400 252066 227412
rect 276382 227400 276388 227412
rect 276440 227400 276446 227452
rect 306374 227400 306380 227452
rect 306432 227440 306438 227452
rect 322014 227440 322020 227452
rect 306432 227412 322020 227440
rect 306432 227400 306438 227412
rect 322014 227400 322020 227412
rect 322072 227400 322078 227452
rect 323118 227400 323124 227452
rect 323176 227440 323182 227452
rect 344002 227440 344008 227452
rect 323176 227412 344008 227440
rect 323176 227400 323182 227412
rect 344002 227400 344008 227412
rect 344060 227400 344066 227452
rect 347314 227400 347320 227452
rect 347372 227440 347378 227452
rect 411070 227440 411076 227452
rect 347372 227412 411076 227440
rect 347372 227400 347378 227412
rect 411070 227400 411076 227412
rect 411128 227400 411134 227452
rect 167086 227332 167092 227384
rect 167144 227372 167150 227384
rect 241422 227372 241428 227384
rect 167144 227344 241428 227372
rect 167144 227332 167150 227344
rect 241422 227332 241428 227344
rect 241480 227332 241486 227384
rect 248598 227332 248604 227384
rect 248656 227372 248662 227384
rect 268562 227372 268568 227384
rect 248656 227344 268568 227372
rect 248656 227332 248662 227344
rect 268562 227332 268568 227344
rect 268620 227332 268626 227384
rect 300946 227332 300952 227384
rect 301004 227372 301010 227384
rect 301004 227344 302280 227372
rect 301004 227332 301010 227344
rect 173618 227264 173624 227316
rect 173676 227304 173682 227316
rect 244274 227304 244280 227316
rect 173676 227276 244280 227304
rect 173676 227264 173682 227276
rect 244274 227264 244280 227276
rect 244332 227264 244338 227316
rect 253750 227264 253756 227316
rect 253808 227304 253814 227316
rect 272794 227304 272800 227316
rect 253808 227276 272800 227304
rect 253808 227264 253814 227276
rect 272794 227264 272800 227276
rect 272852 227264 272858 227316
rect 295242 227264 295248 227316
rect 295300 227304 295306 227316
rect 296806 227304 296812 227316
rect 295300 227276 296812 227304
rect 295300 227264 295306 227276
rect 296806 227264 296812 227276
rect 296864 227264 296870 227316
rect 297818 227264 297824 227316
rect 297876 227304 297882 227316
rect 301866 227304 301872 227316
rect 297876 227276 301872 227304
rect 297876 227264 297882 227276
rect 301866 227264 301872 227276
rect 301924 227264 301930 227316
rect 302252 227304 302280 227344
rect 302418 227332 302424 227384
rect 302476 227372 302482 227384
rect 313642 227372 313648 227384
rect 302476 227344 313648 227372
rect 302476 227332 302482 227344
rect 313642 227332 313648 227344
rect 313700 227332 313706 227384
rect 332042 227332 332048 227384
rect 332100 227372 332106 227384
rect 364334 227372 364340 227384
rect 332100 227344 364340 227372
rect 332100 227332 332106 227344
rect 364334 227332 364340 227344
rect 364392 227332 364398 227384
rect 374454 227332 374460 227384
rect 374512 227372 374518 227384
rect 433242 227372 433248 227384
rect 374512 227344 433248 227372
rect 374512 227332 374518 227344
rect 433242 227332 433248 227344
rect 433300 227332 433306 227384
rect 310238 227304 310244 227316
rect 302252 227276 310244 227304
rect 310238 227264 310244 227276
rect 310296 227264 310302 227316
rect 325970 227264 325976 227316
rect 326028 227304 326034 227316
rect 345106 227304 345112 227316
rect 326028 227276 345112 227304
rect 326028 227264 326034 227276
rect 345106 227264 345112 227276
rect 345164 227264 345170 227316
rect 368750 227264 368756 227316
rect 368808 227304 368814 227316
rect 425698 227304 425704 227316
rect 368808 227276 425704 227304
rect 368808 227264 368814 227276
rect 425698 227264 425704 227276
rect 425756 227264 425762 227316
rect 169570 227196 169576 227248
rect 169628 227236 169634 227248
rect 241054 227236 241060 227248
rect 169628 227208 241060 227236
rect 169628 227196 169634 227208
rect 241054 227196 241060 227208
rect 241112 227196 241118 227248
rect 248414 227196 248420 227248
rect 248472 227236 248478 227248
rect 269942 227236 269948 227248
rect 248472 227208 269948 227236
rect 248472 227196 248478 227208
rect 269942 227196 269948 227208
rect 270000 227196 270006 227248
rect 303522 227196 303528 227248
rect 303580 227236 303586 227248
rect 315298 227236 315304 227248
rect 303580 227208 315304 227236
rect 303580 227196 303586 227208
rect 315298 227196 315304 227208
rect 315356 227196 315362 227248
rect 371602 227196 371608 227248
rect 371660 227236 371666 227248
rect 430482 227236 430488 227248
rect 371660 227208 430488 227236
rect 371660 227196 371666 227208
rect 430482 227196 430488 227208
rect 430540 227196 430546 227248
rect 172146 227128 172152 227180
rect 172204 227168 172210 227180
rect 243262 227168 243268 227180
rect 172204 227140 243268 227168
rect 172204 227128 172210 227140
rect 243262 227128 243268 227140
rect 243320 227128 243326 227180
rect 252922 227128 252928 227180
rect 252980 227168 252986 227180
rect 271414 227168 271420 227180
rect 252980 227140 271420 227168
rect 252980 227128 252986 227140
rect 271414 227128 271420 227140
rect 271472 227128 271478 227180
rect 376202 227128 376208 227180
rect 376260 227168 376266 227180
rect 434622 227168 434628 227180
rect 376260 227140 434628 227168
rect 376260 227128 376266 227140
rect 434622 227128 434628 227140
rect 434680 227128 434686 227180
rect 176378 227060 176384 227112
rect 176436 227100 176442 227112
rect 243906 227100 243912 227112
rect 176436 227072 243912 227100
rect 176436 227060 176442 227072
rect 243906 227060 243912 227072
rect 243964 227060 243970 227112
rect 255222 227060 255228 227112
rect 255280 227100 255286 227112
rect 275646 227100 275652 227112
rect 255280 227072 275652 227100
rect 255280 227060 255286 227072
rect 275646 227060 275652 227072
rect 275704 227060 275710 227112
rect 317414 227060 317420 227112
rect 317472 227100 317478 227112
rect 337654 227100 337660 227112
rect 317472 227072 337660 227100
rect 317472 227060 317478 227072
rect 337654 227060 337660 227072
rect 337712 227060 337718 227112
rect 366174 227060 366180 227112
rect 366232 227100 366238 227112
rect 419534 227100 419540 227112
rect 366232 227072 419540 227100
rect 366232 227060 366238 227072
rect 419534 227060 419540 227072
rect 419592 227060 419598 227112
rect 181898 226992 181904 227044
rect 181956 227032 181962 227044
rect 246114 227032 246120 227044
rect 181956 227004 246120 227032
rect 181956 226992 181962 227004
rect 246114 226992 246120 227004
rect 246172 226992 246178 227044
rect 248506 226992 248512 227044
rect 248564 227032 248570 227044
rect 265710 227032 265716 227044
rect 248564 227004 265716 227032
rect 248564 226992 248570 227004
rect 265710 226992 265716 227004
rect 265768 226992 265774 227044
rect 312078 226992 312084 227044
rect 312136 227032 312142 227044
rect 335538 227032 335544 227044
rect 312136 227004 335544 227032
rect 312136 226992 312142 227004
rect 335538 226992 335544 227004
rect 335596 226992 335602 227044
rect 361574 226992 361580 227044
rect 361632 227032 361638 227044
rect 418890 227032 418896 227044
rect 361632 227004 418896 227032
rect 361632 226992 361638 227004
rect 418890 226992 418896 227004
rect 418948 226992 418954 227044
rect 180518 226924 180524 226976
rect 180576 226964 180582 226976
rect 247126 226964 247132 226976
rect 180576 226936 247132 226964
rect 180576 226924 180582 226936
rect 247126 226924 247132 226936
rect 247184 226924 247190 226976
rect 255590 226924 255596 226976
rect 255648 226964 255654 226976
rect 271782 226964 271788 226976
rect 255648 226936 271788 226964
rect 255648 226924 255654 226936
rect 271782 226924 271788 226936
rect 271840 226924 271846 226976
rect 358722 226924 358728 226976
rect 358780 226964 358786 226976
rect 411990 226964 411996 226976
rect 358780 226936 411996 226964
rect 358780 226924 358786 226936
rect 411990 226924 411996 226936
rect 412048 226924 412054 226976
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 248966 226896 248972 226908
rect 185636 226868 248972 226896
rect 185636 226856 185642 226868
rect 248966 226856 248972 226868
rect 249024 226856 249030 226908
rect 258442 226856 258448 226908
rect 258500 226896 258506 226908
rect 274634 226896 274640 226908
rect 258500 226868 274640 226896
rect 258500 226856 258506 226868
rect 274634 226856 274640 226868
rect 274692 226856 274698 226908
rect 300670 226856 300676 226908
rect 300728 226896 300734 226908
rect 308582 226896 308588 226908
rect 300728 226868 308588 226896
rect 300728 226856 300734 226868
rect 308582 226856 308588 226868
rect 308640 226856 308646 226908
rect 355870 226856 355876 226908
rect 355928 226896 355934 226908
rect 408310 226896 408316 226908
rect 355928 226868 408316 226896
rect 355928 226856 355934 226868
rect 408310 226856 408316 226868
rect 408368 226856 408374 226908
rect 408678 226856 408684 226908
rect 408736 226896 408742 226908
rect 449710 226896 449716 226908
rect 408736 226868 449716 226896
rect 408736 226856 408742 226868
rect 449710 226856 449716 226868
rect 449768 226856 449774 226908
rect 190362 226788 190368 226840
rect 190420 226828 190426 226840
rect 251450 226828 251456 226840
rect 190420 226800 251456 226828
rect 190420 226788 190426 226800
rect 251450 226788 251456 226800
rect 251508 226788 251514 226840
rect 255406 226788 255412 226840
rect 255464 226828 255470 226840
rect 270310 226828 270316 226840
rect 255464 226800 270316 226828
rect 255464 226788 255470 226800
rect 270310 226788 270316 226800
rect 270368 226788 270374 226840
rect 299566 226788 299572 226840
rect 299624 226828 299630 226840
rect 306926 226828 306932 226840
rect 299624 226800 306932 226828
rect 299624 226788 299630 226800
rect 306926 226788 306932 226800
rect 306984 226788 306990 226840
rect 323486 226788 323492 226840
rect 323544 226828 323550 226840
rect 362402 226828 362408 226840
rect 323544 226800 362408 226828
rect 323544 226788 323550 226800
rect 362402 226788 362408 226800
rect 362460 226788 362466 226840
rect 366910 226788 366916 226840
rect 366968 226828 366974 226840
rect 408402 226828 408408 226840
rect 366968 226800 408408 226828
rect 366968 226788 366974 226800
rect 408402 226788 408408 226800
rect 408460 226788 408466 226840
rect 409690 226788 409696 226840
rect 409748 226828 409754 226840
rect 448790 226828 448796 226840
rect 409748 226800 448796 226828
rect 409748 226788 409754 226800
rect 448790 226788 448796 226800
rect 448848 226788 448854 226840
rect 186406 226720 186412 226772
rect 186464 226760 186470 226772
rect 248230 226760 248236 226772
rect 186464 226732 248236 226760
rect 186464 226720 186470 226732
rect 248230 226720 248236 226732
rect 248288 226720 248294 226772
rect 299198 226720 299204 226772
rect 299256 226760 299262 226772
rect 305270 226760 305276 226772
rect 299256 226732 305276 226760
rect 299256 226720 299262 226732
rect 305270 226720 305276 226732
rect 305328 226720 305334 226772
rect 345198 226720 345204 226772
rect 345256 226760 345262 226772
rect 376570 226760 376576 226772
rect 345256 226732 376576 226760
rect 345256 226720 345262 226732
rect 376570 226720 376576 226732
rect 376628 226720 376634 226772
rect 379790 226720 379796 226772
rect 379848 226760 379854 226772
rect 391750 226760 391756 226772
rect 379848 226732 391756 226760
rect 379848 226720 379854 226732
rect 391750 226720 391756 226732
rect 391808 226720 391814 226772
rect 402238 226720 402244 226772
rect 402296 226760 402302 226772
rect 441614 226760 441620 226772
rect 402296 226732 441620 226760
rect 402296 226720 402302 226732
rect 441614 226720 441620 226732
rect 441672 226720 441678 226772
rect 42150 226652 42156 226704
rect 42208 226692 42214 226704
rect 43990 226692 43996 226704
rect 42208 226664 43996 226692
rect 42208 226652 42214 226664
rect 43990 226652 43996 226664
rect 44048 226652 44054 226704
rect 192938 226652 192944 226704
rect 192996 226692 193002 226704
rect 251082 226692 251088 226704
rect 192996 226664 251088 226692
rect 192996 226652 193002 226664
rect 251082 226652 251088 226664
rect 251140 226652 251146 226704
rect 259362 226652 259368 226704
rect 259420 226692 259426 226704
rect 273162 226692 273168 226704
rect 259420 226664 273168 226692
rect 259420 226652 259426 226664
rect 273162 226652 273168 226664
rect 273220 226652 273226 226704
rect 298094 226652 298100 226704
rect 298152 226692 298158 226704
rect 303614 226692 303620 226704
rect 298152 226664 303620 226692
rect 298152 226652 298158 226664
rect 303614 226652 303620 226664
rect 303672 226652 303678 226704
rect 361206 226652 361212 226704
rect 361264 226692 361270 226704
rect 383654 226692 383660 226704
rect 361264 226664 383660 226692
rect 361264 226652 361270 226664
rect 383654 226652 383660 226664
rect 383712 226652 383718 226704
rect 399018 226652 399024 226704
rect 399076 226692 399082 226704
rect 436094 226692 436100 226704
rect 399076 226664 436100 226692
rect 399076 226652 399082 226664
rect 436094 226652 436100 226664
rect 436152 226652 436158 226704
rect 234706 226584 234712 226636
rect 234764 226624 234770 226636
rect 256786 226624 256792 226636
rect 234764 226596 256792 226624
rect 234764 226584 234770 226596
rect 256786 226584 256792 226596
rect 256844 226584 256850 226636
rect 300302 226584 300308 226636
rect 300360 226624 300366 226636
rect 306374 226624 306380 226636
rect 300360 226596 306380 226624
rect 300360 226584 300366 226596
rect 306374 226584 306380 226596
rect 306432 226584 306438 226636
rect 371970 226584 371976 226636
rect 372028 226624 372034 226636
rect 397546 226624 397552 226636
rect 372028 226596 397552 226624
rect 372028 226584 372034 226596
rect 397546 226584 397552 226596
rect 397604 226584 397610 226636
rect 404354 226584 404360 226636
rect 404412 226624 404418 226636
rect 438854 226624 438860 226636
rect 404412 226596 438860 226624
rect 404412 226584 404418 226596
rect 438854 226584 438860 226596
rect 438912 226584 438918 226636
rect 247034 226516 247040 226568
rect 247092 226556 247098 226568
rect 264698 226556 264704 226568
rect 247092 226528 264704 226556
rect 247092 226516 247098 226528
rect 264698 226516 264704 226528
rect 264756 226516 264762 226568
rect 301314 226516 301320 226568
rect 301372 226556 301378 226568
rect 307754 226556 307760 226568
rect 301372 226528 307760 226556
rect 301372 226516 301378 226528
rect 307754 226516 307760 226528
rect 307812 226516 307818 226568
rect 374086 226516 374092 226568
rect 374144 226556 374150 226568
rect 402974 226556 402980 226568
rect 374144 226528 402980 226556
rect 374144 226516 374150 226528
rect 402974 226516 402980 226528
rect 403032 226516 403038 226568
rect 197814 226448 197820 226500
rect 197872 226488 197878 226500
rect 207934 226488 207940 226500
rect 197872 226460 207940 226488
rect 197872 226448 197878 226460
rect 207934 226448 207940 226460
rect 207992 226448 207998 226500
rect 245654 226448 245660 226500
rect 245712 226488 245718 226500
rect 258534 226488 258540 226500
rect 245712 226460 258540 226488
rect 245712 226448 245718 226460
rect 258534 226448 258540 226460
rect 258592 226448 258598 226500
rect 303798 226448 303804 226500
rect 303856 226488 303862 226500
rect 317414 226488 317420 226500
rect 303856 226460 317420 226488
rect 303856 226448 303862 226460
rect 317414 226448 317420 226460
rect 317472 226448 317478 226500
rect 330570 226448 330576 226500
rect 330628 226488 330634 226500
rect 379238 226488 379244 226500
rect 330628 226460 379244 226488
rect 330628 226448 330634 226460
rect 379238 226448 379244 226460
rect 379296 226448 379302 226500
rect 395798 226448 395804 226500
rect 395856 226488 395862 226500
rect 422294 226488 422300 226500
rect 395856 226460 422300 226488
rect 395856 226448 395862 226460
rect 422294 226448 422300 226460
rect 422352 226448 422358 226500
rect 304902 226380 304908 226432
rect 304960 226420 304966 226432
rect 318702 226420 318708 226432
rect 304960 226392 318708 226420
rect 304960 226380 304966 226392
rect 318702 226380 318708 226392
rect 318760 226380 318766 226432
rect 373350 226380 373356 226432
rect 373408 226420 373414 226432
rect 397454 226420 397460 226432
rect 373408 226392 397460 226420
rect 373408 226380 373414 226392
rect 397454 226380 397460 226392
rect 397512 226380 397518 226432
rect 254670 226312 254676 226364
rect 254728 226352 254734 226364
rect 268930 226352 268936 226364
rect 254728 226324 268936 226352
rect 254728 226312 254734 226324
rect 268930 226312 268936 226324
rect 268988 226312 268994 226364
rect 299934 226312 299940 226364
rect 299992 226352 299998 226364
rect 304350 226352 304356 226364
rect 299992 226324 304356 226352
rect 299992 226312 299998 226324
rect 304350 226312 304356 226324
rect 304408 226312 304414 226364
rect 309870 226312 309876 226364
rect 309928 226352 309934 226364
rect 327902 226352 327908 226364
rect 309928 226324 327908 226352
rect 309928 226312 309934 226324
rect 327902 226312 327908 226324
rect 327960 226312 327966 226364
rect 331674 226312 331680 226364
rect 331732 226352 331738 226364
rect 347406 226352 347412 226364
rect 331732 226324 347412 226352
rect 331732 226312 331738 226324
rect 347406 226312 347412 226324
rect 347464 226312 347470 226364
rect 368014 226312 368020 226364
rect 368072 226352 368078 226364
rect 369946 226352 369952 226364
rect 368072 226324 369952 226352
rect 368072 226312 368078 226324
rect 369946 226312 369952 226324
rect 370004 226312 370010 226364
rect 389358 226312 389364 226364
rect 389416 226352 389422 226364
rect 411162 226352 411168 226364
rect 389416 226324 411168 226352
rect 389416 226312 389422 226324
rect 411162 226312 411168 226324
rect 411220 226312 411226 226364
rect 411896 226356 411902 226408
rect 411954 226396 411960 226408
rect 485546 226396 485552 226406
rect 411954 226368 485552 226396
rect 411954 226356 411960 226368
rect 485546 226354 485552 226368
rect 485604 226396 485610 226406
rect 485604 226368 485612 226396
rect 485604 226354 485610 226368
rect 154482 226244 154488 226296
rect 154540 226284 154546 226296
rect 235074 226284 235080 226296
rect 154540 226256 235080 226284
rect 154540 226244 154546 226256
rect 235074 226244 235080 226256
rect 235132 226244 235138 226296
rect 354122 226244 354128 226296
rect 354180 226284 354186 226296
rect 432230 226284 432236 226296
rect 354180 226256 432236 226284
rect 354180 226244 354186 226256
rect 432230 226244 432236 226256
rect 432288 226244 432294 226296
rect 434806 226284 434812 226296
rect 433076 226256 434812 226284
rect 144362 226176 144368 226228
rect 144420 226216 144426 226228
rect 230750 226216 230756 226228
rect 144420 226188 230756 226216
rect 144420 226176 144426 226188
rect 230750 226176 230756 226188
rect 230808 226176 230814 226228
rect 353754 226176 353760 226228
rect 353812 226216 353818 226228
rect 433076 226216 433104 226256
rect 434806 226244 434812 226256
rect 434864 226244 434870 226296
rect 435634 226216 435640 226228
rect 353812 226188 433104 226216
rect 433168 226188 435640 226216
rect 353812 226176 353818 226188
rect 147766 226108 147772 226160
rect 147824 226148 147830 226160
rect 232222 226148 232228 226160
rect 147824 226120 232228 226148
rect 147824 226108 147830 226120
rect 232222 226108 232228 226120
rect 232280 226108 232286 226160
rect 352282 226108 352288 226160
rect 352340 226148 352346 226160
rect 431402 226148 431408 226160
rect 352340 226120 431408 226148
rect 352340 226108 352346 226120
rect 431402 226108 431408 226120
rect 431460 226108 431466 226160
rect 141050 226040 141056 226092
rect 141108 226080 141114 226092
rect 229370 226080 229376 226092
rect 141108 226052 229376 226080
rect 141108 226040 141114 226052
rect 229370 226040 229376 226052
rect 229428 226040 229434 226092
rect 355502 226040 355508 226092
rect 355560 226080 355566 226092
rect 433168 226080 433196 226188
rect 435634 226176 435640 226188
rect 435692 226176 435698 226228
rect 466362 226176 466368 226228
rect 466420 226216 466426 226228
rect 487798 226216 487804 226228
rect 466420 226188 487804 226216
rect 466420 226176 466426 226188
rect 487798 226176 487804 226188
rect 487856 226176 487862 226228
rect 433242 226108 433248 226160
rect 433300 226148 433306 226160
rect 480990 226148 480996 226160
rect 433300 226120 480996 226148
rect 433300 226108 433306 226120
rect 480990 226108 480996 226120
rect 481048 226108 481054 226160
rect 355560 226052 433196 226080
rect 355560 226040 355566 226052
rect 434622 226040 434628 226092
rect 434680 226080 434686 226092
rect 487154 226080 487160 226092
rect 434680 226052 487160 226080
rect 434680 226040 434686 226052
rect 487154 226040 487160 226052
rect 487212 226040 487218 226092
rect 137646 225972 137652 226024
rect 137704 226012 137710 226024
rect 227898 226012 227904 226024
rect 137704 225984 227904 226012
rect 137704 225972 137710 225984
rect 227898 225972 227904 225984
rect 227956 225972 227962 226024
rect 340230 225972 340236 226024
rect 340288 226012 340294 226024
rect 370222 226012 370228 226024
rect 340288 225984 370228 226012
rect 340288 225972 340294 225984
rect 370222 225972 370228 225984
rect 370280 225972 370286 226024
rect 397454 225972 397460 226024
rect 397512 226012 397518 226024
rect 480346 226012 480352 226024
rect 397512 225984 480352 226012
rect 397512 225972 397518 225984
rect 480346 225972 480352 225984
rect 480404 225972 480410 226024
rect 130930 225904 130936 225956
rect 130988 225944 130994 225956
rect 225046 225944 225052 225956
rect 130988 225916 225052 225944
rect 130988 225904 130994 225916
rect 225046 225904 225052 225916
rect 225104 225904 225110 225956
rect 356606 225904 356612 225956
rect 356664 225944 356670 225956
rect 441706 225944 441712 225956
rect 356664 225916 441712 225944
rect 356664 225904 356670 225916
rect 441706 225904 441712 225916
rect 441764 225904 441770 225956
rect 480254 225904 480260 225956
rect 480312 225944 480318 225956
rect 502334 225944 502340 225956
rect 480312 225916 502340 225944
rect 480312 225904 480318 225916
rect 502334 225904 502340 225916
rect 502392 225904 502398 225956
rect 134242 225836 134248 225888
rect 134300 225876 134306 225888
rect 226518 225876 226524 225888
rect 134300 225848 226524 225876
rect 134300 225836 134306 225848
rect 226518 225836 226524 225848
rect 226576 225836 226582 225888
rect 360838 225836 360844 225888
rect 360896 225876 360902 225888
rect 451550 225876 451556 225888
rect 360896 225848 451556 225876
rect 360896 225836 360902 225848
rect 451550 225836 451556 225848
rect 451608 225836 451614 225888
rect 472066 225836 472072 225888
rect 472124 225876 472130 225888
rect 523954 225876 523960 225888
rect 472124 225848 523960 225876
rect 472124 225836 472130 225848
rect 523954 225836 523960 225848
rect 524012 225836 524018 225888
rect 127526 225768 127532 225820
rect 127584 225808 127590 225820
rect 223666 225808 223672 225820
rect 127584 225780 223672 225808
rect 127584 225768 127590 225780
rect 223666 225768 223672 225780
rect 223724 225768 223730 225820
rect 362310 225768 362316 225820
rect 362368 225808 362374 225820
rect 454954 225808 454960 225820
rect 362368 225780 454960 225808
rect 362368 225768 362374 225780
rect 454954 225768 454960 225780
rect 455012 225768 455018 225820
rect 458174 225768 458180 225820
rect 458232 225808 458238 225820
rect 507946 225808 507952 225820
rect 458232 225780 507952 225808
rect 458232 225768 458238 225780
rect 507946 225768 507952 225780
rect 508004 225768 508010 225820
rect 119154 225700 119160 225752
rect 119212 225740 119218 225752
rect 219710 225740 219716 225752
rect 119212 225712 219716 225740
rect 119212 225700 119218 225712
rect 219710 225700 219716 225712
rect 219768 225700 219774 225752
rect 220630 225700 220636 225752
rect 220688 225740 220694 225752
rect 249610 225740 249616 225752
rect 220688 225712 249616 225740
rect 220688 225700 220694 225712
rect 249610 225700 249616 225712
rect 249668 225700 249674 225752
rect 362678 225700 362684 225752
rect 362736 225740 362742 225752
rect 452654 225740 452660 225752
rect 362736 225712 452660 225740
rect 362736 225700 362742 225712
rect 452654 225700 452660 225712
rect 452712 225700 452718 225752
rect 453850 225700 453856 225752
rect 453908 225740 453914 225752
rect 503162 225740 503168 225752
rect 453908 225712 503168 225740
rect 453908 225700 453914 225712
rect 503162 225700 503168 225712
rect 503220 225700 503226 225752
rect 124122 225632 124128 225684
rect 124180 225672 124186 225684
rect 222194 225672 222200 225684
rect 124180 225644 222200 225672
rect 124180 225632 124186 225644
rect 222194 225632 222200 225644
rect 222252 225632 222258 225684
rect 231854 225632 231860 225684
rect 231912 225672 231918 225684
rect 253934 225672 253940 225684
rect 231912 225644 253940 225672
rect 231912 225632 231918 225644
rect 253934 225632 253940 225644
rect 253992 225632 253998 225684
rect 363690 225632 363696 225684
rect 363748 225672 363754 225684
rect 458450 225672 458456 225684
rect 363748 225644 458456 225672
rect 363748 225632 363754 225644
rect 458450 225632 458456 225644
rect 458508 225632 458514 225684
rect 460934 225632 460940 225684
rect 460992 225672 460998 225684
rect 513466 225672 513472 225684
rect 460992 225644 513472 225672
rect 460992 225632 460998 225644
rect 513466 225632 513472 225644
rect 513524 225632 513530 225684
rect 42426 225564 42432 225616
rect 42484 225604 42490 225616
rect 48682 225604 48688 225616
rect 42484 225576 48688 225604
rect 42484 225564 42490 225576
rect 48682 225564 48688 225576
rect 48740 225564 48746 225616
rect 114094 225564 114100 225616
rect 114152 225604 114158 225616
rect 217962 225604 217968 225616
rect 114152 225576 217968 225604
rect 114152 225564 114158 225576
rect 217962 225564 217968 225576
rect 218020 225564 218026 225616
rect 228450 225564 228456 225616
rect 228508 225604 228514 225616
rect 266446 225604 266452 225616
rect 228508 225576 266452 225604
rect 228508 225564 228514 225576
rect 266446 225564 266452 225576
rect 266504 225564 266510 225616
rect 365162 225564 365168 225616
rect 365220 225604 365226 225616
rect 461670 225604 461676 225616
rect 365220 225576 461676 225604
rect 365220 225564 365226 225576
rect 461670 225564 461676 225576
rect 461728 225564 461734 225616
rect 474734 225564 474740 225616
rect 474792 225604 474798 225616
rect 529014 225604 529020 225616
rect 474792 225576 529020 225604
rect 474792 225564 474798 225576
rect 529014 225564 529020 225576
rect 529072 225564 529078 225616
rect 117498 225496 117504 225548
rect 117556 225536 117562 225548
rect 219342 225536 219348 225548
rect 117556 225508 219348 225536
rect 117556 225496 117562 225508
rect 219342 225496 219348 225508
rect 219400 225496 219406 225548
rect 262122 225536 262128 225548
rect 219452 225508 262128 225536
rect 105722 225428 105728 225480
rect 105780 225468 105786 225480
rect 214006 225468 214012 225480
rect 105780 225440 214012 225468
rect 105780 225428 105786 225440
rect 214006 225428 214012 225440
rect 214064 225428 214070 225480
rect 218422 225428 218428 225480
rect 218480 225468 218486 225480
rect 219452 225468 219480 225508
rect 262122 225496 262128 225508
rect 262180 225496 262186 225548
rect 343082 225496 343088 225548
rect 343140 225536 343146 225548
rect 368198 225536 368204 225548
rect 343140 225508 368204 225536
rect 343140 225496 343146 225508
rect 368198 225496 368204 225508
rect 368256 225496 368262 225548
rect 369762 225496 369768 225548
rect 369820 225536 369826 225548
rect 468386 225536 468392 225548
rect 369820 225508 468392 225536
rect 369820 225496 369826 225508
rect 468386 225496 468392 225508
rect 468444 225496 468450 225548
rect 469122 225496 469128 225548
rect 469180 225536 469186 225548
rect 518894 225536 518900 225548
rect 469180 225508 518900 225536
rect 469180 225496 469186 225508
rect 518894 225496 518900 225508
rect 518952 225496 518958 225548
rect 218480 225440 219480 225468
rect 218480 225428 218486 225440
rect 221734 225428 221740 225480
rect 221792 225468 221798 225480
rect 263594 225468 263600 225480
rect 221792 225440 263600 225468
rect 221792 225428 221798 225440
rect 263594 225428 263600 225440
rect 263652 225428 263658 225480
rect 366542 225428 366548 225480
rect 366600 225468 366606 225480
rect 465074 225468 465080 225480
rect 366600 225440 465080 225468
rect 366600 225428 366606 225440
rect 465074 225428 465080 225440
rect 465132 225428 465138 225480
rect 474826 225428 474832 225480
rect 474884 225468 474890 225480
rect 533982 225468 533988 225480
rect 474884 225440 533988 225468
rect 474884 225428 474890 225440
rect 533982 225428 533988 225440
rect 534040 225428 534046 225480
rect 107378 225360 107384 225412
rect 107436 225400 107442 225412
rect 215110 225400 215116 225412
rect 107436 225372 215116 225400
rect 107436 225360 107442 225372
rect 215110 225360 215116 225372
rect 215168 225360 215174 225412
rect 225138 225360 225144 225412
rect 225196 225400 225202 225412
rect 264974 225400 264980 225412
rect 225196 225372 264980 225400
rect 225196 225360 225202 225372
rect 264974 225360 264980 225372
rect 265032 225360 265038 225412
rect 339862 225360 339868 225412
rect 339920 225400 339926 225412
rect 369578 225400 369584 225412
rect 339920 225372 369584 225400
rect 339920 225360 339926 225372
rect 369578 225360 369584 225372
rect 369636 225360 369642 225412
rect 369670 225360 369676 225412
rect 369728 225400 369734 225412
rect 469214 225400 469220 225412
rect 369728 225372 469220 225400
rect 369728 225360 369734 225372
rect 469214 225360 469220 225372
rect 469272 225360 469278 225412
rect 477494 225360 477500 225412
rect 477552 225400 477558 225412
rect 539042 225400 539048 225412
rect 477552 225372 539048 225400
rect 477552 225360 477558 225372
rect 539042 225360 539048 225372
rect 539100 225360 539106 225412
rect 90542 225292 90548 225344
rect 90600 225332 90606 225344
rect 197814 225332 197820 225344
rect 90600 225304 197820 225332
rect 90600 225292 90606 225304
rect 197814 225292 197820 225304
rect 197872 225292 197878 225344
rect 198182 225292 198188 225344
rect 198240 225332 198246 225344
rect 253566 225332 253572 225344
rect 198240 225304 253572 225332
rect 198240 225292 198246 225304
rect 253566 225292 253572 225304
rect 253624 225292 253630 225344
rect 355134 225292 355140 225344
rect 355192 225332 355198 225344
rect 355192 225304 436048 225332
rect 355192 225292 355198 225304
rect 103974 225224 103980 225276
rect 104032 225264 104038 225276
rect 213638 225264 213644 225276
rect 104032 225236 213644 225264
rect 104032 225224 104038 225236
rect 213638 225224 213644 225236
rect 213696 225224 213702 225276
rect 215018 225224 215024 225276
rect 215076 225264 215082 225276
rect 260742 225264 260748 225276
rect 215076 225236 260748 225264
rect 215076 225224 215082 225236
rect 260742 225224 260748 225236
rect 260800 225224 260806 225276
rect 313458 225224 313464 225276
rect 313516 225264 313522 225276
rect 338850 225264 338856 225276
rect 313516 225236 338856 225264
rect 313516 225224 313522 225236
rect 338850 225224 338856 225236
rect 338908 225224 338914 225276
rect 358354 225224 358360 225276
rect 358412 225264 358418 225276
rect 429102 225264 429108 225276
rect 358412 225236 429108 225264
rect 358412 225224 358418 225236
rect 429102 225224 429108 225236
rect 429160 225224 429166 225276
rect 436020 225264 436048 225304
rect 436094 225292 436100 225344
rect 436152 225332 436158 225344
rect 541434 225332 541440 225344
rect 436152 225304 541440 225332
rect 436152 225292 436158 225304
rect 541434 225292 541440 225304
rect 541492 225292 541498 225344
rect 438118 225264 438124 225276
rect 436020 225236 438124 225264
rect 438118 225224 438124 225236
rect 438176 225224 438182 225276
rect 441614 225224 441620 225276
rect 441672 225264 441678 225276
rect 546494 225264 546500 225276
rect 441672 225236 546500 225264
rect 441672 225224 441678 225236
rect 546494 225224 546500 225236
rect 546552 225224 546558 225276
rect 100662 225156 100668 225208
rect 100720 225196 100726 225208
rect 197446 225196 197452 225208
rect 100720 225168 197452 225196
rect 100720 225156 100726 225168
rect 197446 225156 197452 225168
rect 197504 225156 197510 225208
rect 208302 225156 208308 225208
rect 208360 225196 208366 225208
rect 208360 225168 209820 225196
rect 208360 225156 208366 225168
rect 95602 225088 95608 225140
rect 95660 225128 95666 225140
rect 209682 225128 209688 225140
rect 95660 225100 209688 225128
rect 95660 225088 95666 225100
rect 209682 225088 209688 225100
rect 209740 225088 209746 225140
rect 209792 225128 209820 225168
rect 211706 225156 211712 225208
rect 211764 225196 211770 225208
rect 259270 225196 259276 225208
rect 211764 225168 259276 225196
rect 211764 225156 211770 225168
rect 259270 225156 259276 225168
rect 259328 225156 259334 225208
rect 314930 225156 314936 225208
rect 314988 225196 314994 225208
rect 342438 225196 342444 225208
rect 314988 225168 342444 225196
rect 314988 225156 314994 225168
rect 342438 225156 342444 225168
rect 342496 225156 342502 225208
rect 349798 225156 349804 225208
rect 349856 225196 349862 225208
rect 422202 225196 422208 225208
rect 349856 225168 422208 225196
rect 349856 225156 349862 225168
rect 422202 225156 422208 225168
rect 422260 225156 422266 225208
rect 422294 225156 422300 225208
rect 422352 225196 422358 225208
rect 532786 225196 532792 225208
rect 422352 225168 532792 225196
rect 422352 225156 422358 225168
rect 532786 225156 532792 225168
rect 532844 225156 532850 225208
rect 257890 225128 257896 225140
rect 209792 225100 257896 225128
rect 257890 225088 257896 225100
rect 257948 225088 257954 225140
rect 317782 225088 317788 225140
rect 317840 225128 317846 225140
rect 348970 225128 348976 225140
rect 317840 225100 348976 225128
rect 317840 225088 317846 225100
rect 348970 225088 348976 225100
rect 349028 225088 349034 225140
rect 356974 225088 356980 225140
rect 357032 225128 357038 225140
rect 438762 225128 438768 225140
rect 357032 225100 438768 225128
rect 357032 225088 357038 225100
rect 438762 225088 438768 225100
rect 438820 225088 438826 225140
rect 438854 225088 438860 225140
rect 438912 225128 438918 225140
rect 554314 225128 554320 225140
rect 438912 225100 554320 225128
rect 438912 225088 438918 225100
rect 554314 225088 554320 225100
rect 554372 225088 554378 225140
rect 88886 225020 88892 225072
rect 88944 225060 88950 225072
rect 206738 225060 206744 225072
rect 88944 225032 206744 225060
rect 88944 225020 88950 225032
rect 206738 225020 206744 225032
rect 206796 225020 206802 225072
rect 206922 225020 206928 225072
rect 206980 225060 206986 225072
rect 256418 225060 256424 225072
rect 206980 225032 256424 225060
rect 206980 225020 206986 225032
rect 256418 225020 256424 225032
rect 256476 225020 256482 225072
rect 316310 225020 316316 225072
rect 316368 225060 316374 225072
rect 345566 225060 345572 225072
rect 316368 225032 345572 225060
rect 316368 225020 316374 225032
rect 345566 225020 345572 225032
rect 345624 225020 345630 225072
rect 357986 225020 357992 225072
rect 358044 225060 358050 225072
rect 444834 225060 444840 225072
rect 358044 225032 444840 225060
rect 358044 225020 358050 225032
rect 444834 225020 444840 225032
rect 444892 225020 444898 225072
rect 449710 225020 449716 225072
rect 449768 225060 449774 225072
rect 563698 225060 563704 225072
rect 449768 225032 563704 225060
rect 449768 225020 449774 225032
rect 563698 225020 563704 225032
rect 563756 225020 563762 225072
rect 73706 224952 73712 225004
rect 73764 224992 73770 225004
rect 200850 224992 200856 225004
rect 73764 224964 200856 224992
rect 73764 224952 73770 224964
rect 200850 224952 200856 224964
rect 200908 224952 200914 225004
rect 255038 224992 255044 225004
rect 206848 224964 255044 224992
rect 60274 224884 60280 224936
rect 60332 224924 60338 224936
rect 195146 224924 195152 224936
rect 60332 224896 195152 224924
rect 60332 224884 60338 224896
rect 195146 224884 195152 224896
rect 195204 224884 195210 224936
rect 201402 224884 201408 224936
rect 201460 224924 201466 224936
rect 206848 224924 206876 224964
rect 255038 224952 255044 224964
rect 255096 224952 255102 225004
rect 319162 224952 319168 225004
rect 319220 224992 319226 225004
rect 352374 224992 352380 225004
rect 319220 224964 352380 224992
rect 319220 224952 319226 224964
rect 352374 224952 352380 224964
rect 352432 224952 352438 225004
rect 359458 224952 359464 225004
rect 359516 224992 359522 225004
rect 448238 224992 448244 225004
rect 359516 224964 448244 224992
rect 359516 224952 359522 224964
rect 448238 224952 448244 224964
rect 448296 224952 448302 225004
rect 448790 224952 448796 225004
rect 448848 224992 448854 225004
rect 565998 224992 566004 225004
rect 448848 224964 566004 224992
rect 448848 224952 448854 224964
rect 565998 224952 566004 224964
rect 566056 224952 566062 225004
rect 201460 224896 206876 224924
rect 201460 224884 201466 224896
rect 207014 224884 207020 224936
rect 207072 224924 207078 224936
rect 252186 224924 252192 224936
rect 207072 224896 252192 224924
rect 207072 224884 207078 224896
rect 252186 224884 252192 224896
rect 252244 224884 252250 224936
rect 335170 224884 335176 224936
rect 335228 224924 335234 224936
rect 391014 224924 391020 224936
rect 335228 224896 391020 224924
rect 335228 224884 335234 224896
rect 391014 224884 391020 224896
rect 391072 224884 391078 224936
rect 406470 224884 406476 224936
rect 406528 224924 406534 224936
rect 559098 224924 559104 224936
rect 406528 224896 559104 224924
rect 406528 224884 406534 224896
rect 559098 224884 559104 224896
rect 559156 224884 559162 224936
rect 151078 224816 151084 224868
rect 151136 224856 151142 224868
rect 233602 224856 233608 224868
rect 151136 224828 233608 224856
rect 151136 224816 151142 224828
rect 233602 224816 233608 224828
rect 233660 224816 233666 224868
rect 350902 224816 350908 224868
rect 350960 224856 350966 224868
rect 427998 224856 428004 224868
rect 350960 224828 428004 224856
rect 350960 224816 350966 224828
rect 427998 224816 428004 224828
rect 428056 224816 428062 224868
rect 430482 224816 430488 224868
rect 430540 224856 430546 224868
rect 474274 224856 474280 224868
rect 430540 224828 474280 224856
rect 430540 224816 430546 224828
rect 474274 224816 474280 224828
rect 474332 224816 474338 224868
rect 157794 224748 157800 224800
rect 157852 224788 157858 224800
rect 236454 224788 236460 224800
rect 157852 224760 236460 224788
rect 157852 224748 157858 224760
rect 236454 224748 236460 224760
rect 236512 224748 236518 224800
rect 349430 224748 349436 224800
rect 349488 224788 349494 224800
rect 425054 224788 425060 224800
rect 349488 224760 425060 224788
rect 349488 224748 349494 224760
rect 425054 224748 425060 224760
rect 425112 224748 425118 224800
rect 425698 224748 425704 224800
rect 425756 224788 425762 224800
rect 467558 224788 467564 224800
rect 425756 224760 467564 224788
rect 425756 224748 425762 224760
rect 467558 224748 467564 224760
rect 467616 224748 467622 224800
rect 161198 224680 161204 224732
rect 161256 224720 161262 224732
rect 237926 224720 237932 224732
rect 161256 224692 237932 224720
rect 161256 224680 161262 224692
rect 237926 224680 237932 224692
rect 237984 224680 237990 224732
rect 352650 224680 352656 224732
rect 352708 224720 352714 224732
rect 428918 224720 428924 224732
rect 352708 224692 428924 224720
rect 352708 224680 352714 224692
rect 428918 224680 428924 224692
rect 428976 224680 428982 224732
rect 429102 224680 429108 224732
rect 429160 224720 429166 224732
rect 442350 224720 442356 224732
rect 429160 224692 442356 224720
rect 429160 224680 429166 224692
rect 442350 224680 442356 224692
rect 442408 224680 442414 224732
rect 167914 224612 167920 224664
rect 167972 224652 167978 224664
rect 240778 224652 240784 224664
rect 167972 224624 240784 224652
rect 167972 224612 167978 224624
rect 240778 224612 240784 224624
rect 240836 224612 240842 224664
rect 380894 224612 380900 224664
rect 380952 224652 380958 224664
rect 402790 224652 402796 224664
rect 380952 224624 402796 224652
rect 380952 224612 380958 224624
rect 402790 224612 402796 224624
rect 402848 224612 402854 224664
rect 402974 224612 402980 224664
rect 403032 224652 403038 224664
rect 479334 224652 479340 224664
rect 403032 224624 479340 224652
rect 403032 224612 403038 224624
rect 479334 224612 479340 224624
rect 479392 224612 479398 224664
rect 164602 224544 164608 224596
rect 164660 224584 164666 224596
rect 239306 224584 239312 224596
rect 164660 224556 239312 224584
rect 164660 224544 164666 224556
rect 239306 224544 239312 224556
rect 239364 224544 239370 224596
rect 351270 224544 351276 224596
rect 351328 224584 351334 224596
rect 425514 224584 425520 224596
rect 351328 224556 425520 224584
rect 351328 224544 351334 224556
rect 425514 224544 425520 224556
rect 425572 224544 425578 224596
rect 170950 224476 170956 224528
rect 171008 224516 171014 224528
rect 242158 224516 242164 224528
rect 171008 224488 242164 224516
rect 171008 224476 171014 224488
rect 242158 224476 242164 224488
rect 242216 224476 242222 224528
rect 348050 224476 348056 224528
rect 348108 224516 348114 224528
rect 348108 224488 408908 224516
rect 348108 224476 348114 224488
rect 174630 224408 174636 224460
rect 174688 224448 174694 224460
rect 243354 224448 243360 224460
rect 174688 224420 243360 224448
rect 174688 224408 174694 224420
rect 243354 224408 243360 224420
rect 243412 224408 243418 224460
rect 346578 224408 346584 224460
rect 346636 224448 346642 224460
rect 346636 224420 402744 224448
rect 346636 224408 346642 224420
rect 181346 224340 181352 224392
rect 181404 224380 181410 224392
rect 246482 224380 246488 224392
rect 181404 224352 246488 224380
rect 181404 224340 181410 224352
rect 246482 224340 246488 224352
rect 246540 224340 246546 224392
rect 348418 224340 348424 224392
rect 348476 224380 348482 224392
rect 402606 224380 402612 224392
rect 348476 224352 402612 224380
rect 348476 224340 348482 224352
rect 402606 224340 402612 224352
rect 402664 224340 402670 224392
rect 402716 224380 402744 224420
rect 402790 224408 402796 224460
rect 402848 224448 402854 224460
rect 404446 224448 404452 224460
rect 402848 224420 404452 224448
rect 402848 224408 402854 224420
rect 404446 224408 404452 224420
rect 404504 224408 404510 224460
rect 408880 224448 408908 224488
rect 419534 224476 419540 224528
rect 419592 224516 419598 224528
rect 460934 224516 460940 224528
rect 419592 224488 460940 224516
rect 419592 224476 419598 224488
rect 460934 224476 460940 224488
rect 460992 224476 460998 224528
rect 408880 224420 419534 224448
rect 417970 224380 417976 224392
rect 402716 224352 417976 224380
rect 417970 224340 417976 224352
rect 418028 224340 418034 224392
rect 419506 224380 419534 224420
rect 421282 224380 421288 224392
rect 419506 224352 421288 224380
rect 421282 224340 421288 224352
rect 421340 224340 421346 224392
rect 178034 224272 178040 224324
rect 178092 224312 178098 224324
rect 245010 224312 245016 224324
rect 178092 224284 245016 224312
rect 178092 224272 178098 224284
rect 245010 224272 245016 224284
rect 245068 224272 245074 224324
rect 346946 224272 346952 224324
rect 347004 224312 347010 224324
rect 415394 224312 415400 224324
rect 347004 224284 415400 224312
rect 347004 224272 347010 224284
rect 415394 224272 415400 224284
rect 415452 224272 415458 224324
rect 418890 224272 418896 224324
rect 418948 224312 418954 224324
rect 450722 224312 450728 224324
rect 418948 224284 450728 224312
rect 418948 224272 418954 224284
rect 450722 224272 450728 224284
rect 450780 224272 450786 224324
rect 184750 224204 184756 224256
rect 184808 224244 184814 224256
rect 247862 224244 247868 224256
rect 184808 224216 247868 224244
rect 184808 224204 184814 224216
rect 247862 224204 247868 224216
rect 247920 224204 247926 224256
rect 344094 224204 344100 224256
rect 344152 224244 344158 224256
rect 408678 224244 408684 224256
rect 344152 224216 408684 224244
rect 344152 224204 344158 224216
rect 408678 224204 408684 224216
rect 408736 224204 408742 224256
rect 411990 224204 411996 224256
rect 412048 224244 412054 224256
rect 444374 224244 444380 224256
rect 412048 224216 444380 224244
rect 412048 224204 412054 224216
rect 444374 224204 444380 224216
rect 444432 224204 444438 224256
rect 188154 224136 188160 224188
rect 188212 224176 188218 224188
rect 249334 224176 249340 224188
rect 188212 224148 249340 224176
rect 188212 224136 188218 224148
rect 249334 224136 249340 224148
rect 249392 224136 249398 224188
rect 345658 224136 345664 224188
rect 345716 224176 345722 224188
rect 412082 224176 412088 224188
rect 345716 224148 412088 224176
rect 345716 224136 345722 224148
rect 412082 224136 412088 224148
rect 412140 224136 412146 224188
rect 191466 224068 191472 224120
rect 191524 224108 191530 224120
rect 250714 224108 250720 224120
rect 191524 224080 250720 224108
rect 191524 224068 191530 224080
rect 250714 224068 250720 224080
rect 250772 224068 250778 224120
rect 383654 224068 383660 224120
rect 383712 224108 383718 224120
rect 449066 224108 449072 224120
rect 383712 224080 449072 224108
rect 383712 224068 383718 224080
rect 449066 224068 449072 224080
rect 449124 224068 449130 224120
rect 155402 224000 155408 224052
rect 155460 224040 155466 224052
rect 155460 224012 190224 224040
rect 155460 224000 155466 224012
rect 190196 223836 190224 224012
rect 197446 224000 197452 224052
rect 197504 224040 197510 224052
rect 212258 224040 212264 224052
rect 197504 224012 212264 224040
rect 197504 224000 197510 224012
rect 212258 224000 212264 224012
rect 212316 224000 212322 224052
rect 214282 224000 214288 224052
rect 214340 224040 214346 224052
rect 245378 224040 245384 224052
rect 214340 224012 245384 224040
rect 214340 224000 214346 224012
rect 245378 224000 245384 224012
rect 245436 224000 245442 224052
rect 378226 224000 378232 224052
rect 378284 224040 378290 224052
rect 407850 224040 407856 224052
rect 378284 224012 407856 224040
rect 378284 224000 378290 224012
rect 407850 224000 407856 224012
rect 407908 224000 407914 224052
rect 408402 224000 408408 224052
rect 408460 224040 408466 224052
rect 462498 224040 462504 224052
rect 408460 224012 462504 224040
rect 408460 224000 408466 224012
rect 462498 224000 462504 224012
rect 462556 224000 462562 224052
rect 204254 223932 204260 223984
rect 204312 223972 204318 223984
rect 252462 223972 252468 223984
rect 204312 223944 252468 223972
rect 204312 223932 204318 223944
rect 252462 223932 252468 223944
rect 252520 223932 252526 223984
rect 376570 223932 376576 223984
rect 376628 223972 376634 223984
rect 414566 223972 414572 223984
rect 376628 223944 414572 223972
rect 376628 223932 376634 223944
rect 414566 223932 414572 223944
rect 414624 223932 414630 223984
rect 190270 223864 190276 223916
rect 190328 223904 190334 223916
rect 232498 223904 232504 223916
rect 190328 223876 232504 223904
rect 190328 223864 190334 223876
rect 232498 223864 232504 223876
rect 232556 223864 232562 223916
rect 378134 223864 378140 223916
rect 378192 223904 378198 223916
rect 411254 223904 411260 223916
rect 378192 223876 411260 223904
rect 378192 223864 378198 223876
rect 411254 223864 411260 223876
rect 411312 223864 411318 223916
rect 209406 223836 209412 223848
rect 190196 223808 209412 223836
rect 209406 223796 209412 223808
rect 209464 223796 209470 223848
rect 216214 223796 216220 223848
rect 216272 223836 216278 223848
rect 246758 223836 246764 223848
rect 216272 223808 246764 223836
rect 216272 223796 216278 223808
rect 246758 223796 246764 223808
rect 246816 223796 246822 223848
rect 380986 223796 380992 223848
rect 381044 223836 381050 223848
rect 405734 223836 405740 223848
rect 381044 223808 405740 223836
rect 381044 223796 381050 223808
rect 405734 223796 405740 223808
rect 405792 223796 405798 223848
rect 171042 223728 171048 223780
rect 171100 223768 171106 223780
rect 206554 223768 206560 223780
rect 171100 223740 206560 223768
rect 171100 223728 171106 223740
rect 206554 223728 206560 223740
rect 206612 223728 206618 223780
rect 209682 223728 209688 223780
rect 209740 223768 209746 223780
rect 236822 223768 236828 223780
rect 209740 223740 236828 223768
rect 209740 223728 209746 223740
rect 236822 223728 236828 223740
rect 236880 223728 236886 223780
rect 402606 223728 402612 223780
rect 402664 223768 402670 223780
rect 418798 223768 418804 223780
rect 402664 223740 418804 223768
rect 402664 223728 402670 223740
rect 418798 223728 418804 223740
rect 418856 223728 418862 223780
rect 194870 223660 194876 223712
rect 194928 223700 194934 223712
rect 206922 223700 206928 223712
rect 194928 223672 206928 223700
rect 194928 223660 194934 223672
rect 206922 223660 206928 223672
rect 206980 223660 206986 223712
rect 215202 223660 215208 223712
rect 215260 223700 215266 223712
rect 242526 223700 242532 223712
rect 215260 223672 242532 223700
rect 215260 223660 215266 223672
rect 242526 223660 242532 223672
rect 242584 223660 242590 223712
rect 57974 223592 57980 223644
rect 58032 223632 58038 223644
rect 63494 223632 63500 223644
rect 58032 223604 63500 223632
rect 58032 223592 58038 223604
rect 63494 223592 63500 223604
rect 63552 223592 63558 223644
rect 169662 223592 169668 223644
rect 169720 223632 169726 223644
rect 180702 223632 180708 223644
rect 169720 223604 180708 223632
rect 169720 223592 169726 223604
rect 180702 223592 180708 223604
rect 180760 223592 180766 223644
rect 182174 223592 182180 223644
rect 182232 223632 182238 223644
rect 192294 223632 192300 223644
rect 182232 223604 192300 223632
rect 182232 223592 182238 223604
rect 192294 223592 192300 223604
rect 192352 223592 192358 223644
rect 411070 223592 411076 223644
rect 411128 223632 411134 223644
rect 417142 223632 417148 223644
rect 411128 223604 417148 223632
rect 411128 223592 411134 223604
rect 417142 223592 417148 223604
rect 417200 223592 417206 223644
rect 488442 223592 488448 223644
rect 488500 223632 488506 223644
rect 489730 223632 489736 223644
rect 488500 223604 489736 223632
rect 488500 223592 488506 223604
rect 489730 223592 489736 223604
rect 489788 223592 489794 223644
rect 153654 223524 153660 223576
rect 153712 223564 153718 223576
rect 222102 223564 222108 223576
rect 153712 223536 222108 223564
rect 153712 223524 153718 223536
rect 222102 223524 222108 223536
rect 222160 223524 222166 223576
rect 224402 223524 224408 223576
rect 224460 223564 224466 223576
rect 232866 223564 232872 223576
rect 224460 223536 232872 223564
rect 224460 223524 224466 223536
rect 232866 223524 232872 223536
rect 232924 223524 232930 223576
rect 241146 223524 241152 223576
rect 241204 223564 241210 223576
rect 253750 223564 253756 223576
rect 241204 223536 253756 223564
rect 241204 223524 241210 223536
rect 253750 223524 253756 223536
rect 253808 223524 253814 223576
rect 278682 223524 278688 223576
rect 278740 223564 278746 223576
rect 287790 223564 287796 223576
rect 278740 223536 287796 223564
rect 278740 223524 278746 223536
rect 287790 223524 287796 223536
rect 287848 223524 287854 223576
rect 324130 223524 324136 223576
rect 324188 223564 324194 223576
rect 361758 223564 361764 223576
rect 324188 223536 361764 223564
rect 324188 223524 324194 223536
rect 361758 223524 361764 223536
rect 361816 223524 361822 223576
rect 364334 223524 364340 223576
rect 364392 223564 364398 223576
rect 365898 223564 365904 223576
rect 364392 223536 365904 223564
rect 364392 223524 364398 223536
rect 365898 223524 365904 223536
rect 365956 223524 365962 223576
rect 494054 223524 494060 223576
rect 494112 223564 494118 223576
rect 607582 223564 607588 223576
rect 494112 223536 607588 223564
rect 494112 223524 494118 223536
rect 607582 223524 607588 223536
rect 607640 223524 607646 223576
rect 87138 223456 87144 223508
rect 87196 223496 87202 223508
rect 171042 223496 171048 223508
rect 87196 223468 171048 223496
rect 87196 223456 87202 223468
rect 171042 223456 171048 223468
rect 171100 223456 171106 223508
rect 175458 223456 175464 223508
rect 175516 223496 175522 223508
rect 244642 223496 244648 223508
rect 175516 223468 244648 223496
rect 175516 223456 175522 223468
rect 244642 223456 244648 223468
rect 244700 223456 244706 223508
rect 322382 223456 322388 223508
rect 322440 223496 322446 223508
rect 360746 223496 360752 223508
rect 322440 223468 360752 223496
rect 322440 223456 322446 223468
rect 360746 223456 360752 223468
rect 360804 223456 360810 223508
rect 387610 223456 387616 223508
rect 387668 223496 387674 223508
rect 513834 223496 513840 223508
rect 387668 223468 513840 223496
rect 387668 223456 387674 223468
rect 513834 223456 513840 223468
rect 513892 223456 513898 223508
rect 535454 223456 535460 223508
rect 535512 223496 535518 223508
rect 536098 223496 536104 223508
rect 535512 223468 536104 223496
rect 535512 223456 535518 223468
rect 536098 223456 536104 223468
rect 536156 223496 536162 223508
rect 615034 223496 615040 223508
rect 536156 223468 615040 223496
rect 536156 223456 536162 223468
rect 615034 223456 615040 223468
rect 615092 223456 615098 223508
rect 148594 223388 148600 223440
rect 148652 223428 148658 223440
rect 223850 223428 223856 223440
rect 148652 223400 223856 223428
rect 148652 223388 148658 223400
rect 223850 223388 223856 223400
rect 223908 223388 223914 223440
rect 227438 223388 227444 223440
rect 227496 223428 227502 223440
rect 242894 223428 242900 223440
rect 227496 223400 242900 223428
rect 227496 223388 227502 223400
rect 242894 223388 242900 223400
rect 242952 223388 242958 223440
rect 323762 223388 323768 223440
rect 323820 223428 323826 223440
rect 364334 223428 364340 223440
rect 323820 223400 364340 223428
rect 323820 223388 323826 223400
rect 364334 223388 364340 223400
rect 364392 223388 364398 223440
rect 499482 223388 499488 223440
rect 499540 223428 499546 223440
rect 608042 223428 608048 223440
rect 499540 223400 608048 223428
rect 499540 223388 499546 223400
rect 608042 223388 608048 223400
rect 608100 223388 608106 223440
rect 146938 223320 146944 223372
rect 146996 223360 147002 223372
rect 224126 223360 224132 223372
rect 146996 223332 224132 223360
rect 146996 223320 147002 223332
rect 224126 223320 224132 223332
rect 224184 223320 224190 223372
rect 230382 223360 230388 223372
rect 224236 223332 230388 223360
rect 141878 223252 141884 223304
rect 141936 223292 141942 223304
rect 224236 223292 224264 223332
rect 230382 223320 230388 223332
rect 230440 223320 230446 223372
rect 237742 223320 237748 223372
rect 237800 223360 237806 223372
rect 252922 223360 252928 223372
rect 237800 223332 252928 223360
rect 237800 223320 237806 223332
rect 252922 223320 252928 223332
rect 252980 223320 252986 223372
rect 273070 223320 273076 223372
rect 273128 223360 273134 223372
rect 286042 223360 286048 223372
rect 273128 223332 286048 223360
rect 273128 223320 273134 223332
rect 286042 223320 286048 223332
rect 286100 223320 286106 223372
rect 324498 223320 324504 223372
rect 324556 223360 324562 223372
rect 363230 223360 363236 223372
rect 324556 223332 363236 223360
rect 324556 223320 324562 223332
rect 363230 223320 363236 223332
rect 363288 223320 363294 223372
rect 388714 223320 388720 223372
rect 388772 223360 388778 223372
rect 516410 223360 516416 223372
rect 388772 223332 516416 223360
rect 388772 223320 388778 223332
rect 516410 223320 516416 223332
rect 516468 223320 516474 223372
rect 541434 223320 541440 223372
rect 541492 223360 541498 223372
rect 615954 223360 615960 223372
rect 541492 223332 615960 223360
rect 541492 223320 541498 223332
rect 615954 223320 615960 223332
rect 616012 223320 616018 223372
rect 141936 223264 224264 223292
rect 141936 223252 141942 223264
rect 227622 223252 227628 223304
rect 227680 223292 227686 223304
rect 249978 223292 249984 223304
rect 227680 223264 249984 223292
rect 227680 223252 227686 223264
rect 249978 223252 249984 223264
rect 250036 223252 250042 223304
rect 325602 223252 325608 223304
rect 325660 223292 325666 223304
rect 364978 223292 364984 223304
rect 325660 223264 364984 223292
rect 325660 223252 325666 223264
rect 364978 223252 364984 223264
rect 365036 223252 365042 223304
rect 390830 223252 390836 223304
rect 390888 223292 390894 223304
rect 521654 223292 521660 223304
rect 390888 223264 521660 223292
rect 390888 223252 390894 223264
rect 521654 223252 521660 223264
rect 521712 223252 521718 223304
rect 538858 223252 538864 223304
rect 538916 223292 538922 223304
rect 539318 223292 539324 223304
rect 538916 223264 539324 223292
rect 538916 223252 538922 223264
rect 539318 223252 539324 223264
rect 539376 223292 539382 223304
rect 615494 223292 615500 223304
rect 539376 223264 615500 223292
rect 539376 223252 539382 223264
rect 615494 223252 615500 223264
rect 615552 223252 615558 223304
rect 140130 223184 140136 223236
rect 140188 223224 140194 223236
rect 230014 223224 230020 223236
rect 140188 223196 230020 223224
rect 140188 223184 140194 223196
rect 230014 223184 230020 223196
rect 230072 223184 230078 223236
rect 239398 223184 239404 223236
rect 239456 223224 239462 223236
rect 255590 223224 255596 223236
rect 239456 223196 255596 223224
rect 239456 223184 239462 223196
rect 255590 223184 255596 223196
rect 255648 223184 255654 223236
rect 326982 223184 326988 223236
rect 327040 223224 327046 223236
rect 368290 223224 368296 223236
rect 327040 223196 368296 223224
rect 327040 223184 327046 223196
rect 368290 223184 368296 223196
rect 368348 223184 368354 223236
rect 392946 223184 392952 223236
rect 393004 223224 393010 223236
rect 526438 223224 526444 223236
rect 393004 223196 526444 223224
rect 393004 223184 393010 223196
rect 526438 223184 526444 223196
rect 526496 223184 526502 223236
rect 546494 223184 546500 223236
rect 546552 223224 546558 223236
rect 548610 223224 548616 223236
rect 546552 223196 548616 223224
rect 546552 223184 546558 223196
rect 548610 223184 548616 223196
rect 548668 223224 548674 223236
rect 617334 223224 617340 223236
rect 548668 223196 617340 223224
rect 548668 223184 548674 223196
rect 617334 223184 617340 223196
rect 617392 223184 617398 223236
rect 135162 223116 135168 223168
rect 135220 223156 135226 223168
rect 227530 223156 227536 223168
rect 135220 223128 227536 223156
rect 135220 223116 135226 223128
rect 227530 223116 227536 223128
rect 227588 223116 227594 223168
rect 227806 223116 227812 223168
rect 227864 223156 227870 223168
rect 235718 223156 235724 223168
rect 227864 223128 235724 223156
rect 227864 223116 227870 223128
rect 235718 223116 235724 223128
rect 235776 223116 235782 223168
rect 242802 223116 242808 223168
rect 242860 223156 242866 223168
rect 259362 223156 259368 223168
rect 242860 223128 259368 223156
rect 242860 223116 242866 223128
rect 259362 223116 259368 223128
rect 259420 223116 259426 223168
rect 274726 223116 274732 223168
rect 274784 223156 274790 223168
rect 287054 223156 287060 223168
rect 274784 223128 287060 223156
rect 274784 223116 274790 223128
rect 287054 223116 287060 223128
rect 287112 223116 287118 223168
rect 328454 223116 328460 223168
rect 328512 223156 328518 223168
rect 371694 223156 371700 223168
rect 328512 223128 371700 223156
rect 328512 223116 328518 223128
rect 371694 223116 371700 223128
rect 371752 223116 371758 223168
rect 395062 223116 395068 223168
rect 395120 223156 395126 223168
rect 531498 223156 531504 223168
rect 395120 223128 531504 223156
rect 395120 223116 395126 223128
rect 531498 223116 531504 223128
rect 531556 223116 531562 223168
rect 557442 223116 557448 223168
rect 557500 223156 557506 223168
rect 618714 223156 618720 223168
rect 557500 223128 618720 223156
rect 557500 223116 557506 223128
rect 618714 223116 618720 223128
rect 618772 223116 618778 223168
rect 133414 223048 133420 223100
rect 133472 223088 133478 223100
rect 227162 223088 227168 223100
rect 133472 223060 227168 223088
rect 133472 223048 133478 223060
rect 227162 223048 227168 223060
rect 227220 223048 227226 223100
rect 231026 223048 231032 223100
rect 231084 223088 231090 223100
rect 248598 223088 248604 223100
rect 231084 223060 248604 223088
rect 231084 223048 231090 223060
rect 248598 223048 248604 223060
rect 248656 223048 248662 223100
rect 271414 223048 271420 223100
rect 271472 223088 271478 223100
rect 271472 223060 281166 223088
rect 271472 223048 271478 223060
rect 128354 222980 128360 223032
rect 128412 223020 128418 223032
rect 224678 223020 224684 223032
rect 128412 222992 224684 223020
rect 128412 222980 128418 222992
rect 224678 222980 224684 222992
rect 224736 222980 224742 223032
rect 233234 223020 233240 223032
rect 224788 222992 233240 223020
rect 77938 222912 77944 222964
rect 77996 222952 78002 222964
rect 121178 222952 121184 222964
rect 77996 222924 121184 222952
rect 77996 222912 78002 222924
rect 121178 222912 121184 222924
rect 121236 222912 121242 222964
rect 126698 222912 126704 222964
rect 126756 222952 126762 222964
rect 224034 222952 224040 222964
rect 126756 222924 224040 222952
rect 126756 222912 126762 222924
rect 224034 222912 224040 222924
rect 224092 222912 224098 222964
rect 224788 222952 224816 222992
rect 233234 222980 233240 222992
rect 233292 222980 233298 223032
rect 236086 222980 236092 223032
rect 236144 223020 236150 223032
rect 255406 223020 255412 223032
rect 236144 222992 255412 223020
rect 236144 222980 236150 222992
rect 255406 222980 255412 222992
rect 255464 222980 255470 223032
rect 224144 222924 224816 222952
rect 116578 222844 116584 222896
rect 116636 222884 116642 222896
rect 220078 222884 220084 222896
rect 116636 222856 220084 222884
rect 116636 222844 116642 222856
rect 220078 222844 220084 222856
rect 220136 222844 220142 222896
rect 223850 222844 223856 222896
rect 223908 222884 223914 222896
rect 224144 222884 224172 222924
rect 232682 222912 232688 222964
rect 232740 222952 232746 222964
rect 254670 222952 254676 222964
rect 232740 222924 254676 222952
rect 232740 222912 232746 222924
rect 254670 222912 254676 222924
rect 254728 222912 254734 222964
rect 263778 222912 263784 222964
rect 263836 222952 263842 222964
rect 280982 222952 280988 222964
rect 263836 222924 280988 222952
rect 263836 222912 263842 222924
rect 280982 222912 280988 222924
rect 281040 222912 281046 222964
rect 223908 222856 224172 222884
rect 223908 222844 223914 222856
rect 224310 222844 224316 222896
rect 224368 222884 224374 222896
rect 248506 222884 248512 222896
rect 224368 222856 248512 222884
rect 224368 222844 224374 222856
rect 248506 222844 248512 222856
rect 248564 222844 248570 222896
rect 257062 222844 257068 222896
rect 257120 222884 257126 222896
rect 278130 222884 278136 222896
rect 257120 222856 278136 222884
rect 257120 222844 257126 222856
rect 278130 222844 278136 222856
rect 278188 222844 278194 222896
rect 281138 222884 281166 223060
rect 326338 223048 326344 223100
rect 326396 223088 326402 223100
rect 369118 223088 369124 223100
rect 326396 223060 369124 223088
rect 326396 223048 326402 223060
rect 369118 223048 369124 223060
rect 369176 223048 369182 223100
rect 395430 223048 395436 223100
rect 395488 223088 395494 223100
rect 532694 223088 532700 223100
rect 395488 223060 532700 223088
rect 395488 223048 395494 223060
rect 532694 223048 532700 223060
rect 532752 223048 532758 223100
rect 565998 223048 566004 223100
rect 566056 223088 566062 223100
rect 620554 223088 620560 223100
rect 566056 223060 620560 223088
rect 566056 223048 566062 223060
rect 620554 223048 620560 223060
rect 620612 223048 620618 223100
rect 324866 222980 324872 223032
rect 324924 223020 324930 223032
rect 365806 223020 365812 223032
rect 324924 222992 365812 223020
rect 324924 222980 324930 222992
rect 365806 222980 365812 222992
rect 365864 222980 365870 223032
rect 365898 222980 365904 223032
rect 365956 223020 365962 223032
rect 382642 223020 382648 223032
rect 365956 222992 382648 223020
rect 365956 222980 365962 222992
rect 382642 222980 382648 222992
rect 382700 222980 382706 223032
rect 397270 222980 397276 223032
rect 397328 223020 397334 223032
rect 536558 223020 536564 223032
rect 397328 222992 536564 223020
rect 397328 222980 397334 222992
rect 536558 222980 536564 222992
rect 536616 222980 536622 223032
rect 326614 222912 326620 222964
rect 326672 222952 326678 222964
rect 370866 222952 370872 222964
rect 326672 222924 370872 222952
rect 326672 222912 326678 222924
rect 370866 222912 370872 222924
rect 370924 222912 370930 222964
rect 399386 222912 399392 222964
rect 399444 222952 399450 222964
rect 541618 222952 541624 222964
rect 399444 222924 541624 222952
rect 399444 222912 399450 222924
rect 541618 222912 541624 222924
rect 541676 222912 541682 222964
rect 285674 222884 285680 222896
rect 281138 222856 285680 222884
rect 285674 222844 285680 222856
rect 285732 222844 285738 222896
rect 327350 222844 327356 222896
rect 327408 222884 327414 222896
rect 370038 222884 370044 222896
rect 327408 222856 370044 222884
rect 327408 222844 327414 222856
rect 370038 222844 370044 222856
rect 370096 222844 370102 222896
rect 370222 222844 370228 222896
rect 370280 222884 370286 222896
rect 400398 222884 400404 222896
rect 370280 222856 400404 222884
rect 370280 222844 370286 222856
rect 400398 222844 400404 222856
rect 400456 222844 400462 222896
rect 400766 222844 400772 222896
rect 400824 222884 400830 222896
rect 545114 222884 545120 222896
rect 400824 222856 545120 222884
rect 400824 222844 400830 222856
rect 545114 222844 545120 222856
rect 545172 222844 545178 222896
rect 568574 222844 568580 222896
rect 568632 222884 568638 222896
rect 621014 222884 621020 222896
rect 568632 222856 621020 222884
rect 568632 222844 568638 222856
rect 621014 222844 621020 222856
rect 621072 222844 621078 222896
rect 119982 222776 119988 222828
rect 120040 222816 120046 222828
rect 221458 222816 221464 222828
rect 120040 222788 221464 222816
rect 120040 222776 120046 222788
rect 221458 222776 221464 222788
rect 221516 222776 221522 222828
rect 222562 222776 222568 222828
rect 222620 222816 222626 222828
rect 256970 222816 256976 222828
rect 222620 222788 256976 222816
rect 222620 222776 222626 222788
rect 256970 222776 256976 222788
rect 257028 222776 257034 222828
rect 261294 222776 261300 222828
rect 261352 222816 261358 222828
rect 281350 222816 281356 222828
rect 261352 222788 281356 222816
rect 261352 222776 261358 222788
rect 281350 222776 281356 222788
rect 281408 222776 281414 222828
rect 325234 222776 325240 222828
rect 325292 222816 325298 222828
rect 367462 222816 367468 222828
rect 325292 222788 367468 222816
rect 325292 222776 325298 222788
rect 367462 222776 367468 222788
rect 367520 222776 367526 222828
rect 369578 222776 369584 222828
rect 369636 222816 369642 222828
rect 398558 222816 398564 222828
rect 369636 222788 398564 222816
rect 369636 222776 369642 222788
rect 398558 222776 398564 222788
rect 398616 222776 398622 222828
rect 400122 222776 400128 222828
rect 400180 222816 400186 222828
rect 543642 222816 543648 222828
rect 400180 222788 543648 222816
rect 400180 222776 400186 222788
rect 543642 222776 543648 222788
rect 543700 222776 543706 222828
rect 545758 222776 545764 222828
rect 545816 222816 545822 222828
rect 616874 222816 616880 222828
rect 545816 222788 616880 222816
rect 545816 222776 545822 222788
rect 616874 222776 616880 222788
rect 616932 222776 616938 222828
rect 91370 222708 91376 222760
rect 91428 222748 91434 222760
rect 197262 222748 197268 222760
rect 91428 222720 197268 222748
rect 91428 222708 91434 222720
rect 197262 222708 197268 222720
rect 197320 222708 197326 222760
rect 207474 222708 207480 222760
rect 207532 222748 207538 222760
rect 245654 222748 245660 222760
rect 207532 222720 245660 222748
rect 207532 222708 207538 222720
rect 245654 222708 245660 222720
rect 245712 222708 245718 222760
rect 266354 222708 266360 222760
rect 266412 222748 266418 222760
rect 283190 222748 283196 222760
rect 266412 222720 283196 222748
rect 266412 222708 266418 222720
rect 283190 222708 283196 222720
rect 283248 222708 283254 222760
rect 328086 222708 328092 222760
rect 328144 222748 328150 222760
rect 374178 222748 374184 222760
rect 328144 222720 374184 222748
rect 328144 222708 328150 222720
rect 374178 222708 374184 222720
rect 374236 222708 374242 222760
rect 401502 222708 401508 222760
rect 401560 222748 401566 222760
rect 546678 222748 546684 222760
rect 401560 222720 546684 222748
rect 401560 222708 401566 222720
rect 546678 222708 546684 222720
rect 546736 222708 546742 222760
rect 85482 222640 85488 222692
rect 85540 222680 85546 222692
rect 192846 222680 192852 222692
rect 85540 222652 192852 222680
rect 85540 222640 85546 222652
rect 192846 222640 192852 222652
rect 192904 222640 192910 222692
rect 203978 222680 203984 222692
rect 193048 222652 203984 222680
rect 82170 222572 82176 222624
rect 82228 222612 82234 222624
rect 193048 222612 193076 222652
rect 203978 222640 203984 222652
rect 204036 222640 204042 222692
rect 215846 222640 215852 222692
rect 215904 222680 215910 222692
rect 256694 222680 256700 222692
rect 215904 222652 256700 222680
rect 215904 222640 215910 222652
rect 256694 222640 256700 222652
rect 256752 222640 256758 222692
rect 260466 222640 260472 222692
rect 260524 222680 260530 222692
rect 279602 222680 279608 222692
rect 260524 222652 279608 222680
rect 260524 222640 260530 222652
rect 279602 222640 279608 222652
rect 279660 222640 279666 222692
rect 329466 222640 329472 222692
rect 329524 222680 329530 222692
rect 377582 222680 377588 222692
rect 329524 222652 377588 222680
rect 329524 222640 329530 222652
rect 377582 222640 377588 222652
rect 377640 222640 377646 222692
rect 403342 222640 403348 222692
rect 403400 222680 403406 222692
rect 549346 222680 549352 222692
rect 403400 222652 549352 222680
rect 403400 222640 403406 222652
rect 549346 222640 549352 222652
rect 549404 222640 549410 222692
rect 563698 222640 563704 222692
rect 563756 222680 563762 222692
rect 620094 222680 620100 222692
rect 563756 222652 620100 222680
rect 563756 222640 563762 222652
rect 620094 222640 620100 222652
rect 620152 222640 620158 222692
rect 82228 222584 193076 222612
rect 82228 222572 82234 222584
rect 193122 222572 193128 222624
rect 193180 222612 193186 222624
rect 201310 222612 201316 222624
rect 193180 222584 201316 222612
rect 193180 222572 193186 222584
rect 201310 222572 201316 222584
rect 201368 222572 201374 222624
rect 209130 222572 209136 222624
rect 209188 222612 209194 222624
rect 258902 222612 258908 222624
rect 209188 222584 258908 222612
rect 209188 222572 209194 222584
rect 258902 222572 258908 222584
rect 258960 222572 258966 222624
rect 262950 222572 262956 222624
rect 263008 222612 263014 222624
rect 281718 222612 281724 222624
rect 263008 222584 281724 222612
rect 263008 222572 263014 222584
rect 281718 222572 281724 222584
rect 281776 222572 281782 222624
rect 284938 222612 284944 222624
rect 281828 222584 284944 222612
rect 75362 222504 75368 222556
rect 75420 222544 75426 222556
rect 201126 222544 201132 222556
rect 75420 222516 201132 222544
rect 75420 222504 75426 222516
rect 201126 222504 201132 222516
rect 201184 222504 201190 222556
rect 205818 222504 205824 222556
rect 205876 222544 205882 222556
rect 257522 222544 257528 222556
rect 205876 222516 257528 222544
rect 205876 222504 205882 222516
rect 257522 222504 257528 222516
rect 257580 222504 257586 222556
rect 262122 222504 262128 222556
rect 262180 222544 262186 222556
rect 280706 222544 280712 222556
rect 262180 222516 280712 222544
rect 262180 222504 262186 222516
rect 280706 222504 280712 222516
rect 280764 222504 280770 222556
rect 72878 222436 72884 222488
rect 72936 222476 72942 222488
rect 193122 222476 193128 222488
rect 72936 222448 193128 222476
rect 72936 222436 72942 222448
rect 193122 222436 193128 222448
rect 193180 222436 193186 222488
rect 193214 222436 193220 222488
rect 193272 222476 193278 222488
rect 195790 222476 195796 222488
rect 193272 222448 195796 222476
rect 193272 222436 193278 222448
rect 195790 222436 195796 222448
rect 195848 222436 195854 222488
rect 202414 222436 202420 222488
rect 202472 222476 202478 222488
rect 256050 222476 256056 222488
rect 202472 222448 256056 222476
rect 202472 222436 202478 222448
rect 256050 222436 256056 222448
rect 256108 222436 256114 222488
rect 257890 222436 257896 222488
rect 257948 222476 257954 222488
rect 279970 222476 279976 222488
rect 257948 222448 279976 222476
rect 257948 222436 257954 222448
rect 279970 222436 279976 222448
rect 280028 222436 280034 222488
rect 68646 222368 68652 222420
rect 68704 222408 68710 222420
rect 198274 222408 198280 222420
rect 68704 222380 198280 222408
rect 68704 222368 68710 222380
rect 198274 222368 198280 222380
rect 198332 222368 198338 222420
rect 200758 222368 200764 222420
rect 200816 222408 200822 222420
rect 255682 222408 255688 222420
rect 200816 222380 255688 222408
rect 200816 222368 200822 222380
rect 255682 222368 255688 222380
rect 255740 222368 255746 222420
rect 272242 222368 272248 222420
rect 272300 222408 272306 222420
rect 281828 222408 281856 222584
rect 284938 222572 284944 222584
rect 284996 222572 285002 222624
rect 329834 222572 329840 222624
rect 329892 222612 329898 222624
rect 375374 222612 375380 222624
rect 329892 222584 375380 222612
rect 329892 222572 329898 222584
rect 375374 222572 375380 222584
rect 375432 222572 375438 222624
rect 376662 222572 376668 222624
rect 376720 222612 376726 222624
rect 394694 222612 394700 222624
rect 376720 222584 394700 222612
rect 376720 222572 376726 222584
rect 394694 222572 394700 222584
rect 394752 222572 394758 222624
rect 403250 222572 403256 222624
rect 403308 222612 403314 222624
rect 549990 222612 549996 222624
rect 403308 222584 549996 222612
rect 403308 222572 403314 222584
rect 549990 222572 549996 222584
rect 550048 222572 550054 222624
rect 553762 222572 553768 222624
rect 553820 222612 553826 222624
rect 553820 222584 554360 222612
rect 553820 222572 553826 222584
rect 554332 222556 554360 222584
rect 561214 222572 561220 222624
rect 561272 222612 561278 222624
rect 619634 222612 619640 222624
rect 561272 222584 619640 222612
rect 561272 222572 561278 222584
rect 619634 222572 619640 222584
rect 619692 222572 619698 222624
rect 283190 222504 283196 222556
rect 283248 222544 283254 222556
rect 290274 222544 290280 222556
rect 283248 222516 290280 222544
rect 283248 222504 283254 222516
rect 290274 222504 290280 222516
rect 290332 222504 290338 222556
rect 331582 222504 331588 222556
rect 331640 222544 331646 222556
rect 378410 222544 378416 222556
rect 331640 222516 378416 222544
rect 331640 222504 331646 222516
rect 378410 222504 378416 222516
rect 378468 222504 378474 222556
rect 404722 222504 404728 222556
rect 404780 222544 404786 222556
rect 554222 222544 554228 222556
rect 404780 222516 554228 222544
rect 404780 222504 404786 222516
rect 554222 222504 554228 222516
rect 554280 222504 554286 222556
rect 554314 222504 554320 222556
rect 554372 222544 554378 222556
rect 618254 222544 618260 222556
rect 554372 222516 618260 222544
rect 554372 222504 554378 222516
rect 618254 222504 618260 222516
rect 618312 222504 618318 222556
rect 327718 222436 327724 222488
rect 327776 222476 327782 222488
rect 372614 222476 372620 222488
rect 327776 222448 372620 222476
rect 327776 222436 327782 222448
rect 372614 222436 372620 222448
rect 372672 222436 372678 222488
rect 373902 222436 373908 222488
rect 373960 222476 373966 222488
rect 397730 222476 397736 222488
rect 373960 222448 397736 222476
rect 373960 222436 373966 222448
rect 397730 222436 397736 222448
rect 397788 222436 397794 222488
rect 405826 222436 405832 222488
rect 405884 222476 405890 222488
rect 556706 222476 556712 222488
rect 405884 222448 556712 222476
rect 405884 222436 405890 222448
rect 556706 222436 556712 222448
rect 556764 222436 556770 222488
rect 559098 222436 559104 222488
rect 559156 222476 559162 222488
rect 619174 222476 619180 222488
rect 559156 222448 619180 222476
rect 559156 222436 559162 222448
rect 619174 222436 619180 222448
rect 619232 222436 619238 222488
rect 272300 222380 281856 222408
rect 272300 222368 272306 222380
rect 332686 222368 332692 222420
rect 332744 222408 332750 222420
rect 351914 222408 351920 222420
rect 332744 222380 351920 222408
rect 332744 222368 332750 222380
rect 351914 222368 351920 222380
rect 351972 222368 351978 222420
rect 352006 222368 352012 222420
rect 352064 222408 352070 222420
rect 376754 222408 376760 222420
rect 352064 222380 376760 222408
rect 352064 222368 352070 222380
rect 376754 222368 376760 222380
rect 376812 222368 376818 222420
rect 376846 222368 376852 222420
rect 376904 222408 376910 222420
rect 401134 222408 401140 222420
rect 376904 222380 401140 222408
rect 376904 222368 376910 222380
rect 401134 222368 401140 222380
rect 401192 222368 401198 222420
rect 405090 222368 405096 222420
rect 405148 222408 405154 222420
rect 555050 222408 555056 222420
rect 405148 222380 555056 222408
rect 405148 222368 405154 222380
rect 555050 222368 555056 222380
rect 555108 222368 555114 222420
rect 562870 222368 562876 222420
rect 562928 222408 562934 222420
rect 634538 222408 634544 222420
rect 562928 222380 634544 222408
rect 562928 222368 562934 222380
rect 634538 222368 634544 222380
rect 634596 222368 634602 222420
rect 53558 222300 53564 222352
rect 53616 222340 53622 222352
rect 182174 222340 182180 222352
rect 53616 222312 182180 222340
rect 53616 222300 53622 222312
rect 182174 222300 182180 222312
rect 182232 222300 182238 222352
rect 187234 222300 187240 222352
rect 187292 222340 187298 222352
rect 227622 222340 227628 222352
rect 187292 222312 227628 222340
rect 187292 222300 187298 222312
rect 227622 222300 227628 222312
rect 227680 222300 227686 222352
rect 259362 222300 259368 222352
rect 259420 222340 259426 222352
rect 280338 222340 280344 222352
rect 259420 222312 280344 222340
rect 259420 222300 259426 222312
rect 280338 222300 280344 222312
rect 280396 222300 280402 222352
rect 310974 222300 310980 222352
rect 311032 222340 311038 222352
rect 333974 222340 333980 222352
rect 311032 222312 333980 222340
rect 311032 222300 311038 222312
rect 333974 222300 333980 222312
rect 334032 222300 334038 222352
rect 334158 222300 334164 222352
rect 334216 222340 334222 222352
rect 385126 222340 385132 222352
rect 334216 222312 385132 222340
rect 334216 222300 334222 222312
rect 385126 222300 385132 222312
rect 385184 222300 385190 222352
rect 405458 222300 405464 222352
rect 405516 222340 405522 222352
rect 556246 222340 556252 222352
rect 405516 222312 556252 222340
rect 405516 222300 405522 222312
rect 556246 222300 556252 222312
rect 556304 222340 556310 222352
rect 557442 222340 557448 222352
rect 556304 222312 557448 222340
rect 556304 222300 556310 222312
rect 557442 222300 557448 222312
rect 557500 222300 557506 222352
rect 557626 222300 557632 222352
rect 557684 222340 557690 222352
rect 633618 222340 633624 222352
rect 557684 222312 633624 222340
rect 557684 222300 557690 222312
rect 633618 222300 633624 222312
rect 633676 222300 633682 222352
rect 61930 222232 61936 222284
rect 61988 222272 61994 222284
rect 195422 222272 195428 222284
rect 61988 222244 195428 222272
rect 61988 222232 61994 222244
rect 195422 222232 195428 222244
rect 195480 222232 195486 222284
rect 195698 222232 195704 222284
rect 195756 222272 195762 222284
rect 253198 222272 253204 222284
rect 195756 222244 253204 222272
rect 195756 222232 195762 222244
rect 253198 222232 253204 222244
rect 253256 222232 253262 222284
rect 254578 222232 254584 222284
rect 254636 222272 254642 222284
rect 278498 222272 278504 222284
rect 254636 222244 278504 222272
rect 254636 222232 254642 222244
rect 278498 222232 278504 222244
rect 278556 222232 278562 222284
rect 337378 222232 337384 222284
rect 337436 222272 337442 222284
rect 337436 222244 351868 222272
rect 337436 222232 337442 222244
rect 59446 222164 59452 222216
rect 59504 222204 59510 222216
rect 193214 222204 193220 222216
rect 59504 222176 193220 222204
rect 59504 222164 59510 222176
rect 193214 222164 193220 222176
rect 193272 222164 193278 222216
rect 194042 222164 194048 222216
rect 194100 222204 194106 222216
rect 252830 222204 252836 222216
rect 194100 222176 252836 222204
rect 194100 222164 194106 222176
rect 252830 222164 252836 222176
rect 252888 222164 252894 222216
rect 255406 222164 255412 222216
rect 255464 222204 255470 222216
rect 277854 222204 277860 222216
rect 255464 222176 277860 222204
rect 255464 222164 255470 222176
rect 277854 222164 277860 222176
rect 277912 222164 277918 222216
rect 314194 222164 314200 222216
rect 314252 222204 314258 222216
rect 338022 222204 338028 222216
rect 314252 222176 338028 222204
rect 314252 222164 314258 222176
rect 338022 222164 338028 222176
rect 338080 222164 338086 222216
rect 338114 222164 338120 222216
rect 338172 222204 338178 222216
rect 343082 222204 343088 222216
rect 338172 222176 343088 222204
rect 338172 222164 338178 222176
rect 343082 222164 343088 222176
rect 343140 222164 343146 222216
rect 351840 222204 351868 222244
rect 351914 222232 351920 222284
rect 351972 222272 351978 222284
rect 381814 222272 381820 222284
rect 351972 222244 381820 222272
rect 351972 222232 351978 222244
rect 381814 222232 381820 222244
rect 381872 222232 381878 222284
rect 396166 222232 396172 222284
rect 396224 222272 396230 222284
rect 401962 222272 401968 222284
rect 396224 222244 401968 222272
rect 396224 222232 396230 222244
rect 401962 222232 401968 222244
rect 402020 222232 402026 222284
rect 409322 222232 409328 222284
rect 409380 222272 409386 222284
rect 565170 222272 565176 222284
rect 409380 222244 565176 222272
rect 409380 222232 409386 222244
rect 565170 222232 565176 222244
rect 565228 222232 565234 222284
rect 393590 222204 393596 222216
rect 351840 222176 393596 222204
rect 393590 222164 393596 222176
rect 393648 222164 393654 222216
rect 400030 222164 400036 222216
rect 400088 222204 400094 222216
rect 403618 222204 403624 222216
rect 400088 222176 403624 222204
rect 400088 222164 400094 222176
rect 403618 222164 403624 222176
rect 403676 222164 403682 222216
rect 543642 222164 543648 222216
rect 543700 222204 543706 222216
rect 616414 222204 616420 222216
rect 543700 222176 616420 222204
rect 543700 222164 543706 222176
rect 616414 222164 616420 222176
rect 616472 222164 616478 222216
rect 155310 222096 155316 222148
rect 155368 222136 155374 222148
rect 219986 222136 219992 222148
rect 155368 222108 219992 222136
rect 155368 222096 155374 222108
rect 219986 222096 219992 222108
rect 220044 222096 220050 222148
rect 220078 222096 220084 222148
rect 220136 222136 220142 222148
rect 234614 222136 234620 222148
rect 220136 222108 234620 222136
rect 220136 222096 220142 222108
rect 234614 222096 234620 222108
rect 234672 222096 234678 222148
rect 269666 222096 269672 222148
rect 269724 222136 269730 222148
rect 284570 222136 284576 222148
rect 269724 222108 284576 222136
rect 269724 222096 269730 222108
rect 284570 222096 284576 222108
rect 284628 222096 284634 222148
rect 320910 222096 320916 222148
rect 320968 222136 320974 222148
rect 357342 222136 357348 222148
rect 320968 222108 357348 222136
rect 320968 222096 320974 222108
rect 357342 222096 357348 222108
rect 357400 222096 357406 222148
rect 384022 222096 384028 222148
rect 384080 222136 384086 222148
rect 505738 222136 505744 222148
rect 384080 222108 505744 222136
rect 384080 222096 384086 222108
rect 505738 222096 505744 222108
rect 505796 222096 505802 222148
rect 532786 222096 532792 222148
rect 532844 222136 532850 222148
rect 533430 222136 533436 222148
rect 532844 222108 533436 222136
rect 532844 222096 532850 222108
rect 533430 222096 533436 222108
rect 533488 222136 533494 222148
rect 614574 222136 614580 222148
rect 533488 222108 614580 222136
rect 533488 222096 533494 222108
rect 614574 222096 614580 222108
rect 614632 222096 614638 222148
rect 93762 222028 93768 222080
rect 93820 222068 93826 222080
rect 155402 222068 155408 222080
rect 93820 222040 155408 222068
rect 93820 222028 93826 222040
rect 155402 222028 155408 222040
rect 155460 222028 155466 222080
rect 160370 222028 160376 222080
rect 160428 222068 160434 222080
rect 238294 222068 238300 222080
rect 160428 222040 238300 222068
rect 160428 222028 160434 222040
rect 238294 222028 238300 222040
rect 238352 222028 238358 222080
rect 244458 222028 244464 222080
rect 244516 222068 244522 222080
rect 256142 222068 256148 222080
rect 244516 222040 256148 222068
rect 244516 222028 244522 222040
rect 256142 222028 256148 222040
rect 256200 222028 256206 222080
rect 319806 222028 319812 222080
rect 319864 222068 319870 222080
rect 354030 222068 354036 222080
rect 319864 222040 354036 222068
rect 319864 222028 319870 222040
rect 354030 222028 354036 222040
rect 354088 222028 354094 222080
rect 383378 222028 383384 222080
rect 383436 222068 383442 222080
rect 503714 222068 503720 222080
rect 383436 222040 503720 222068
rect 383436 222028 383442 222040
rect 503714 222028 503720 222040
rect 503772 222028 503778 222080
rect 552566 222028 552572 222080
rect 552624 222068 552630 222080
rect 553210 222068 553216 222080
rect 552624 222040 553216 222068
rect 552624 222028 552630 222040
rect 553210 222028 553216 222040
rect 553268 222068 553274 222080
rect 632698 222068 632704 222080
rect 553268 222040 632704 222068
rect 553268 222028 553274 222040
rect 632698 222028 632704 222040
rect 632756 222028 632762 222080
rect 162026 221960 162032 222012
rect 162084 222000 162090 222012
rect 238938 222000 238944 222012
rect 162084 221972 238944 222000
rect 162084 221960 162090 221972
rect 238938 221960 238944 221972
rect 238996 221960 239002 222012
rect 322750 221960 322756 222012
rect 322808 222000 322814 222012
rect 358262 222000 358268 222012
rect 322808 221972 358268 222000
rect 322808 221960 322814 221972
rect 358262 221960 358268 221972
rect 358320 221960 358326 222012
rect 381906 221960 381912 222012
rect 381964 222000 381970 222012
rect 501046 222000 501052 222012
rect 381964 221972 501052 222000
rect 381964 221960 381970 221972
rect 501046 221960 501052 221972
rect 501104 221960 501110 222012
rect 547782 221960 547788 222012
rect 547840 222000 547846 222012
rect 631778 222000 631784 222012
rect 547840 221972 631784 222000
rect 547840 221960 547846 221972
rect 631778 221960 631784 221972
rect 631836 221960 631842 222012
rect 170490 221892 170496 221944
rect 170548 221932 170554 221944
rect 227438 221932 227444 221944
rect 170548 221904 227444 221932
rect 170548 221892 170554 221904
rect 227438 221892 227444 221904
rect 227496 221892 227502 221944
rect 241790 221932 241796 221944
rect 227548 221904 241796 221932
rect 168742 221824 168748 221876
rect 168800 221864 168806 221876
rect 227548 221864 227576 221904
rect 241790 221892 241796 221904
rect 241848 221892 241854 221944
rect 275554 221892 275560 221944
rect 275612 221932 275618 221944
rect 286410 221932 286416 221944
rect 275612 221904 286416 221932
rect 275612 221892 275618 221904
rect 286410 221892 286416 221904
rect 286468 221892 286474 221944
rect 316678 221892 316684 221944
rect 316736 221932 316742 221944
rect 347314 221932 347320 221944
rect 316736 221904 347320 221932
rect 316736 221892 316742 221904
rect 347314 221892 347320 221904
rect 347372 221892 347378 221944
rect 347406 221892 347412 221944
rect 347464 221932 347470 221944
rect 380066 221932 380072 221944
rect 347464 221904 380072 221932
rect 347464 221892 347470 221904
rect 380066 221892 380072 221904
rect 380124 221892 380130 221944
rect 382274 221892 382280 221944
rect 382332 221932 382338 221944
rect 501230 221932 501236 221944
rect 382332 221904 501236 221932
rect 382332 221892 382338 221904
rect 501230 221892 501236 221904
rect 501288 221892 501294 221944
rect 530670 221892 530676 221944
rect 530728 221932 530734 221944
rect 614022 221932 614028 221944
rect 530728 221904 614028 221932
rect 530728 221892 530734 221904
rect 614022 221892 614028 221904
rect 614080 221892 614086 221944
rect 239674 221864 239680 221876
rect 168800 221836 227576 221864
rect 227640 221836 239680 221864
rect 168800 221824 168806 221836
rect 166258 221756 166264 221808
rect 166316 221796 166322 221808
rect 227640 221796 227668 221836
rect 239674 221824 239680 221836
rect 239732 221824 239738 221876
rect 321278 221824 321284 221876
rect 321336 221864 321342 221876
rect 354858 221864 354864 221876
rect 321336 221836 354864 221864
rect 321336 221824 321342 221836
rect 354858 221824 354864 221836
rect 354916 221824 354922 221876
rect 380526 221824 380532 221876
rect 380584 221864 380590 221876
rect 497366 221864 497372 221876
rect 380584 221836 497372 221864
rect 380584 221824 380590 221836
rect 497366 221824 497372 221836
rect 497424 221864 497430 221876
rect 499482 221864 499488 221876
rect 497424 221836 499488 221864
rect 497424 221824 497430 221836
rect 499482 221824 499488 221836
rect 499540 221824 499546 221876
rect 528094 221824 528100 221876
rect 528152 221864 528158 221876
rect 613562 221864 613568 221876
rect 528152 221836 613568 221864
rect 528152 221824 528158 221836
rect 613562 221824 613568 221836
rect 613620 221824 613626 221876
rect 166316 221768 227668 221796
rect 166316 221756 166322 221768
rect 234338 221756 234344 221808
rect 234396 221796 234402 221808
rect 248414 221796 248420 221808
rect 234396 221768 248420 221796
rect 234396 221756 234402 221768
rect 248414 221756 248420 221768
rect 248472 221756 248478 221808
rect 278130 221756 278136 221808
rect 278188 221796 278194 221808
rect 288526 221796 288532 221808
rect 278188 221768 288532 221796
rect 278188 221756 278194 221768
rect 288526 221756 288532 221768
rect 288584 221756 288590 221808
rect 319898 221756 319904 221808
rect 319956 221796 319962 221808
rect 351454 221796 351460 221808
rect 319956 221768 351460 221796
rect 319956 221756 319962 221768
rect 351454 221756 351460 221768
rect 351512 221756 351518 221808
rect 377950 221756 377956 221808
rect 378008 221796 378014 221808
rect 491294 221796 491300 221808
rect 378008 221768 491300 221796
rect 378008 221756 378014 221768
rect 491294 221756 491300 221768
rect 491352 221756 491358 221808
rect 542722 221756 542728 221808
rect 542780 221796 542786 221808
rect 630858 221796 630864 221808
rect 542780 221768 630864 221796
rect 542780 221756 542786 221768
rect 630858 221756 630864 221768
rect 630916 221756 630922 221808
rect 177206 221688 177212 221740
rect 177264 221728 177270 221740
rect 245746 221728 245752 221740
rect 177264 221700 245752 221728
rect 177264 221688 177270 221700
rect 245746 221688 245752 221700
rect 245804 221688 245810 221740
rect 281442 221688 281448 221740
rect 281500 221728 281506 221740
rect 289906 221728 289912 221740
rect 281500 221700 289912 221728
rect 281500 221688 281506 221700
rect 289906 221688 289912 221700
rect 289964 221688 289970 221740
rect 318058 221688 318064 221740
rect 318116 221728 318122 221740
rect 350626 221728 350632 221740
rect 318116 221700 350632 221728
rect 318116 221688 318122 221700
rect 350626 221688 350632 221700
rect 350684 221688 350690 221740
rect 380802 221688 380808 221740
rect 380860 221728 380866 221740
rect 497826 221728 497832 221740
rect 380860 221700 497832 221728
rect 380860 221688 380866 221700
rect 497826 221688 497832 221700
rect 497884 221688 497890 221740
rect 538306 221688 538312 221740
rect 538364 221728 538370 221740
rect 540146 221728 540152 221740
rect 538364 221700 540152 221728
rect 538364 221688 538370 221700
rect 540146 221688 540152 221700
rect 540204 221728 540210 221740
rect 630398 221728 630404 221740
rect 540204 221700 630404 221728
rect 540204 221688 540210 221700
rect 630398 221688 630404 221700
rect 630456 221688 630462 221740
rect 183922 221620 183928 221672
rect 183980 221660 183986 221672
rect 248322 221660 248328 221672
rect 183980 221632 248328 221660
rect 183980 221620 183986 221632
rect 248322 221620 248328 221632
rect 248380 221620 248386 221672
rect 264606 221620 264612 221672
rect 264664 221660 264670 221672
rect 282822 221660 282828 221672
rect 264664 221632 282828 221660
rect 264664 221620 264670 221632
rect 282822 221620 282828 221632
rect 282880 221620 282886 221672
rect 317046 221620 317052 221672
rect 317104 221660 317110 221672
rect 345014 221660 345020 221672
rect 317104 221632 345020 221660
rect 317104 221620 317110 221632
rect 345014 221620 345020 221632
rect 345072 221620 345078 221672
rect 345934 221620 345940 221672
rect 345992 221660 345998 221672
rect 373350 221660 373356 221672
rect 345992 221632 373356 221660
rect 345992 221620 345998 221632
rect 373350 221620 373356 221632
rect 373408 221620 373414 221672
rect 377674 221620 377680 221672
rect 377732 221660 377738 221672
rect 490282 221660 490288 221672
rect 377732 221632 490288 221660
rect 377732 221620 377738 221632
rect 490282 221620 490288 221632
rect 490340 221620 490346 221672
rect 534902 221620 534908 221672
rect 534960 221660 534966 221672
rect 629478 221660 629484 221672
rect 534960 221632 629484 221660
rect 534960 221620 534966 221632
rect 629478 221620 629484 221632
rect 629536 221620 629542 221672
rect 182082 221552 182088 221604
rect 182140 221592 182146 221604
rect 182140 221564 235948 221592
rect 182140 221552 182146 221564
rect 188982 221484 188988 221536
rect 189040 221524 189046 221536
rect 189040 221496 219756 221524
rect 189040 221484 189046 221496
rect 159542 221416 159548 221468
rect 159600 221456 159606 221468
rect 209682 221456 209688 221468
rect 159600 221428 209688 221456
rect 159600 221416 159606 221428
rect 209682 221416 209688 221428
rect 209740 221416 209746 221468
rect 178862 221348 178868 221400
rect 178920 221388 178926 221400
rect 181898 221388 181904 221400
rect 178920 221360 181904 221388
rect 178920 221348 178926 221360
rect 181898 221348 181904 221360
rect 181956 221348 181962 221400
rect 181990 221348 181996 221400
rect 182048 221388 182054 221400
rect 215202 221388 215208 221400
rect 182048 221360 215208 221388
rect 182048 221348 182054 221360
rect 215202 221348 215208 221360
rect 215260 221348 215266 221400
rect 219728 221388 219756 221496
rect 219986 221484 219992 221536
rect 220044 221524 220050 221536
rect 235810 221524 235816 221536
rect 220044 221496 235816 221524
rect 220044 221484 220050 221496
rect 235810 221484 235816 221496
rect 235868 221484 235874 221536
rect 235920 221524 235948 221564
rect 258810 221552 258816 221604
rect 258868 221592 258874 221604
rect 279234 221592 279240 221604
rect 258868 221564 279240 221592
rect 258868 221552 258874 221564
rect 279234 221552 279240 221564
rect 279292 221552 279298 221604
rect 283926 221552 283932 221604
rect 283984 221592 283990 221604
rect 289538 221592 289544 221604
rect 283984 221564 289544 221592
rect 283984 221552 283990 221564
rect 289538 221552 289544 221564
rect 289596 221552 289602 221604
rect 318426 221552 318432 221604
rect 318484 221592 318490 221604
rect 348142 221592 348148 221604
rect 318484 221564 348148 221592
rect 318484 221552 318490 221564
rect 348142 221552 348148 221564
rect 348200 221552 348206 221604
rect 379054 221552 379060 221604
rect 379112 221592 379118 221604
rect 494054 221592 494060 221604
rect 379112 221564 494060 221592
rect 379112 221552 379118 221564
rect 494054 221552 494060 221564
rect 494112 221552 494118 221604
rect 530118 221552 530124 221604
rect 530176 221592 530182 221604
rect 628466 221592 628472 221604
rect 530176 221564 628472 221592
rect 530176 221552 530182 221564
rect 628466 221552 628472 221564
rect 628524 221552 628530 221604
rect 247494 221524 247500 221536
rect 235920 221496 247500 221524
rect 247494 221484 247500 221496
rect 247552 221484 247558 221536
rect 273898 221484 273904 221536
rect 273956 221524 273962 221536
rect 285306 221524 285312 221536
rect 273956 221496 285312 221524
rect 273956 221484 273962 221496
rect 285306 221484 285312 221496
rect 285364 221484 285370 221536
rect 286502 221484 286508 221536
rect 286560 221524 286566 221536
rect 291746 221524 291752 221536
rect 286560 221496 291752 221524
rect 286560 221484 286566 221496
rect 291746 221484 291752 221496
rect 291804 221484 291810 221536
rect 314562 221484 314568 221536
rect 314620 221524 314626 221536
rect 339678 221524 339684 221536
rect 314620 221496 339684 221524
rect 314620 221484 314626 221496
rect 339678 221484 339684 221496
rect 339736 221484 339742 221536
rect 345106 221484 345112 221536
rect 345164 221524 345170 221536
rect 366634 221524 366640 221536
rect 345164 221496 366640 221524
rect 345164 221484 345170 221496
rect 366634 221484 366640 221496
rect 366692 221484 366698 221536
rect 375098 221484 375104 221536
rect 375156 221524 375162 221536
rect 483566 221524 483572 221536
rect 375156 221496 483572 221524
rect 375156 221484 375162 221496
rect 483566 221484 483572 221496
rect 483624 221484 483630 221536
rect 510614 221484 510620 221536
rect 510672 221524 510678 221536
rect 610342 221524 610348 221536
rect 510672 221496 610348 221524
rect 510672 221484 510678 221496
rect 610342 221484 610348 221496
rect 610400 221484 610406 221536
rect 219894 221416 219900 221468
rect 219952 221456 219958 221468
rect 245838 221456 245844 221468
rect 219952 221428 245844 221456
rect 219952 221416 219958 221428
rect 245838 221416 245844 221428
rect 245896 221416 245902 221468
rect 249518 221416 249524 221468
rect 249576 221456 249582 221468
rect 257706 221456 257712 221468
rect 249576 221428 257712 221456
rect 249576 221416 249582 221428
rect 257706 221416 257712 221428
rect 257764 221416 257770 221468
rect 268838 221416 268844 221468
rect 268896 221456 268902 221468
rect 283558 221456 283564 221468
rect 268896 221428 283564 221456
rect 268896 221416 268902 221428
rect 283558 221416 283564 221428
rect 283616 221416 283622 221468
rect 288250 221416 288256 221468
rect 288308 221456 288314 221468
rect 292758 221456 292764 221468
rect 288308 221428 292764 221456
rect 288308 221416 288314 221428
rect 292758 221416 292764 221428
rect 292816 221416 292822 221468
rect 315206 221416 315212 221468
rect 315264 221456 315270 221468
rect 343910 221456 343916 221468
rect 315264 221428 343916 221456
rect 315264 221416 315270 221428
rect 343910 221416 343916 221428
rect 343968 221416 343974 221468
rect 344002 221416 344008 221468
rect 344060 221456 344066 221468
rect 359918 221456 359924 221468
rect 344060 221428 359924 221456
rect 344060 221416 344066 221428
rect 359918 221416 359924 221428
rect 359976 221416 359982 221468
rect 372982 221416 372988 221468
rect 373040 221456 373046 221468
rect 477770 221456 477776 221468
rect 373040 221428 477776 221456
rect 373040 221416 373046 221428
rect 477770 221416 477776 221428
rect 477828 221416 477834 221468
rect 525058 221416 525064 221468
rect 525116 221456 525122 221468
rect 627546 221456 627552 221468
rect 525116 221428 627552 221456
rect 525116 221416 525122 221428
rect 627546 221416 627552 221428
rect 627604 221416 627610 221468
rect 250070 221388 250076 221400
rect 219728 221360 250076 221388
rect 250070 221348 250076 221360
rect 250128 221348 250134 221400
rect 251082 221348 251088 221400
rect 251140 221388 251146 221400
rect 256602 221388 256608 221400
rect 251140 221360 256608 221388
rect 251140 221348 251146 221360
rect 256602 221348 256608 221360
rect 256660 221348 256666 221400
rect 267182 221348 267188 221400
rect 267240 221388 267246 221400
rect 282454 221388 282460 221400
rect 267240 221360 282460 221388
rect 267240 221348 267246 221360
rect 282454 221348 282460 221360
rect 282512 221348 282518 221400
rect 289078 221348 289084 221400
rect 289136 221388 289142 221400
rect 292114 221388 292120 221400
rect 289136 221360 292120 221388
rect 289136 221348 289142 221360
rect 292114 221348 292120 221360
rect 292172 221348 292178 221400
rect 292390 221348 292396 221400
rect 292448 221388 292454 221400
rect 293494 221388 293500 221400
rect 292448 221360 293500 221388
rect 292448 221348 292454 221360
rect 293494 221348 293500 221360
rect 293552 221348 293558 221400
rect 313826 221348 313832 221400
rect 313884 221388 313890 221400
rect 340598 221388 340604 221400
rect 313884 221360 340604 221388
rect 313884 221348 313890 221360
rect 340598 221348 340604 221360
rect 340656 221348 340662 221400
rect 340690 221348 340696 221400
rect 340748 221388 340754 221400
rect 356514 221388 356520 221400
rect 340748 221360 356520 221388
rect 340748 221348 340754 221360
rect 356514 221348 356520 221360
rect 356572 221348 356578 221400
rect 367278 221348 367284 221400
rect 367336 221388 367342 221400
rect 464246 221388 464252 221400
rect 367336 221360 464252 221388
rect 367336 221348 367342 221360
rect 464246 221348 464252 221360
rect 464304 221348 464310 221400
rect 505738 221348 505744 221400
rect 505796 221388 505802 221400
rect 609422 221388 609428 221400
rect 505796 221360 609428 221388
rect 505796 221348 505802 221360
rect 609422 221348 609428 221360
rect 609480 221348 609486 221400
rect 149422 221280 149428 221332
rect 149480 221320 149486 221332
rect 190270 221320 190276 221332
rect 149480 221292 190276 221320
rect 149480 221280 149486 221292
rect 190270 221280 190276 221292
rect 190328 221280 190334 221332
rect 199930 221280 199936 221332
rect 199988 221320 199994 221332
rect 231854 221320 231860 221332
rect 199988 221292 231860 221320
rect 199988 221280 199994 221292
rect 231854 221280 231860 221292
rect 231912 221280 231918 221332
rect 236914 221280 236920 221332
rect 236972 221320 236978 221332
rect 240318 221320 240324 221332
rect 236972 221292 240324 221320
rect 236972 221280 236978 221292
rect 240318 221280 240324 221292
rect 240376 221280 240382 221332
rect 247862 221280 247868 221332
rect 247920 221320 247926 221332
rect 255222 221320 255228 221332
rect 247920 221292 255228 221320
rect 247920 221280 247926 221292
rect 255222 221280 255228 221292
rect 255280 221280 255286 221332
rect 256234 221280 256240 221332
rect 256292 221320 256298 221332
rect 259638 221320 259644 221332
rect 256292 221292 259644 221320
rect 256292 221280 256298 221292
rect 259638 221280 259644 221292
rect 259696 221280 259702 221332
rect 280614 221280 280620 221332
rect 280672 221320 280678 221332
rect 288158 221320 288164 221332
rect 280672 221292 288164 221320
rect 280672 221280 280678 221292
rect 288158 221280 288164 221292
rect 288216 221280 288222 221332
rect 289722 221280 289728 221332
rect 289780 221320 289786 221332
rect 293126 221320 293132 221332
rect 289780 221292 293132 221320
rect 289780 221280 289786 221292
rect 293126 221280 293132 221292
rect 293184 221280 293190 221332
rect 294966 221280 294972 221332
rect 295024 221320 295030 221332
rect 295610 221320 295616 221332
rect 295024 221292 295616 221320
rect 295024 221280 295030 221292
rect 295610 221280 295616 221292
rect 295668 221280 295674 221332
rect 315574 221280 315580 221332
rect 315632 221320 315638 221332
rect 341426 221320 341432 221332
rect 315632 221292 341432 221320
rect 315632 221280 315638 221292
rect 341426 221280 341432 221292
rect 341484 221280 341490 221332
rect 341518 221280 341524 221332
rect 341576 221320 341582 221332
rect 353294 221320 353300 221332
rect 341576 221292 353300 221320
rect 341576 221280 341582 221292
rect 353294 221280 353300 221292
rect 353352 221280 353358 221332
rect 365990 221280 365996 221332
rect 366048 221320 366054 221332
rect 454126 221320 454132 221332
rect 366048 221292 454132 221320
rect 366048 221280 366054 221292
rect 454126 221280 454132 221292
rect 454184 221280 454190 221332
rect 501046 221280 501052 221332
rect 501104 221320 501110 221332
rect 608502 221320 608508 221332
rect 501104 221292 608508 221320
rect 501104 221280 501110 221292
rect 608502 221280 608508 221292
rect 608560 221280 608566 221332
rect 179690 221212 179696 221264
rect 179748 221252 179754 221264
rect 214282 221252 214288 221264
rect 179748 221224 214288 221252
rect 179748 221212 179754 221224
rect 214282 221212 214288 221224
rect 214340 221212 214346 221264
rect 226794 221212 226800 221264
rect 226852 221252 226858 221264
rect 239858 221252 239864 221264
rect 226852 221224 239864 221252
rect 226852 221212 226858 221224
rect 239858 221212 239864 221224
rect 239916 221212 239922 221264
rect 252922 221212 252928 221264
rect 252980 221252 252986 221264
rect 258258 221252 258264 221264
rect 252980 221224 258264 221252
rect 252980 221212 252986 221224
rect 258258 221212 258264 221224
rect 258316 221212 258322 221264
rect 270402 221212 270408 221264
rect 270460 221252 270466 221264
rect 283834 221252 283840 221264
rect 270460 221224 283840 221252
rect 270460 221212 270466 221224
rect 283834 221212 283840 221224
rect 283892 221212 283898 221264
rect 284846 221212 284852 221264
rect 284904 221252 284910 221264
rect 291378 221252 291384 221264
rect 284904 221224 291384 221252
rect 284904 221212 284910 221224
rect 291378 221212 291384 221224
rect 291436 221212 291442 221264
rect 291562 221212 291568 221264
rect 291620 221252 291626 221264
rect 294230 221252 294236 221264
rect 291620 221224 294236 221252
rect 291620 221212 291626 221224
rect 294230 221212 294236 221224
rect 294288 221212 294294 221264
rect 312354 221212 312360 221264
rect 312412 221252 312418 221264
rect 337194 221252 337200 221264
rect 312412 221224 337200 221252
rect 312412 221212 312418 221224
rect 337194 221212 337200 221224
rect 337252 221212 337258 221264
rect 337654 221212 337660 221264
rect 337712 221252 337718 221264
rect 346486 221252 346492 221264
rect 337712 221224 346492 221252
rect 337712 221212 337718 221224
rect 346486 221212 346492 221224
rect 346544 221212 346550 221264
rect 389910 221212 389916 221264
rect 389968 221252 389974 221264
rect 392670 221252 392676 221264
rect 389968 221224 392676 221252
rect 389968 221212 389974 221224
rect 392670 221212 392676 221224
rect 392728 221212 392734 221264
rect 397546 221212 397552 221264
rect 397604 221252 397610 221264
rect 476850 221252 476856 221264
rect 397604 221224 476856 221252
rect 397604 221212 397610 221224
rect 476850 221212 476856 221224
rect 476908 221212 476914 221264
rect 518986 221212 518992 221264
rect 519044 221252 519050 221264
rect 519998 221252 520004 221264
rect 519044 221224 520004 221252
rect 519044 221212 519050 221224
rect 519998 221212 520004 221224
rect 520056 221252 520062 221264
rect 626626 221252 626632 221264
rect 520056 221224 626632 221252
rect 520056 221212 520062 221224
rect 626626 221212 626632 221224
rect 626684 221212 626690 221264
rect 172974 221144 172980 221196
rect 173032 221184 173038 221196
rect 181990 221184 181996 221196
rect 173032 221156 181996 221184
rect 173032 221144 173038 221156
rect 181990 221144 181996 221156
rect 182048 221144 182054 221196
rect 183094 221144 183100 221196
rect 183152 221184 183158 221196
rect 216214 221184 216220 221196
rect 183152 221156 216220 221184
rect 183152 221144 183158 221156
rect 216214 221144 216220 221156
rect 216272 221144 216278 221196
rect 246114 221144 246120 221196
rect 246172 221184 246178 221196
rect 258442 221184 258448 221196
rect 246172 221156 258448 221184
rect 246172 221144 246178 221156
rect 258442 221144 258448 221156
rect 258500 221144 258506 221196
rect 276474 221144 276480 221196
rect 276532 221184 276538 221196
rect 287422 221184 287428 221196
rect 276532 221156 287428 221184
rect 276532 221144 276538 221156
rect 287422 221144 287428 221156
rect 287480 221144 287486 221196
rect 330202 221144 330208 221196
rect 330260 221184 330266 221196
rect 330260 221156 336872 221184
rect 330260 221144 330266 221156
rect 189810 221076 189816 221128
rect 189868 221116 189874 221128
rect 220630 221116 220636 221128
rect 189868 221088 220636 221116
rect 189868 221076 189874 221088
rect 220630 221076 220636 221088
rect 220688 221076 220694 221128
rect 234706 221116 234712 221128
rect 227640 221088 234712 221116
rect 192294 221008 192300 221060
rect 192352 221048 192358 221060
rect 193030 221048 193036 221060
rect 192352 221020 193036 221048
rect 192352 221008 192358 221020
rect 193030 221008 193036 221020
rect 193088 221008 193094 221060
rect 205450 221048 205456 221060
rect 193140 221020 205456 221048
rect 192846 220940 192852 220992
rect 192904 220980 192910 220992
rect 193140 220980 193168 221020
rect 205450 221008 205456 221020
rect 205508 221008 205514 221060
rect 206646 221008 206652 221060
rect 206704 221048 206710 221060
rect 227640 221048 227668 221088
rect 234706 221076 234712 221088
rect 234764 221076 234770 221128
rect 277302 221076 277308 221128
rect 277360 221116 277366 221128
rect 286686 221116 286692 221128
rect 277360 221088 286692 221116
rect 277360 221076 277366 221088
rect 286686 221076 286692 221088
rect 286744 221076 286750 221128
rect 289262 221116 289268 221128
rect 286796 221088 289268 221116
rect 206704 221020 227668 221048
rect 206704 221008 206710 221020
rect 230198 221008 230204 221060
rect 230256 221048 230262 221060
rect 239950 221048 239956 221060
rect 230256 221020 239956 221048
rect 230256 221008 230262 221020
rect 239950 221008 239956 221020
rect 240008 221008 240014 221060
rect 265526 221008 265532 221060
rect 265584 221048 265590 221060
rect 282086 221048 282092 221060
rect 265584 221020 282092 221048
rect 265584 221008 265590 221020
rect 282086 221008 282092 221020
rect 282144 221008 282150 221060
rect 282362 221008 282368 221060
rect 282420 221048 282426 221060
rect 286796 221048 286824 221088
rect 289262 221076 289268 221088
rect 289320 221076 289326 221128
rect 313090 221076 313096 221128
rect 313148 221116 313154 221128
rect 336734 221116 336740 221128
rect 313148 221088 336740 221116
rect 313148 221076 313154 221088
rect 336734 221076 336740 221088
rect 336792 221076 336798 221128
rect 336844 221116 336872 221156
rect 339586 221144 339592 221196
rect 339644 221184 339650 221196
rect 349798 221184 349804 221196
rect 339644 221156 349804 221184
rect 339644 221144 339650 221156
rect 349798 221144 349804 221156
rect 349856 221144 349862 221196
rect 368198 221144 368204 221196
rect 368256 221184 368262 221196
rect 368256 221156 400214 221184
rect 368256 221144 368262 221156
rect 352006 221116 352012 221128
rect 336844 221088 352012 221116
rect 352006 221076 352012 221088
rect 352064 221076 352070 221128
rect 383746 221076 383752 221128
rect 383804 221116 383810 221128
rect 396074 221116 396080 221128
rect 383804 221088 396080 221116
rect 383804 221076 383810 221088
rect 396074 221076 396080 221088
rect 396132 221076 396138 221128
rect 400186 221116 400214 221156
rect 403710 221144 403716 221196
rect 403768 221184 403774 221196
rect 406194 221184 406200 221196
rect 403768 221156 406200 221184
rect 403768 221144 403774 221156
rect 406194 221144 406200 221156
rect 406252 221144 406258 221196
rect 408310 221144 408316 221196
rect 408368 221184 408374 221196
rect 437290 221184 437296 221196
rect 408368 221156 437296 221184
rect 408368 221144 408374 221156
rect 437290 221144 437296 221156
rect 437348 221144 437354 221196
rect 513374 221144 513380 221196
rect 513432 221184 513438 221196
rect 514938 221184 514944 221196
rect 513432 221156 514944 221184
rect 513432 221144 513438 221156
rect 514938 221144 514944 221156
rect 514996 221184 515002 221196
rect 625706 221184 625712 221196
rect 514996 221156 625712 221184
rect 514996 221144 515002 221156
rect 625706 221144 625712 221156
rect 625764 221144 625770 221196
rect 655790 221144 655796 221196
rect 655848 221184 655854 221196
rect 675938 221184 675944 221196
rect 655848 221156 675944 221184
rect 655848 221144 655854 221156
rect 675938 221144 675944 221156
rect 675996 221144 676002 221196
rect 407022 221116 407028 221128
rect 400186 221088 407028 221116
rect 407022 221076 407028 221088
rect 407080 221076 407086 221128
rect 407942 221076 407948 221128
rect 408000 221116 408006 221128
rect 561766 221116 561772 221128
rect 408000 221088 561772 221116
rect 408000 221076 408006 221088
rect 561766 221076 561772 221088
rect 561824 221076 561830 221128
rect 282420 221020 286824 221048
rect 282420 221008 282426 221020
rect 287330 221008 287336 221060
rect 287388 221048 287394 221060
rect 291010 221048 291016 221060
rect 287388 221020 291016 221048
rect 287388 221008 287394 221020
rect 291010 221008 291016 221020
rect 291068 221008 291074 221060
rect 386230 221008 386236 221060
rect 386288 221048 386294 221060
rect 510614 221048 510620 221060
rect 386288 221020 510620 221048
rect 386288 221008 386294 221020
rect 510614 221008 510620 221020
rect 510672 221008 510678 221060
rect 549346 221008 549352 221060
rect 549404 221048 549410 221060
rect 551094 221048 551100 221060
rect 549404 221020 551100 221048
rect 549404 221008 549410 221020
rect 551094 221008 551100 221020
rect 551152 221048 551158 221060
rect 617794 221048 617800 221060
rect 551152 221020 617800 221048
rect 551152 221008 551158 221020
rect 617794 221008 617800 221020
rect 617852 221008 617858 221060
rect 655606 221008 655612 221060
rect 655664 221048 655670 221060
rect 676030 221048 676036 221060
rect 655664 221020 676036 221048
rect 655664 221008 655670 221020
rect 676030 221008 676036 221020
rect 676088 221008 676094 221060
rect 192904 220952 193168 220980
rect 192904 220940 192910 220952
rect 197262 220940 197268 220992
rect 197320 220980 197326 220992
rect 209038 220980 209044 220992
rect 197320 220952 209044 220980
rect 197320 220940 197326 220952
rect 209038 220940 209044 220952
rect 209096 220940 209102 220992
rect 213362 220940 213368 220992
rect 213420 220980 213426 220992
rect 234798 220980 234804 220992
rect 213420 220952 234804 220980
rect 213420 220940 213426 220952
rect 234798 220940 234804 220952
rect 234856 220940 234862 220992
rect 268010 220940 268016 220992
rect 268068 220980 268074 220992
rect 284202 220980 284208 220992
rect 268068 220952 284208 220980
rect 268068 220940 268074 220952
rect 284202 220940 284208 220952
rect 284260 220940 284266 220992
rect 285674 220940 285680 220992
rect 285732 220980 285738 220992
rect 290642 220980 290648 220992
rect 285732 220952 290648 220980
rect 285732 220940 285738 220952
rect 290642 220940 290648 220952
rect 290700 220940 290706 220992
rect 385494 220940 385500 220992
rect 385552 220980 385558 220992
rect 508774 220980 508780 220992
rect 385552 220952 508780 220980
rect 385552 220940 385558 220952
rect 508774 220940 508780 220952
rect 508832 220940 508838 220992
rect 509602 220940 509608 220992
rect 509660 220980 509666 220992
rect 624786 220980 624792 220992
rect 509660 220952 624792 220980
rect 509660 220940 509666 220952
rect 624786 220940 624792 220952
rect 624844 220940 624850 220992
rect 279786 220872 279792 220924
rect 279844 220912 279850 220924
rect 288894 220912 288900 220924
rect 279844 220884 288900 220912
rect 279844 220872 279850 220884
rect 288894 220872 288900 220884
rect 288952 220872 288958 220924
rect 393774 220872 393780 220924
rect 393832 220912 393838 220924
rect 399478 220912 399484 220924
rect 393832 220884 399484 220912
rect 393832 220872 393838 220884
rect 399478 220872 399484 220884
rect 399536 220872 399542 220924
rect 504818 220872 504824 220924
rect 504876 220912 504882 220924
rect 623866 220912 623872 220924
rect 504876 220884 623872 220912
rect 504876 220872 504882 220884
rect 623866 220872 623872 220884
rect 623924 220872 623930 220924
rect 196526 220804 196532 220856
rect 196584 220844 196590 220856
rect 204254 220844 204260 220856
rect 196584 220816 204260 220844
rect 196584 220804 196590 220816
rect 204254 220804 204260 220816
rect 204312 220804 204318 220856
rect 204898 220804 204904 220856
rect 204956 220844 204962 220856
rect 206830 220844 206836 220856
rect 204956 220816 206836 220844
rect 204956 220804 204962 220816
rect 206830 220804 206836 220816
rect 206888 220804 206894 220856
rect 233510 220804 233516 220856
rect 233568 220844 233574 220856
rect 238478 220844 238484 220856
rect 233568 220816 238484 220844
rect 233568 220804 233574 220816
rect 238478 220804 238484 220816
rect 238536 220804 238542 220856
rect 499298 220804 499304 220856
rect 499356 220844 499362 220856
rect 622946 220844 622952 220856
rect 499356 220816 622952 220844
rect 499356 220804 499362 220816
rect 622946 220804 622952 220816
rect 623004 220804 623010 220856
rect 655514 220804 655520 220856
rect 655572 220844 655578 220856
rect 675846 220844 675852 220856
rect 655572 220816 675852 220844
rect 655572 220804 655578 220816
rect 675846 220804 675852 220816
rect 675904 220804 675910 220856
rect 350534 220736 350540 220788
rect 350592 220776 350598 220788
rect 426342 220776 426348 220788
rect 350592 220748 426348 220776
rect 350592 220736 350598 220748
rect 426342 220736 426348 220748
rect 426400 220736 426406 220788
rect 675202 220736 675208 220788
rect 675260 220776 675266 220788
rect 676030 220776 676036 220788
rect 675260 220748 676036 220776
rect 675260 220736 675266 220748
rect 676030 220736 676036 220748
rect 676088 220736 676094 220788
rect 352098 220668 352104 220720
rect 352156 220708 352162 220720
rect 429746 220708 429752 220720
rect 352156 220680 429752 220708
rect 352156 220668 352162 220680
rect 429746 220668 429752 220680
rect 429804 220668 429810 220720
rect 353386 220600 353392 220652
rect 353444 220640 353450 220652
rect 433334 220640 433340 220652
rect 353444 220612 433340 220640
rect 353444 220600 353450 220612
rect 433334 220600 433340 220612
rect 433392 220600 433398 220652
rect 355042 220532 355048 220584
rect 355100 220572 355106 220584
rect 436462 220572 436468 220584
rect 355100 220544 436468 220572
rect 355100 220532 355106 220544
rect 436462 220532 436468 220544
rect 436520 220532 436526 220584
rect 356238 220464 356244 220516
rect 356296 220504 356302 220516
rect 439774 220504 439780 220516
rect 356296 220476 439780 220504
rect 356296 220464 356302 220476
rect 439774 220464 439780 220476
rect 439832 220464 439838 220516
rect 359366 220396 359372 220448
rect 359424 220436 359430 220448
rect 446582 220436 446588 220448
rect 359424 220408 446588 220436
rect 359424 220396 359430 220408
rect 446582 220396 446588 220408
rect 446640 220396 446646 220448
rect 357710 220328 357716 220380
rect 357768 220368 357774 220380
rect 443178 220368 443184 220380
rect 357768 220340 443184 220368
rect 357768 220328 357774 220340
rect 443178 220328 443184 220340
rect 443236 220328 443242 220380
rect 361942 220260 361948 220312
rect 362000 220300 362006 220312
rect 453298 220300 453304 220312
rect 362000 220272 453304 220300
rect 362000 220260 362006 220272
rect 453298 220260 453304 220272
rect 453356 220260 453362 220312
rect 142706 220192 142712 220244
rect 142764 220232 142770 220244
rect 229646 220232 229652 220244
rect 142764 220204 229652 220232
rect 142764 220192 142770 220204
rect 229646 220192 229652 220204
rect 229704 220192 229710 220244
rect 360562 220192 360568 220244
rect 360620 220232 360626 220244
rect 449894 220232 449900 220244
rect 360620 220204 449900 220232
rect 360620 220192 360626 220204
rect 449894 220192 449900 220204
rect 449952 220192 449958 220244
rect 139302 220124 139308 220176
rect 139360 220164 139366 220176
rect 228266 220164 228272 220176
rect 139360 220136 228272 220164
rect 139360 220124 139366 220136
rect 228266 220124 228272 220136
rect 228324 220124 228330 220176
rect 364794 220124 364800 220176
rect 364852 220164 364858 220176
rect 460014 220164 460020 220176
rect 364852 220136 460020 220164
rect 364852 220124 364858 220136
rect 460014 220124 460020 220136
rect 460072 220124 460078 220176
rect 135990 220056 135996 220108
rect 136048 220096 136054 220108
rect 226610 220096 226616 220108
rect 136048 220068 226616 220096
rect 136048 220056 136054 220068
rect 226610 220056 226616 220068
rect 226668 220056 226674 220108
rect 363414 220056 363420 220108
rect 363472 220096 363478 220108
rect 456610 220096 456616 220108
rect 363472 220068 456616 220096
rect 363472 220056 363478 220068
rect 456610 220056 456616 220068
rect 456668 220056 456674 220108
rect 132402 219988 132408 220040
rect 132460 220028 132466 220040
rect 225414 220028 225420 220040
rect 132460 220000 225420 220028
rect 132460 219988 132466 220000
rect 225414 219988 225420 220000
rect 225472 219988 225478 220040
rect 368382 219988 368388 220040
rect 368440 220028 368446 220040
rect 465902 220028 465908 220040
rect 368440 220000 465908 220028
rect 368440 219988 368446 220000
rect 465902 219988 465908 220000
rect 465960 219988 465966 220040
rect 129274 219920 129280 219972
rect 129332 219960 129338 219972
rect 223758 219960 223764 219972
rect 129332 219932 223764 219960
rect 129332 219920 129338 219932
rect 223758 219920 223764 219932
rect 223816 219920 223822 219972
rect 367646 219920 367652 219972
rect 367704 219960 367710 219972
rect 466730 219960 466736 219972
rect 367704 219932 466736 219960
rect 367704 219920 367710 219932
rect 466730 219920 466736 219932
rect 466788 219920 466794 219972
rect 125870 219852 125876 219904
rect 125928 219892 125934 219904
rect 222286 219892 222292 219904
rect 125928 219864 222292 219892
rect 125928 219852 125934 219864
rect 222286 219852 222292 219864
rect 222344 219852 222350 219904
rect 366266 219852 366272 219904
rect 366324 219892 366330 219904
rect 463694 219892 463700 219904
rect 366324 219864 463700 219892
rect 366324 219852 366330 219864
rect 463694 219852 463700 219864
rect 463752 219852 463758 219904
rect 122466 219784 122472 219836
rect 122524 219824 122530 219836
rect 221090 219824 221096 219836
rect 122524 219796 221096 219824
rect 122524 219784 122530 219796
rect 221090 219784 221096 219796
rect 221148 219784 221154 219836
rect 370498 219784 370504 219836
rect 370556 219824 370562 219836
rect 473446 219824 473452 219836
rect 370556 219796 473452 219824
rect 370556 219784 370562 219796
rect 473446 219784 473452 219796
rect 473504 219784 473510 219836
rect 58618 219716 58624 219768
rect 58676 219756 58682 219768
rect 193766 219756 193772 219768
rect 58676 219728 193772 219756
rect 58676 219716 58682 219728
rect 193766 219716 193772 219728
rect 193824 219716 193830 219768
rect 369302 219716 369308 219768
rect 369360 219756 369366 219768
rect 470134 219756 470140 219768
rect 369360 219728 470140 219756
rect 369360 219716 369366 219728
rect 470134 219716 470140 219728
rect 470192 219716 470198 219768
rect 45462 219648 45468 219700
rect 45520 219688 45526 219700
rect 648522 219688 648528 219700
rect 45520 219660 648528 219688
rect 45520 219648 45526 219660
rect 648522 219648 648528 219660
rect 648580 219648 648586 219700
rect 45554 219580 45560 219632
rect 45612 219620 45618 219632
rect 649902 219620 649908 219632
rect 45612 219592 649908 219620
rect 45612 219580 45618 219592
rect 649902 219580 649908 219592
rect 649960 219580 649966 219632
rect 45738 219512 45744 219564
rect 45796 219552 45802 219564
rect 651282 219552 651288 219564
rect 45796 219524 651288 219552
rect 45796 219512 45802 219524
rect 651282 219512 651288 219524
rect 651340 219512 651346 219564
rect 45830 219444 45836 219496
rect 45888 219484 45894 219496
rect 652754 219484 652760 219496
rect 45888 219456 652760 219484
rect 45888 219444 45894 219456
rect 652754 219444 652760 219456
rect 652812 219444 652818 219496
rect 45922 219376 45928 219428
rect 45980 219416 45986 219428
rect 654134 219416 654140 219428
rect 45980 219388 654140 219416
rect 45980 219376 45986 219388
rect 654134 219376 654140 219388
rect 654192 219376 654198 219428
rect 347682 219308 347688 219360
rect 347740 219348 347746 219360
rect 419718 219348 419724 219360
rect 347740 219320 419724 219348
rect 347740 219308 347746 219320
rect 419718 219308 419724 219320
rect 419776 219308 419782 219360
rect 349154 219240 349160 219292
rect 349212 219280 349218 219292
rect 423030 219280 423036 219292
rect 349212 219252 423036 219280
rect 349212 219240 349218 219252
rect 423030 219240 423036 219252
rect 423088 219240 423094 219292
rect 346302 219172 346308 219224
rect 346360 219212 346366 219224
rect 416222 219212 416228 219224
rect 346360 219184 416228 219212
rect 346360 219172 346366 219184
rect 416222 219172 416228 219184
rect 416280 219172 416286 219224
rect 344830 219104 344836 219156
rect 344888 219144 344894 219156
rect 412910 219144 412916 219156
rect 344888 219116 412916 219144
rect 344888 219104 344894 219116
rect 412910 219104 412916 219116
rect 412968 219104 412974 219156
rect 343450 219036 343456 219088
rect 343508 219076 343514 219088
rect 409506 219076 409512 219088
rect 343508 219048 409512 219076
rect 343508 219036 343514 219048
rect 409506 219036 409512 219048
rect 409564 219036 409570 219088
rect 666554 218560 666560 218612
rect 666612 218600 666618 218612
rect 666830 218600 666836 218612
rect 666612 218572 666836 218600
rect 666612 218560 666618 218572
rect 666830 218560 666836 218572
rect 666888 218560 666894 218612
rect 525794 218424 525800 218476
rect 525852 218464 525858 218476
rect 613102 218464 613108 218476
rect 525852 218436 613108 218464
rect 525852 218424 525858 218436
rect 613102 218424 613108 218436
rect 613160 218424 613166 218476
rect 523402 218356 523408 218408
rect 523460 218396 523466 218408
rect 612642 218396 612648 218408
rect 523460 218368 612648 218396
rect 523460 218356 523466 218368
rect 612642 218356 612648 218368
rect 612700 218356 612706 218408
rect 520826 218288 520832 218340
rect 520884 218328 520890 218340
rect 612182 218328 612188 218340
rect 520884 218300 612188 218328
rect 520884 218288 520890 218300
rect 612182 218288 612188 218300
rect 612240 218288 612246 218340
rect 674558 218288 674564 218340
rect 674616 218328 674622 218340
rect 676030 218328 676036 218340
rect 674616 218300 676036 218328
rect 674616 218288 674622 218300
rect 676030 218288 676036 218300
rect 676088 218288 676094 218340
rect 518618 218220 518624 218272
rect 518676 218260 518682 218272
rect 611722 218260 611728 218272
rect 518676 218232 611728 218260
rect 518676 218220 518682 218232
rect 611722 218220 611728 218232
rect 611780 218220 611786 218272
rect 515490 218152 515496 218204
rect 515548 218192 515554 218204
rect 611262 218192 611268 218204
rect 515548 218164 611268 218192
rect 515548 218152 515554 218164
rect 611262 218152 611268 218164
rect 611320 218152 611326 218204
rect 490282 218084 490288 218136
rect 490340 218124 490346 218136
rect 607122 218124 607128 218136
rect 490340 218096 607128 218124
rect 490340 218084 490346 218096
rect 607122 218084 607128 218096
rect 607180 218084 607186 218136
rect 487154 218016 487160 218068
rect 487212 218056 487218 218068
rect 606662 218056 606668 218068
rect 487212 218028 606668 218056
rect 487212 218016 487218 218028
rect 606662 218016 606668 218028
rect 606720 218016 606726 218068
rect 674834 218016 674840 218068
rect 674892 218056 674898 218068
rect 676030 218056 676036 218068
rect 674892 218028 676036 218056
rect 674892 218016 674898 218028
rect 676030 218016 676036 218028
rect 676088 218016 676094 218068
rect 418154 217948 418160 218000
rect 418212 217988 418218 218000
rect 418614 217988 418620 218000
rect 418212 217960 418620 217988
rect 418212 217948 418218 217960
rect 418614 217948 418620 217960
rect 418672 217948 418678 218000
rect 213868 217608 213874 217660
rect 213926 217648 213932 217660
rect 219894 217648 219900 217660
rect 213926 217620 219900 217648
rect 213926 217608 213932 217620
rect 219894 217608 219900 217620
rect 219952 217608 219958 217660
rect 492260 217540 492266 217592
rect 492318 217580 492324 217592
rect 622026 217580 622032 217592
rect 492318 217552 622032 217580
rect 492318 217540 492324 217552
rect 622026 217540 622032 217552
rect 622084 217540 622090 217592
rect 24946 217472 24952 217524
rect 25004 217512 25010 217524
rect 665726 217512 665732 217524
rect 25004 217484 665732 217512
rect 25004 217472 25010 217484
rect 665726 217472 665732 217484
rect 665784 217472 665790 217524
rect 570874 217404 570880 217456
rect 570932 217444 570938 217456
rect 635918 217444 635924 217456
rect 570932 217416 635924 217444
rect 570932 217404 570938 217416
rect 635918 217404 635924 217416
rect 635976 217404 635982 217456
rect 568298 217336 568304 217388
rect 568356 217376 568362 217388
rect 635458 217376 635464 217388
rect 568356 217348 635464 217376
rect 568356 217336 568362 217348
rect 635458 217336 635464 217348
rect 635516 217336 635522 217388
rect 565630 217268 565636 217320
rect 565688 217308 565694 217320
rect 634998 217308 635004 217320
rect 565688 217280 635004 217308
rect 565688 217268 565694 217280
rect 634998 217268 635004 217280
rect 635056 217268 635062 217320
rect 560754 217200 560760 217252
rect 560812 217240 560818 217252
rect 634078 217240 634084 217252
rect 560812 217212 634084 217240
rect 560812 217200 560818 217212
rect 634078 217200 634084 217212
rect 634136 217200 634142 217252
rect 555694 217132 555700 217184
rect 555752 217172 555758 217184
rect 633158 217172 633164 217184
rect 555752 217144 633164 217172
rect 555752 217132 555758 217144
rect 633158 217132 633164 217144
rect 633216 217132 633222 217184
rect 508590 217064 508596 217116
rect 508648 217104 508654 217116
rect 533062 217104 533068 217116
rect 508648 217076 533068 217104
rect 508648 217064 508654 217076
rect 533062 217064 533068 217076
rect 533120 217064 533126 217116
rect 550450 217064 550456 217116
rect 550508 217104 550514 217116
rect 632238 217104 632244 217116
rect 550508 217076 632244 217104
rect 550508 217064 550514 217076
rect 632238 217064 632244 217076
rect 632296 217064 632302 217116
rect 418522 216996 418528 217048
rect 418580 217036 418586 217048
rect 639690 217036 639696 217048
rect 418580 217008 639696 217036
rect 418580 216996 418586 217008
rect 639690 216996 639696 217008
rect 639748 216996 639754 217048
rect 418614 216928 418620 216980
rect 418672 216968 418678 216980
rect 640150 216968 640156 216980
rect 418672 216940 640156 216968
rect 418672 216928 418678 216940
rect 640150 216928 640156 216940
rect 640208 216928 640214 216980
rect 418430 216860 418436 216912
rect 418488 216900 418494 216912
rect 640610 216900 640616 216912
rect 418488 216872 640616 216900
rect 418488 216860 418494 216872
rect 640610 216860 640616 216872
rect 640668 216860 640674 216912
rect 52178 216792 52184 216844
rect 52236 216832 52242 216844
rect 57974 216832 57980 216844
rect 52236 216804 57980 216832
rect 52236 216792 52242 216804
rect 57974 216792 57980 216804
rect 58032 216792 58038 216844
rect 417878 216792 417884 216844
rect 417936 216832 417942 216844
rect 641070 216832 641076 216844
rect 417936 216804 641076 216832
rect 417936 216792 417942 216804
rect 641070 216792 641076 216804
rect 641128 216792 641134 216844
rect 52270 216724 52276 216776
rect 52328 216764 52334 216776
rect 169662 216764 169668 216776
rect 52328 216736 169668 216764
rect 52328 216724 52334 216736
rect 169662 216724 169668 216736
rect 169720 216724 169726 216776
rect 187602 216724 187608 216776
rect 187660 216764 187666 216776
rect 603442 216764 603448 216776
rect 187660 216736 603448 216764
rect 187660 216724 187666 216736
rect 603442 216724 603448 216736
rect 603500 216724 603506 216776
rect 46290 216656 46296 216708
rect 46348 216696 46354 216708
rect 664806 216696 664812 216708
rect 46348 216668 664812 216696
rect 46348 216656 46354 216668
rect 664806 216656 664812 216668
rect 664864 216656 664870 216708
rect 673822 216656 673828 216708
rect 673880 216696 673886 216708
rect 676030 216696 676036 216708
rect 673880 216668 676036 216696
rect 673880 216656 673886 216668
rect 676030 216656 676036 216668
rect 676088 216656 676094 216708
rect 45646 216588 45652 216640
rect 45704 216628 45710 216640
rect 664346 216628 664352 216640
rect 45704 216600 664352 216628
rect 45704 216588 45710 216600
rect 664346 216588 664352 216600
rect 664404 216588 664410 216640
rect 503530 216520 503536 216572
rect 503588 216560 503594 216572
rect 524046 216560 524052 216572
rect 503588 216532 524052 216560
rect 503588 216520 503594 216532
rect 524046 216520 524052 216532
rect 524104 216520 524110 216572
rect 532970 216520 532976 216572
rect 533028 216560 533034 216572
rect 533028 216532 537340 216560
rect 533028 216520 533034 216532
rect 502702 216452 502708 216504
rect 502760 216492 502766 216504
rect 502760 216464 512684 216492
rect 502760 216452 502766 216464
rect 486694 216384 486700 216436
rect 486752 216384 486758 216436
rect 490098 216384 490104 216436
rect 490156 216384 490162 216436
rect 493226 216384 493232 216436
rect 493284 216424 493290 216436
rect 493284 216396 496814 216424
rect 493284 216384 493290 216396
rect 486712 215540 486740 216384
rect 490116 215608 490144 216384
rect 496786 215676 496814 216396
rect 507762 216384 507768 216436
rect 507820 216384 507826 216436
rect 507780 215812 507808 216384
rect 512656 215880 512684 216464
rect 517624 216464 536788 216492
rect 512822 216384 512828 216436
rect 512880 216384 512886 216436
rect 513650 216384 513656 216436
rect 513708 216424 513714 216436
rect 517624 216424 517652 216464
rect 513708 216396 517652 216424
rect 513708 216384 513714 216396
rect 517882 216384 517888 216436
rect 517940 216424 517946 216436
rect 517940 216396 520688 216424
rect 517940 216384 517946 216396
rect 512840 216356 512868 216384
rect 512840 216328 517284 216356
rect 517256 215948 517284 216328
rect 520660 216016 520688 216396
rect 522850 216384 522856 216436
rect 522908 216424 522914 216436
rect 522908 216396 524000 216424
rect 522908 216384 522914 216396
rect 523972 216084 524000 216396
rect 524046 216384 524052 216436
rect 524104 216384 524110 216436
rect 527910 216384 527916 216436
rect 527968 216424 527974 216436
rect 527968 216396 530072 216424
rect 527968 216384 527974 216396
rect 524064 216152 524092 216384
rect 530044 216220 530072 216396
rect 533062 216384 533068 216436
rect 533120 216384 533126 216436
rect 533080 216288 533108 216384
rect 536760 216356 536788 216464
rect 537312 216424 537340 216532
rect 545574 216520 545580 216572
rect 545632 216560 545638 216572
rect 631318 216560 631324 216572
rect 545632 216532 631324 216560
rect 545632 216520 545638 216532
rect 631318 216520 631324 216532
rect 631376 216520 631382 216572
rect 538030 216452 538036 216504
rect 538088 216492 538094 216504
rect 629938 216492 629944 216504
rect 538088 216464 629944 216492
rect 538088 216452 538094 216464
rect 629938 216452 629944 216464
rect 629996 216452 630002 216504
rect 628926 216424 628932 216436
rect 537312 216396 628932 216424
rect 628926 216384 628932 216396
rect 628984 216384 628990 216436
rect 610802 216356 610808 216368
rect 536760 216328 610808 216356
rect 610802 216316 610808 216328
rect 610860 216316 610866 216368
rect 609882 216288 609888 216300
rect 533080 216260 609888 216288
rect 609882 216248 609888 216260
rect 609940 216248 609946 216300
rect 673546 216248 673552 216300
rect 673604 216288 673610 216300
rect 675938 216288 675944 216300
rect 673604 216260 675944 216288
rect 673604 216248 673610 216260
rect 675938 216248 675944 216260
rect 675996 216248 676002 216300
rect 628006 216220 628012 216232
rect 530044 216192 628012 216220
rect 628006 216180 628012 216192
rect 628064 216180 628070 216232
rect 608962 216152 608968 216164
rect 524064 216124 608968 216152
rect 608962 216112 608968 216124
rect 609020 216112 609026 216164
rect 627086 216084 627092 216096
rect 523972 216056 627092 216084
rect 627086 216044 627092 216056
rect 627144 216044 627150 216096
rect 626166 216016 626172 216028
rect 520660 215988 626172 216016
rect 626166 215976 626172 215988
rect 626224 215976 626230 216028
rect 625246 215948 625252 215960
rect 517256 215920 625252 215948
rect 625246 215908 625252 215920
rect 625304 215908 625310 215960
rect 623406 215880 623412 215892
rect 512656 215852 623412 215880
rect 623406 215840 623412 215852
rect 623464 215840 623470 215892
rect 624326 215812 624332 215824
rect 507780 215784 624332 215812
rect 624326 215772 624332 215784
rect 624384 215772 624390 215824
rect 580902 215704 580908 215756
rect 580960 215744 580966 215756
rect 638770 215744 638776 215756
rect 580960 215716 638776 215744
rect 580960 215704 580966 215716
rect 638770 215704 638776 215716
rect 638828 215704 638834 215756
rect 636930 215676 636936 215688
rect 496786 215648 636936 215676
rect 636930 215636 636936 215648
rect 636988 215636 636994 215688
rect 636378 215608 636384 215620
rect 490116 215580 636384 215608
rect 636378 215568 636384 215580
rect 636436 215568 636442 215620
rect 638310 215540 638316 215552
rect 486712 215512 638316 215540
rect 638310 215500 638316 215512
rect 638368 215500 638374 215552
rect 673454 215500 673460 215552
rect 673512 215540 673518 215552
rect 675570 215540 675576 215552
rect 673512 215512 675576 215540
rect 673512 215500 673518 215512
rect 675570 215500 675576 215512
rect 675628 215500 675634 215552
rect 25130 215432 25136 215484
rect 25188 215472 25194 215484
rect 666186 215472 666192 215484
rect 25188 215444 666192 215472
rect 25188 215432 25194 215444
rect 666186 215432 666192 215444
rect 666244 215432 666250 215484
rect 674466 215432 674472 215484
rect 674524 215472 674530 215484
rect 675846 215472 675852 215484
rect 674524 215444 675852 215472
rect 674524 215432 674530 215444
rect 675846 215432 675852 215444
rect 675904 215432 675910 215484
rect 24854 215364 24860 215416
rect 24912 215404 24918 215416
rect 665266 215404 665272 215416
rect 24912 215376 665272 215404
rect 24912 215364 24918 215376
rect 665266 215364 665272 215376
rect 665324 215364 665330 215416
rect 674650 215364 674656 215416
rect 674708 215404 674714 215416
rect 675938 215404 675944 215416
rect 674708 215376 675944 215404
rect 674708 215364 674714 215376
rect 675938 215364 675944 215376
rect 675996 215364 676002 215416
rect 582282 215296 582288 215348
rect 582340 215336 582346 215348
rect 599854 215336 599860 215348
rect 582340 215308 599860 215336
rect 582340 215296 582346 215308
rect 599854 215296 599860 215308
rect 599912 215296 599918 215348
rect 603442 215296 603448 215348
rect 603500 215336 603506 215348
rect 604362 215336 604368 215348
rect 603500 215308 604368 215336
rect 603500 215296 603506 215308
rect 604362 215296 604368 215308
rect 604420 215336 604426 215348
rect 639230 215336 639236 215348
rect 604420 215308 639236 215336
rect 604420 215296 604426 215308
rect 639230 215296 639236 215308
rect 639288 215296 639294 215348
rect 674926 215296 674932 215348
rect 674984 215336 674990 215348
rect 676030 215336 676036 215348
rect 674984 215308 676036 215336
rect 674984 215296 674990 215308
rect 676030 215296 676036 215308
rect 676088 215296 676094 215348
rect 51816 215172 579138 215200
rect 41506 215092 41512 215144
rect 41564 215132 41570 215144
rect 46198 215132 46204 215144
rect 41564 215104 46204 215132
rect 41564 215092 41570 215104
rect 46198 215092 46204 215104
rect 46256 215092 46262 215144
rect 41506 214684 41512 214736
rect 41564 214724 41570 214736
rect 46106 214724 46112 214736
rect 41564 214696 46112 214724
rect 41564 214684 41570 214696
rect 46106 214684 46112 214696
rect 46164 214684 46170 214736
rect 41506 214276 41512 214328
rect 41564 214316 41570 214328
rect 50982 214316 50988 214328
rect 41564 214288 50988 214316
rect 41564 214276 41570 214288
rect 50982 214276 50988 214288
rect 51040 214276 51046 214328
rect 41506 214072 41512 214124
rect 41564 214112 41570 214124
rect 43530 214112 43536 214124
rect 41564 214084 43536 214112
rect 41564 214072 41570 214084
rect 43530 214072 43536 214084
rect 43588 214072 43594 214124
rect 33042 213596 33048 213648
rect 33100 213636 33106 213648
rect 51816 213636 51844 215172
rect 33100 213608 51844 213636
rect 51884 215104 579070 215132
rect 33100 213596 33106 213608
rect 32950 213528 32956 213580
rect 33008 213568 33014 213580
rect 51884 213568 51912 215104
rect 33008 213540 51912 213568
rect 51952 215036 579002 215064
rect 33008 213528 33014 213540
rect 32858 213460 32864 213512
rect 32916 213500 32922 213512
rect 51952 213500 51980 215036
rect 32916 213472 51980 213500
rect 52020 214968 578934 214996
rect 32916 213460 32922 213472
rect 41506 213392 41512 213444
rect 41564 213432 41570 213444
rect 52020 213432 52048 214968
rect 41564 213404 52048 213432
rect 578906 213432 578934 214968
rect 578974 213500 579002 215036
rect 579042 213568 579070 215104
rect 579110 213636 579138 215172
rect 659654 215092 659660 215144
rect 659712 215132 659718 215144
rect 660758 215132 660764 215144
rect 659712 215104 660764 215132
rect 659712 215092 659718 215104
rect 660758 215092 660764 215104
rect 660816 215092 660822 215144
rect 673730 214616 673736 214668
rect 673788 214656 673794 214668
rect 676030 214656 676036 214668
rect 673788 214628 676036 214656
rect 673788 214616 673794 214628
rect 676030 214616 676036 214628
rect 676088 214616 676094 214668
rect 673638 213800 673644 213852
rect 673696 213840 673702 213852
rect 675938 213840 675944 213852
rect 673696 213812 675944 213840
rect 673696 213800 673702 213812
rect 675938 213800 675944 213812
rect 675996 213800 676002 213852
rect 670878 213636 670884 213648
rect 579110 213608 670884 213636
rect 670878 213596 670884 213608
rect 670936 213596 670942 213648
rect 671798 213568 671804 213580
rect 579042 213540 671804 213568
rect 671798 213528 671804 213540
rect 671856 213528 671862 213580
rect 673086 213500 673092 213512
rect 578974 213472 673092 213500
rect 673086 213460 673092 213472
rect 673144 213460 673150 213512
rect 671890 213432 671896 213444
rect 578906 213404 671896 213432
rect 41564 213392 41570 213404
rect 671890 213392 671896 213404
rect 671948 213392 671954 213444
rect 580166 212576 580172 212628
rect 580224 212616 580230 212628
rect 598934 212616 598940 212628
rect 580224 212588 598940 212616
rect 580224 212576 580230 212588
rect 598934 212576 598940 212588
rect 598992 212576 598998 212628
rect 674282 212576 674288 212628
rect 674340 212616 674346 212628
rect 675938 212616 675944 212628
rect 674340 212588 675944 212616
rect 674340 212576 674346 212588
rect 675938 212576 675944 212588
rect 675996 212576 676002 212628
rect 580442 212508 580448 212560
rect 580500 212548 580506 212560
rect 599946 212548 599952 212560
rect 580500 212520 599952 212548
rect 580500 212508 580506 212520
rect 599946 212508 599952 212520
rect 600004 212508 600010 212560
rect 674742 212508 674748 212560
rect 674800 212548 674806 212560
rect 676030 212548 676036 212560
rect 674800 212520 676036 212548
rect 674800 212508 674806 212520
rect 676030 212508 676036 212520
rect 676088 212508 676094 212560
rect 655422 212440 655428 212492
rect 655480 212480 655486 212492
rect 669682 212480 669688 212492
rect 655480 212452 669688 212480
rect 655480 212440 655486 212452
rect 669682 212440 669688 212452
rect 669740 212440 669746 212492
rect 41506 212236 41512 212288
rect 41564 212276 41570 212288
rect 43162 212276 43168 212288
rect 41564 212248 43168 212276
rect 41564 212236 41570 212248
rect 43162 212236 43168 212248
rect 43220 212236 43226 212288
rect 41506 212100 41512 212152
rect 41564 212140 41570 212152
rect 43622 212140 43628 212152
rect 41564 212112 43628 212140
rect 41564 212100 41570 212112
rect 43622 212100 43628 212112
rect 43680 212100 43686 212152
rect 672994 212032 673000 212084
rect 673052 212072 673058 212084
rect 676030 212072 676036 212084
rect 673052 212044 676036 212072
rect 673052 212032 673058 212044
rect 676030 212032 676036 212044
rect 676088 212032 676094 212084
rect 662690 210060 662696 210112
rect 662748 210100 662754 210112
rect 663518 210100 663524 210112
rect 662748 210072 663524 210100
rect 662748 210060 662754 210072
rect 663518 210060 663524 210072
rect 663576 210060 663582 210112
rect 582282 209856 582288 209908
rect 582340 209896 582346 209908
rect 599118 209896 599124 209908
rect 582340 209868 599124 209896
rect 582340 209856 582346 209868
rect 599118 209856 599124 209868
rect 599176 209856 599182 209908
rect 580074 209788 580080 209840
rect 580132 209828 580138 209840
rect 601142 209828 601148 209840
rect 580132 209800 601148 209828
rect 580132 209788 580138 209800
rect 601142 209788 601148 209800
rect 601200 209788 601206 209840
rect 641806 209788 641812 209840
rect 641864 209828 641870 209840
rect 642082 209828 642088 209840
rect 641864 209800 642088 209828
rect 641864 209788 641870 209800
rect 642082 209788 642088 209800
rect 642140 209788 642146 209840
rect 644658 209788 644664 209840
rect 644716 209828 644722 209840
rect 644934 209828 644940 209840
rect 644716 209800 644940 209828
rect 644716 209788 644722 209800
rect 644934 209788 644940 209800
rect 644992 209788 644998 209840
rect 647418 209788 647424 209840
rect 647476 209828 647482 209840
rect 647694 209828 647700 209840
rect 647476 209800 647700 209828
rect 647476 209788 647482 209800
rect 647694 209788 647700 209800
rect 647752 209788 647758 209840
rect 675018 208360 675024 208412
rect 675076 208400 675082 208412
rect 675294 208400 675300 208412
rect 675076 208372 675300 208400
rect 675076 208360 675082 208372
rect 675294 208360 675300 208372
rect 675352 208360 675358 208412
rect 675110 208292 675116 208344
rect 675168 208332 675174 208344
rect 675386 208332 675392 208344
rect 675168 208304 675392 208332
rect 675168 208292 675174 208304
rect 675386 208292 675392 208304
rect 675444 208292 675450 208344
rect 41506 208224 41512 208276
rect 41564 208264 41570 208276
rect 43346 208264 43352 208276
rect 41564 208236 43352 208264
rect 41564 208224 41570 208236
rect 43346 208224 43352 208236
rect 43404 208224 43410 208276
rect 674834 208224 674840 208276
rect 674892 208264 674898 208276
rect 675294 208264 675300 208276
rect 674892 208236 675300 208264
rect 674892 208224 674898 208236
rect 675294 208224 675300 208236
rect 675352 208224 675358 208276
rect 41506 207272 41512 207324
rect 41564 207312 41570 207324
rect 43438 207312 43444 207324
rect 41564 207284 43444 207312
rect 41564 207272 41570 207284
rect 43438 207272 43444 207284
rect 43496 207272 43502 207324
rect 41782 207136 41788 207188
rect 41840 207176 41846 207188
rect 43714 207176 43720 207188
rect 41840 207148 43720 207176
rect 41840 207136 41846 207148
rect 43714 207136 43720 207148
rect 43772 207136 43778 207188
rect 582282 207068 582288 207120
rect 582340 207108 582346 207120
rect 601510 207108 601516 207120
rect 582340 207080 601516 207108
rect 582340 207068 582346 207080
rect 601510 207068 601516 207080
rect 601568 207068 601574 207120
rect 579798 207000 579804 207052
rect 579856 207040 579862 207052
rect 600958 207040 600964 207052
rect 579856 207012 600964 207040
rect 579856 207000 579862 207012
rect 600958 207000 600964 207012
rect 601016 207000 601022 207052
rect 666922 206932 666928 206984
rect 666980 206972 666986 206984
rect 675386 206972 675392 206984
rect 666980 206944 675392 206972
rect 666980 206932 666986 206944
rect 675386 206932 675392 206944
rect 675444 206932 675450 206984
rect 674834 206252 674840 206304
rect 674892 206292 674898 206304
rect 675754 206292 675760 206304
rect 674892 206264 675760 206292
rect 674892 206252 674898 206264
rect 675754 206252 675760 206264
rect 675812 206252 675818 206304
rect 673362 206184 673368 206236
rect 673420 206224 673426 206236
rect 675478 206224 675484 206236
rect 673420 206196 675484 206224
rect 673420 206184 673426 206196
rect 675478 206184 675484 206196
rect 675536 206184 675542 206236
rect 675662 206184 675668 206236
rect 675720 206184 675726 206236
rect 674558 205164 674564 205216
rect 674616 205204 674622 205216
rect 675294 205204 675300 205216
rect 674616 205176 675300 205204
rect 674616 205164 674622 205176
rect 675294 205164 675300 205176
rect 675352 205164 675358 205216
rect 674558 205028 674564 205080
rect 674616 205068 674622 205080
rect 675680 205068 675708 206184
rect 674616 205040 675708 205068
rect 674616 205028 674622 205040
rect 674926 204960 674932 205012
rect 674984 205000 674990 205012
rect 675386 205000 675392 205012
rect 674984 204972 675392 205000
rect 674984 204960 674990 204972
rect 675386 204960 675392 204972
rect 675444 204960 675450 205012
rect 581454 204280 581460 204332
rect 581512 204320 581518 204332
rect 599946 204320 599952 204332
rect 581512 204292 599952 204320
rect 581512 204280 581518 204292
rect 599946 204280 599952 204292
rect 600004 204280 600010 204332
rect 675110 203872 675116 203924
rect 675168 203912 675174 203924
rect 675294 203912 675300 203924
rect 675168 203884 675300 203912
rect 675168 203872 675174 203884
rect 675294 203872 675300 203884
rect 675352 203872 675358 203924
rect 674834 203804 674840 203856
rect 674892 203844 674898 203856
rect 674892 203816 675156 203844
rect 674892 203804 674898 203816
rect 675128 203788 675156 203816
rect 675110 203736 675116 203788
rect 675168 203736 675174 203788
rect 674282 203668 674288 203720
rect 674340 203708 674346 203720
rect 674834 203708 674840 203720
rect 674340 203680 674840 203708
rect 674340 203668 674346 203680
rect 674834 203668 674840 203680
rect 674892 203668 674898 203720
rect 673822 202716 673828 202768
rect 673880 202756 673886 202768
rect 675386 202756 675392 202768
rect 673880 202728 675392 202756
rect 673880 202716 673886 202728
rect 675386 202716 675392 202728
rect 675444 202716 675450 202768
rect 674650 202036 674656 202088
rect 674708 202076 674714 202088
rect 675386 202076 675392 202088
rect 674708 202048 675392 202076
rect 674708 202036 674714 202048
rect 675386 202036 675392 202048
rect 675444 202036 675450 202088
rect 582282 201560 582288 201612
rect 582340 201600 582346 201612
rect 599946 201600 599952 201612
rect 582340 201572 599952 201600
rect 582340 201560 582346 201572
rect 599946 201560 599952 201572
rect 600004 201560 600010 201612
rect 580626 201492 580632 201544
rect 580684 201532 580690 201544
rect 598934 201532 598940 201544
rect 580684 201504 598940 201532
rect 580684 201492 580690 201504
rect 598934 201492 598940 201504
rect 598992 201492 598998 201544
rect 674466 201492 674472 201544
rect 674524 201532 674530 201544
rect 675386 201532 675392 201544
rect 674524 201504 675392 201532
rect 674524 201492 674530 201504
rect 675386 201492 675392 201504
rect 675444 201492 675450 201544
rect 38010 201424 38016 201476
rect 38068 201464 38074 201476
rect 43530 201464 43536 201476
rect 38068 201436 43536 201464
rect 38068 201424 38074 201436
rect 43530 201424 43536 201436
rect 43588 201424 43594 201476
rect 41414 201356 41420 201408
rect 41472 201396 41478 201408
rect 43070 201396 43076 201408
rect 41472 201368 43076 201396
rect 41472 201356 41478 201368
rect 43070 201356 43076 201368
rect 43128 201356 43134 201408
rect 674742 200880 674748 200932
rect 674800 200920 674806 200932
rect 675386 200920 675392 200932
rect 674800 200892 675392 200920
rect 674800 200880 674806 200892
rect 675386 200880 675392 200892
rect 675444 200880 675450 200932
rect 673546 200744 673552 200796
rect 673604 200784 673610 200796
rect 674742 200784 674748 200796
rect 673604 200756 674748 200784
rect 673604 200744 673610 200756
rect 674742 200744 674748 200756
rect 674800 200744 674806 200796
rect 30190 200608 30196 200660
rect 30248 200648 30254 200660
rect 42702 200648 42708 200660
rect 30248 200620 42708 200648
rect 30248 200608 30254 200620
rect 42702 200608 42708 200620
rect 42760 200608 42766 200660
rect 30282 200472 30288 200524
rect 30340 200512 30346 200524
rect 42242 200512 42248 200524
rect 30340 200484 42248 200512
rect 30340 200472 30346 200484
rect 42242 200472 42248 200484
rect 42300 200472 42306 200524
rect 582282 200064 582288 200116
rect 582340 200104 582346 200116
rect 599946 200104 599952 200116
rect 582340 200076 599952 200104
rect 582340 200064 582346 200076
rect 599946 200064 599952 200076
rect 600004 200064 600010 200116
rect 41598 199112 41604 199164
rect 41656 199152 41662 199164
rect 43162 199152 43168 199164
rect 41656 199124 43168 199152
rect 41656 199112 41662 199124
rect 43162 199112 43168 199124
rect 43220 199112 43226 199164
rect 41690 198976 41696 199028
rect 41748 199016 41754 199028
rect 43254 199016 43260 199028
rect 41748 198988 43260 199016
rect 41748 198976 41754 198988
rect 43254 198976 43260 198988
rect 43312 198976 43318 199028
rect 41782 198908 41788 198960
rect 41840 198948 41846 198960
rect 43622 198948 43628 198960
rect 41840 198920 43628 198948
rect 41840 198908 41846 198920
rect 43622 198908 43628 198920
rect 43680 198908 43686 198960
rect 41506 198772 41512 198824
rect 41564 198812 41570 198824
rect 42334 198812 42340 198824
rect 41564 198784 42340 198812
rect 41564 198772 41570 198784
rect 42334 198772 42340 198784
rect 42392 198772 42398 198824
rect 581086 198704 581092 198756
rect 581144 198744 581150 198756
rect 599118 198744 599124 198756
rect 581144 198716 599124 198744
rect 581144 198704 581150 198716
rect 599118 198704 599124 198716
rect 599176 198704 599182 198756
rect 673454 198364 673460 198416
rect 673512 198404 673518 198416
rect 675386 198404 675392 198416
rect 673512 198376 675392 198404
rect 673512 198364 673518 198376
rect 675386 198364 675392 198376
rect 675444 198364 675450 198416
rect 673638 197752 673644 197804
rect 673696 197792 673702 197804
rect 675478 197792 675484 197804
rect 673696 197764 675484 197792
rect 673696 197752 673702 197764
rect 675478 197752 675484 197764
rect 675536 197752 675542 197804
rect 582282 197344 582288 197396
rect 582340 197384 582346 197396
rect 599302 197384 599308 197396
rect 582340 197356 599308 197384
rect 582340 197344 582346 197356
rect 599302 197344 599308 197356
rect 599360 197344 599366 197396
rect 580718 197276 580724 197328
rect 580776 197316 580782 197328
rect 599946 197316 599952 197328
rect 580776 197288 599952 197316
rect 580776 197276 580782 197288
rect 599946 197276 599952 197288
rect 600004 197276 600010 197328
rect 673730 197004 673736 197056
rect 673788 197044 673794 197056
rect 675386 197044 675392 197056
rect 673788 197016 675392 197044
rect 673788 197004 673794 197016
rect 675386 197004 675392 197016
rect 675444 197004 675450 197056
rect 42242 196528 42248 196580
rect 42300 196568 42306 196580
rect 42702 196568 42708 196580
rect 42300 196540 42708 196568
rect 42300 196528 42306 196540
rect 42702 196528 42708 196540
rect 42760 196528 42766 196580
rect 674834 196528 674840 196580
rect 674892 196568 674898 196580
rect 675386 196568 675392 196580
rect 674892 196540 675392 196568
rect 674892 196528 674898 196540
rect 675386 196528 675392 196540
rect 675444 196528 675450 196580
rect 673546 195304 673552 195356
rect 673604 195344 673610 195356
rect 675386 195344 675392 195356
rect 673604 195316 675392 195344
rect 673604 195304 673610 195316
rect 675386 195304 675392 195316
rect 675444 195304 675450 195356
rect 582190 194624 582196 194676
rect 582248 194664 582254 194676
rect 599118 194664 599124 194676
rect 582248 194636 599124 194664
rect 582248 194624 582254 194636
rect 599118 194624 599124 194636
rect 599176 194624 599182 194676
rect 582282 194556 582288 194608
rect 582340 194596 582346 194608
rect 599946 194596 599952 194608
rect 582340 194568 599952 194596
rect 582340 194556 582346 194568
rect 599946 194556 599952 194568
rect 600004 194556 600010 194608
rect 42058 193468 42064 193520
rect 42116 193508 42122 193520
rect 43070 193508 43076 193520
rect 42116 193480 43076 193508
rect 42116 193468 42122 193480
rect 43070 193468 43076 193480
rect 43128 193468 43134 193520
rect 674466 192788 674472 192840
rect 674524 192828 674530 192840
rect 675294 192828 675300 192840
rect 674524 192800 675300 192828
rect 674524 192788 674530 192800
rect 675294 192788 675300 192800
rect 675352 192788 675358 192840
rect 582190 191836 582196 191888
rect 582248 191876 582254 191888
rect 599118 191876 599124 191888
rect 582248 191848 599124 191876
rect 582248 191836 582254 191848
rect 599118 191836 599124 191848
rect 599176 191836 599182 191888
rect 582282 191768 582288 191820
rect 582340 191808 582346 191820
rect 599946 191808 599952 191820
rect 582340 191780 599952 191808
rect 582340 191768 582346 191780
rect 599946 191768 599952 191780
rect 600004 191768 600010 191820
rect 42334 191632 42340 191684
rect 42392 191672 42398 191684
rect 43162 191672 43168 191684
rect 42392 191644 43168 191672
rect 42392 191632 42398 191644
rect 43162 191632 43168 191644
rect 43220 191632 43226 191684
rect 674742 191632 674748 191684
rect 674800 191672 674806 191684
rect 675386 191672 675392 191684
rect 674800 191644 675392 191672
rect 674800 191632 674806 191644
rect 675386 191632 675392 191644
rect 675444 191632 675450 191684
rect 42058 191428 42064 191480
rect 42116 191468 42122 191480
rect 43254 191468 43260 191480
rect 42116 191440 43260 191468
rect 42116 191428 42122 191440
rect 43254 191428 43260 191440
rect 43312 191428 43318 191480
rect 581362 190408 581368 190460
rect 581420 190448 581426 190460
rect 599854 190448 599860 190460
rect 581420 190420 599860 190448
rect 581420 190408 581426 190420
rect 599854 190408 599860 190420
rect 599912 190408 599918 190460
rect 42242 190136 42248 190188
rect 42300 190176 42306 190188
rect 43438 190176 43444 190188
rect 42300 190148 43444 190176
rect 42300 190136 42306 190148
rect 43438 190136 43444 190148
rect 43496 190136 43502 190188
rect 42150 190068 42156 190120
rect 42208 190108 42214 190120
rect 43530 190108 43536 190120
rect 42208 190080 43536 190108
rect 42208 190068 42214 190080
rect 43530 190068 43536 190080
rect 43588 190068 43594 190120
rect 42426 189116 42432 189168
rect 42484 189156 42490 189168
rect 43346 189156 43352 189168
rect 42484 189128 43352 189156
rect 42484 189116 42490 189128
rect 43346 189116 43352 189128
rect 43404 189116 43410 189168
rect 42150 187824 42156 187876
rect 42208 187864 42214 187876
rect 43622 187864 43628 187876
rect 42208 187836 43628 187864
rect 42208 187824 42214 187836
rect 43622 187824 43628 187836
rect 43680 187824 43686 187876
rect 582190 187620 582196 187672
rect 582248 187660 582254 187672
rect 601602 187660 601608 187672
rect 582248 187632 601608 187660
rect 582248 187620 582254 187632
rect 601602 187620 601608 187632
rect 601660 187620 601666 187672
rect 582282 187552 582288 187604
rect 582340 187592 582346 187604
rect 600958 187592 600964 187604
rect 582340 187564 600964 187592
rect 582340 187552 582346 187564
rect 600958 187552 600964 187564
rect 601016 187552 601022 187604
rect 42150 187144 42156 187196
rect 42208 187184 42214 187196
rect 43714 187184 43720 187196
rect 42208 187156 43720 187184
rect 42208 187144 42214 187156
rect 43714 187144 43720 187156
rect 43772 187144 43778 187196
rect 579798 184832 579804 184884
rect 579856 184872 579862 184884
rect 599946 184872 599952 184884
rect 579856 184844 599952 184872
rect 579856 184832 579862 184844
rect 599946 184832 599952 184844
rect 600004 184832 600010 184884
rect 582282 184764 582288 184816
rect 582340 184804 582346 184816
rect 601510 184804 601516 184816
rect 582340 184776 601516 184804
rect 582340 184764 582346 184776
rect 601510 184764 601516 184776
rect 601568 184764 601574 184816
rect 42150 182112 42156 182164
rect 42208 182152 42214 182164
rect 48498 182152 48504 182164
rect 42208 182124 48504 182152
rect 42208 182112 42214 182124
rect 48498 182112 48504 182124
rect 48556 182112 48562 182164
rect 580166 182112 580172 182164
rect 580224 182152 580230 182164
rect 599854 182152 599860 182164
rect 580224 182124 599860 182152
rect 580224 182112 580230 182124
rect 599854 182112 599860 182124
rect 599912 182112 599918 182164
rect 582282 182044 582288 182096
rect 582340 182084 582346 182096
rect 600038 182084 600044 182096
rect 582340 182056 600044 182084
rect 582340 182044 582346 182056
rect 600038 182044 600044 182056
rect 600096 182044 600102 182096
rect 580534 179324 580540 179376
rect 580592 179364 580598 179376
rect 599762 179364 599768 179376
rect 580592 179336 599768 179364
rect 580592 179324 580598 179336
rect 599762 179324 599768 179336
rect 599820 179324 599826 179376
rect 580258 179256 580264 179308
rect 580316 179296 580322 179308
rect 599946 179296 599952 179308
rect 580316 179268 599952 179296
rect 580316 179256 580322 179268
rect 599946 179256 599952 179268
rect 600004 179256 600010 179308
rect 669406 178780 669412 178832
rect 669464 178820 669470 178832
rect 676214 178820 676220 178832
rect 669464 178792 676220 178820
rect 669464 178780 669470 178792
rect 676214 178780 676220 178792
rect 676272 178780 676278 178832
rect 675202 178576 675208 178628
rect 675260 178616 675266 178628
rect 676030 178616 676036 178628
rect 675260 178588 676036 178616
rect 675260 178576 675266 178588
rect 676030 178576 676036 178588
rect 676088 178576 676094 178628
rect 669498 178100 669504 178152
rect 669556 178140 669562 178152
rect 675938 178140 675944 178152
rect 669556 178112 675944 178140
rect 669556 178100 669562 178112
rect 675938 178100 675944 178112
rect 675996 178100 676002 178152
rect 669590 177692 669596 177744
rect 669648 177732 669654 177744
rect 675938 177732 675944 177744
rect 669648 177704 675944 177732
rect 669648 177692 669654 177704
rect 675938 177692 675944 177704
rect 675996 177692 676002 177744
rect 671706 176808 671712 176860
rect 671764 176848 671770 176860
rect 676030 176848 676036 176860
rect 671764 176820 676036 176848
rect 671764 176808 671770 176820
rect 676030 176808 676036 176820
rect 676088 176808 676094 176860
rect 581270 176672 581276 176724
rect 581328 176712 581334 176724
rect 598934 176712 598940 176724
rect 581328 176684 598940 176712
rect 581328 176672 581334 176684
rect 598934 176672 598940 176684
rect 598992 176672 598998 176724
rect 580534 176604 580540 176656
rect 580592 176644 580598 176656
rect 599854 176644 599860 176656
rect 580592 176616 599860 176644
rect 580592 176604 580598 176616
rect 599854 176604 599860 176616
rect 599912 176604 599918 176656
rect 675110 176604 675116 176656
rect 675168 176644 675174 176656
rect 676030 176644 676036 176656
rect 675168 176616 676036 176644
rect 675168 176604 675174 176616
rect 676030 176604 676036 176616
rect 676088 176604 676094 176656
rect 580810 176536 580816 176588
rect 580868 176576 580874 176588
rect 600130 176576 600136 176588
rect 580868 176548 600136 176576
rect 580868 176536 580874 176548
rect 600130 176536 600136 176548
rect 600188 176536 600194 176588
rect 675018 176332 675024 176384
rect 675076 176372 675082 176384
rect 676030 176372 676036 176384
rect 675076 176344 676036 176372
rect 675076 176332 675082 176344
rect 676030 176332 676036 176344
rect 676088 176332 676094 176384
rect 673178 175992 673184 176044
rect 673236 176032 673242 176044
rect 675938 176032 675944 176044
rect 673236 176004 675944 176032
rect 673236 175992 673242 176004
rect 675938 175992 675944 176004
rect 675996 175992 676002 176044
rect 673270 175176 673276 175228
rect 673328 175216 673334 175228
rect 675938 175216 675944 175228
rect 673328 175188 675944 175216
rect 673328 175176 673334 175188
rect 675938 175176 675944 175188
rect 675996 175176 676002 175228
rect 673362 174360 673368 174412
rect 673420 174400 673426 174412
rect 676030 174400 676036 174412
rect 673420 174372 676036 174400
rect 673420 174360 673426 174372
rect 676030 174360 676036 174372
rect 676088 174360 676094 174412
rect 580994 173884 581000 173936
rect 581052 173924 581058 173936
rect 599946 173924 599952 173936
rect 581052 173896 599952 173924
rect 581052 173884 581058 173896
rect 599946 173884 599952 173896
rect 600004 173884 600010 173936
rect 674558 173884 674564 173936
rect 674616 173924 674622 173936
rect 676030 173924 676036 173936
rect 674616 173896 676036 173924
rect 674616 173884 674622 173896
rect 676030 173884 676036 173896
rect 676088 173884 676094 173936
rect 582282 173816 582288 173868
rect 582340 173856 582346 173868
rect 599670 173856 599676 173868
rect 582340 173828 599676 173856
rect 582340 173816 582346 173828
rect 599670 173816 599676 173828
rect 599728 173816 599734 173868
rect 582190 173748 582196 173800
rect 582248 173788 582254 173800
rect 600038 173788 600044 173800
rect 582248 173760 600044 173788
rect 582248 173748 582254 173760
rect 600038 173748 600044 173760
rect 600096 173748 600102 173800
rect 673546 172864 673552 172916
rect 673604 172904 673610 172916
rect 676030 172904 676036 172916
rect 673604 172876 676036 172904
rect 673604 172864 673610 172876
rect 676030 172864 676036 172876
rect 676088 172864 676094 172916
rect 673730 172048 673736 172100
rect 673788 172088 673794 172100
rect 675938 172088 675944 172100
rect 673788 172060 675944 172088
rect 673788 172048 673794 172060
rect 675938 172048 675944 172060
rect 675996 172048 676002 172100
rect 674742 171640 674748 171692
rect 674800 171680 674806 171692
rect 675938 171680 675944 171692
rect 674800 171652 675944 171680
rect 674800 171640 674806 171652
rect 675938 171640 675944 171652
rect 675996 171640 676002 171692
rect 582006 171164 582012 171216
rect 582064 171204 582070 171216
rect 599946 171204 599952 171216
rect 582064 171176 599952 171204
rect 582064 171164 582070 171176
rect 599946 171164 599952 171176
rect 600004 171164 600010 171216
rect 674926 171164 674932 171216
rect 674984 171204 674990 171216
rect 675938 171204 675944 171216
rect 674984 171176 675944 171204
rect 674984 171164 674990 171176
rect 675938 171164 675944 171176
rect 675996 171164 676002 171216
rect 579890 171096 579896 171148
rect 579948 171136 579954 171148
rect 599854 171136 599860 171148
rect 579948 171108 599860 171136
rect 579948 171096 579954 171108
rect 599854 171096 599860 171108
rect 599912 171096 599918 171148
rect 675018 171096 675024 171148
rect 675076 171136 675082 171148
rect 676030 171136 676036 171148
rect 675076 171108 676036 171136
rect 675076 171096 675082 171108
rect 676030 171096 676036 171108
rect 676088 171096 676094 171148
rect 582282 171028 582288 171080
rect 582340 171068 582346 171080
rect 599762 171068 599768 171080
rect 582340 171040 599768 171068
rect 582340 171028 582346 171040
rect 599762 171028 599768 171040
rect 599820 171028 599826 171080
rect 674282 169600 674288 169652
rect 674340 169640 674346 169652
rect 675938 169640 675944 169652
rect 674340 169612 675944 169640
rect 674340 169600 674346 169612
rect 675938 169600 675944 169612
rect 675996 169600 676002 169652
rect 673638 169192 673644 169244
rect 673696 169232 673702 169244
rect 675846 169232 675852 169244
rect 673696 169204 675852 169232
rect 673696 169192 673702 169204
rect 675846 169192 675852 169204
rect 675904 169192 675910 169244
rect 673822 168580 673828 168632
rect 673880 168620 673886 168632
rect 675754 168620 675760 168632
rect 673880 168592 675760 168620
rect 673880 168580 673886 168592
rect 675754 168580 675760 168592
rect 675812 168580 675818 168632
rect 579798 168512 579804 168564
rect 579856 168552 579862 168564
rect 599946 168552 599952 168564
rect 579856 168524 599952 168552
rect 579856 168512 579862 168524
rect 599946 168512 599952 168524
rect 600004 168512 600010 168564
rect 674466 168512 674472 168564
rect 674524 168552 674530 168564
rect 675846 168552 675852 168564
rect 674524 168524 675852 168552
rect 674524 168512 674530 168524
rect 675846 168512 675852 168524
rect 675904 168512 675910 168564
rect 581730 168444 581736 168496
rect 581788 168484 581794 168496
rect 599026 168484 599032 168496
rect 581788 168456 599032 168484
rect 581788 168444 581794 168456
rect 599026 168444 599032 168456
rect 599084 168444 599090 168496
rect 674834 168444 674840 168496
rect 674892 168484 674898 168496
rect 675938 168484 675944 168496
rect 674892 168456 675944 168484
rect 674892 168444 674898 168456
rect 675938 168444 675944 168456
rect 675996 168444 676002 168496
rect 579706 168376 579712 168428
rect 579764 168416 579770 168428
rect 599854 168416 599860 168428
rect 579764 168388 599860 168416
rect 579764 168376 579770 168388
rect 599854 168376 599860 168388
rect 599912 168376 599918 168428
rect 675202 168376 675208 168428
rect 675260 168416 675266 168428
rect 676030 168416 676036 168428
rect 675260 168388 676036 168416
rect 675260 168376 675266 168388
rect 676030 168376 676036 168388
rect 676088 168376 676094 168428
rect 581454 168308 581460 168360
rect 581512 168348 581518 168360
rect 600314 168348 600320 168360
rect 581512 168320 600320 168348
rect 581512 168308 581518 168320
rect 600314 168308 600320 168320
rect 600372 168308 600378 168360
rect 671982 167016 671988 167068
rect 672040 167056 672046 167068
rect 676030 167056 676036 167068
rect 672040 167028 676036 167056
rect 672040 167016 672046 167028
rect 676030 167016 676036 167028
rect 676088 167016 676094 167068
rect 666554 165928 666560 165980
rect 666612 165968 666618 165980
rect 666922 165968 666928 165980
rect 666612 165940 666928 165968
rect 666612 165928 666618 165940
rect 666922 165928 666928 165940
rect 666980 165928 666986 165980
rect 582282 165724 582288 165776
rect 582340 165764 582346 165776
rect 599854 165764 599860 165776
rect 582340 165736 599860 165764
rect 582340 165724 582346 165736
rect 599854 165724 599860 165736
rect 599912 165724 599918 165776
rect 581914 165656 581920 165708
rect 581972 165696 581978 165708
rect 600038 165696 600044 165708
rect 581972 165668 600044 165696
rect 581972 165656 581978 165668
rect 600038 165656 600044 165668
rect 600096 165656 600102 165708
rect 581822 165588 581828 165640
rect 581880 165628 581886 165640
rect 599946 165628 599952 165640
rect 581880 165600 599952 165628
rect 581880 165588 581886 165600
rect 599946 165588 599952 165600
rect 600004 165588 600010 165640
rect 580258 165520 580264 165572
rect 580316 165560 580322 165572
rect 600130 165560 600136 165572
rect 580316 165532 600136 165560
rect 580316 165520 580322 165532
rect 600130 165520 600136 165532
rect 600188 165520 600194 165572
rect 582098 162936 582104 162988
rect 582156 162976 582162 162988
rect 599854 162976 599860 162988
rect 582156 162948 599860 162976
rect 582156 162936 582162 162948
rect 599854 162936 599860 162948
rect 599912 162936 599918 162988
rect 581454 162868 581460 162920
rect 581512 162908 581518 162920
rect 599946 162908 599952 162920
rect 581512 162880 599952 162908
rect 581512 162868 581518 162880
rect 599946 162868 599952 162880
rect 600004 162868 600010 162920
rect 675110 160488 675116 160540
rect 675168 160528 675174 160540
rect 675386 160528 675392 160540
rect 675168 160500 675392 160528
rect 675168 160488 675174 160500
rect 675386 160488 675392 160500
rect 675444 160488 675450 160540
rect 675018 160352 675024 160404
rect 675076 160352 675082 160404
rect 581270 160216 581276 160268
rect 581328 160256 581334 160268
rect 599854 160256 599860 160268
rect 581328 160228 599860 160256
rect 581328 160216 581334 160228
rect 599854 160216 599860 160228
rect 599912 160216 599918 160268
rect 580994 160148 581000 160200
rect 581052 160188 581058 160200
rect 599946 160188 599952 160200
rect 581052 160160 599952 160188
rect 581052 160148 581058 160160
rect 599946 160148 599952 160160
rect 600004 160148 600010 160200
rect 674742 160148 674748 160200
rect 674800 160188 674806 160200
rect 675036 160188 675064 160352
rect 675294 160188 675300 160200
rect 674800 160160 674972 160188
rect 675036 160160 675300 160188
rect 674800 160148 674806 160160
rect 674944 160132 674972 160160
rect 675294 160148 675300 160160
rect 675352 160148 675358 160200
rect 581362 160080 581368 160132
rect 581420 160120 581426 160132
rect 599302 160120 599308 160132
rect 581420 160092 599308 160120
rect 581420 160080 581426 160092
rect 599302 160080 599308 160092
rect 599360 160080 599366 160132
rect 674926 160080 674932 160132
rect 674984 160080 674990 160132
rect 675018 160012 675024 160064
rect 675076 160052 675082 160064
rect 675386 160052 675392 160064
rect 675076 160024 675392 160052
rect 675076 160012 675082 160024
rect 675386 160012 675392 160024
rect 675444 160012 675450 160064
rect 674926 159984 674932 159996
rect 674852 159956 674932 159984
rect 674852 159792 674880 159956
rect 674926 159944 674932 159956
rect 674984 159944 674990 159996
rect 674834 159740 674840 159792
rect 674892 159740 674898 159792
rect 674558 159536 674564 159588
rect 674616 159576 674622 159588
rect 675478 159576 675484 159588
rect 674616 159548 675484 159576
rect 674616 159536 674622 159548
rect 675478 159536 675484 159548
rect 675536 159536 675542 159588
rect 581546 157496 581552 157548
rect 581604 157536 581610 157548
rect 599946 157536 599952 157548
rect 581604 157508 599952 157536
rect 581604 157496 581610 157508
rect 599946 157496 599952 157508
rect 600004 157496 600010 157548
rect 581086 157428 581092 157480
rect 581144 157468 581150 157480
rect 600038 157468 600044 157480
rect 581144 157440 600044 157468
rect 581144 157428 581150 157440
rect 600038 157428 600044 157440
rect 600096 157428 600102 157480
rect 580718 157360 580724 157412
rect 580776 157400 580782 157412
rect 599854 157400 599860 157412
rect 580776 157372 599860 157400
rect 580776 157360 580782 157372
rect 599854 157360 599860 157372
rect 599912 157360 599918 157412
rect 666830 157292 666836 157344
rect 666888 157332 666894 157344
rect 675110 157332 675116 157344
rect 666888 157304 675116 157332
rect 666888 157292 666894 157304
rect 675110 157292 675116 157304
rect 675168 157292 675174 157344
rect 674466 155252 674472 155304
rect 674524 155292 674530 155304
rect 675110 155292 675116 155304
rect 674524 155264 675116 155292
rect 674524 155252 674530 155264
rect 675110 155252 675116 155264
rect 675168 155252 675174 155304
rect 673730 155184 673736 155236
rect 673788 155224 673794 155236
rect 675202 155224 675208 155236
rect 673788 155196 675208 155224
rect 673788 155184 673794 155196
rect 675202 155184 675208 155196
rect 675260 155184 675266 155236
rect 581178 154640 581184 154692
rect 581236 154680 581242 154692
rect 599946 154680 599952 154692
rect 581236 154652 599952 154680
rect 581236 154640 581242 154652
rect 599946 154640 599952 154652
rect 600004 154640 600010 154692
rect 580442 154572 580448 154624
rect 580500 154612 580506 154624
rect 599854 154612 599860 154624
rect 580500 154584 599860 154612
rect 580500 154572 580506 154584
rect 599854 154572 599860 154584
rect 599912 154572 599918 154624
rect 674282 152192 674288 152244
rect 674340 152232 674346 152244
rect 675110 152232 675116 152244
rect 674340 152204 675116 152232
rect 674340 152192 674346 152204
rect 675110 152192 675116 152204
rect 675168 152192 675174 152244
rect 673822 152124 673828 152176
rect 673880 152164 673886 152176
rect 675202 152164 675208 152176
rect 673880 152136 675208 152164
rect 673880 152124 673886 152136
rect 675202 152124 675208 152136
rect 675260 152124 675266 152176
rect 673638 152056 673644 152108
rect 673696 152096 673702 152108
rect 675294 152096 675300 152108
rect 673696 152068 675300 152096
rect 673696 152056 673702 152068
rect 675294 152056 675300 152068
rect 675352 152056 675358 152108
rect 582190 151920 582196 151972
rect 582248 151960 582254 151972
rect 599302 151960 599308 151972
rect 582248 151932 599308 151960
rect 582248 151920 582254 151932
rect 599302 151920 599308 151932
rect 599360 151920 599366 151972
rect 580810 151852 580816 151904
rect 580868 151892 580874 151904
rect 599946 151892 599952 151904
rect 580868 151864 599952 151892
rect 580868 151852 580874 151864
rect 599946 151852 599952 151864
rect 600004 151852 600010 151904
rect 580626 151784 580632 151836
rect 580684 151824 580690 151836
rect 599854 151824 599860 151836
rect 580684 151796 599860 151824
rect 580684 151784 580690 151796
rect 599854 151784 599860 151796
rect 599912 151784 599918 151836
rect 582006 149200 582012 149252
rect 582064 149240 582070 149252
rect 599762 149240 599768 149252
rect 582064 149212 599768 149240
rect 582064 149200 582070 149212
rect 599762 149200 599768 149212
rect 599820 149200 599826 149252
rect 582282 149132 582288 149184
rect 582340 149172 582346 149184
rect 598934 149172 598940 149184
rect 582340 149144 598940 149172
rect 582340 149132 582346 149144
rect 598934 149132 598940 149144
rect 598992 149132 598998 149184
rect 581822 149064 581828 149116
rect 581880 149104 581886 149116
rect 599946 149104 599952 149116
rect 581880 149076 599952 149104
rect 581880 149064 581886 149076
rect 599946 149064 599952 149076
rect 600004 149064 600010 149116
rect 673546 148452 673552 148504
rect 673604 148492 673610 148504
rect 675386 148492 675392 148504
rect 673604 148464 675392 148492
rect 673604 148452 673610 148464
rect 675386 148452 675392 148464
rect 675444 148452 675450 148504
rect 581638 146344 581644 146396
rect 581696 146384 581702 146396
rect 599946 146384 599952 146396
rect 581696 146356 599952 146384
rect 581696 146344 581702 146356
rect 599946 146344 599952 146356
rect 600004 146344 600010 146396
rect 580534 146276 580540 146328
rect 580592 146316 580598 146328
rect 599854 146316 599860 146328
rect 580592 146288 599860 146316
rect 580592 146276 580598 146288
rect 599854 146276 599860 146288
rect 599912 146276 599918 146328
rect 582098 143692 582104 143744
rect 582156 143732 582162 143744
rect 600038 143732 600044 143744
rect 582156 143704 600044 143732
rect 582156 143692 582162 143704
rect 600038 143692 600044 143704
rect 600096 143692 600102 143744
rect 581730 143624 581736 143676
rect 581788 143664 581794 143676
rect 599854 143664 599860 143676
rect 581788 143636 599860 143664
rect 581788 143624 581794 143636
rect 599854 143624 599860 143636
rect 599912 143624 599918 143676
rect 581454 143556 581460 143608
rect 581512 143596 581518 143608
rect 599946 143596 599952 143608
rect 581512 143568 599952 143596
rect 581512 143556 581518 143568
rect 599946 143556 599952 143568
rect 600004 143556 600010 143608
rect 581914 140904 581920 140956
rect 581972 140944 581978 140956
rect 599854 140944 599860 140956
rect 581972 140916 599860 140944
rect 581972 140904 581978 140916
rect 599854 140904 599860 140916
rect 599912 140904 599918 140956
rect 581270 140836 581276 140888
rect 581328 140876 581334 140888
rect 599946 140876 599952 140888
rect 581328 140848 599952 140876
rect 581328 140836 581334 140848
rect 599946 140836 599952 140848
rect 600004 140836 600010 140888
rect 580994 140768 581000 140820
rect 581052 140808 581058 140820
rect 599302 140808 599308 140820
rect 581052 140780 599308 140808
rect 581052 140768 581058 140780
rect 599302 140768 599308 140780
rect 599360 140768 599366 140820
rect 581546 138116 581552 138168
rect 581604 138156 581610 138168
rect 599854 138156 599860 138168
rect 581604 138128 599860 138156
rect 581604 138116 581610 138128
rect 599854 138116 599860 138128
rect 599912 138116 599918 138168
rect 581086 138048 581092 138100
rect 581144 138088 581150 138100
rect 599946 138088 599952 138100
rect 581144 138060 599952 138088
rect 581144 138048 581150 138060
rect 599946 138048 599952 138060
rect 600004 138048 600010 138100
rect 579890 137980 579896 138032
rect 579948 138020 579954 138032
rect 600038 138020 600044 138032
rect 579948 137992 600044 138020
rect 579948 137980 579954 137992
rect 600038 137980 600044 137992
rect 600096 137980 600102 138032
rect 581362 135328 581368 135380
rect 581420 135368 581426 135380
rect 599854 135368 599860 135380
rect 581420 135340 599860 135368
rect 581420 135328 581426 135340
rect 599854 135328 599860 135340
rect 599912 135328 599918 135380
rect 579982 135260 579988 135312
rect 580040 135300 580046 135312
rect 599946 135300 599952 135312
rect 580040 135272 599952 135300
rect 580040 135260 580046 135272
rect 599946 135260 599952 135272
rect 600004 135260 600010 135312
rect 669682 132880 669688 132932
rect 669740 132920 669746 132932
rect 676030 132920 676036 132932
rect 669740 132892 676036 132920
rect 669740 132880 669746 132892
rect 676030 132880 676036 132892
rect 676088 132880 676094 132932
rect 669314 132744 669320 132796
rect 669372 132784 669378 132796
rect 676214 132784 676220 132796
rect 669372 132756 676220 132784
rect 669372 132744 669378 132756
rect 676214 132744 676220 132756
rect 676272 132744 676278 132796
rect 580902 132608 580908 132660
rect 580960 132648 580966 132660
rect 599854 132648 599860 132660
rect 580960 132620 599860 132648
rect 580960 132608 580966 132620
rect 599854 132608 599860 132620
rect 599912 132608 599918 132660
rect 669222 132608 669228 132660
rect 669280 132648 669286 132660
rect 676122 132648 676128 132660
rect 669280 132620 676128 132648
rect 669280 132608 669286 132620
rect 676122 132608 676128 132620
rect 676180 132608 676186 132660
rect 580442 132540 580448 132592
rect 580500 132580 580506 132592
rect 599946 132580 599952 132592
rect 580500 132552 599952 132580
rect 580500 132540 580506 132552
rect 599946 132540 599952 132552
rect 600004 132540 600010 132592
rect 579798 132472 579804 132524
rect 579856 132512 579862 132524
rect 600038 132512 600044 132524
rect 579856 132484 600044 132512
rect 579856 132472 579862 132484
rect 600038 132472 600044 132484
rect 600096 132472 600102 132524
rect 671706 132268 671712 132320
rect 671764 132308 671770 132320
rect 676214 132308 676220 132320
rect 671764 132280 676220 132308
rect 671764 132268 671770 132280
rect 676214 132268 676220 132280
rect 676272 132268 676278 132320
rect 671890 131656 671896 131708
rect 671948 131696 671954 131708
rect 672166 131696 672172 131708
rect 671948 131668 672172 131696
rect 671948 131656 671954 131668
rect 672166 131656 672172 131668
rect 672224 131696 672230 131708
rect 676030 131696 676036 131708
rect 672224 131668 676036 131696
rect 672224 131656 672230 131668
rect 676030 131656 676036 131668
rect 676088 131656 676094 131708
rect 673178 131452 673184 131504
rect 673236 131492 673242 131504
rect 676214 131492 676220 131504
rect 673236 131464 676220 131492
rect 673236 131452 673242 131464
rect 676214 131452 676220 131464
rect 676272 131452 676278 131504
rect 672258 130840 672264 130892
rect 672316 130880 672322 130892
rect 676030 130880 676036 130892
rect 672316 130852 676036 130880
rect 672316 130840 672322 130852
rect 676030 130840 676036 130852
rect 676088 130840 676094 130892
rect 673270 130636 673276 130688
rect 673328 130676 673334 130688
rect 676214 130676 676220 130688
rect 673328 130648 676220 130676
rect 673328 130636 673334 130648
rect 676214 130636 676220 130648
rect 676272 130636 676278 130688
rect 671798 130024 671804 130076
rect 671856 130064 671862 130076
rect 672074 130064 672080 130076
rect 671856 130036 672080 130064
rect 671856 130024 671862 130036
rect 672074 130024 672080 130036
rect 672132 130064 672138 130076
rect 676030 130064 676036 130076
rect 672132 130036 676036 130064
rect 672132 130024 672138 130036
rect 676030 130024 676036 130036
rect 676088 130024 676094 130076
rect 581178 129888 581184 129940
rect 581236 129928 581242 129940
rect 599946 129928 599952 129940
rect 581236 129900 599952 129928
rect 581236 129888 581242 129900
rect 599946 129888 599952 129900
rect 600004 129888 600010 129940
rect 580626 129820 580632 129872
rect 580684 129860 580690 129872
rect 599762 129860 599768 129872
rect 580684 129832 599768 129860
rect 580684 129820 580690 129832
rect 599762 129820 599768 129832
rect 599820 129820 599826 129872
rect 580074 129752 580080 129804
rect 580132 129792 580138 129804
rect 598934 129792 598940 129804
rect 580132 129764 598940 129792
rect 580132 129752 580138 129764
rect 598934 129752 598940 129764
rect 598992 129752 598998 129804
rect 673362 129684 673368 129736
rect 673420 129724 673426 129736
rect 676030 129724 676036 129736
rect 673420 129696 676036 129724
rect 673420 129684 673426 129696
rect 676030 129684 676036 129696
rect 676088 129684 676094 129736
rect 672350 129412 672356 129464
rect 672408 129452 672414 129464
rect 673086 129452 673092 129464
rect 672408 129424 673092 129452
rect 672408 129412 672414 129424
rect 673086 129412 673092 129424
rect 673144 129452 673150 129464
rect 676214 129452 676220 129464
rect 673144 129424 676220 129452
rect 673144 129412 673150 129424
rect 676214 129412 676220 129424
rect 676272 129412 676278 129464
rect 674650 127712 674656 127764
rect 674708 127752 674714 127764
rect 676030 127752 676036 127764
rect 674708 127724 676036 127752
rect 674708 127712 674714 127724
rect 676030 127712 676036 127724
rect 676088 127712 676094 127764
rect 673546 127304 673552 127356
rect 673604 127344 673610 127356
rect 675938 127344 675944 127356
rect 673604 127316 675944 127344
rect 673604 127304 673610 127316
rect 675938 127304 675944 127316
rect 675996 127304 676002 127356
rect 582190 127032 582196 127084
rect 582248 127072 582254 127084
rect 599854 127072 599860 127084
rect 582248 127044 599860 127072
rect 582248 127032 582254 127044
rect 599854 127032 599860 127044
rect 599912 127032 599918 127084
rect 673822 127032 673828 127084
rect 673880 127072 673886 127084
rect 675938 127072 675944 127084
rect 673880 127044 675944 127072
rect 673880 127032 673886 127044
rect 675938 127032 675944 127044
rect 675996 127032 676002 127084
rect 580258 126964 580264 127016
rect 580316 127004 580322 127016
rect 599946 127004 599952 127016
rect 580316 126976 599952 127004
rect 580316 126964 580322 126976
rect 599946 126964 599952 126976
rect 600004 126964 600010 127016
rect 674742 126964 674748 127016
rect 674800 127004 674806 127016
rect 676030 127004 676036 127016
rect 674800 126976 676036 127004
rect 674800 126964 674806 126976
rect 676030 126964 676036 126976
rect 676088 126964 676094 127016
rect 674558 126080 674564 126132
rect 674616 126120 674622 126132
rect 676030 126120 676036 126132
rect 674616 126092 676036 126120
rect 674616 126080 674622 126092
rect 676030 126080 676036 126092
rect 676088 126080 676094 126132
rect 673638 124584 673644 124636
rect 673696 124624 673702 124636
rect 676122 124624 676128 124636
rect 673696 124596 676128 124624
rect 673696 124584 673702 124596
rect 676122 124584 676128 124596
rect 676180 124584 676186 124636
rect 674926 124448 674932 124500
rect 674984 124488 674990 124500
rect 676030 124488 676036 124500
rect 674984 124460 676036 124488
rect 674984 124448 674990 124460
rect 676030 124448 676036 124460
rect 676088 124448 676094 124500
rect 580718 124312 580724 124364
rect 580776 124352 580782 124364
rect 599946 124352 599952 124364
rect 580776 124324 599952 124352
rect 580776 124312 580782 124324
rect 599946 124312 599952 124324
rect 600004 124312 600010 124364
rect 673730 124312 673736 124364
rect 673788 124352 673794 124364
rect 676122 124352 676128 124364
rect 673788 124324 676128 124352
rect 673788 124312 673794 124324
rect 676122 124312 676128 124324
rect 676180 124312 676186 124364
rect 580350 124244 580356 124296
rect 580408 124284 580414 124296
rect 599854 124284 599860 124296
rect 580408 124256 599860 124284
rect 580408 124244 580414 124256
rect 599854 124244 599860 124256
rect 599912 124244 599918 124296
rect 674834 124244 674840 124296
rect 674892 124284 674898 124296
rect 675938 124284 675944 124296
rect 674892 124256 675944 124284
rect 674892 124244 674898 124256
rect 675938 124244 675944 124256
rect 675996 124244 676002 124296
rect 580166 124176 580172 124228
rect 580224 124216 580230 124228
rect 600038 124216 600044 124228
rect 580224 124188 600044 124216
rect 580224 124176 580230 124188
rect 600038 124176 600044 124188
rect 600096 124176 600102 124228
rect 675202 124176 675208 124228
rect 675260 124216 675266 124228
rect 676030 124216 676036 124228
rect 675260 124188 676036 124216
rect 675260 124176 675266 124188
rect 676030 124176 676036 124188
rect 676088 124176 676094 124228
rect 674282 123632 674288 123684
rect 674340 123672 674346 123684
rect 676030 123672 676036 123684
rect 674340 123644 676036 123672
rect 674340 123632 674346 123644
rect 676030 123632 676036 123644
rect 676088 123632 676094 123684
rect 582006 121592 582012 121644
rect 582064 121632 582070 121644
rect 599578 121632 599584 121644
rect 582064 121604 599584 121632
rect 582064 121592 582070 121604
rect 599578 121592 599584 121604
rect 599636 121592 599642 121644
rect 672442 121592 672448 121644
rect 672500 121632 672506 121644
rect 676214 121632 676220 121644
rect 672500 121604 676220 121632
rect 672500 121592 672506 121604
rect 676214 121592 676220 121604
rect 676272 121592 676278 121644
rect 580810 121524 580816 121576
rect 580868 121564 580874 121576
rect 599946 121564 599952 121576
rect 580868 121536 599952 121564
rect 580868 121524 580874 121536
rect 599946 121524 599952 121536
rect 600004 121524 600010 121576
rect 580534 121456 580540 121508
rect 580592 121496 580598 121508
rect 599854 121496 599860 121508
rect 580592 121468 599860 121496
rect 580592 121456 580598 121468
rect 599854 121456 599860 121468
rect 599912 121456 599918 121508
rect 675018 121456 675024 121508
rect 675076 121496 675082 121508
rect 676030 121496 676036 121508
rect 675076 121468 676036 121496
rect 675076 121456 675082 121468
rect 676030 121456 676036 121468
rect 676088 121456 676094 121508
rect 586422 118804 586428 118856
rect 586480 118844 586486 118856
rect 599854 118844 599860 118856
rect 586480 118816 599860 118844
rect 586480 118804 586486 118816
rect 599854 118804 599860 118816
rect 599912 118804 599918 118856
rect 583662 118736 583668 118788
rect 583720 118776 583726 118788
rect 599946 118776 599952 118788
rect 583720 118748 599952 118776
rect 583720 118736 583726 118748
rect 599946 118736 599952 118748
rect 600004 118736 600010 118788
rect 582282 118668 582288 118720
rect 582340 118708 582346 118720
rect 600038 118708 600044 118720
rect 582340 118680 600044 118708
rect 582340 118668 582346 118680
rect 600038 118668 600044 118680
rect 600096 118668 600102 118720
rect 582098 116016 582104 116068
rect 582156 116056 582162 116068
rect 599854 116056 599860 116068
rect 582156 116028 599860 116056
rect 582156 116016 582162 116028
rect 599854 116016 599860 116028
rect 599912 116016 599918 116068
rect 581822 115948 581828 116000
rect 581880 115988 581886 116000
rect 599946 115988 599952 116000
rect 581880 115960 599952 115988
rect 581880 115948 581886 115960
rect 599946 115948 599952 115960
rect 600004 115948 600010 116000
rect 666738 115880 666744 115932
rect 666796 115920 666802 115932
rect 675386 115920 675392 115932
rect 666796 115892 675392 115920
rect 666796 115880 666802 115892
rect 675386 115880 675392 115892
rect 675444 115880 675450 115932
rect 674650 114316 674656 114368
rect 674708 114356 674714 114368
rect 675202 114356 675208 114368
rect 674708 114328 675208 114356
rect 674708 114316 674714 114328
rect 675202 114316 675208 114328
rect 675260 114316 675266 114368
rect 674742 113704 674748 113756
rect 674800 113744 674806 113756
rect 675202 113744 675208 113756
rect 674800 113716 675208 113744
rect 674800 113704 674806 113716
rect 675202 113704 675208 113716
rect 675260 113704 675266 113756
rect 581914 113296 581920 113348
rect 581972 113336 581978 113348
rect 600038 113336 600044 113348
rect 581972 113308 600044 113336
rect 581972 113296 581978 113308
rect 600038 113296 600044 113308
rect 600096 113296 600102 113348
rect 581638 113228 581644 113280
rect 581696 113268 581702 113280
rect 599946 113268 599952 113280
rect 581696 113240 599952 113268
rect 581696 113228 581702 113240
rect 599946 113228 599952 113240
rect 600004 113228 600010 113280
rect 581730 113160 581736 113212
rect 581788 113200 581794 113212
rect 599854 113200 599860 113212
rect 581788 113172 599860 113200
rect 581788 113160 581794 113172
rect 599854 113160 599860 113172
rect 599912 113160 599918 113212
rect 674926 111868 674932 111920
rect 674984 111908 674990 111920
rect 675202 111908 675208 111920
rect 674984 111880 675208 111908
rect 674984 111868 674990 111880
rect 675202 111868 675208 111880
rect 675260 111868 675266 111920
rect 674834 111120 674840 111172
rect 674892 111160 674898 111172
rect 675386 111160 675392 111172
rect 674892 111132 675392 111160
rect 674892 111120 674898 111132
rect 675386 111120 675392 111132
rect 675444 111120 675450 111172
rect 581270 110508 581276 110560
rect 581328 110548 581334 110560
rect 599946 110548 599952 110560
rect 581328 110520 599952 110548
rect 581328 110508 581334 110520
rect 599946 110508 599952 110520
rect 600004 110508 600010 110560
rect 581454 110440 581460 110492
rect 581512 110480 581518 110492
rect 598934 110480 598940 110492
rect 581512 110452 598940 110480
rect 581512 110440 581518 110452
rect 598934 110440 598940 110452
rect 598992 110440 598998 110492
rect 673730 110032 673736 110084
rect 673788 110072 673794 110084
rect 675110 110072 675116 110084
rect 673788 110044 675116 110072
rect 673788 110032 673794 110044
rect 675110 110032 675116 110044
rect 675168 110032 675174 110084
rect 673822 108196 673828 108248
rect 673880 108236 673886 108248
rect 675386 108236 675392 108248
rect 673880 108208 675392 108236
rect 673880 108196 673886 108208
rect 675386 108196 675392 108208
rect 675444 108196 675450 108248
rect 581546 107720 581552 107772
rect 581604 107760 581610 107772
rect 599854 107760 599860 107772
rect 581604 107732 599860 107760
rect 581604 107720 581610 107732
rect 599854 107720 599860 107732
rect 599912 107720 599918 107772
rect 580994 107652 581000 107704
rect 581052 107692 581058 107704
rect 599946 107692 599952 107704
rect 581052 107664 599952 107692
rect 581052 107652 581058 107664
rect 599946 107652 599952 107664
rect 600004 107652 600010 107704
rect 674282 107516 674288 107568
rect 674340 107556 674346 107568
rect 675386 107556 675392 107568
rect 674340 107528 675392 107556
rect 674340 107516 674346 107528
rect 675386 107516 675392 107528
rect 675444 107516 675450 107568
rect 673638 105680 673644 105732
rect 673696 105720 673702 105732
rect 675110 105720 675116 105732
rect 673696 105692 675116 105720
rect 673696 105680 673702 105692
rect 675110 105680 675116 105692
rect 675168 105680 675174 105732
rect 581362 104932 581368 104984
rect 581420 104972 581426 104984
rect 599854 104972 599860 104984
rect 581420 104944 599860 104972
rect 581420 104932 581426 104944
rect 599854 104932 599860 104944
rect 599912 104932 599918 104984
rect 581086 104864 581092 104916
rect 581144 104904 581150 104916
rect 599946 104904 599952 104916
rect 581144 104876 599952 104904
rect 581144 104864 581150 104876
rect 599946 104864 599952 104876
rect 600004 104864 600010 104916
rect 673546 104524 673552 104576
rect 673604 104564 673610 104576
rect 675110 104564 675116 104576
rect 673604 104536 675116 104564
rect 673604 104524 673610 104536
rect 675110 104524 675116 104536
rect 675168 104524 675174 104576
rect 657722 99764 657728 99816
rect 657780 99804 657786 99816
rect 660896 99804 660902 99816
rect 657780 99776 660902 99804
rect 657780 99764 657786 99776
rect 660896 99764 660902 99776
rect 660954 99764 660960 99816
rect 580902 99356 580908 99408
rect 580960 99396 580966 99408
rect 599946 99396 599952 99408
rect 580960 99368 599952 99396
rect 580960 99356 580966 99368
rect 599946 99356 599952 99368
rect 600004 99356 600010 99408
rect 633802 96568 633808 96620
rect 633860 96608 633866 96620
rect 636378 96608 636384 96620
rect 633860 96580 636384 96608
rect 633860 96568 633866 96580
rect 636378 96568 636384 96580
rect 636436 96568 636442 96620
rect 637022 96568 637028 96620
rect 637080 96608 637086 96620
rect 642174 96608 642180 96620
rect 637080 96580 642180 96608
rect 637080 96568 637086 96580
rect 642174 96568 642180 96580
rect 642232 96568 642238 96620
rect 655974 96568 655980 96620
rect 656032 96608 656038 96620
rect 659562 96608 659568 96620
rect 656032 96580 659568 96608
rect 656032 96568 656038 96580
rect 659562 96568 659568 96580
rect 659620 96568 659626 96620
rect 661862 96568 661868 96620
rect 661920 96608 661926 96620
rect 663058 96608 663064 96620
rect 661920 96580 663064 96608
rect 661920 96568 661926 96580
rect 663058 96568 663064 96580
rect 663116 96568 663122 96620
rect 634446 96500 634452 96552
rect 634504 96540 634510 96552
rect 637574 96540 637580 96552
rect 634504 96512 637580 96540
rect 634504 96500 634510 96512
rect 637574 96500 637580 96512
rect 637632 96500 637638 96552
rect 654686 96500 654692 96552
rect 654744 96540 654750 96552
rect 658274 96540 658280 96552
rect 654744 96512 658280 96540
rect 654744 96500 654750 96512
rect 658274 96500 658280 96512
rect 658332 96500 658338 96552
rect 659102 96500 659108 96552
rect 659160 96540 659166 96552
rect 662506 96540 662512 96552
rect 659160 96512 662512 96540
rect 659160 96500 659166 96512
rect 662506 96500 662512 96512
rect 662564 96500 662570 96552
rect 635734 96432 635740 96484
rect 635792 96472 635798 96484
rect 639874 96472 639880 96484
rect 635792 96444 639880 96472
rect 635792 96432 635798 96444
rect 639874 96432 639880 96444
rect 639932 96432 639938 96484
rect 652018 96432 652024 96484
rect 652076 96472 652082 96484
rect 661954 96472 661960 96484
rect 652076 96444 661960 96472
rect 652076 96432 652082 96444
rect 661954 96432 661960 96444
rect 662012 96432 662018 96484
rect 636286 96364 636292 96416
rect 636344 96404 636350 96416
rect 640978 96404 640984 96416
rect 636344 96376 640984 96404
rect 636344 96364 636350 96376
rect 640978 96364 640984 96376
rect 641036 96364 641042 96416
rect 633066 96296 633072 96348
rect 633124 96336 633130 96348
rect 635274 96336 635280 96348
rect 633124 96308 635280 96336
rect 633124 96296 633130 96308
rect 635274 96296 635280 96308
rect 635332 96296 635338 96348
rect 640334 96228 640340 96280
rect 640392 96268 640398 96280
rect 641714 96268 641720 96280
rect 640392 96240 641720 96268
rect 640392 96228 640398 96240
rect 641714 96228 641720 96240
rect 641772 96228 641778 96280
rect 638954 96160 638960 96212
rect 639012 96200 639018 96212
rect 646222 96200 646228 96212
rect 639012 96172 646228 96200
rect 639012 96160 639018 96172
rect 646222 96160 646228 96172
rect 646280 96160 646286 96212
rect 622026 96092 622032 96144
rect 622084 96132 622090 96144
rect 642818 96132 642824 96144
rect 622084 96104 642824 96132
rect 622084 96092 622090 96104
rect 642818 96092 642824 96104
rect 642876 96092 642882 96144
rect 631134 96024 631140 96076
rect 631192 96064 631198 96076
rect 632100 96064 632106 96076
rect 631192 96036 632106 96064
rect 631192 96024 631198 96036
rect 632100 96024 632106 96036
rect 632158 96024 632164 96076
rect 632422 96024 632428 96076
rect 632480 96064 632486 96076
rect 634400 96064 634406 96076
rect 632480 96036 634406 96064
rect 632480 96024 632486 96036
rect 634400 96024 634406 96036
rect 634458 96024 634464 96076
rect 635090 96024 635096 96076
rect 635148 96064 635154 96076
rect 639000 96064 639006 96076
rect 635148 96036 639006 96064
rect 635148 96024 635154 96036
rect 639000 96024 639006 96036
rect 639058 96024 639064 96076
rect 640058 95956 640064 96008
rect 640116 95996 640122 96008
rect 646038 95996 646044 96008
rect 640116 95968 646044 95996
rect 640116 95956 640122 95968
rect 646038 95956 646044 95968
rect 646096 95956 646102 96008
rect 631778 95888 631784 95940
rect 631836 95928 631842 95940
rect 632974 95928 632980 95940
rect 631836 95900 632980 95928
rect 631836 95888 631842 95900
rect 632974 95888 632980 95900
rect 633032 95888 633038 95940
rect 639598 95888 639604 95940
rect 639656 95928 639662 95940
rect 645946 95928 645952 95940
rect 639656 95900 645952 95928
rect 639656 95888 639662 95900
rect 645946 95888 645952 95900
rect 646004 95888 646010 95940
rect 623682 95820 623688 95872
rect 623740 95860 623746 95872
rect 642910 95860 642916 95872
rect 623740 95832 642916 95860
rect 623740 95820 623746 95832
rect 642910 95820 642916 95832
rect 642968 95820 642974 95872
rect 647510 95820 647516 95872
rect 647568 95860 647574 95872
rect 651558 95860 651564 95872
rect 647568 95832 651564 95860
rect 647568 95820 647574 95832
rect 651558 95820 651564 95832
rect 651616 95820 651622 95872
rect 621382 95752 621388 95804
rect 621440 95792 621446 95804
rect 643002 95792 643008 95804
rect 621440 95764 643008 95792
rect 621440 95752 621446 95764
rect 643002 95752 643008 95764
rect 643060 95752 643066 95804
rect 626534 95684 626540 95736
rect 626592 95724 626598 95736
rect 640334 95724 640340 95736
rect 626592 95696 640340 95724
rect 626592 95684 626598 95696
rect 640334 95684 640340 95696
rect 640392 95684 640398 95736
rect 640886 95684 640892 95736
rect 640944 95724 640950 95736
rect 645854 95724 645860 95736
rect 640944 95696 645860 95724
rect 640944 95684 640950 95696
rect 645854 95684 645860 95696
rect 645912 95684 645918 95736
rect 596174 95616 596180 95668
rect 596232 95656 596238 95668
rect 607674 95656 607680 95668
rect 596232 95628 607680 95656
rect 596232 95616 596238 95628
rect 607674 95616 607680 95628
rect 607732 95616 607738 95668
rect 638310 95616 638316 95668
rect 638368 95656 638374 95668
rect 642634 95656 642640 95668
rect 638368 95628 642640 95656
rect 638368 95616 638374 95628
rect 642634 95616 642640 95628
rect 642692 95616 642698 95668
rect 652662 95616 652668 95668
rect 652720 95656 652726 95668
rect 663794 95656 663800 95668
rect 652720 95628 663800 95656
rect 652720 95616 652726 95628
rect 663794 95616 663800 95628
rect 663852 95616 663858 95668
rect 607490 95548 607496 95600
rect 607548 95588 607554 95600
rect 608962 95588 608968 95600
rect 607548 95560 608968 95588
rect 607548 95548 607554 95560
rect 608962 95548 608968 95560
rect 609020 95548 609026 95600
rect 610342 95548 610348 95600
rect 610400 95588 610406 95600
rect 611538 95588 611544 95600
rect 610400 95560 611544 95588
rect 610400 95548 610406 95560
rect 611538 95548 611544 95560
rect 611596 95548 611602 95600
rect 616138 95548 616144 95600
rect 616196 95588 616202 95600
rect 623222 95588 623228 95600
rect 616196 95560 623228 95588
rect 616196 95548 616202 95560
rect 623222 95548 623228 95560
rect 623280 95548 623286 95600
rect 623774 95548 623780 95600
rect 623832 95588 623838 95600
rect 624602 95588 624608 95600
rect 623832 95560 624608 95588
rect 623832 95548 623838 95560
rect 624602 95548 624608 95560
rect 624660 95548 624666 95600
rect 637482 95548 637488 95600
rect 637540 95548 637546 95600
rect 641622 95548 641628 95600
rect 641680 95588 641686 95600
rect 643094 95588 643100 95600
rect 641680 95560 643100 95588
rect 641680 95548 641686 95560
rect 643094 95548 643100 95560
rect 643152 95548 643158 95600
rect 656986 95548 656992 95600
rect 657044 95588 657050 95600
rect 659194 95588 659200 95600
rect 657044 95560 659200 95588
rect 657044 95548 657050 95560
rect 659194 95548 659200 95560
rect 659252 95548 659258 95600
rect 619358 95480 619364 95532
rect 619416 95520 619422 95532
rect 621198 95520 621204 95532
rect 619416 95492 621204 95520
rect 619416 95480 619422 95492
rect 621198 95480 621204 95492
rect 621256 95480 621262 95532
rect 637500 95520 637528 95548
rect 642726 95520 642732 95532
rect 637500 95492 642732 95520
rect 642726 95480 642732 95492
rect 642784 95480 642790 95532
rect 660574 95480 660580 95532
rect 660632 95520 660638 95532
rect 661402 95520 661408 95532
rect 660632 95492 661408 95520
rect 660632 95480 660638 95492
rect 661402 95480 661408 95492
rect 661460 95480 661466 95532
rect 620002 95412 620008 95464
rect 620060 95452 620066 95464
rect 623498 95452 623504 95464
rect 620060 95424 623504 95452
rect 620060 95412 620066 95424
rect 623498 95412 623504 95424
rect 623556 95412 623562 95464
rect 642818 95412 642824 95464
rect 642876 95452 642882 95464
rect 642876 95424 642956 95452
rect 642876 95412 642882 95424
rect 588078 95344 588084 95396
rect 588136 95384 588142 95396
rect 610894 95384 610900 95396
rect 588136 95356 610900 95384
rect 588136 95344 588142 95356
rect 610894 95344 610900 95356
rect 610952 95344 610958 95396
rect 581178 95276 581184 95328
rect 581236 95316 581242 95328
rect 612182 95316 612188 95328
rect 581236 95288 612188 95316
rect 581236 95276 581242 95288
rect 612182 95276 612188 95288
rect 612240 95276 612246 95328
rect 620738 95276 620744 95328
rect 620796 95316 620802 95328
rect 642818 95316 642824 95328
rect 620796 95288 642824 95316
rect 620796 95276 620802 95288
rect 642818 95276 642824 95288
rect 642876 95276 642882 95328
rect 575658 95208 575664 95260
rect 575716 95248 575722 95260
rect 606386 95248 606392 95260
rect 575716 95220 606392 95248
rect 575716 95208 575722 95220
rect 606386 95208 606392 95220
rect 606444 95208 606450 95260
rect 622670 95208 622676 95260
rect 622728 95248 622734 95260
rect 623682 95248 623688 95260
rect 622728 95220 623688 95248
rect 622728 95208 622734 95220
rect 623682 95208 623688 95220
rect 623740 95208 623746 95260
rect 617426 95072 617432 95124
rect 617484 95112 617490 95124
rect 621934 95112 621940 95124
rect 617484 95084 621940 95112
rect 617484 95072 617490 95084
rect 621934 95072 621940 95084
rect 621992 95072 621998 95124
rect 614850 94936 614856 94988
rect 614908 94976 614914 94988
rect 615402 94976 615408 94988
rect 614908 94948 615408 94976
rect 614908 94936 614914 94948
rect 615402 94936 615408 94948
rect 615460 94936 615466 94988
rect 618714 94936 618720 94988
rect 618772 94976 618778 94988
rect 623314 94976 623320 94988
rect 618772 94948 623320 94976
rect 618772 94936 618778 94948
rect 623314 94936 623320 94948
rect 623372 94936 623378 94988
rect 616782 94868 616788 94920
rect 616840 94908 616846 94920
rect 622486 94908 622492 94920
rect 616840 94880 622492 94908
rect 616840 94868 616846 94880
rect 622486 94868 622492 94880
rect 622544 94868 622550 94920
rect 642928 94784 642956 95424
rect 646774 95276 646780 95328
rect 646832 95316 646838 95328
rect 663334 95316 663340 95328
rect 646832 95288 663340 95316
rect 646832 95276 646838 95288
rect 663334 95276 663340 95288
rect 663392 95276 663398 95328
rect 657078 95208 657084 95260
rect 657136 95248 657142 95260
rect 657906 95248 657912 95260
rect 657136 95220 657912 95248
rect 657136 95208 657142 95220
rect 657906 95208 657912 95220
rect 657964 95208 657970 95260
rect 646130 95140 646136 95192
rect 646188 95180 646194 95192
rect 663426 95180 663432 95192
rect 646188 95152 663432 95180
rect 646188 95140 646194 95152
rect 663426 95140 663432 95152
rect 663484 95140 663490 95192
rect 643462 95072 643468 95124
rect 643520 95112 643526 95124
rect 644842 95112 644848 95124
rect 643520 95084 644848 95112
rect 643520 95072 643526 95084
rect 644842 95072 644848 95084
rect 644900 95072 644906 95124
rect 648614 94936 648620 94988
rect 648672 94976 648678 94988
rect 650730 94976 650736 94988
rect 648672 94948 650736 94976
rect 648672 94936 648678 94948
rect 650730 94936 650736 94948
rect 650788 94936 650794 94988
rect 646038 94868 646044 94920
rect 646096 94908 646102 94920
rect 646222 94908 646228 94920
rect 646096 94880 646228 94908
rect 646096 94868 646102 94880
rect 646222 94868 646228 94880
rect 646280 94868 646286 94920
rect 648706 94800 648712 94852
rect 648764 94840 648770 94852
rect 649442 94840 649448 94852
rect 648764 94812 649448 94840
rect 648764 94800 648770 94812
rect 649442 94800 649448 94812
rect 649500 94800 649506 94852
rect 642910 94732 642916 94784
rect 642968 94732 642974 94784
rect 653306 94732 653312 94784
rect 653364 94772 653370 94784
rect 663702 94772 663708 94784
rect 653364 94744 663708 94772
rect 653364 94732 653370 94744
rect 663702 94732 663708 94744
rect 663760 94732 663766 94784
rect 647510 94664 647516 94716
rect 647568 94704 647574 94716
rect 648154 94704 648160 94716
rect 647568 94676 648160 94704
rect 647568 94664 647574 94676
rect 648154 94664 648160 94676
rect 648212 94664 648218 94716
rect 651834 94664 651840 94716
rect 651892 94704 651898 94716
rect 653398 94704 653404 94716
rect 651892 94676 653404 94704
rect 651892 94664 651898 94676
rect 653398 94664 653404 94676
rect 653456 94664 653462 94716
rect 656618 94664 656624 94716
rect 656676 94704 656682 94716
rect 663886 94704 663892 94716
rect 656676 94676 663892 94704
rect 656676 94664 656682 94676
rect 663886 94664 663892 94676
rect 663944 94664 663950 94716
rect 657262 94596 657268 94648
rect 657320 94636 657326 94648
rect 663518 94636 663524 94648
rect 657320 94608 663524 94636
rect 657320 94596 657326 94608
rect 663518 94596 663524 94608
rect 663576 94596 663582 94648
rect 618070 94528 618076 94580
rect 618128 94568 618134 94580
rect 623130 94568 623136 94580
rect 618128 94540 623136 94568
rect 618128 94528 618134 94540
rect 623130 94528 623136 94540
rect 623188 94528 623194 94580
rect 648798 94528 648804 94580
rect 648856 94568 648862 94580
rect 650086 94568 650092 94580
rect 648856 94540 650092 94568
rect 648856 94528 648862 94540
rect 650086 94528 650092 94540
rect 650144 94528 650150 94580
rect 656894 94528 656900 94580
rect 656952 94568 656958 94580
rect 658550 94568 658556 94580
rect 656952 94540 658556 94568
rect 656952 94528 656958 94540
rect 658550 94528 658556 94540
rect 658608 94528 658614 94580
rect 648062 94460 648068 94512
rect 648120 94500 648126 94512
rect 659838 94500 659844 94512
rect 648120 94472 659844 94500
rect 648120 94460 648126 94472
rect 659838 94460 659844 94472
rect 659896 94460 659902 94512
rect 660390 94460 660396 94512
rect 660448 94460 660454 94512
rect 643554 94188 643560 94240
rect 643612 94228 643618 94240
rect 660408 94228 660436 94460
rect 643612 94200 660436 94228
rect 643612 94188 643618 94200
rect 644750 94120 644756 94172
rect 644808 94160 644814 94172
rect 652754 94160 652760 94172
rect 644808 94132 652760 94160
rect 644808 94120 644814 94132
rect 652754 94120 652760 94132
rect 652812 94120 652818 94172
rect 644198 94052 644204 94104
rect 644256 94092 644262 94104
rect 654042 94092 654048 94104
rect 644256 94064 654048 94092
rect 644256 94052 644262 94064
rect 654042 94052 654048 94064
rect 654100 94052 654106 94104
rect 607214 93848 607220 93900
rect 607272 93888 607278 93900
rect 613562 93888 613568 93900
rect 607272 93860 613568 93888
rect 607272 93848 607278 93860
rect 613562 93848 613568 93860
rect 613620 93848 613626 93900
rect 649350 93848 649356 93900
rect 649408 93888 649414 93900
rect 656894 93888 656900 93900
rect 649408 93860 656900 93888
rect 649408 93848 649414 93860
rect 656894 93848 656900 93860
rect 656952 93848 656958 93900
rect 585134 89632 585140 89684
rect 585192 89672 585198 89684
rect 607214 89672 607220 89684
rect 585192 89644 607220 89672
rect 585192 89632 585198 89644
rect 607214 89632 607220 89644
rect 607272 89632 607278 89684
rect 657078 88816 657084 88868
rect 657136 88856 657142 88868
rect 657998 88856 658004 88868
rect 657136 88828 658004 88856
rect 657136 88816 657142 88828
rect 657998 88816 658004 88828
rect 658056 88816 658062 88868
rect 659470 88816 659476 88868
rect 659528 88856 659534 88868
rect 663610 88856 663616 88868
rect 659528 88828 663616 88856
rect 659528 88816 659534 88828
rect 663610 88816 663616 88828
rect 663668 88816 663674 88868
rect 582190 88340 582196 88392
rect 582248 88380 582254 88392
rect 588078 88380 588084 88392
rect 582248 88352 588084 88380
rect 582248 88340 582254 88352
rect 588078 88340 588084 88352
rect 588136 88340 588142 88392
rect 591942 85960 591948 86012
rect 592000 86000 592006 86012
rect 596174 86000 596180 86012
rect 592000 85972 596180 86000
rect 592000 85960 592006 85972
rect 596174 85960 596180 85972
rect 596232 85960 596238 86012
rect 648798 85484 648804 85536
rect 648856 85524 648862 85536
rect 657722 85524 657728 85536
rect 648856 85496 657728 85524
rect 648856 85484 648862 85496
rect 657722 85484 657728 85496
rect 657780 85484 657786 85536
rect 651834 85416 651840 85468
rect 651892 85456 651898 85468
rect 658826 85456 658832 85468
rect 651892 85428 658832 85456
rect 651892 85416 651898 85428
rect 658826 85416 658832 85428
rect 658884 85416 658890 85468
rect 648706 85348 648712 85400
rect 648764 85388 648770 85400
rect 660666 85388 660672 85400
rect 648764 85360 660672 85388
rect 648764 85348 648770 85360
rect 660666 85348 660672 85360
rect 660724 85348 660730 85400
rect 648614 85280 648620 85332
rect 648672 85320 648678 85332
rect 657170 85320 657176 85332
rect 648672 85292 657176 85320
rect 648672 85280 648678 85292
rect 657170 85280 657176 85292
rect 657228 85280 657234 85332
rect 643462 85212 643468 85264
rect 643520 85252 643526 85264
rect 660114 85252 660120 85264
rect 643520 85224 660120 85252
rect 643520 85212 643526 85224
rect 660114 85212 660120 85224
rect 660172 85212 660178 85264
rect 647510 85144 647516 85196
rect 647568 85184 647574 85196
rect 661402 85184 661408 85196
rect 647568 85156 661408 85184
rect 647568 85144 647574 85156
rect 661402 85144 661408 85156
rect 661460 85144 661466 85196
rect 583754 84396 583760 84448
rect 583812 84436 583818 84448
rect 600498 84436 600504 84448
rect 583812 84408 600504 84436
rect 583812 84396 583818 84408
rect 600498 84396 600504 84408
rect 600556 84396 600562 84448
rect 583846 84328 583852 84380
rect 583904 84368 583910 84380
rect 600682 84368 600688 84380
rect 583904 84340 600688 84368
rect 583904 84328 583910 84340
rect 600682 84328 600688 84340
rect 600740 84328 600746 84380
rect 580810 84260 580816 84312
rect 580868 84300 580874 84312
rect 600314 84300 600320 84312
rect 580868 84272 600320 84300
rect 580868 84260 580874 84272
rect 600314 84260 600320 84272
rect 600372 84260 600378 84312
rect 580718 84192 580724 84244
rect 580776 84232 580782 84244
rect 600222 84232 600228 84244
rect 580776 84204 600228 84232
rect 580776 84192 580782 84204
rect 600222 84192 600228 84204
rect 600280 84192 600286 84244
rect 580626 84124 580632 84176
rect 580684 84164 580690 84176
rect 600406 84164 600412 84176
rect 580684 84136 600412 84164
rect 580684 84124 580690 84136
rect 600406 84124 600412 84136
rect 600464 84124 600470 84176
rect 602982 82832 602988 82884
rect 603040 82872 603046 82884
rect 610158 82872 610164 82884
rect 603040 82844 610164 82872
rect 603040 82832 603046 82844
rect 610158 82832 610164 82844
rect 610216 82832 610222 82884
rect 579982 82764 579988 82816
rect 580040 82804 580046 82816
rect 586422 82804 586428 82816
rect 580040 82776 586428 82804
rect 580040 82764 580046 82776
rect 586422 82764 586428 82776
rect 586480 82764 586486 82816
rect 579614 82288 579620 82340
rect 579672 82328 579678 82340
rect 583662 82328 583668 82340
rect 579672 82300 583668 82328
rect 579672 82288 579678 82300
rect 583662 82288 583668 82300
rect 583720 82288 583726 82340
rect 604362 81268 604368 81320
rect 604420 81308 604426 81320
rect 631318 81308 631324 81320
rect 604420 81280 631324 81308
rect 604420 81268 604426 81280
rect 631318 81268 631324 81280
rect 631376 81268 631382 81320
rect 628558 81200 628564 81252
rect 628616 81240 628622 81252
rect 637022 81240 637028 81252
rect 628616 81212 637028 81240
rect 628616 81200 628622 81212
rect 637022 81200 637028 81212
rect 637080 81200 637086 81252
rect 575750 80112 575756 80164
rect 575808 80152 575814 80164
rect 585134 80152 585140 80164
rect 575808 80124 585140 80152
rect 575808 80112 575814 80124
rect 585134 80112 585140 80124
rect 585192 80112 585198 80164
rect 629202 80044 629208 80096
rect 629260 80084 629266 80096
rect 639874 80084 639880 80096
rect 629260 80056 639880 80084
rect 629260 80044 629266 80056
rect 639874 80044 639880 80056
rect 639932 80044 639938 80096
rect 615310 77188 615316 77240
rect 615368 77228 615374 77240
rect 640334 77228 640340 77240
rect 615368 77200 640340 77228
rect 615368 77188 615374 77200
rect 640334 77188 640340 77200
rect 640392 77188 640398 77240
rect 623682 75964 623688 76016
rect 623740 76004 623746 76016
rect 641070 76004 641076 76016
rect 623740 75976 641076 76004
rect 623740 75964 623746 75976
rect 641070 75964 641076 75976
rect 641128 75964 641134 76016
rect 623590 75828 623596 75880
rect 623648 75868 623654 75880
rect 640978 75868 640984 75880
rect 623648 75840 640984 75868
rect 623648 75828 623654 75840
rect 640978 75828 640984 75840
rect 641036 75828 641042 75880
rect 612734 75760 612740 75812
rect 612792 75800 612798 75812
rect 623084 75800 623090 75812
rect 612792 75772 623090 75800
rect 612792 75760 612798 75772
rect 623084 75760 623090 75772
rect 623142 75800 623148 75812
rect 631502 75800 631508 75812
rect 623142 75772 631508 75800
rect 623142 75760 623148 75772
rect 631502 75760 631508 75772
rect 631560 75760 631566 75812
rect 625614 74984 625620 74996
rect 593386 74956 625620 74984
rect 578142 74740 578148 74792
rect 578200 74780 578206 74792
rect 593386 74780 593414 74956
rect 625614 74944 625620 74956
rect 625672 74984 625678 74996
rect 638954 74984 638960 74996
rect 625672 74956 638960 74984
rect 625672 74944 625678 74956
rect 638954 74944 638960 74956
rect 639012 74944 639018 74996
rect 578200 74752 593414 74780
rect 578200 74740 578206 74752
rect 598934 66444 598940 66496
rect 598992 66484 598998 66496
rect 612734 66484 612740 66496
rect 598992 66456 612740 66484
rect 598992 66444 598998 66456
rect 612734 66444 612740 66456
rect 612792 66444 612798 66496
rect 579614 60392 579620 60444
rect 579672 60432 579678 60444
rect 583754 60432 583760 60444
rect 579672 60404 583760 60432
rect 579672 60392 579678 60404
rect 583754 60392 583760 60404
rect 583812 60392 583818 60444
rect 597462 58352 597468 58404
rect 597520 58392 597526 58404
rect 602982 58392 602988 58404
rect 597520 58364 602988 58392
rect 597520 58352 597526 58364
rect 602982 58352 602988 58364
rect 603040 58352 603046 58404
rect 579614 58284 579620 58336
rect 579672 58324 579678 58336
rect 583846 58324 583852 58336
rect 579672 58296 583852 58324
rect 579672 58284 579678 58296
rect 583846 58284 583852 58296
rect 583904 58284 583910 58336
rect 594794 57944 594800 57996
rect 594852 57984 594858 57996
rect 598934 57984 598940 57996
rect 594852 57956 598940 57984
rect 594852 57944 594858 57956
rect 598934 57944 598940 57956
rect 598992 57944 598998 57996
rect 52178 53864 52184 53916
rect 52236 53904 52242 53916
rect 582190 53904 582196 53916
rect 52236 53876 331168 53904
rect 52236 53864 52242 53876
rect 145392 53808 322934 53836
rect 145392 53632 145420 53808
rect 145374 53580 145380 53632
rect 145432 53580 145438 53632
rect 322906 53532 322934 53808
rect 331140 53668 331168 53876
rect 546466 53876 582196 53904
rect 342226 53808 516134 53836
rect 331140 53640 339448 53668
rect 339420 53612 339448 53640
rect 339402 53560 339408 53612
rect 339460 53560 339466 53612
rect 342226 53532 342254 53808
rect 516106 53768 516134 53808
rect 516106 53740 527174 53768
rect 527146 53632 527174 53740
rect 546466 53736 546494 53876
rect 582190 53864 582196 53876
rect 582248 53864 582254 53916
rect 594794 53836 594800 53848
rect 554746 53808 594800 53836
rect 554746 53768 554774 53808
rect 594794 53796 594800 53808
rect 594852 53796 594858 53848
rect 543752 53708 546494 53736
rect 546606 53740 554774 53768
rect 527146 53604 543518 53632
rect 322906 53504 342254 53532
rect 543490 53532 543518 53604
rect 543642 53560 543648 53612
rect 543700 53600 543706 53612
rect 543752 53600 543780 53708
rect 543700 53572 543780 53600
rect 543700 53560 543706 53572
rect 546606 53532 546634 53740
rect 543490 53504 546634 53532
rect 600038 52436 600044 52488
rect 600096 52476 600102 52488
rect 613010 52476 613016 52488
rect 600096 52448 613016 52476
rect 600096 52436 600102 52448
rect 613010 52436 613016 52448
rect 613068 52436 613074 52488
rect 52270 52368 52276 52420
rect 52328 52408 52334 52420
rect 149974 52408 149980 52420
rect 52328 52380 149980 52408
rect 52328 52368 52334 52380
rect 149974 52368 149980 52380
rect 150032 52368 150038 52420
rect 568574 51008 568580 51060
rect 568632 51048 568638 51060
rect 581178 51048 581184 51060
rect 568632 51020 581184 51048
rect 568632 51008 568638 51020
rect 581178 51008 581184 51020
rect 581236 51008 581242 51060
rect 150342 49648 150348 49700
rect 150400 49688 150406 49700
rect 184934 49688 184940 49700
rect 150400 49660 184940 49688
rect 150400 49648 150406 49660
rect 184934 49648 184940 49660
rect 184992 49648 184998 49700
rect 649994 49620 650000 49632
rect 632026 49592 650000 49620
rect 615402 49512 615408 49564
rect 615460 49552 615466 49564
rect 632026 49552 632054 49592
rect 649994 49580 650000 49592
rect 650052 49580 650058 49632
rect 615460 49524 632054 49552
rect 615460 49512 615466 49524
rect 478138 48424 478144 48476
rect 478196 48464 478202 48476
rect 526162 48464 526168 48476
rect 478196 48436 526168 48464
rect 478196 48424 478202 48436
rect 526162 48424 526168 48436
rect 526220 48424 526226 48476
rect 412634 48356 412640 48408
rect 412692 48396 412698 48408
rect 506382 48396 506388 48408
rect 412692 48368 506388 48396
rect 412692 48356 412698 48368
rect 506382 48356 506388 48368
rect 506440 48356 506446 48408
rect 281442 48288 281448 48340
rect 281500 48328 281506 48340
rect 507854 48328 507860 48340
rect 281500 48300 507860 48328
rect 281500 48288 281506 48300
rect 507854 48288 507860 48300
rect 507912 48288 507918 48340
rect 660960 47376 660988 47581
rect 661034 47376 661040 47388
rect 660960 47348 661040 47376
rect 661034 47336 661040 47348
rect 661092 47336 661098 47388
rect 658348 47243 658406 47249
rect 658348 47240 658360 47243
rect 657372 47212 658360 47240
rect 649994 46928 650000 46980
rect 650052 46968 650058 46980
rect 657372 46968 657400 47212
rect 658348 47209 658360 47212
rect 658394 47209 658406 47243
rect 658348 47203 658406 47209
rect 650052 46940 657400 46968
rect 650052 46928 650058 46940
rect 460658 45772 460664 45824
rect 460716 45812 460722 45824
rect 610342 45812 610348 45824
rect 460716 45784 610348 45812
rect 460716 45772 460722 45784
rect 610342 45772 610348 45784
rect 610400 45772 610406 45824
rect 367094 45704 367100 45756
rect 367152 45744 367158 45756
rect 607398 45744 607404 45756
rect 367152 45716 607404 45744
rect 367152 45704 367158 45716
rect 607398 45704 607404 45716
rect 607456 45704 607462 45756
rect 312814 45636 312820 45688
rect 312872 45676 312878 45688
rect 607582 45676 607588 45688
rect 312872 45648 607588 45676
rect 312872 45636 312878 45648
rect 607582 45636 607588 45648
rect 607640 45636 607646 45688
rect 85114 45568 85120 45620
rect 85172 45608 85178 45620
rect 475562 45608 475568 45620
rect 85172 45580 475568 45608
rect 85172 45568 85178 45580
rect 475562 45568 475568 45580
rect 475620 45568 475626 45620
rect 187326 45500 187332 45552
rect 187384 45540 187390 45552
rect 578142 45540 578148 45552
rect 187384 45512 578148 45540
rect 187384 45500 187390 45512
rect 578142 45500 578148 45512
rect 578200 45500 578206 45552
rect 312814 44180 312820 44192
rect 310440 44152 312820 44180
rect 310440 44124 310468 44152
rect 312814 44140 312820 44152
rect 312872 44140 312878 44192
rect 367094 44180 367100 44192
rect 365180 44152 367100 44180
rect 365180 44124 365208 44152
rect 367094 44140 367100 44152
rect 367152 44140 367158 44192
rect 310422 44072 310428 44124
rect 310480 44072 310486 44124
rect 365162 44072 365168 44124
rect 365220 44072 365226 44124
rect 390186 43120 390192 43172
rect 390244 43160 390250 43172
rect 575658 43160 575664 43172
rect 390244 43132 575664 43160
rect 390244 43120 390250 43132
rect 575658 43120 575664 43132
rect 575716 43120 575722 43172
rect 223574 43052 223580 43104
rect 223632 43092 223638 43104
rect 661454 43092 661460 43104
rect 223632 43064 661460 43092
rect 223632 43052 223638 43064
rect 661454 43052 661460 43064
rect 661512 43052 661518 43104
rect 475470 42616 475476 42628
rect 474490 42588 475476 42616
rect 475470 42576 475476 42588
rect 475528 42576 475534 42628
rect 513282 41964 513288 42016
rect 513340 42004 513346 42016
rect 518526 42004 518532 42016
rect 513340 41976 518532 42004
rect 513340 41964 513346 41976
rect 518526 41964 518532 41976
rect 518584 41964 518590 42016
rect 405826 41896 405832 41948
rect 405884 41936 405890 41948
rect 420638 41936 420644 41948
rect 405884 41908 420644 41936
rect 405884 41896 405890 41908
rect 420638 41896 420644 41908
rect 420696 41896 420702 41948
rect 514018 41896 514024 41948
rect 514076 41936 514082 41948
rect 514846 41936 514852 41948
rect 514076 41908 514852 41936
rect 514076 41896 514082 41908
rect 514846 41896 514852 41908
rect 514904 41896 514910 41948
rect 529658 41896 529664 41948
rect 529716 41936 529722 41948
rect 530486 41936 530492 41948
rect 529716 41908 530492 41936
rect 529716 41896 529722 41908
rect 530486 41896 530492 41908
rect 530544 41896 530550 41948
rect 420656 41772 430574 41800
rect 420656 41744 420684 41772
rect 420638 41692 420644 41744
rect 420696 41692 420702 41744
rect 430546 41460 430574 41772
rect 607490 41460 607496 41472
rect 430546 41432 607496 41460
rect 607490 41420 607496 41432
rect 607548 41420 607554 41472
rect 506382 41352 506388 41404
rect 506440 41392 506446 41404
rect 513282 41392 513288 41404
rect 506440 41364 513288 41392
rect 506440 41352 506446 41364
rect 513282 41352 513288 41364
rect 513340 41352 513346 41404
rect 530302 41352 530308 41404
rect 530360 41392 530366 41404
rect 610250 41392 610256 41404
rect 530360 41364 610256 41392
rect 530360 41352 530366 41364
rect 610250 41352 610256 41364
rect 610308 41352 610314 41404
rect 507854 41284 507860 41336
rect 507912 41324 507918 41336
rect 513190 41324 513196 41336
rect 507912 41296 513196 41324
rect 507912 41284 507918 41296
rect 513190 41284 513196 41296
rect 513248 41284 513254 41336
rect 530394 41284 530400 41336
rect 530452 41324 530458 41336
rect 575750 41324 575756 41336
rect 530452 41296 575756 41324
rect 530452 41284 530458 41296
rect 575750 41284 575756 41296
rect 575808 41284 575814 41336
rect 475562 38564 475568 38616
rect 475620 38604 475626 38616
rect 514018 38604 514024 38616
rect 475620 38576 514024 38604
rect 475620 38564 475626 38576
rect 514018 38564 514024 38576
rect 514076 38564 514082 38616
rect 530486 38564 530492 38616
rect 530544 38604 530550 38616
rect 542998 38604 543004 38616
rect 530544 38576 543004 38604
rect 530544 38564 530550 38576
rect 542998 38564 543004 38576
rect 543056 38564 543062 38616
<< via1 >>
rect 655428 896996 655480 897048
rect 676036 896996 676088 897048
rect 673368 894616 673420 894668
rect 675944 894616 675996 894668
rect 655612 894344 655664 894396
rect 676036 894344 676088 894396
rect 655520 894276 655572 894328
rect 676128 894276 676180 894328
rect 673276 892984 673328 893036
rect 676036 892984 676088 893036
rect 674748 891488 674800 891540
rect 676036 891488 676088 891540
rect 674932 890672 674984 890724
rect 676036 890672 676088 890724
rect 675024 889040 675076 889092
rect 676036 889040 676088 889092
rect 675208 888700 675260 888752
rect 676036 888700 676088 888752
rect 673736 887816 673788 887868
rect 676036 887816 676088 887868
rect 674288 887408 674340 887460
rect 676036 887408 676088 887460
rect 674196 885980 674248 886032
rect 676036 885980 676088 886032
rect 671988 884960 672040 885012
rect 678980 884960 679032 885012
rect 655704 883260 655756 883312
rect 675392 883260 675444 883312
rect 674472 880676 674524 880728
rect 675208 880676 675260 880728
rect 674840 880608 674892 880660
rect 680268 880608 680320 880660
rect 675208 880540 675260 880592
rect 679164 880540 679216 880592
rect 675300 880472 675352 880524
rect 679440 880472 679492 880524
rect 675116 878772 675168 878824
rect 679256 878772 679308 878824
rect 674564 878636 674616 878688
rect 679532 878636 679584 878688
rect 674656 878568 674708 878620
rect 679716 878568 679768 878620
rect 674932 878500 674984 878552
rect 679072 878500 679124 878552
rect 674840 877208 674892 877260
rect 675392 877208 675444 877260
rect 674380 875848 674432 875900
rect 674840 875848 674892 875900
rect 674656 874284 674708 874336
rect 675116 874284 675168 874336
rect 673736 874148 673788 874200
rect 674656 874148 674708 874200
rect 674564 873740 674616 873792
rect 675116 873740 675168 873792
rect 675024 872720 675076 872772
rect 675024 872516 675076 872568
rect 674748 872448 674800 872500
rect 675208 872448 675260 872500
rect 655796 872176 655848 872228
rect 675116 872176 675168 872228
rect 674288 869932 674340 869984
rect 675208 869932 675260 869984
rect 674196 869388 674248 869440
rect 675208 869388 675260 869440
rect 674656 869320 674708 869372
rect 675300 869320 675352 869372
rect 674472 867552 674524 867604
rect 675116 867552 675168 867604
rect 674748 865716 674800 865768
rect 675208 865716 675260 865768
rect 656808 863812 656860 863864
rect 675116 863812 675168 863864
rect 41788 817640 41840 817692
rect 50988 817640 51040 817692
rect 41788 817232 41840 817284
rect 48228 817232 48280 817284
rect 41788 816824 41840 816876
rect 45560 816824 45612 816876
rect 41788 815668 41840 815720
rect 43812 815668 43864 815720
rect 41788 814512 41840 814564
rect 43628 814512 43680 814564
rect 41788 814376 41840 814428
rect 43536 814376 43588 814428
rect 41788 813288 41840 813340
rect 43352 813288 43404 813340
rect 41788 812880 41840 812932
rect 42800 812880 42852 812932
rect 41788 812744 41840 812796
rect 42708 812744 42760 812796
rect 41788 811452 41840 811504
rect 43444 811452 43496 811504
rect 41788 810092 41840 810144
rect 43904 810092 43956 810144
rect 41880 808800 41932 808852
rect 44088 808800 44140 808852
rect 41788 808664 41840 808716
rect 43260 808664 43312 808716
rect 41788 807984 41840 808036
rect 43076 807984 43128 808036
rect 41788 806012 41840 806064
rect 42984 806012 43036 806064
rect 42064 805944 42116 805996
rect 45468 805944 45520 805996
rect 41880 803088 41932 803140
rect 42892 803088 42944 803140
rect 41972 803020 42024 803072
rect 43168 803020 43220 803072
rect 42340 800436 42392 800488
rect 58256 800436 58308 800488
rect 42340 798940 42392 798992
rect 42800 798940 42852 798992
rect 42156 798124 42208 798176
rect 42708 798124 42760 798176
rect 42708 797988 42760 798040
rect 43168 797988 43220 798040
rect 43536 797920 43588 797972
rect 43168 797852 43220 797904
rect 43352 797852 43404 797904
rect 43352 797716 43404 797768
rect 43720 797784 43772 797836
rect 43720 797648 43772 797700
rect 42340 796696 42392 796748
rect 43260 796696 43312 796748
rect 42248 795880 42300 795932
rect 43260 795880 43312 795932
rect 42248 794996 42300 795048
rect 42984 794996 43036 795048
rect 42248 794452 42300 794504
rect 42708 794452 42760 794504
rect 43628 794044 43680 794096
rect 43812 794044 43864 794096
rect 42156 793772 42208 793824
rect 43076 793772 43128 793824
rect 42340 792208 42392 792260
rect 42708 792208 42760 792260
rect 655520 792140 655572 792192
rect 675392 792140 675444 792192
rect 42156 790644 42208 790696
rect 42892 790644 42944 790696
rect 42248 789488 42300 789540
rect 43720 789488 43772 789540
rect 42432 789352 42484 789404
rect 58164 789352 58216 789404
rect 42708 789284 42760 789336
rect 58532 789284 58584 789336
rect 42156 789216 42208 789268
rect 44088 789216 44140 789268
rect 45560 789216 45612 789268
rect 58440 789216 58492 789268
rect 42340 789148 42392 789200
rect 43260 789148 43312 789200
rect 48228 786564 48280 786616
rect 58440 786564 58492 786616
rect 50988 786496 51040 786548
rect 58532 786496 58584 786548
rect 42340 786428 42392 786480
rect 43444 786428 43496 786480
rect 42064 786224 42116 786276
rect 43904 786224 43956 786276
rect 673828 784728 673880 784780
rect 675116 784728 675168 784780
rect 656532 783844 656584 783896
rect 675116 783844 675168 783896
rect 674564 780444 674616 780496
rect 675484 780444 675536 780496
rect 674288 779968 674340 780020
rect 675484 779968 675536 780020
rect 673644 779764 673696 779816
rect 675208 779764 675260 779816
rect 673736 778744 673788 778796
rect 675484 778744 675536 778796
rect 674472 778540 674524 778592
rect 675208 778540 675260 778592
rect 674656 777316 674708 777368
rect 675392 777316 675444 777368
rect 675024 776840 675076 776892
rect 675024 776636 675076 776688
rect 654968 775480 655020 775532
rect 675116 775480 675168 775532
rect 41788 774392 41840 774444
rect 50988 774392 51040 774444
rect 41512 774256 41564 774308
rect 43628 774256 43680 774308
rect 41420 773848 41472 773900
rect 48228 773848 48280 773900
rect 41788 773576 41840 773628
rect 45744 773576 45796 773628
rect 675024 773372 675076 773424
rect 675668 773372 675720 773424
rect 674748 773304 674800 773356
rect 675760 773304 675812 773356
rect 41880 772828 41932 772880
rect 44088 772828 44140 772880
rect 41788 772760 41840 772812
rect 43352 772760 43404 772812
rect 41512 772692 41564 772744
rect 43536 772692 43588 772744
rect 41788 771468 41840 771520
rect 43168 771468 43220 771520
rect 41420 770992 41472 771044
rect 43168 770992 43220 771044
rect 41512 770312 41564 770364
rect 42432 770312 42484 770364
rect 41512 769496 41564 769548
rect 43260 769496 43312 769548
rect 41512 769360 41564 769412
rect 43076 769360 43128 769412
rect 41512 768952 41564 769004
rect 43720 768952 43772 769004
rect 41512 768272 41564 768324
rect 43444 768272 43496 768324
rect 41512 768136 41564 768188
rect 43352 768136 43404 768188
rect 41512 767388 41564 767440
rect 43536 767388 43588 767440
rect 42708 767320 42760 767372
rect 45652 767320 45704 767372
rect 674656 767320 674708 767372
rect 674932 767320 674984 767372
rect 43536 766300 43588 766352
rect 43996 766300 44048 766352
rect 41512 766096 41564 766148
rect 42432 766096 42484 766148
rect 43352 765824 43404 765876
rect 43628 765824 43680 765876
rect 41512 765688 41564 765740
rect 43352 765688 43404 765740
rect 41512 764872 41564 764924
rect 43812 764872 43864 764924
rect 41512 764532 41564 764584
rect 42708 764532 42760 764584
rect 41512 762832 41564 762884
rect 45560 762832 45612 762884
rect 41788 761744 41840 761796
rect 42248 761744 42300 761796
rect 42340 760928 42392 760980
rect 43628 760928 43680 760980
rect 42340 760792 42392 760844
rect 43076 760792 43128 760844
rect 42432 760656 42484 760708
rect 43076 760656 43128 760708
rect 41604 759296 41656 759348
rect 43904 759296 43956 759348
rect 41420 759024 41472 759076
rect 44180 759024 44232 759076
rect 43352 757800 43404 757852
rect 43536 757664 43588 757716
rect 43168 757460 43220 757512
rect 43352 757460 43404 757512
rect 43444 757460 43496 757512
rect 674656 757596 674708 757648
rect 675300 757596 675352 757648
rect 43352 757324 43404 757376
rect 43720 757324 43772 757376
rect 43720 757188 43772 757240
rect 42248 756236 42300 756288
rect 59268 756236 59320 756288
rect 42156 754876 42208 754928
rect 42340 754876 42392 754928
rect 42340 754264 42392 754316
rect 42708 754264 42760 754316
rect 42156 753312 42208 753364
rect 42708 753312 42760 753364
rect 42156 753040 42208 753092
rect 43076 753040 43128 753092
rect 42340 751204 42392 751256
rect 43444 751204 43496 751256
rect 43536 751136 43588 751188
rect 43536 750932 43588 750984
rect 42064 750592 42116 750644
rect 43812 750592 43864 750644
rect 42340 750524 42392 750576
rect 43904 750524 43956 750576
rect 42248 750456 42300 750508
rect 43720 750456 43772 750508
rect 43812 750456 43864 750508
rect 44180 750456 44232 750508
rect 42708 750388 42760 750440
rect 43904 750388 43956 750440
rect 43076 750320 43128 750372
rect 43720 750320 43772 750372
rect 655980 747940 656032 747992
rect 675392 747940 675444 747992
rect 43904 747872 43956 747924
rect 58440 747872 58492 747924
rect 42340 746920 42392 746972
rect 43812 746920 43864 746972
rect 42248 745560 42300 745612
rect 43536 745560 43588 745612
rect 42340 745220 42392 745272
rect 58440 745220 58492 745272
rect 45744 745152 45796 745204
rect 58532 745152 58584 745204
rect 42248 745084 42300 745136
rect 43168 745084 43220 745136
rect 673460 744200 673512 744252
rect 675760 744200 675812 744252
rect 673552 744132 673604 744184
rect 675668 744132 675720 744184
rect 42248 743248 42300 743300
rect 43352 743248 43404 743300
rect 42156 743044 42208 743096
rect 43996 743044 44048 743096
rect 48228 742364 48280 742416
rect 58440 742364 58492 742416
rect 50988 742296 51040 742348
rect 57980 742296 58032 742348
rect 673736 738352 673788 738404
rect 674656 738352 674708 738404
rect 654324 736992 654376 737044
rect 675208 736992 675260 737044
rect 656072 736924 656124 736976
rect 675300 736924 675352 736976
rect 674748 735632 674800 735684
rect 675392 735632 675444 735684
rect 674840 734952 674892 735004
rect 675392 734952 675444 735004
rect 674288 734136 674340 734188
rect 675392 734136 675444 734188
rect 675300 733728 675352 733780
rect 675392 733728 675444 733780
rect 675300 733388 675352 733440
rect 675208 733320 675260 733372
rect 673276 732436 673328 732488
rect 673460 732436 673512 732488
rect 673460 732300 673512 732352
rect 675392 732300 675444 732352
rect 675208 732096 675260 732148
rect 674840 731960 674892 732012
rect 675208 731960 675260 732012
rect 674840 731824 674892 731876
rect 41512 731008 41564 731060
rect 50988 731008 51040 731060
rect 41788 730736 41840 730788
rect 43444 730736 43496 730788
rect 41512 730600 41564 730652
rect 48228 730600 48280 730652
rect 41880 730464 41932 730516
rect 44088 730464 44140 730516
rect 41512 730192 41564 730244
rect 45836 730192 45888 730244
rect 41512 729104 41564 729156
rect 43996 729104 44048 729156
rect 673552 728832 673604 728884
rect 673276 728764 673328 728816
rect 675208 728764 675260 728816
rect 674840 728628 674892 728680
rect 41512 728560 41564 728612
rect 43260 728560 43312 728612
rect 673460 728560 673512 728612
rect 673736 728560 673788 728612
rect 675392 728628 675444 728680
rect 674932 728492 674984 728544
rect 41512 727880 41564 727932
rect 43720 727880 43772 727932
rect 41512 726520 41564 726572
rect 43168 726520 43220 726572
rect 41788 726180 41840 726232
rect 43076 726180 43128 726232
rect 41512 726112 41564 726164
rect 43352 726112 43404 726164
rect 41788 725976 41840 726028
rect 43720 725976 43772 726028
rect 674472 724752 674524 724804
rect 675116 724752 675168 724804
rect 41512 724208 41564 724260
rect 43904 724208 43956 724260
rect 41788 723392 41840 723444
rect 44088 723392 44140 723444
rect 41512 723256 41564 723308
rect 43536 723256 43588 723308
rect 673184 723188 673236 723240
rect 679072 723188 679124 723240
rect 41788 723120 41840 723172
rect 42708 723120 42760 723172
rect 673368 723120 673420 723172
rect 678980 723120 679032 723172
rect 41512 722032 41564 722084
rect 43444 722032 43496 722084
rect 41604 720672 41656 720724
rect 43812 720672 43864 720724
rect 41512 720400 41564 720452
rect 43260 720400 43312 720452
rect 41512 719584 41564 719636
rect 45744 719584 45796 719636
rect 30288 716252 30340 716304
rect 43628 716252 43680 716304
rect 655796 715232 655848 715284
rect 675944 715232 675996 715284
rect 655612 715096 655664 715148
rect 676036 715096 676088 715148
rect 655428 714960 655480 715012
rect 675852 714960 675904 715012
rect 41696 714892 41748 714944
rect 44272 714892 44324 714944
rect 673276 714892 673328 714944
rect 676036 714892 676088 714944
rect 42340 714824 42392 714876
rect 59360 714824 59412 714876
rect 674656 714756 674708 714808
rect 676036 714756 676088 714808
rect 674564 714688 674616 714740
rect 675760 714688 675812 714740
rect 673828 714620 673880 714672
rect 675668 714620 675720 714672
rect 673460 714552 673512 714604
rect 676128 714552 676180 714604
rect 673184 714008 673236 714060
rect 675944 714008 675996 714060
rect 41972 713872 42024 713924
rect 44364 713872 44416 713924
rect 41880 713804 41932 713856
rect 673368 713192 673420 713244
rect 675944 713192 675996 713244
rect 42248 712920 42300 712972
rect 673092 712376 673144 712428
rect 675944 712376 675996 712428
rect 44088 712104 44140 712156
rect 59268 712104 59320 712156
rect 675116 712036 675168 712088
rect 675944 712036 675996 712088
rect 675024 711968 675076 712020
rect 675852 711968 675904 712020
rect 42156 711696 42208 711748
rect 43352 711696 43404 711748
rect 42156 710880 42208 710932
rect 42340 710880 42392 710932
rect 673552 710676 673604 710728
rect 674656 710676 674708 710728
rect 42340 710404 42392 710456
rect 42708 710404 42760 710456
rect 42708 710268 42760 710320
rect 43260 710268 43312 710320
rect 43260 710132 43312 710184
rect 43904 710132 43956 710184
rect 43904 709996 43956 710048
rect 44364 709996 44416 710048
rect 42248 709928 42300 709980
rect 42340 709724 42392 709776
rect 44088 709656 44140 709708
rect 42248 709384 42300 709436
rect 44088 709384 44140 709436
rect 43720 709316 43772 709368
rect 675208 709248 675260 709300
rect 676036 709248 676088 709300
rect 674840 709180 674892 709232
rect 675760 709180 675812 709232
rect 673644 708636 673696 708688
rect 676036 708636 676088 708688
rect 42156 708568 42208 708620
rect 43812 708568 43864 708620
rect 42156 708024 42208 708076
rect 42340 708024 42392 708076
rect 42156 707208 42208 707260
rect 42708 707208 42760 707260
rect 42156 706732 42208 706784
rect 43720 706732 43772 706784
rect 672080 705100 672132 705152
rect 676036 705100 676088 705152
rect 42064 704216 42116 704268
rect 43352 704216 43404 704268
rect 655980 703876 656032 703928
rect 675392 703876 675444 703928
rect 42340 703808 42392 703860
rect 58532 703808 58584 703860
rect 42156 703536 42208 703588
rect 44088 703536 44140 703588
rect 42064 703060 42116 703112
rect 43628 703060 43680 703112
rect 42064 702380 42116 702432
rect 43260 702380 43312 702432
rect 45836 700952 45888 701004
rect 58256 700952 58308 701004
rect 50988 700884 51040 700936
rect 58532 700884 58584 700936
rect 42156 700544 42208 700596
rect 43812 700544 43864 700596
rect 42156 700000 42208 700052
rect 43536 700000 43588 700052
rect 48228 698232 48280 698284
rect 58532 698232 58584 698284
rect 654232 692860 654284 692912
rect 675024 692860 675076 692912
rect 654140 690004 654192 690056
rect 675116 690004 675168 690056
rect 673828 689324 673880 689376
rect 675484 689324 675536 689376
rect 675024 688916 675076 688968
rect 675484 688916 675536 688968
rect 675024 688576 675076 688628
rect 675392 688576 675444 688628
rect 41788 688032 41840 688084
rect 50988 688032 51040 688084
rect 41788 687624 41840 687676
rect 48228 687624 48280 687676
rect 41788 687284 41840 687336
rect 45928 687284 45980 687336
rect 674564 687284 674616 687336
rect 675392 687284 675444 687336
rect 41788 687148 41840 687200
rect 43996 687148 44048 687200
rect 675116 687012 675168 687064
rect 675484 687012 675536 687064
rect 41788 686128 41840 686180
rect 43996 686128 44048 686180
rect 41788 685992 41840 686044
rect 43444 685992 43496 686044
rect 675116 685448 675168 685500
rect 675392 685448 675444 685500
rect 41788 684428 41840 684480
rect 43904 684428 43956 684480
rect 41788 683680 41840 683732
rect 43536 683680 43588 683732
rect 675024 683612 675076 683664
rect 675392 683612 675444 683664
rect 41696 682456 41748 682508
rect 43628 682456 43680 682508
rect 41696 682184 41748 682236
rect 43720 682184 43772 682236
rect 41788 681708 41840 681760
rect 43444 681708 43496 681760
rect 673276 681436 673328 681488
rect 679164 681436 679216 681488
rect 673092 680824 673144 680876
rect 679256 680824 679308 680876
rect 673184 680756 673236 680808
rect 679072 680756 679124 680808
rect 41788 680008 41840 680060
rect 43904 680008 43956 680060
rect 41788 679872 41840 679924
rect 43812 679872 43864 679924
rect 41696 679328 41748 679380
rect 44088 679328 44140 679380
rect 41696 676608 41748 676660
rect 43352 676608 43404 676660
rect 41696 676472 41748 676524
rect 45836 676472 45888 676524
rect 41788 676200 41840 676252
rect 42708 676200 42760 676252
rect 674564 673820 674616 673872
rect 674932 673820 674984 673872
rect 30288 672188 30340 672240
rect 43076 672188 43128 672240
rect 27528 672120 27580 672172
rect 43168 672120 43220 672172
rect 27436 672052 27488 672104
rect 43260 672052 43312 672104
rect 655888 670896 655940 670948
rect 676220 670896 676272 670948
rect 42432 670828 42484 670880
rect 60648 670828 60700 670880
rect 655520 670760 655572 670812
rect 676036 670760 676088 670812
rect 42064 670692 42116 670744
rect 43536 670692 43588 670744
rect 43168 670624 43220 670676
rect 43720 670624 43772 670676
rect 44272 670624 44324 670676
rect 43628 670556 43680 670608
rect 43904 670488 43956 670540
rect 44364 670488 44416 670540
rect 42708 670352 42760 670404
rect 43076 670352 43128 670404
rect 42432 670216 42484 670268
rect 42708 670216 42760 670268
rect 42248 669944 42300 669996
rect 42340 669740 42392 669792
rect 673552 668992 673604 669044
rect 676036 668992 676088 669044
rect 673368 668652 673420 668704
rect 676220 668652 676272 668704
rect 655704 668040 655756 668092
rect 678980 668040 679032 668092
rect 674932 667972 674984 668024
rect 676036 667972 676088 668024
rect 42340 667904 42392 667956
rect 42708 667904 42760 667956
rect 674748 667836 674800 667888
rect 676036 667836 676088 667888
rect 42708 667768 42760 667820
rect 44180 667768 44232 667820
rect 42340 667224 42392 667276
rect 43812 667224 43864 667276
rect 43812 667088 43864 667140
rect 44272 667088 44324 667140
rect 42248 665388 42300 665440
rect 43076 665388 43128 665440
rect 42156 665184 42208 665236
rect 43352 665184 43404 665236
rect 675208 665116 675260 665168
rect 676036 665116 676088 665168
rect 43352 665048 43404 665100
rect 44364 665048 44416 665100
rect 674656 664708 674708 664760
rect 676036 664708 676088 664760
rect 42156 664640 42208 664692
rect 42708 664640 42760 664692
rect 42248 663552 42300 663604
rect 43168 663552 43220 663604
rect 674288 663076 674340 663128
rect 676036 663076 676088 663128
rect 42248 663008 42300 663060
rect 43720 663008 43772 663060
rect 673736 662328 673788 662380
rect 676036 662328 676088 662380
rect 42156 661036 42208 661088
rect 43628 661036 43680 661088
rect 42432 659676 42484 659728
rect 58440 659676 58492 659728
rect 672172 659676 672224 659728
rect 678980 659676 679032 659728
rect 42340 659608 42392 659660
rect 58532 659608 58584 659660
rect 45928 659540 45980 659592
rect 58624 659540 58676 659592
rect 42340 659472 42392 659524
rect 43260 659472 43312 659524
rect 42340 659200 42392 659252
rect 43352 659200 43404 659252
rect 42156 658996 42208 659048
rect 43812 658996 43864 659048
rect 42156 657364 42208 657416
rect 43904 657364 43956 657416
rect 655704 656888 655756 656940
rect 675392 656888 675444 656940
rect 48228 656820 48280 656872
rect 58072 656820 58124 656872
rect 50988 656752 51040 656804
rect 58440 656752 58492 656804
rect 42156 656140 42208 656192
rect 43076 656140 43128 656192
rect 674656 649544 674708 649596
rect 675392 649544 675444 649596
rect 654416 648592 654468 648644
rect 674748 648592 674800 648644
rect 674288 647844 674340 647896
rect 674932 647844 674984 647896
rect 674932 647708 674984 647760
rect 675392 647708 675444 647760
rect 673460 646144 673512 646196
rect 675208 646144 675260 646196
rect 656440 645872 656492 645924
rect 675300 645872 675352 645924
rect 673736 645192 673788 645244
rect 675392 645192 675444 645244
rect 41512 644648 41564 644700
rect 50988 644648 51040 644700
rect 673644 644580 673696 644632
rect 675392 644580 675444 644632
rect 41512 644240 41564 644292
rect 48228 644240 48280 644292
rect 673184 644240 673236 644292
rect 673552 644240 673604 644292
rect 673552 644104 673604 644156
rect 675392 644104 675444 644156
rect 41788 644036 41840 644088
rect 46020 644036 46072 644088
rect 41512 643968 41564 644020
rect 43996 643968 44048 644020
rect 675208 643900 675260 643952
rect 675300 643832 675352 643884
rect 674748 643492 674800 643544
rect 674748 643356 674800 643408
rect 675300 643424 675352 643476
rect 675392 643356 675444 643408
rect 41788 643220 41840 643272
rect 43812 643220 43864 643272
rect 41512 643016 41564 643068
rect 43536 643016 43588 643068
rect 41512 642812 41564 642864
rect 43444 642812 43496 642864
rect 41788 642676 41840 642728
rect 44088 642676 44140 642728
rect 673276 642200 673328 642252
rect 674288 642200 674340 642252
rect 674288 642064 674340 642116
rect 675392 642064 675444 642116
rect 41512 640568 41564 640620
rect 43720 640568 43772 640620
rect 41788 640500 41840 640552
rect 43260 640500 43312 640552
rect 41788 640364 41840 640416
rect 42708 640364 42760 640416
rect 41604 640296 41656 640348
rect 43352 640296 43404 640348
rect 41512 639072 41564 639124
rect 43628 639072 43680 639124
rect 674748 639208 674800 639260
rect 674748 639072 674800 639124
rect 675300 639072 675352 639124
rect 41788 638460 41840 638512
rect 43444 638460 43496 638512
rect 675300 638664 675352 638716
rect 675300 638392 675352 638444
rect 674840 638188 674892 638240
rect 674932 638188 674984 638240
rect 675576 638188 675628 638240
rect 674656 638120 674708 638172
rect 675484 638120 675536 638172
rect 41512 637984 41564 638036
rect 43168 637984 43220 638036
rect 673736 637984 673788 638036
rect 674656 637984 674708 638036
rect 41512 637712 41564 637764
rect 43076 637712 43128 637764
rect 674840 637508 674892 637560
rect 679256 637508 679308 637560
rect 673368 637440 673420 637492
rect 679348 637440 679400 637492
rect 673276 637372 673328 637424
rect 679164 637372 679216 637424
rect 673184 637304 673236 637356
rect 679072 637304 679124 637356
rect 41604 635400 41656 635452
rect 43904 635400 43956 635452
rect 675116 635400 675168 635452
rect 41604 635128 41656 635180
rect 44088 635128 44140 635180
rect 675116 635060 675168 635112
rect 41512 634856 41564 634908
rect 43536 634856 43588 634908
rect 41604 634788 41656 634840
rect 43996 634788 44048 634840
rect 41512 633224 41564 633276
rect 45928 633224 45980 633276
rect 43168 632000 43220 632052
rect 43076 631932 43128 631984
rect 38108 631864 38160 631916
rect 43168 631864 43220 631916
rect 38200 631796 38252 631848
rect 43076 631796 43128 631848
rect 43996 631796 44048 631848
rect 44088 631728 44140 631780
rect 42432 629688 42484 629740
rect 43904 629688 43956 629740
rect 43444 629552 43496 629604
rect 43904 629552 43956 629604
rect 41880 629416 41932 629468
rect 43444 629416 43496 629468
rect 42248 626696 42300 626748
rect 42708 626696 42760 626748
rect 42708 626560 42760 626612
rect 58532 626560 58584 626612
rect 42156 625268 42208 625320
rect 42340 625268 42392 625320
rect 42340 624452 42392 624504
rect 42708 624452 42760 624504
rect 42248 624248 42300 624300
rect 42708 624248 42760 624300
rect 655796 624112 655848 624164
rect 676220 624112 676272 624164
rect 655612 623976 655664 624028
rect 678980 623976 679032 624028
rect 673368 623908 673420 623960
rect 676036 623908 676088 623960
rect 655428 623840 655480 623892
rect 676128 623840 676180 623892
rect 675116 623704 675168 623756
rect 676036 623704 676088 623756
rect 42156 623432 42208 623484
rect 43536 623432 43588 623484
rect 43536 623296 43588 623348
rect 44180 623296 44232 623348
rect 42156 622820 42208 622872
rect 42340 622820 42392 622872
rect 673276 621936 673328 621988
rect 676220 621936 676272 621988
rect 673460 621324 673512 621376
rect 676036 621324 676088 621376
rect 674840 620916 674892 620968
rect 676036 620916 676088 620968
rect 42064 620780 42116 620832
rect 43536 620780 43588 620832
rect 42064 620304 42116 620356
rect 43904 620304 43956 620356
rect 42432 619148 42484 619200
rect 43076 619148 43128 619200
rect 42340 618196 42392 618248
rect 58164 618196 58216 618248
rect 674472 618196 674524 618248
rect 676036 618196 676088 618248
rect 673828 618128 673880 618180
rect 676128 618128 676180 618180
rect 674564 618060 674616 618112
rect 676036 618060 676088 618112
rect 42432 617312 42484 617364
rect 43168 617312 43220 617364
rect 42432 616700 42484 616752
rect 43444 616700 43496 616752
rect 42432 616020 42484 616072
rect 43996 616020 44048 616072
rect 42340 615476 42392 615528
rect 58532 615476 58584 615528
rect 46020 615408 46072 615460
rect 58164 615408 58216 615460
rect 672264 614592 672316 614644
rect 678980 614592 679032 614644
rect 42156 614184 42208 614236
rect 42708 614184 42760 614236
rect 42248 614048 42300 614100
rect 43628 614048 43680 614100
rect 42156 613436 42208 613488
rect 44088 613436 44140 613488
rect 655428 612824 655480 612876
rect 675668 612824 675720 612876
rect 48228 612688 48280 612740
rect 58348 612688 58400 612740
rect 50988 612620 51040 612672
rect 58532 612620 58584 612672
rect 674564 609084 674616 609136
rect 675760 609084 675812 609136
rect 673736 609016 673788 609068
rect 675484 609016 675536 609068
rect 674472 608948 674524 609000
rect 675576 608948 675628 609000
rect 673828 606908 673880 606960
rect 675300 606908 675352 606960
rect 655244 601740 655296 601792
rect 675116 601740 675168 601792
rect 41788 601672 41840 601724
rect 50988 601672 51040 601724
rect 655612 601672 655664 601724
rect 675024 601672 675076 601724
rect 41788 601264 41840 601316
rect 48228 601264 48280 601316
rect 41512 600992 41564 601044
rect 43812 600992 43864 601044
rect 41788 600856 41840 600908
rect 46112 600856 46164 600908
rect 41512 600312 41564 600364
rect 43352 600312 43404 600364
rect 673552 599768 673604 599820
rect 675484 599768 675536 599820
rect 41788 599020 41840 599072
rect 43996 599020 44048 599072
rect 41512 598952 41564 599004
rect 43352 598952 43404 599004
rect 41788 598884 41840 598936
rect 43260 598884 43312 598936
rect 675116 598680 675168 598732
rect 675392 598680 675444 598732
rect 673460 598544 673512 598596
rect 675484 598544 675536 598596
rect 41512 598476 41564 598528
rect 43720 598476 43772 598528
rect 674564 598476 674616 598528
rect 675116 598476 675168 598528
rect 674564 598340 674616 598392
rect 675300 598340 675352 598392
rect 675024 598068 675076 598120
rect 675300 598068 675352 598120
rect 673184 597252 673236 597304
rect 673828 597252 673880 597304
rect 673828 597116 673880 597168
rect 675392 597116 675444 597168
rect 41512 597048 41564 597100
rect 44088 597048 44140 597100
rect 675116 597048 675168 597100
rect 675208 596844 675260 596896
rect 41512 596640 41564 596692
rect 43812 596640 43864 596692
rect 41512 596368 41564 596420
rect 43628 596368 43680 596420
rect 674472 596300 674524 596352
rect 675300 596300 675352 596352
rect 41512 595416 41564 595468
rect 43444 595416 43496 595468
rect 674472 595280 674524 595332
rect 675392 595280 675444 595332
rect 41512 594600 41564 594652
rect 43536 594600 43588 594652
rect 41512 594056 41564 594108
rect 43168 594056 43220 594108
rect 41788 593512 41840 593564
rect 43076 593512 43128 593564
rect 673552 593512 673604 593564
rect 673736 593444 673788 593496
rect 673184 593376 673236 593428
rect 673552 593376 673604 593428
rect 675668 593376 675720 593428
rect 675208 593172 675260 593224
rect 41512 592152 41564 592204
rect 43720 592152 43772 592204
rect 42340 591880 42392 591932
rect 43536 591880 43588 591932
rect 41512 591744 41564 591796
rect 43536 591744 43588 591796
rect 41512 591200 41564 591252
rect 43260 591200 43312 591252
rect 41512 589976 41564 590028
rect 46020 589976 46072 590028
rect 42156 588480 42208 588532
rect 43904 588480 43956 588532
rect 673276 587936 673328 587988
rect 679072 587936 679124 587988
rect 673368 587868 673420 587920
rect 678980 587868 679032 587920
rect 38016 587800 38068 587852
rect 42708 587800 42760 587852
rect 38108 587732 38160 587784
rect 41420 587732 41472 587784
rect 41420 585216 41472 585268
rect 44180 585216 44232 585268
rect 42340 585148 42392 585200
rect 58532 585148 58584 585200
rect 42432 584196 42484 584248
rect 43904 583856 43956 583908
rect 42708 583720 42760 583772
rect 43168 583720 43220 583772
rect 674472 583856 674524 583908
rect 673460 583720 673512 583772
rect 674472 583720 674524 583772
rect 44088 583652 44140 583704
rect 675392 583652 675444 583704
rect 43168 583584 43220 583636
rect 42248 582564 42300 582616
rect 59268 582564 59320 582616
rect 673552 582292 673604 582344
rect 676036 582292 676088 582344
rect 42156 582088 42208 582140
rect 43628 582088 43680 582140
rect 43168 581952 43220 582004
rect 43628 581952 43680 582004
rect 42248 581272 42300 581324
rect 42248 581068 42300 581120
rect 42156 580252 42208 580304
rect 43076 580252 43128 580304
rect 43076 580116 43128 580168
rect 43812 580116 43864 580168
rect 656072 580048 656124 580100
rect 676220 580048 676272 580100
rect 655888 579912 655940 579964
rect 676128 579912 676180 579964
rect 655520 579776 655572 579828
rect 676312 579776 676364 579828
rect 42248 578960 42300 579012
rect 43536 578960 43588 579012
rect 43536 578824 43588 578876
rect 44088 578824 44140 578876
rect 42156 578756 42208 578808
rect 43260 578756 43312 578808
rect 42156 578416 42208 578468
rect 43720 578416 43772 578468
rect 674840 576920 674892 576972
rect 676036 576920 676088 576972
rect 675116 576784 675168 576836
rect 676036 576784 676088 576836
rect 674748 576716 674800 576768
rect 675944 576716 675996 576768
rect 673828 576648 673880 576700
rect 675116 576648 675168 576700
rect 674656 575220 674708 575272
rect 676036 575220 676088 575272
rect 674932 574812 674984 574864
rect 676036 574812 676088 574864
rect 42340 574132 42392 574184
rect 43168 574132 43220 574184
rect 42432 574064 42484 574116
rect 60648 574064 60700 574116
rect 42156 573792 42208 573844
rect 44088 573792 44140 573844
rect 674288 573588 674340 573640
rect 676036 573588 676088 573640
rect 673644 572772 673696 572824
rect 676036 572772 676088 572824
rect 42064 572636 42116 572688
rect 43444 572636 43496 572688
rect 42248 571956 42300 572008
rect 42708 571956 42760 572008
rect 46112 571276 46164 571328
rect 58072 571276 58124 571328
rect 50988 571208 51040 571260
rect 58348 571208 58400 571260
rect 42064 570936 42116 570988
rect 43076 570936 43128 570988
rect 42064 569576 42116 569628
rect 43536 569576 43588 569628
rect 674288 568760 674340 568812
rect 675392 568760 675444 568812
rect 655888 568624 655940 568676
rect 675392 568624 675444 568676
rect 672356 568556 672408 568608
rect 678980 568556 679032 568608
rect 48228 568488 48280 568540
rect 58256 568488 58308 568540
rect 673644 559512 673696 559564
rect 675484 559512 675536 559564
rect 41512 558288 41564 558340
rect 50988 558288 51040 558340
rect 673460 558220 673512 558272
rect 675392 558220 675444 558272
rect 41512 557880 41564 557932
rect 48320 557880 48372 557932
rect 41512 557540 41564 557592
rect 46112 557540 46164 557592
rect 654232 557540 654284 557592
rect 674748 557540 674800 557592
rect 673552 557472 673604 557524
rect 675392 557472 675444 557524
rect 41788 557268 41840 557320
rect 43996 557268 44048 557320
rect 41788 556792 41840 556844
rect 43352 556792 43404 556844
rect 41512 556656 41564 556708
rect 43628 556656 43680 556708
rect 674656 555024 674708 555076
rect 675392 555024 675444 555076
rect 673828 554888 673880 554940
rect 675300 554888 675352 554940
rect 38568 554752 38620 554804
rect 43904 554752 43956 554804
rect 654140 554752 654192 554804
rect 675300 554752 675352 554804
rect 674288 553732 674340 553784
rect 675392 553732 675444 553784
rect 673368 553528 673420 553580
rect 673644 553528 673696 553580
rect 674748 553460 674800 553512
rect 675392 553460 675444 553512
rect 673644 553392 673696 553444
rect 675484 553392 675536 553444
rect 41512 552304 41564 552356
rect 43260 552304 43312 552356
rect 674748 551896 674800 551948
rect 675392 551896 675444 551948
rect 41420 549720 41472 549772
rect 43352 549720 43404 549772
rect 41512 549584 41564 549636
rect 43076 549584 43128 549636
rect 41512 549312 41564 549364
rect 43444 549312 43496 549364
rect 41512 548632 41564 548684
rect 43904 548632 43956 548684
rect 675668 548224 675720 548276
rect 674656 547952 674708 548004
rect 674840 547952 674892 548004
rect 675300 547884 675352 547936
rect 674288 547816 674340 547868
rect 674656 547816 674708 547868
rect 673736 547680 673788 547732
rect 673828 547680 673880 547732
rect 674288 547680 674340 547732
rect 673736 547476 673788 547528
rect 41512 547000 41564 547052
rect 43168 547000 43220 547052
rect 41512 546864 41564 546916
rect 48228 546864 48280 546916
rect 674932 543736 674984 543788
rect 679348 543736 679400 543788
rect 43168 541288 43220 541340
rect 43352 541288 43404 541340
rect 43076 541016 43128 541068
rect 59268 541016 59320 541068
rect 42708 540948 42760 541000
rect 59452 540948 59504 541000
rect 674288 539452 674340 539504
rect 675576 539452 675628 539504
rect 42064 538908 42116 538960
rect 43260 538908 43312 538960
rect 42248 538432 42300 538484
rect 43076 538432 43128 538484
rect 42156 538228 42208 538280
rect 42708 538228 42760 538280
rect 42064 537072 42116 537124
rect 43168 537072 43220 537124
rect 673460 537072 673512 537124
rect 674288 537072 674340 537124
rect 673460 536732 673512 536784
rect 673644 536732 673696 536784
rect 674840 536732 674892 536784
rect 675300 536732 675352 536784
rect 673460 536596 673512 536648
rect 675392 536596 675444 536648
rect 655980 535712 656032 535764
rect 676036 535712 676088 535764
rect 42156 535576 42208 535628
rect 43352 535576 43404 535628
rect 655704 535576 655756 535628
rect 676220 535576 676272 535628
rect 42064 535032 42116 535084
rect 43444 535032 43496 535084
rect 42156 534420 42208 534472
rect 43904 534420 43956 534472
rect 42156 533944 42208 533996
rect 43076 533944 43128 533996
rect 655796 532856 655848 532908
rect 679164 532856 679216 532908
rect 675024 532652 675076 532704
rect 676036 532652 676088 532704
rect 42156 531428 42208 531480
rect 43536 531428 43588 531480
rect 42156 530884 42208 530936
rect 42708 530884 42760 530936
rect 42432 530068 42484 530120
rect 42248 529592 42300 529644
rect 42432 529932 42484 529984
rect 58532 529932 58584 529984
rect 46112 529864 46164 529916
rect 58348 529864 58400 529916
rect 675208 529864 675260 529916
rect 676036 529864 676088 529916
rect 675116 529456 675168 529508
rect 676036 529456 676088 529508
rect 674564 527824 674616 527876
rect 676036 527824 676088 527876
rect 42156 527756 42208 527808
rect 43168 527756 43220 527808
rect 48320 527076 48372 527128
rect 58072 527076 58124 527128
rect 674472 527076 674524 527128
rect 676036 527076 676088 527128
rect 50988 527008 51040 527060
rect 57980 527008 58032 527060
rect 673736 527008 673788 527060
rect 675944 527008 675996 527060
rect 42340 526600 42392 526652
rect 43076 526600 43128 526652
rect 672448 524424 672500 524476
rect 679072 524424 679124 524476
rect 676128 521568 676180 521620
rect 678980 521568 679032 521620
rect 677396 521500 677448 521552
rect 679164 521500 679216 521552
rect 677304 521432 677356 521484
rect 679348 521432 679400 521484
rect 677488 521364 677540 521416
rect 679256 521364 679308 521416
rect 655612 491648 655664 491700
rect 676036 491648 676088 491700
rect 655520 491512 655572 491564
rect 676036 491512 676088 491564
rect 655428 491376 655480 491428
rect 675944 491376 675996 491428
rect 676220 491240 676272 491292
rect 677304 491240 677356 491292
rect 676220 490764 676272 490816
rect 677488 490764 677540 490816
rect 676220 489948 676272 490000
rect 677396 489948 677448 490000
rect 676036 489336 676088 489388
rect 676128 489132 676180 489184
rect 674932 488452 674984 488504
rect 676036 488452 676088 488504
rect 674288 488384 674340 488436
rect 675852 488384 675904 488436
rect 673460 488316 673512 488368
rect 675484 488316 675536 488368
rect 674840 485732 674892 485784
rect 676036 485732 676088 485784
rect 673644 485664 673696 485716
rect 675852 485664 675904 485716
rect 674748 485460 674800 485512
rect 676036 485460 676088 485512
rect 674656 483828 674708 483880
rect 676036 483828 676088 483880
rect 673552 483420 673604 483472
rect 676036 483420 676088 483472
rect 673828 482944 673880 482996
rect 676036 482944 676088 482996
rect 672540 480700 672592 480752
rect 676036 480700 676088 480752
rect 41788 430856 41840 430908
rect 50988 430856 51040 430908
rect 41788 430448 41840 430500
rect 48412 430448 48464 430500
rect 41788 430040 41840 430092
rect 46112 430040 46164 430092
rect 41788 429904 41840 429956
rect 43352 429904 43404 429956
rect 41788 429020 41840 429072
rect 43904 429020 43956 429072
rect 41788 428884 41840 428936
rect 43720 428884 43772 428936
rect 41788 426504 41840 426556
rect 43720 426504 43772 426556
rect 41788 426368 41840 426420
rect 43812 426368 43864 426420
rect 41788 425416 41840 425468
rect 42708 425416 42760 425468
rect 41788 425144 41840 425196
rect 43260 425144 43312 425196
rect 41880 423648 41932 423700
rect 43536 423648 43588 423700
rect 41880 423512 41932 423564
rect 43076 423512 43128 423564
rect 41880 422900 41932 422952
rect 43628 422900 43680 422952
rect 41880 422628 41932 422680
rect 43444 422628 43496 422680
rect 41788 422424 41840 422476
rect 43996 422424 44048 422476
rect 41788 422288 41840 422340
rect 44088 422288 44140 422340
rect 41788 421540 41840 421592
rect 43352 421540 43404 421592
rect 41788 419432 41840 419484
rect 48320 419432 48372 419484
rect 41880 416304 41932 416356
rect 43168 416304 43220 416356
rect 43996 413924 44048 413976
rect 44272 413924 44324 413976
rect 44088 413856 44140 413908
rect 44180 413856 44232 413908
rect 42064 413788 42116 413840
rect 43996 413788 44048 413840
rect 42432 413720 42484 413772
rect 44088 413720 44140 413772
rect 41972 413380 42024 413432
rect 42248 412972 42300 413024
rect 43260 411272 43312 411324
rect 43904 411272 43956 411324
rect 43904 411136 43956 411188
rect 44180 411136 44232 411188
rect 42156 409708 42208 409760
rect 42340 409708 42392 409760
rect 42156 409436 42208 409488
rect 43444 409436 43496 409488
rect 43076 409300 43128 409352
rect 43444 409300 43496 409352
rect 42156 407872 42208 407924
rect 43076 407872 43128 407924
rect 42248 407532 42300 407584
rect 43904 407532 43956 407584
rect 42064 406988 42116 407040
rect 43168 406988 43220 407040
rect 42248 406920 42300 406972
rect 44272 406920 44324 406972
rect 42340 405628 42392 405680
rect 58440 405628 58492 405680
rect 42340 405492 42392 405544
rect 43352 405492 43404 405544
rect 42432 405152 42484 405204
rect 42708 405152 42760 405204
rect 42340 403316 42392 403368
rect 43628 403316 43680 403368
rect 655704 403112 655756 403164
rect 676128 403112 676180 403164
rect 655520 403044 655572 403096
rect 676220 403044 676272 403096
rect 655428 402976 655480 403028
rect 676128 402976 676180 403028
rect 43076 402908 43128 402960
rect 58532 402908 58584 402960
rect 42248 402568 42300 402620
rect 43536 402568 43588 402620
rect 42156 402500 42208 402552
rect 43444 402500 43496 402552
rect 42156 401820 42208 401872
rect 43168 401820 43220 401872
rect 42156 400188 42208 400240
rect 43812 400188 43864 400240
rect 46112 400120 46164 400172
rect 58440 400120 58492 400172
rect 48412 400052 48464 400104
rect 58348 400052 58400 400104
rect 50988 399984 51040 400036
rect 58532 399984 58584 400036
rect 674288 399440 674340 399492
rect 676036 399440 676088 399492
rect 674564 398216 674616 398268
rect 676036 398216 676088 398268
rect 675024 397604 675076 397656
rect 675944 397604 675996 397656
rect 673644 397536 673696 397588
rect 676128 397536 676180 397588
rect 674656 397468 674708 397520
rect 676036 397468 676088 397520
rect 674472 396992 674524 397044
rect 676036 396992 676088 397044
rect 673460 395360 673512 395412
rect 675668 395360 675720 395412
rect 674748 394952 674800 395004
rect 675944 394952 675996 395004
rect 673552 394884 673604 394936
rect 675668 394884 675720 394936
rect 674840 394816 674892 394868
rect 676128 394816 676180 394868
rect 675116 394748 675168 394800
rect 675944 394748 675996 394800
rect 675208 394680 675260 394732
rect 676036 394680 676088 394732
rect 42156 394612 42208 394664
rect 60372 394612 60424 394664
rect 673736 394136 673788 394188
rect 676036 394136 676088 394188
rect 672632 392028 672684 392080
rect 678980 392028 679032 392080
rect 673828 391960 673880 392012
rect 676036 391960 676088 392012
rect 674932 390532 674984 390584
rect 675760 390532 675812 390584
rect 41512 388016 41564 388068
rect 43260 388016 43312 388068
rect 41420 387472 41472 387524
rect 50988 387472 51040 387524
rect 41420 387064 41472 387116
rect 48504 387064 48556 387116
rect 41788 386792 41840 386844
rect 46112 386792 46164 386844
rect 675760 386588 675812 386640
rect 41788 386316 41840 386368
rect 43720 386316 43772 386368
rect 675024 386112 675076 386164
rect 41512 386044 41564 386096
rect 44088 386044 44140 386096
rect 41512 385772 41564 385824
rect 43996 385772 44048 385824
rect 675024 385976 675076 386028
rect 675392 385976 675444 386028
rect 675760 385976 675812 386028
rect 675208 385568 675260 385620
rect 675392 385568 675444 385620
rect 674288 384956 674340 385008
rect 675208 384956 675260 385008
rect 674288 384820 674340 384872
rect 674564 384752 674616 384804
rect 675392 384752 675444 384804
rect 41880 383732 41932 383784
rect 44088 383732 44140 383784
rect 41512 383664 41564 383716
rect 43812 383664 43864 383716
rect 674656 383120 674708 383172
rect 675392 383120 675444 383172
rect 41512 382712 41564 382764
rect 43720 382712 43772 382764
rect 674840 382440 674892 382492
rect 675392 382440 675444 382492
rect 41512 381896 41564 381948
rect 42708 381896 42760 381948
rect 674748 381896 674800 381948
rect 675392 381896 675444 381948
rect 41512 381760 41564 381812
rect 43076 381760 43128 381812
rect 41512 381216 41564 381268
rect 43628 381216 43680 381268
rect 675116 381216 675168 381268
rect 674932 381080 674984 381132
rect 675116 381080 675168 381132
rect 675392 381080 675444 381132
rect 673644 381012 673696 381064
rect 673644 380876 673696 380928
rect 674288 380876 674340 380928
rect 674472 380876 674524 380928
rect 41512 380128 41564 380180
rect 43628 380128 43680 380180
rect 41512 379448 41564 379500
rect 43996 379448 44048 379500
rect 41420 378904 41472 378956
rect 43352 378904 43404 378956
rect 673644 378768 673696 378820
rect 675392 378768 675444 378820
rect 41512 378496 41564 378548
rect 43168 378496 43220 378548
rect 41604 378224 41656 378276
rect 43444 378224 43496 378276
rect 673736 377952 673788 378004
rect 675484 377952 675536 378004
rect 673552 377408 673604 377460
rect 675392 377408 675444 377460
rect 673828 376932 673880 376984
rect 675484 376932 675536 376984
rect 41420 376048 41472 376100
rect 48412 376048 48464 376100
rect 673460 375708 673512 375760
rect 675392 375708 675444 375760
rect 42432 374892 42484 374944
rect 44088 374892 44140 374944
rect 674472 373872 674524 373924
rect 675392 373872 675444 373924
rect 654508 372512 654560 372564
rect 675024 372512 675076 372564
rect 674656 372036 674708 372088
rect 675392 372036 675444 372088
rect 41512 371968 41564 372020
rect 43260 371968 43312 372020
rect 43628 371356 43680 371408
rect 43628 371220 43680 371272
rect 43812 371220 43864 371272
rect 43904 370948 43956 371000
rect 675208 370744 675260 370796
rect 675668 370744 675720 370796
rect 675116 370676 675168 370728
rect 675760 370676 675812 370728
rect 41328 370540 41380 370592
rect 41972 370200 42024 370252
rect 42340 369860 42392 369912
rect 42340 369316 42392 369368
rect 42708 369316 42760 369368
rect 42708 369180 42760 369232
rect 42156 368092 42208 368144
rect 42340 368092 42392 368144
rect 42708 366664 42760 366716
rect 42156 366528 42208 366580
rect 42708 366528 42760 366580
rect 42156 366256 42208 366308
rect 43168 366256 43220 366308
rect 43168 366120 43220 366172
rect 42340 365032 42392 365084
rect 42248 364828 42300 364880
rect 42248 364692 42300 364744
rect 43352 364692 43404 364744
rect 43352 364556 43404 364608
rect 43996 364556 44048 364608
rect 43168 364284 43220 364336
rect 43904 364284 43956 364336
rect 42156 363808 42208 363860
rect 43260 363808 43312 363860
rect 42156 363128 42208 363180
rect 43536 363128 43588 363180
rect 42432 361904 42484 361956
rect 43076 361904 43128 361956
rect 42708 361496 42760 361548
rect 58164 361496 58216 361548
rect 42340 361292 42392 361344
rect 58532 361292 58584 361344
rect 42340 360884 42392 360936
rect 43536 360884 43588 360936
rect 42340 360136 42392 360188
rect 43996 360136 44048 360188
rect 42156 359932 42208 359984
rect 43352 359932 43404 359984
rect 46112 358708 46164 358760
rect 58532 358708 58584 358760
rect 42432 358300 42484 358352
rect 43904 358300 43956 358352
rect 655520 356396 655572 356448
rect 676036 356396 676088 356448
rect 655428 356260 655480 356312
rect 675852 356260 675904 356312
rect 655612 356192 655664 356244
rect 675944 356192 675996 356244
rect 673368 356124 673420 356176
rect 676036 356124 676088 356176
rect 48504 355988 48556 356040
rect 58440 355988 58492 356040
rect 50988 355920 51040 355972
rect 58532 355920 58584 355972
rect 674656 353472 674708 353524
rect 676036 353472 676088 353524
rect 674932 353268 674984 353320
rect 676036 353268 676088 353320
rect 674564 352248 674616 352300
rect 675944 352248 675996 352300
rect 674840 351840 674892 351892
rect 676036 351840 676088 351892
rect 673644 351432 673696 351484
rect 675944 351432 675996 351484
rect 673552 350752 673604 350804
rect 675668 350752 675720 350804
rect 674288 350684 674340 350736
rect 675852 350684 675904 350736
rect 674748 350616 674800 350668
rect 675944 350616 675996 350668
rect 675024 350548 675076 350600
rect 676036 350548 676088 350600
rect 42156 350480 42208 350532
rect 57980 350480 58032 350532
rect 673828 349800 673880 349852
rect 676036 349800 676088 349852
rect 673460 347896 673512 347948
rect 675852 347896 675904 347948
rect 673736 347828 673788 347880
rect 675944 347828 675996 347880
rect 674472 347760 674524 347812
rect 676036 347760 676088 347812
rect 672724 347216 672776 347268
rect 676036 347216 676088 347268
rect 41880 344972 41932 345024
rect 44088 344972 44140 345024
rect 41512 344224 41564 344276
rect 50988 344224 51040 344276
rect 41788 344088 41840 344140
rect 43812 344088 43864 344140
rect 41512 343816 41564 343868
rect 48504 343816 48556 343868
rect 41512 343408 41564 343460
rect 46112 343408 46164 343460
rect 41512 342592 41564 342644
rect 43904 342592 43956 342644
rect 673276 342524 673328 342576
rect 673552 342524 673604 342576
rect 673460 342456 673512 342508
rect 673460 342252 673512 342304
rect 673644 342252 673696 342304
rect 674564 342252 674616 342304
rect 41512 341844 41564 341896
rect 43628 341844 43680 341896
rect 41512 341436 41564 341488
rect 43720 341436 43772 341488
rect 674564 341436 674616 341488
rect 675760 341436 675812 341488
rect 41788 341368 41840 341420
rect 43536 341368 43588 341420
rect 675116 341368 675168 341420
rect 675392 341368 675444 341420
rect 674932 340960 674984 341012
rect 675484 340960 675536 341012
rect 675024 340892 675076 340944
rect 675024 340620 675076 340672
rect 675116 340620 675168 340672
rect 675392 340620 675444 340672
rect 675024 340212 675076 340264
rect 675392 340212 675444 340264
rect 673276 340076 673328 340128
rect 675024 340076 675076 340128
rect 674656 339532 674708 339584
rect 675484 339532 675536 339584
rect 41788 339464 41840 339516
rect 43352 339464 43404 339516
rect 674840 337900 674892 337952
rect 675484 337900 675536 337952
rect 674748 337084 674800 337136
rect 675392 337084 675444 337136
rect 674288 336540 674340 336592
rect 675392 336540 675444 336592
rect 674472 336064 674524 336116
rect 675484 336064 675536 336116
rect 655980 335316 656032 335368
rect 675116 335316 675168 335368
rect 673644 333548 673696 333600
rect 675392 333548 675444 333600
rect 41880 333072 41932 333124
rect 48596 333072 48648 333124
rect 673736 332732 673788 332784
rect 675392 332732 675444 332784
rect 675116 332528 675168 332580
rect 675300 332528 675352 332580
rect 674564 332392 674616 332444
rect 675300 332392 675352 332444
rect 673828 332188 673880 332240
rect 675392 332188 675444 332240
rect 673460 331576 673512 331628
rect 675392 331576 675444 331628
rect 41512 331168 41564 331220
rect 42708 331168 42760 331220
rect 41420 331100 41472 331152
rect 43168 331100 43220 331152
rect 41696 330896 41748 330948
rect 43444 330896 43496 330948
rect 675024 330556 675076 330608
rect 675392 330556 675444 330608
rect 30288 330284 30340 330336
rect 42248 330284 42300 330336
rect 33048 330216 33100 330268
rect 42340 330216 42392 330268
rect 30196 330012 30248 330064
rect 43628 330012 43680 330064
rect 41788 329400 41840 329452
rect 43260 329400 43312 329452
rect 41604 329332 41656 329384
rect 43076 329332 43128 329384
rect 674932 328720 674984 328772
rect 675392 328720 675444 328772
rect 673552 326884 673604 326936
rect 675392 326884 675444 326936
rect 42064 323076 42116 323128
rect 42708 323076 42760 323128
rect 42708 322940 42760 322992
rect 43076 323144 43128 323196
rect 42248 321988 42300 322040
rect 43260 321988 43312 322040
rect 42248 321784 42300 321836
rect 43168 321784 43220 321836
rect 42156 321580 42208 321632
rect 43444 321580 43496 321632
rect 42248 320560 42300 320612
rect 43076 320560 43128 320612
rect 42248 319948 42300 320000
rect 43628 319948 43680 320000
rect 42432 318724 42484 318776
rect 42708 318724 42760 318776
rect 43260 318724 43312 318776
rect 58532 318724 58584 318776
rect 42340 317364 42392 317416
rect 58072 317364 58124 317416
rect 46112 314576 46164 314628
rect 58532 314576 58584 314628
rect 675208 314576 675260 314628
rect 676036 314576 676088 314628
rect 50988 314508 51040 314560
rect 58164 314508 58216 314560
rect 655428 312060 655480 312112
rect 676220 312060 676272 312112
rect 655704 311992 655756 312044
rect 676312 311992 676364 312044
rect 655520 311924 655572 311976
rect 676128 311924 676180 311976
rect 673000 311856 673052 311908
rect 676220 311856 676272 311908
rect 48504 311788 48556 311840
rect 58532 311788 58584 311840
rect 673368 311652 673420 311704
rect 676036 311652 676088 311704
rect 675116 311516 675168 311568
rect 676036 311516 676088 311568
rect 673276 311040 673328 311092
rect 676220 311040 676272 311092
rect 673184 310224 673236 310276
rect 676220 310224 676272 310276
rect 673092 309408 673144 309460
rect 676220 309408 676272 309460
rect 674656 309136 674708 309188
rect 676036 309136 676088 309188
rect 673552 308048 673604 308100
rect 676036 308048 676088 308100
rect 674932 307232 674984 307284
rect 676036 307232 676088 307284
rect 674840 306824 674892 306876
rect 676036 306824 676088 306876
rect 674288 306416 674340 306468
rect 676128 306416 676180 306468
rect 675024 306348 675076 306400
rect 676036 306348 676088 306400
rect 42064 306280 42116 306332
rect 58348 306280 58400 306332
rect 673828 305056 673880 305108
rect 676128 305056 676180 305108
rect 675116 304784 675168 304836
rect 676036 304784 676088 304836
rect 673736 304308 673788 304360
rect 676128 304308 676180 304360
rect 675208 304172 675260 304224
rect 676036 304172 676088 304224
rect 674472 303900 674524 303952
rect 676128 303900 676180 303952
rect 673644 303696 673696 303748
rect 676036 303696 676088 303748
rect 672816 300840 672868 300892
rect 678980 300840 679032 300892
rect 674840 300160 674892 300212
rect 41788 300092 41840 300144
rect 43904 300092 43956 300144
rect 675024 300024 675076 300076
rect 41788 299956 41840 300008
rect 43536 299956 43588 300008
rect 674840 299956 674892 300008
rect 675024 299820 675076 299872
rect 42064 299344 42116 299396
rect 43260 299344 43312 299396
rect 41788 299072 41840 299124
rect 43352 299072 43404 299124
rect 655060 298120 655112 298172
rect 675392 298120 675444 298172
rect 41788 297304 41840 297356
rect 43628 297304 43680 297356
rect 41788 296216 41840 296268
rect 43812 296216 43864 296268
rect 675024 295400 675076 295452
rect 675300 295400 675352 295452
rect 42340 295332 42392 295384
rect 58532 295332 58584 295384
rect 674748 294720 674800 294772
rect 675300 294720 675352 294772
rect 674656 294516 674708 294568
rect 675392 294516 675444 294568
rect 42064 293632 42116 293684
rect 43996 293632 44048 293684
rect 42064 293428 42116 293480
rect 44088 293428 44140 293480
rect 43536 292612 43588 292664
rect 58440 292612 58492 292664
rect 41972 292476 42024 292528
rect 57980 292476 58032 292528
rect 41880 292408 41932 292460
rect 58532 292408 58584 292460
rect 41880 292272 41932 292324
rect 43076 292272 43128 292324
rect 674932 291524 674984 291576
rect 675392 291524 675444 291576
rect 41788 291048 41840 291100
rect 51080 291048 51132 291100
rect 41788 290640 41840 290692
rect 51172 290640 51224 290692
rect 674472 290436 674524 290488
rect 675116 290436 675168 290488
rect 41788 289824 41840 289876
rect 48780 289824 48832 289876
rect 27528 289756 27580 289808
rect 57980 289756 58032 289808
rect 674288 288600 674340 288652
rect 675392 288600 675444 288652
rect 654508 288532 654560 288584
rect 666836 288532 666888 288584
rect 673736 287376 673788 287428
rect 675116 287376 675168 287428
rect 48688 287104 48740 287156
rect 58164 287104 58216 287156
rect 656808 287104 656860 287156
rect 669412 287104 669464 287156
rect 46296 287036 46348 287088
rect 58532 287036 58584 287088
rect 654876 287036 654928 287088
rect 669504 287036 669556 287088
rect 35808 286968 35860 287020
rect 42248 286968 42300 287020
rect 42156 286900 42208 286952
rect 43444 286900 43496 286952
rect 41972 286832 42024 286884
rect 43352 286832 43404 286884
rect 673828 286764 673880 286816
rect 675116 286764 675168 286816
rect 673644 286560 673696 286612
rect 675392 286560 675444 286612
rect 42064 286152 42116 286204
rect 43168 286152 43220 286204
rect 41696 285744 41748 285796
rect 43812 285744 43864 285796
rect 42432 285608 42484 285660
rect 43720 285608 43772 285660
rect 655428 284928 655480 284980
rect 669596 284928 669648 284980
rect 56508 284792 56560 284844
rect 57980 284792 58032 284844
rect 654876 284656 654928 284708
rect 666744 284656 666796 284708
rect 51264 284316 51316 284368
rect 58532 284316 58584 284368
rect 43996 284248 44048 284300
rect 44272 284248 44324 284300
rect 43076 284112 43128 284164
rect 43996 284112 44048 284164
rect 41880 283772 41932 283824
rect 673552 283704 673604 283756
rect 675484 283704 675536 283756
rect 41880 283568 41932 283620
rect 43076 281596 43128 281648
rect 44272 281596 44324 281648
rect 50988 281596 51040 281648
rect 58256 281596 58308 281648
rect 656808 281596 656860 281648
rect 669228 281596 669280 281648
rect 48504 281528 48556 281580
rect 58532 281528 58584 281580
rect 42340 280440 42392 280492
rect 43352 280440 43404 280492
rect 42248 280372 42300 280424
rect 43536 280372 43588 280424
rect 654692 280168 654744 280220
rect 669320 280168 669372 280220
rect 42156 279828 42208 279880
rect 43168 279828 43220 279880
rect 654876 278944 654928 278996
rect 666652 278944 666704 278996
rect 46204 278808 46256 278860
rect 58164 278808 58216 278860
rect 46112 278740 46164 278792
rect 58256 278740 58308 278792
rect 42064 278400 42116 278452
rect 42708 278400 42760 278452
rect 42156 277856 42208 277908
rect 43444 277856 43496 277908
rect 45652 277312 45704 277364
rect 666560 277312 666612 277364
rect 42340 276768 42392 276820
rect 43812 276768 43864 276820
rect 342536 275952 342588 276004
rect 464160 275952 464212 276004
rect 345112 275884 345164 275936
rect 471244 275884 471296 275936
rect 347780 275816 347832 275868
rect 478328 275816 478380 275868
rect 346400 275748 346452 275800
rect 474832 275748 474884 275800
rect 351644 275680 351696 275732
rect 489000 275680 489052 275732
rect 353208 275612 353260 275664
rect 492588 275612 492640 275664
rect 42432 275544 42484 275596
rect 43996 275544 44048 275596
rect 357072 275544 357124 275596
rect 503168 275544 503220 275596
rect 358452 275476 358504 275528
rect 506756 275476 506808 275528
rect 361120 275408 361172 275460
rect 513840 275408 513892 275460
rect 363788 275340 363840 275392
rect 520924 275340 520976 275392
rect 366456 275272 366508 275324
rect 528008 275272 528060 275324
rect 371792 275204 371844 275256
rect 375288 275136 375340 275188
rect 390652 275204 390704 275256
rect 535092 275204 535144 275256
rect 377772 275068 377824 275120
rect 542176 275136 542228 275188
rect 550456 275068 550508 275120
rect 557540 275000 557592 275052
rect 380348 274932 380400 274984
rect 564624 274932 564676 274984
rect 383292 274864 383344 274916
rect 571708 274864 571760 274916
rect 317512 274796 317564 274848
rect 398012 274796 398064 274848
rect 320180 274728 320232 274780
rect 390468 274728 390520 274780
rect 397644 274728 397696 274780
rect 610716 274796 610768 274848
rect 402980 274728 403032 274780
rect 624976 274728 625028 274780
rect 321008 274660 321060 274712
rect 407488 274660 407540 274712
rect 409236 274660 409288 274712
rect 322572 274592 322624 274644
rect 410984 274592 411036 274644
rect 429108 274660 429160 274712
rect 634360 274660 634412 274712
rect 641444 274592 641496 274644
rect 341064 274524 341116 274576
rect 460664 274524 460716 274576
rect 338396 274456 338448 274508
rect 453580 274456 453632 274508
rect 337108 274388 337160 274440
rect 449992 274388 450044 274440
rect 336096 274320 336148 274372
rect 446496 274320 446548 274372
rect 334348 274252 334400 274304
rect 351920 274252 351972 274304
rect 439320 274252 439372 274304
rect 333060 274116 333112 274168
rect 351736 274116 351788 274168
rect 351828 274116 351880 274168
rect 330392 274048 330444 274100
rect 442908 274116 442960 274168
rect 331680 273980 331732 274032
rect 433432 274048 433484 274100
rect 327724 273912 327776 273964
rect 425152 273912 425204 273964
rect 432236 273980 432288 274032
rect 435824 273912 435876 273964
rect 329012 273844 329064 273896
rect 428740 273844 428792 273896
rect 325056 273776 325108 273828
rect 418068 273776 418120 273828
rect 42432 273708 42484 273760
rect 44088 273708 44140 273760
rect 325516 273708 325568 273760
rect 419264 273708 419316 273760
rect 326344 273640 326396 273692
rect 421656 273640 421708 273692
rect 323676 273572 323728 273624
rect 414572 273572 414624 273624
rect 330852 273504 330904 273556
rect 351828 273504 351880 273556
rect 390468 273504 390520 273556
rect 405096 273504 405148 273556
rect 406568 273504 406620 273556
rect 429108 273504 429160 273556
rect 369124 273436 369176 273488
rect 390652 273436 390704 273488
rect 154488 273164 154540 273216
rect 211068 273164 211120 273216
rect 42432 273096 42484 273148
rect 43076 273096 43128 273148
rect 176844 273096 176896 273148
rect 210976 273096 211028 273148
rect 152188 273028 152240 273080
rect 224500 273164 224552 273216
rect 263232 273164 263284 273216
rect 266728 273164 266780 273216
rect 292120 273164 292172 273216
rect 330576 273164 330628 273216
rect 352656 273164 352708 273216
rect 491392 273164 491444 273216
rect 491484 273164 491536 273216
rect 507952 273164 508004 273216
rect 260932 273096 260984 273148
rect 265808 273096 265860 273148
rect 293868 273096 293920 273148
rect 335360 273096 335412 273148
rect 344928 273096 344980 273148
rect 470140 273096 470192 273148
rect 471980 273096 472032 273148
rect 614304 273096 614356 273148
rect 211252 273028 211304 273080
rect 217968 273028 218020 273080
rect 243176 273028 243228 273080
rect 259184 273028 259236 273080
rect 259736 273028 259788 273080
rect 265440 273028 265492 273080
rect 296076 273028 296128 273080
rect 341248 273028 341300 273080
rect 356060 273028 356112 273080
rect 358820 273028 358872 273080
rect 358912 273028 358964 273080
rect 497280 273028 497332 273080
rect 497924 273028 497976 273080
rect 600136 273028 600188 273080
rect 147404 272960 147456 273012
rect 222660 272960 222712 273012
rect 240784 272960 240836 273012
rect 258264 272960 258316 273012
rect 301872 272960 301924 273012
rect 356612 272960 356664 273012
rect 360568 272960 360620 273012
rect 511448 272960 511500 273012
rect 149796 272892 149848 272944
rect 214748 272892 214800 272944
rect 214840 272892 214892 272944
rect 220452 272892 220504 272944
rect 234896 272892 234948 272944
rect 256056 272892 256108 272944
rect 303528 272892 303580 272944
rect 360200 272892 360252 272944
rect 363144 272892 363196 272944
rect 518532 272892 518584 272944
rect 146208 272824 146260 272876
rect 223028 272824 223080 272876
rect 233700 272824 233752 272876
rect 255596 272824 255648 272876
rect 294880 272824 294932 272876
rect 337752 272824 337804 272876
rect 347504 272824 347556 272876
rect 477224 272824 477276 272876
rect 477316 272824 477368 272876
rect 632060 272824 632112 272876
rect 139124 272756 139176 272808
rect 220360 272756 220412 272808
rect 236092 272756 236144 272808
rect 256424 272756 256476 272808
rect 295064 272756 295116 272808
rect 338856 272756 338908 272808
rect 342168 272756 342220 272808
rect 462964 272756 463016 272808
rect 463332 272756 463384 272808
rect 621388 272756 621440 272808
rect 141516 272688 141568 272740
rect 221188 272688 221240 272740
rect 232504 272688 232556 272740
rect 255136 272688 255188 272740
rect 324228 272688 324280 272740
rect 362500 272688 362552 272740
rect 362592 272688 362644 272740
rect 370780 272688 370832 272740
rect 375656 272688 375708 272740
rect 381452 272688 381504 272740
rect 391940 272688 391992 272740
rect 555240 272688 555292 272740
rect 119068 272620 119120 272672
rect 126152 272552 126204 272604
rect 140320 272620 140372 272672
rect 219992 272620 220044 272672
rect 306748 272620 306800 272672
rect 369584 272620 369636 272672
rect 369676 272620 369728 272672
rect 532700 272620 532752 272672
rect 187700 272484 187752 272536
rect 89536 272416 89588 272468
rect 177120 272416 177172 272468
rect 193496 272552 193548 272604
rect 203616 272552 203668 272604
rect 214748 272552 214800 272604
rect 224408 272552 224460 272604
rect 293408 272552 293460 272604
rect 334164 272552 334216 272604
rect 336648 272552 336700 272604
rect 448796 272552 448848 272604
rect 448888 272552 448940 272604
rect 628472 272552 628524 272604
rect 197268 272484 197320 272536
rect 206836 272416 206888 272468
rect 211068 272484 211120 272536
rect 225328 272484 225380 272536
rect 229008 272484 229060 272536
rect 253756 272484 253808 272536
rect 307208 272484 307260 272536
rect 232044 272416 232096 272468
rect 237288 272416 237340 272468
rect 256884 272416 256936 272468
rect 306288 272416 306340 272468
rect 322296 272484 322348 272536
rect 367284 272484 367336 272536
rect 379336 272484 379388 272536
rect 562324 272484 562376 272536
rect 111984 272348 112036 272400
rect 201592 272348 201644 272400
rect 288164 272348 288216 272400
rect 319996 272348 320048 272400
rect 362592 272416 362644 272468
rect 362868 272416 362920 272468
rect 384948 272416 385000 272468
rect 386420 272416 386472 272468
rect 569408 272416 569460 272468
rect 322296 272348 322348 272400
rect 322848 272348 322900 272400
rect 383844 272348 383896 272400
rect 384672 272348 384724 272400
rect 576492 272348 576544 272400
rect 117872 272280 117924 272332
rect 88340 272212 88392 272264
rect 184940 272212 184992 272264
rect 185216 272212 185268 272264
rect 197268 272212 197320 272264
rect 102508 272144 102560 272196
rect 201500 272144 201552 272196
rect 210976 272280 211028 272332
rect 227076 272280 227128 272332
rect 230204 272280 230256 272332
rect 254216 272280 254268 272332
rect 309324 272280 309376 272332
rect 309876 272280 309928 272332
rect 377864 272280 377916 272332
rect 390008 272280 390060 272332
rect 590660 272280 590712 272332
rect 209688 272212 209740 272264
rect 238484 272212 238536 272264
rect 257252 272212 257304 272264
rect 284208 272212 284260 272264
rect 292580 272212 292632 272264
rect 331772 272212 331824 272264
rect 205364 272144 205416 272196
rect 244924 272144 244976 272196
rect 285864 272144 285916 272196
rect 314108 272144 314160 272196
rect 331312 272144 331364 272196
rect 434628 272212 434680 272264
rect 436100 272212 436152 272264
rect 639144 272212 639196 272264
rect 97816 272076 97868 272128
rect 198832 272076 198884 272128
rect 204168 272076 204220 272128
rect 240140 272076 240192 272128
rect 288532 272076 288584 272128
rect 321192 272076 321244 272128
rect 362868 272144 362920 272196
rect 367100 272144 367152 272196
rect 387340 272144 387392 272196
rect 392768 272144 392820 272196
rect 597744 272144 597796 272196
rect 96620 272008 96672 272060
rect 198740 272008 198792 272060
rect 202972 272008 203024 272060
rect 244004 272008 244056 272060
rect 286692 272008 286744 272060
rect 316408 272008 316460 272060
rect 317328 272008 317380 272060
rect 332324 272076 332376 272128
rect 390928 272076 390980 272128
rect 398104 272076 398156 272128
rect 611912 272076 611964 272128
rect 332232 272008 332284 272060
rect 392124 272008 392176 272060
rect 406108 272008 406160 272060
rect 77668 271940 77720 271992
rect 193220 271940 193272 271992
rect 198280 271940 198332 271992
rect 242256 271940 242308 271992
rect 244372 271940 244424 271992
rect 259552 271940 259604 271992
rect 262128 271940 262180 271992
rect 266268 271940 266320 271992
rect 286600 271940 286652 271992
rect 315212 271940 315264 271992
rect 320548 271940 320600 271992
rect 156880 271872 156932 271924
rect 176844 271872 176896 271924
rect 176936 271872 176988 271924
rect 193128 271872 193180 271924
rect 194692 271872 194744 271924
rect 240876 271872 240928 271924
rect 289176 271872 289228 271924
rect 322388 271872 322440 271924
rect 332140 271940 332192 271992
rect 399208 271940 399260 271992
rect 409604 271940 409656 271992
rect 413836 272008 413888 272060
rect 618996 272008 619048 272060
rect 406292 271872 406344 271924
rect 411444 271872 411496 271924
rect 633256 271940 633308 271992
rect 42432 271804 42484 271856
rect 59268 271804 59320 271856
rect 67088 271804 67140 271856
rect 127348 271736 127400 271788
rect 189908 271736 189960 271788
rect 191196 271804 191248 271856
rect 239496 271804 239548 271856
rect 247868 271804 247920 271856
rect 260932 271804 260984 271856
rect 264428 271804 264480 271856
rect 267188 271804 267240 271856
rect 289636 271804 289688 271856
rect 323492 271804 323544 271856
rect 323584 271804 323636 271856
rect 413376 271804 413428 271856
rect 642640 271872 642692 271924
rect 647424 271804 647476 271856
rect 192484 271736 192536 271788
rect 200580 271736 200632 271788
rect 243268 271736 243320 271788
rect 249064 271736 249116 271788
rect 261392 271736 261444 271788
rect 292028 271736 292080 271788
rect 329472 271736 329524 271788
rect 352196 271736 352248 271788
rect 490196 271736 490248 271788
rect 159272 271668 159324 271720
rect 227536 271668 227588 271720
rect 239588 271668 239640 271720
rect 163964 271600 164016 271652
rect 229744 271600 229796 271652
rect 245568 271600 245620 271652
rect 251180 271600 251232 271652
rect 161572 271532 161624 271584
rect 227996 271532 228048 271584
rect 171048 271464 171100 271516
rect 229284 271464 229336 271516
rect 241980 271464 242032 271516
rect 251272 271464 251324 271516
rect 251456 271668 251508 271720
rect 262220 271668 262272 271720
rect 291200 271668 291252 271720
rect 328276 271668 328328 271720
rect 350172 271668 350224 271720
rect 484308 271668 484360 271720
rect 485688 271668 485740 271720
rect 607220 271668 607272 271720
rect 253848 271600 253900 271652
rect 263140 271600 263192 271652
rect 290280 271600 290332 271652
rect 325884 271600 325936 271652
rect 349620 271600 349672 271652
rect 483112 271600 483164 271652
rect 257344 271532 257396 271584
rect 264520 271532 264572 271584
rect 290740 271532 290792 271584
rect 327080 271532 327132 271584
rect 346860 271532 346912 271584
rect 476028 271532 476080 271584
rect 257804 271464 257856 271516
rect 258540 271464 258592 271516
rect 264888 271464 264940 271516
rect 266820 271464 266872 271516
rect 268016 271464 268068 271516
rect 289820 271464 289872 271516
rect 324688 271464 324740 271516
rect 344192 271464 344244 271516
rect 468944 271464 468996 271516
rect 168748 271396 168800 271448
rect 230388 271396 230440 271448
rect 166356 271328 166408 271380
rect 224040 271328 224092 271380
rect 227812 271328 227864 271380
rect 253388 271396 253440 271448
rect 254952 271396 255004 271448
rect 263600 271396 263652 271448
rect 287612 271396 287664 271448
rect 318800 271396 318852 271448
rect 322664 271396 322716 271448
rect 332324 271396 332376 271448
rect 342076 271396 342128 271448
rect 252652 271328 252704 271380
rect 262864 271328 262916 271380
rect 285404 271328 285456 271380
rect 312912 271328 312964 271380
rect 315212 271328 315264 271380
rect 332232 271328 332284 271380
rect 339224 271328 339276 271380
rect 452660 271396 452712 271448
rect 458272 271396 458324 271448
rect 173440 271260 173492 271312
rect 227628 271260 227680 271312
rect 231308 271260 231360 271312
rect 178132 271192 178184 271244
rect 231860 271192 231912 271244
rect 250260 271260 250312 271312
rect 261852 271260 261904 271312
rect 287152 271260 287204 271312
rect 317604 271260 317656 271312
rect 317880 271260 317932 271312
rect 332140 271260 332192 271312
rect 337476 271260 337528 271312
rect 254676 271192 254728 271244
rect 304080 271192 304132 271244
rect 324228 271192 324280 271244
rect 333980 271192 334032 271244
rect 441712 271192 441764 271244
rect 175832 271124 175884 271176
rect 229100 271124 229152 271176
rect 246764 271124 246816 271176
rect 260472 271124 260524 271176
rect 334808 271124 334860 271176
rect 444104 271124 444156 271176
rect 461860 271260 461912 271312
rect 455880 271192 455932 271244
rect 451188 271124 451240 271176
rect 186412 271056 186464 271108
rect 231952 271056 232004 271108
rect 251272 271056 251324 271108
rect 258724 271056 258776 271108
rect 329472 271056 329524 271108
rect 429936 271056 429988 271108
rect 442540 271056 442592 271108
rect 454684 271056 454736 271108
rect 180524 270988 180576 271040
rect 227812 270988 227864 271040
rect 251180 270988 251232 271040
rect 260012 270988 260064 271040
rect 328644 270988 328696 271040
rect 427544 270988 427596 271040
rect 187608 270920 187660 270972
rect 230756 270920 230808 270972
rect 325976 270920 326028 270972
rect 420460 270920 420512 270972
rect 420828 270920 420880 270972
rect 447600 270920 447652 270972
rect 184112 270852 184164 270904
rect 227444 270852 227496 270904
rect 325792 270852 325844 270904
rect 376760 270852 376812 270904
rect 385684 270852 385736 270904
rect 437020 270852 437072 270904
rect 190000 270784 190052 270836
rect 229836 270784 229888 270836
rect 325700 270784 325752 270836
rect 179328 270716 179380 270768
rect 184112 270716 184164 270768
rect 187700 270716 187752 270768
rect 71780 270648 71832 270700
rect 194600 270648 194652 270700
rect 189908 270580 189960 270632
rect 197176 270580 197228 270632
rect 199476 270716 199528 270768
rect 242624 270716 242676 270768
rect 317236 270716 317288 270768
rect 345940 270716 345992 270768
rect 201776 270648 201828 270700
rect 243544 270648 243596 270700
rect 256148 270648 256200 270700
rect 264060 270648 264112 270700
rect 319904 270648 319956 270700
rect 349528 270648 349580 270700
rect 354864 270784 354916 270836
rect 358912 270784 358964 270836
rect 381360 270784 381412 270836
rect 422852 270784 422904 270836
rect 360844 270716 360896 270768
rect 373172 270716 373224 270768
rect 375564 270716 375616 270768
rect 408592 270716 408644 270768
rect 366088 270648 366140 270700
rect 369860 270648 369912 270700
rect 401508 270648 401560 270700
rect 207664 270580 207716 270632
rect 207756 270580 207808 270632
rect 215208 270580 215260 270632
rect 218336 270580 218388 270632
rect 223396 270580 223448 270632
rect 226616 270580 226668 270632
rect 252928 270580 252980 270632
rect 313188 270580 313240 270632
rect 342444 270580 342496 270632
rect 375380 270580 375432 270632
rect 394424 270580 394476 270632
rect 400772 270580 400824 270632
rect 413836 270580 413888 270632
rect 150992 270512 151044 270564
rect 192392 270512 192444 270564
rect 239956 270512 240008 270564
rect 364340 270512 364392 270564
rect 380256 270512 380308 270564
rect 207572 270444 207624 270496
rect 207664 270444 207716 270496
rect 214656 270444 214708 270496
rect 227628 270444 227680 270496
rect 232872 270444 232924 270496
rect 265624 270444 265676 270496
rect 267556 270444 267608 270496
rect 269396 270444 269448 270496
rect 270316 270444 270368 270496
rect 270684 270444 270736 270496
rect 273904 270444 273956 270496
rect 274272 270444 274324 270496
rect 283380 270444 283432 270496
rect 294328 270444 294380 270496
rect 336556 270444 336608 270496
rect 351276 270444 351328 270496
rect 148600 270376 148652 270428
rect 223212 270376 223264 270428
rect 229284 270376 229336 270428
rect 232412 270376 232464 270428
rect 271144 270376 271196 270428
rect 275100 270376 275152 270428
rect 277492 270376 277544 270428
rect 291568 270376 291620 270428
rect 295616 270376 295668 270428
rect 340052 270376 340104 270428
rect 349068 270376 349120 270428
rect 356060 270376 356112 270428
rect 145104 270308 145156 270360
rect 222200 270308 222252 270360
rect 224224 270308 224276 270360
rect 252008 270308 252060 270360
rect 271604 270308 271656 270360
rect 276204 270308 276256 270360
rect 277860 270308 277912 270360
rect 143908 270240 143960 270292
rect 221280 270240 221332 270292
rect 225420 270240 225472 270292
rect 252468 270240 252520 270292
rect 272064 270240 272116 270292
rect 277400 270240 277452 270292
rect 278688 270240 278740 270292
rect 135628 270172 135680 270224
rect 219072 270172 219124 270224
rect 219532 270172 219584 270224
rect 250260 270172 250312 270224
rect 272524 270172 272576 270224
rect 278596 270172 278648 270224
rect 279148 270172 279200 270224
rect 142712 270104 142764 270156
rect 221740 270104 221792 270156
rect 221924 270104 221976 270156
rect 251088 270104 251140 270156
rect 272984 270104 273036 270156
rect 279792 270104 279844 270156
rect 136824 270036 136876 270088
rect 218612 270036 218664 270088
rect 223396 270036 223448 270088
rect 249800 270036 249852 270088
rect 273720 270036 273772 270088
rect 280988 270036 281040 270088
rect 137928 269968 137980 270020
rect 219532 269968 219584 270020
rect 220728 269968 220780 270020
rect 250720 269968 250772 270020
rect 273812 269968 273864 270020
rect 282184 269968 282236 270020
rect 297456 270308 297508 270360
rect 344836 270308 344888 270360
rect 350908 270308 350960 270360
rect 362868 270444 362920 270496
rect 480720 270444 480772 270496
rect 358912 270376 358964 270428
rect 491484 270376 491536 270428
rect 282552 270240 282604 270292
rect 290464 270240 290516 270292
rect 296996 270240 297048 270292
rect 343640 270240 343692 270292
rect 487804 270308 487856 270360
rect 486608 270240 486660 270292
rect 292764 270172 292816 270224
rect 298284 270172 298336 270224
rect 347136 270172 347188 270224
rect 348608 270172 348660 270224
rect 351920 270172 351972 270224
rect 353576 270172 353628 270224
rect 493692 270172 493744 270224
rect 295156 270104 295208 270156
rect 298836 270104 298888 270156
rect 348332 270104 348384 270156
rect 348792 270104 348844 270156
rect 355416 270104 355468 270156
rect 282368 270036 282420 270088
rect 293960 270036 294012 270088
rect 300584 270036 300636 270088
rect 353116 270036 353168 270088
rect 353944 270036 353996 270088
rect 494888 270104 494940 270156
rect 356244 270036 356296 270088
rect 500868 270036 500920 270088
rect 296352 269968 296404 270020
rect 300124 269968 300176 270020
rect 351552 269968 351604 270020
rect 130844 269900 130896 269952
rect 216864 269900 216916 269952
rect 223120 269900 223172 269952
rect 251548 269900 251600 269952
rect 279608 269900 279660 269952
rect 297548 269900 297600 269952
rect 301412 269900 301464 269952
rect 348792 269900 348844 269952
rect 129648 269832 129700 269884
rect 215852 269832 215904 269884
rect 220452 269832 220504 269884
rect 248420 269832 248472 269884
rect 278320 269832 278372 269884
rect 282368 269832 282420 269884
rect 282460 269832 282512 269884
rect 286876 269832 286928 269884
rect 308220 269832 308272 269884
rect 360844 269968 360896 270020
rect 361580 269968 361632 270020
rect 515036 269968 515088 270020
rect 128544 269764 128596 269816
rect 216404 269764 216456 269816
rect 217968 269764 218020 269816
rect 247132 269764 247184 269816
rect 280528 269764 280580 269816
rect 299848 269764 299900 269816
rect 302792 269764 302844 269816
rect 349068 269764 349120 269816
rect 122564 269696 122616 269748
rect 213276 269696 213328 269748
rect 215944 269696 215996 269748
rect 248880 269696 248932 269748
rect 280068 269696 280120 269748
rect 298744 269696 298796 269748
rect 310796 269696 310848 269748
rect 364340 269900 364392 269952
rect 364708 269900 364760 269952
rect 523316 269900 523368 269952
rect 351920 269832 351972 269884
rect 362868 269832 362920 269884
rect 367376 269832 367428 269884
rect 530400 269832 530452 269884
rect 370044 269764 370096 269816
rect 537484 269764 537536 269816
rect 101312 269628 101364 269680
rect 205272 269628 205324 269680
rect 215208 269628 215260 269680
rect 245752 269628 245804 269680
rect 281816 269628 281868 269680
rect 303436 269628 303488 269680
rect 313464 269628 313516 269680
rect 351828 269628 351880 269680
rect 115480 269560 115532 269612
rect 210608 269560 210660 269612
rect 217140 269560 217192 269612
rect 249340 269560 249392 269612
rect 281448 269560 281500 269612
rect 302240 269560 302292 269612
rect 304540 269560 304592 269612
rect 363696 269696 363748 269748
rect 372712 269696 372764 269748
rect 544568 269696 544620 269748
rect 352012 269628 352064 269680
rect 367100 269628 367152 269680
rect 375472 269628 375524 269680
rect 551652 269628 551704 269680
rect 352472 269560 352524 269612
rect 361672 269560 361724 269612
rect 362868 269560 362920 269612
rect 385684 269560 385736 269612
rect 100116 269492 100168 269544
rect 205732 269492 205784 269544
rect 212448 269492 212500 269544
rect 247592 269492 247644 269544
rect 280988 269492 281040 269544
rect 301044 269492 301096 269544
rect 316132 269492 316184 269544
rect 375380 269492 375432 269544
rect 377864 269492 377916 269544
rect 558736 269560 558788 269612
rect 94228 269424 94280 269476
rect 202604 269424 202656 269476
rect 210056 269424 210108 269476
rect 246672 269424 246724 269476
rect 275652 269424 275704 269476
rect 282460 269424 282512 269476
rect 282736 269424 282788 269476
rect 305828 269424 305880 269476
rect 308588 269424 308640 269476
rect 374368 269424 374420 269476
rect 91836 269356 91888 269408
rect 202144 269356 202196 269408
rect 208860 269356 208912 269408
rect 246212 269356 246264 269408
rect 282276 269356 282328 269408
rect 304632 269356 304684 269408
rect 311256 269356 311308 269408
rect 375656 269356 375708 269408
rect 386052 269356 386104 269408
rect 579988 269492 580040 269544
rect 82452 269288 82504 269340
rect 198556 269288 198608 269340
rect 206560 269288 206612 269340
rect 229008 269288 229060 269340
rect 229100 269288 229152 269340
rect 233332 269288 233384 269340
rect 276940 269288 276992 269340
rect 282552 269288 282604 269340
rect 283656 269288 283708 269340
rect 308128 269288 308180 269340
rect 313924 269288 313976 269340
rect 388536 269288 388588 269340
rect 388720 269288 388772 269340
rect 587072 269424 587124 269476
rect 391388 269356 391440 269408
rect 594248 269356 594300 269408
rect 394056 269288 394108 269340
rect 601332 269288 601384 269340
rect 75368 269220 75420 269272
rect 195428 269220 195480 269272
rect 203616 269220 203668 269272
rect 240416 269220 240468 269272
rect 283196 269220 283248 269272
rect 307024 269220 307076 269272
rect 319260 269220 319312 269272
rect 197084 269152 197136 269204
rect 241796 269152 241848 269204
rect 284944 269152 284996 269204
rect 311716 269152 311768 269204
rect 65892 269084 65944 269136
rect 192392 269084 192444 269136
rect 195888 269084 195940 269136
rect 241336 269084 241388 269136
rect 284576 269084 284628 269136
rect 310520 269084 310572 269136
rect 153384 269016 153436 269068
rect 225788 269016 225840 269068
rect 229008 269016 229060 269068
rect 245292 269016 245344 269068
rect 292948 269016 293000 269068
rect 332968 269152 333020 269204
rect 333152 269220 333204 269272
rect 395620 269220 395672 269272
rect 396724 269220 396776 269272
rect 608416 269220 608468 269272
rect 321928 269084 321980 269136
rect 401324 269084 401376 269136
rect 402060 269152 402112 269204
rect 622584 269152 622636 269204
rect 402704 269084 402756 269136
rect 410064 269084 410116 269136
rect 643836 269084 643888 269136
rect 332600 269016 332652 269068
rect 351736 269016 351788 269068
rect 361672 269016 361724 269068
rect 479524 269016 479576 269068
rect 158076 268948 158128 269000
rect 226616 268948 226668 269000
rect 232044 268948 232096 269000
rect 237748 268948 237800 269000
rect 305460 268948 305512 269000
rect 325700 268948 325752 269000
rect 345480 268948 345532 269000
rect 472440 268948 472492 269000
rect 155684 268880 155736 268932
rect 226156 268880 226208 268932
rect 299204 268880 299256 268932
rect 319904 268880 319956 268932
rect 329932 268880 329984 268932
rect 351920 268880 351972 268932
rect 160468 268812 160520 268864
rect 228456 268812 228508 268864
rect 297916 268812 297968 268864
rect 317236 268812 317288 268864
rect 345940 268812 345992 268864
rect 473636 268880 473688 268932
rect 352104 268812 352156 268864
rect 466552 268812 466604 268864
rect 165160 268744 165212 268796
rect 229284 268744 229336 268796
rect 316592 268744 316644 268796
rect 333152 268744 333204 268796
rect 348240 268744 348292 268796
rect 352472 268744 352524 268796
rect 352564 268744 352616 268796
rect 465356 268744 465408 268796
rect 162768 268676 162820 268728
rect 228824 268676 228876 268728
rect 229836 268676 229888 268728
rect 238668 268676 238720 268728
rect 296536 268676 296588 268728
rect 313188 268676 313240 268728
rect 340604 268676 340656 268728
rect 459468 268676 459520 268728
rect 167552 268608 167604 268660
rect 231124 268608 231176 268660
rect 231952 268608 232004 268660
rect 237288 268608 237340 268660
rect 312084 268608 312136 268660
rect 322848 268608 322900 268660
rect 340144 268608 340196 268660
rect 452660 268608 452712 268660
rect 169852 268540 169904 268592
rect 231492 268540 231544 268592
rect 240140 268540 240192 268592
rect 244464 268540 244516 268592
rect 337936 268540 337988 268592
rect 452384 268540 452436 268592
rect 172244 268472 172296 268524
rect 231952 268472 232004 268524
rect 269856 268472 269908 268524
rect 271512 268472 271564 268524
rect 312544 268472 312596 268524
rect 317328 268472 317380 268524
rect 335268 268472 335320 268524
rect 445300 268472 445352 268524
rect 174636 268404 174688 268456
rect 233792 268404 233844 268456
rect 338856 268404 338908 268456
rect 442540 268404 442592 268456
rect 181720 268336 181772 268388
rect 236460 268336 236512 268388
rect 276480 268336 276532 268388
rect 289268 268336 289320 268388
rect 332140 268336 332192 268388
rect 348148 268336 348200 268388
rect 351736 268336 351788 268388
rect 438216 268336 438268 268388
rect 184112 268268 184164 268320
rect 234620 268268 234672 268320
rect 274732 268268 274784 268320
rect 284484 268268 284536 268320
rect 336464 268268 336516 268320
rect 351828 268268 351880 268320
rect 351920 268268 351972 268320
rect 431132 268268 431184 268320
rect 193220 268200 193272 268252
rect 196348 268200 196400 268252
rect 182916 268132 182968 268184
rect 197268 268132 197320 268184
rect 188804 268064 188856 268116
rect 239128 268200 239180 268252
rect 275192 268200 275244 268252
rect 285680 268200 285732 268252
rect 309416 268200 309468 268252
rect 325792 268200 325844 268252
rect 327264 268200 327316 268252
rect 423956 268200 424008 268252
rect 198832 268064 198884 268116
rect 203892 268064 203944 268116
rect 177120 267996 177172 268048
rect 200764 267996 200816 268048
rect 201500 267996 201552 268048
rect 206192 267996 206244 268048
rect 74172 267928 74224 267980
rect 195888 267928 195940 267980
rect 197268 267928 197320 267980
rect 236000 268132 236052 268184
rect 270316 268132 270368 268184
rect 272708 268132 272760 268184
rect 324596 268132 324648 268184
rect 234160 268064 234212 268116
rect 321468 268064 321520 268116
rect 206560 267996 206612 268048
rect 215484 267996 215536 268048
rect 193128 267860 193180 267912
rect 209228 267928 209280 267980
rect 209688 267928 209740 267980
rect 212356 267928 212408 267980
rect 213644 267928 213696 267980
rect 248052 267996 248104 268048
rect 343272 268064 343324 268116
rect 351736 268064 351788 268116
rect 351828 268064 351880 268116
rect 375564 267996 375616 268048
rect 382004 267996 382056 268048
rect 386420 267996 386472 268048
rect 227812 267928 227864 267980
rect 235540 267928 235592 267980
rect 326804 267928 326856 267980
rect 381360 267928 381412 267980
rect 401324 268132 401376 268184
rect 409788 268132 409840 268184
rect 416872 267996 416924 268048
rect 420828 268064 420880 268116
rect 656256 268064 656308 268116
rect 676220 268064 676272 268116
rect 656072 267928 656124 267980
rect 676036 267928 676088 267980
rect 201592 267792 201644 267844
rect 206836 267860 206888 267912
rect 211896 267860 211948 267912
rect 227444 267860 227496 267912
rect 236920 267860 236972 267912
rect 276296 267860 276348 267912
rect 288072 267860 288124 267912
rect 348148 267860 348200 267912
rect 362868 267860 362920 267912
rect 368204 267860 368256 267912
rect 369676 267860 369728 267912
rect 206744 267792 206796 267844
rect 208860 267792 208912 267844
rect 231860 267792 231912 267844
rect 235080 267792 235132 267844
rect 318800 267792 318852 267844
rect 369860 267792 369912 267844
rect 376668 267792 376720 267844
rect 391940 267792 391992 267844
rect 197176 267724 197228 267776
rect 206560 267724 206612 267776
rect 207572 267724 207624 267776
rect 223948 267724 224000 267776
rect 224040 267724 224092 267776
rect 230204 267724 230256 267776
rect 230756 267724 230808 267776
rect 238208 267724 238260 267776
rect 314844 267724 314896 267776
rect 322664 267724 322716 267776
rect 342812 267724 342864 267776
rect 352564 267724 352616 267776
rect 655888 267724 655940 267776
rect 676128 267724 676180 267776
rect 367744 267656 367796 267708
rect 531596 267656 531648 267708
rect 370504 267588 370556 267640
rect 538680 267588 538732 267640
rect 373172 267520 373224 267572
rect 545764 267520 545816 267572
rect 373540 267452 373592 267504
rect 546960 267452 547012 267504
rect 673000 267452 673052 267504
rect 676036 267452 676088 267504
rect 374460 267384 374512 267436
rect 549260 267384 549312 267436
rect 376208 267316 376260 267368
rect 554044 267316 554096 267368
rect 375840 267248 375892 267300
rect 552848 267248 552900 267300
rect 299664 267180 299716 267232
rect 350724 267180 350776 267232
rect 377128 267180 377180 267232
rect 556344 267180 556396 267232
rect 300952 267112 301004 267164
rect 354220 267112 354272 267164
rect 378508 267112 378560 267164
rect 559932 267112 559984 267164
rect 302332 267044 302384 267096
rect 357808 267044 357860 267096
rect 378876 267044 378928 267096
rect 561128 267044 561180 267096
rect 303712 266976 303764 267028
rect 361396 266976 361448 267028
rect 379796 266976 379848 267028
rect 563428 266976 563480 267028
rect 305000 266908 305052 266960
rect 364892 266908 364944 266960
rect 381636 266908 381688 266960
rect 568212 266908 568264 266960
rect 306380 266840 306432 266892
rect 368480 266840 368532 266892
rect 381176 266840 381228 266892
rect 567016 266840 567068 266892
rect 307668 266772 307720 266824
rect 371976 266772 372028 266824
rect 382464 266772 382516 266824
rect 570604 266772 570656 266824
rect 309048 266704 309100 266756
rect 375748 266704 375800 266756
rect 384304 266704 384356 266756
rect 575296 266704 575348 266756
rect 310336 266636 310388 266688
rect 379060 266636 379112 266688
rect 383844 266636 383896 266688
rect 574100 266636 574152 266688
rect 673276 266636 673328 266688
rect 676036 266636 676088 266688
rect 123760 266568 123812 266620
rect 214196 266568 214248 266620
rect 311716 266568 311768 266620
rect 382648 266568 382700 266620
rect 385132 266568 385184 266620
rect 577688 266568 577740 266620
rect 116676 266500 116728 266552
rect 211528 266500 211580 266552
rect 313004 266500 313056 266552
rect 386144 266500 386196 266552
rect 386512 266500 386564 266552
rect 581184 266500 581236 266552
rect 72976 266432 73028 266484
rect 195060 266432 195112 266484
rect 389180 266432 389232 266484
rect 588268 266432 588320 266484
rect 113180 266364 113232 266416
rect 210148 266364 210200 266416
rect 315672 266364 315724 266416
rect 68192 266296 68244 266348
rect 193220 266296 193272 266348
rect 317052 266296 317104 266348
rect 386880 266296 386932 266348
rect 392308 266364 392360 266416
rect 596548 266364 596600 266416
rect 393228 266296 393280 266348
rect 395804 266296 395856 266348
rect 606024 266296 606076 266348
rect 365076 266228 365128 266280
rect 524512 266228 524564 266280
rect 362408 266160 362460 266212
rect 517336 266160 517388 266212
rect 359740 266092 359792 266144
rect 510252 266092 510304 266144
rect 355784 266024 355836 266076
rect 499672 266024 499724 266076
rect 354404 265956 354456 266008
rect 496084 265956 496136 266008
rect 350264 265888 350316 265940
rect 485504 265888 485556 265940
rect 349068 265820 349120 265872
rect 481916 265820 481968 265872
rect 673184 265820 673236 265872
rect 676036 265820 676088 265872
rect 343732 265752 343784 265804
rect 467748 265752 467800 265804
rect 339776 265684 339828 265736
rect 457076 265684 457128 265736
rect 333520 265616 333572 265668
rect 440516 265616 440568 265668
rect 328184 265548 328236 265600
rect 426348 265548 426400 265600
rect 324136 265480 324188 265532
rect 415768 265480 415820 265532
rect 322848 265412 322900 265464
rect 412180 265412 412232 265464
rect 319720 265344 319772 265396
rect 403900 265344 403952 265396
rect 404268 265344 404320 265396
rect 448888 265344 448940 265396
rect 318340 265276 318392 265328
rect 400312 265276 400364 265328
rect 401600 265276 401652 265328
rect 463332 265276 463384 265328
rect 314384 265208 314436 265260
rect 386880 265208 386932 265260
rect 396816 265208 396868 265260
rect 389732 265140 389784 265192
rect 673092 264936 673144 264988
rect 676220 264936 676272 264988
rect 674288 264256 674340 264308
rect 676036 264256 676088 264308
rect 674472 263032 674524 263084
rect 676036 263032 676088 263084
rect 674932 262352 674984 262404
rect 675944 262352 675996 262404
rect 673644 262284 673696 262336
rect 676128 262284 676180 262336
rect 674564 262216 674616 262268
rect 676036 262216 676088 262268
rect 673828 261400 673880 261452
rect 676036 261400 676088 261452
rect 673460 260176 673512 260228
rect 675944 260176 675996 260228
rect 675024 259768 675076 259820
rect 676036 259768 676088 259820
rect 673552 259564 673604 259616
rect 675944 259564 675996 259616
rect 674748 259496 674800 259548
rect 676128 259496 676180 259548
rect 674840 259428 674892 259480
rect 676036 259428 676088 259480
rect 41788 258816 41840 258868
rect 43260 258816 43312 258868
rect 41880 257660 41932 257712
rect 51264 257660 51316 257712
rect 41604 257524 41656 257576
rect 46296 257524 46348 257576
rect 672908 256844 672960 256896
rect 678980 256844 679032 256896
rect 673736 256776 673788 256828
rect 676128 256776 676180 256828
rect 41512 256708 41564 256760
rect 56508 256708 56560 256760
rect 674656 256708 674708 256760
rect 676036 256708 676088 256760
rect 41512 256300 41564 256352
rect 43720 256300 43772 256352
rect 41512 255688 41564 255740
rect 43628 255688 43680 255740
rect 675116 255280 675168 255332
rect 675760 255280 675812 255332
rect 41512 254872 41564 254924
rect 43904 254872 43956 254924
rect 41880 254124 41932 254176
rect 43904 254124 43956 254176
rect 41880 253988 41932 254040
rect 43628 253988 43680 254040
rect 41788 253920 41840 253972
rect 43168 253920 43220 253972
rect 675484 251336 675536 251388
rect 675760 251336 675812 251388
rect 416780 251200 416832 251252
rect 567108 251200 567160 251252
rect 673368 250928 673420 250980
rect 674932 250928 674984 250980
rect 675392 250928 675444 250980
rect 674932 250792 674984 250844
rect 675484 250792 675536 250844
rect 675760 250180 675812 250232
rect 674472 249568 674524 249620
rect 675392 249568 675444 249620
rect 673828 249432 673880 249484
rect 674472 249432 674524 249484
rect 673368 249296 673420 249348
rect 673828 249296 673880 249348
rect 416780 248412 416832 248464
rect 567292 248412 567344 248464
rect 674564 247868 674616 247920
rect 675392 247868 675444 247920
rect 41512 247664 41564 247716
rect 46296 247664 46348 247716
rect 41512 247256 41564 247308
rect 45652 247256 45704 247308
rect 675024 247256 675076 247308
rect 674656 247120 674708 247172
rect 675024 247120 675076 247172
rect 675392 247052 675444 247104
rect 674748 246508 674800 246560
rect 675392 246508 675444 246560
rect 41512 246440 41564 246492
rect 48872 246440 48924 246492
rect 180708 246440 180760 246492
rect 184848 246440 184900 246492
rect 673644 246372 673696 246424
rect 674748 246372 674800 246424
rect 673644 246236 673696 246288
rect 673828 246236 673880 246288
rect 674288 246100 674340 246152
rect 675208 246100 675260 246152
rect 674840 246032 674892 246084
rect 675392 246032 675444 246084
rect 416780 245624 416832 245676
rect 564348 245624 564400 245676
rect 41696 245556 41748 245608
rect 42708 245556 42760 245608
rect 655704 245556 655756 245608
rect 674932 245556 674984 245608
rect 41880 245080 41932 245132
rect 43536 245080 43588 245132
rect 41788 244604 41840 244656
rect 43352 244604 43404 244656
rect 673644 243584 673696 243636
rect 675392 243584 675444 243636
rect 41328 242836 41380 242888
rect 43260 242836 43312 242888
rect 41420 242768 41472 242820
rect 43076 242768 43128 242820
rect 675024 242768 675076 242820
rect 675392 242768 675444 242820
rect 41236 242700 41288 242752
rect 42248 242700 42300 242752
rect 41604 242632 41656 242684
rect 43444 242632 43496 242684
rect 38568 242564 38620 242616
rect 43720 242564 43772 242616
rect 38476 242496 38528 242548
rect 43812 242496 43864 242548
rect 35808 242428 35860 242480
rect 43996 242428 44048 242480
rect 673552 242156 673604 242208
rect 675392 242156 675444 242208
rect 673736 241748 673788 241800
rect 675392 241748 675444 241800
rect 41144 240932 41196 240984
rect 673460 240524 673512 240576
rect 675392 240524 675444 240576
rect 41788 240320 41840 240372
rect 674748 238688 674800 238740
rect 675392 238688 675444 238740
rect 42156 238484 42208 238536
rect 42708 238484 42760 238536
rect 43536 237940 43588 237992
rect 43904 237940 43956 237992
rect 177948 237328 178000 237380
rect 184940 237396 184992 237448
rect 674472 236852 674524 236904
rect 675392 236852 675444 236904
rect 42248 236036 42300 236088
rect 43260 236036 43312 236088
rect 675024 235560 675076 235612
rect 675760 235560 675812 235612
rect 42340 234200 42392 234252
rect 43076 234200 43128 234252
rect 42156 233316 42208 233368
rect 43352 233316 43404 233368
rect 74448 232500 74500 232552
rect 177948 232500 178000 232552
rect 42432 232296 42484 232348
rect 43444 232296 43496 232348
rect 46020 230936 46072 230988
rect 654140 230936 654192 230988
rect 48320 230868 48372 230920
rect 656992 230868 657044 230920
rect 48228 230800 48280 230852
rect 656900 230800 656952 230852
rect 48596 230732 48648 230784
rect 659660 230732 659712 230784
rect 51172 230664 51224 230716
rect 662788 230664 662840 230716
rect 51080 230596 51132 230648
rect 662880 230596 662932 230648
rect 42432 230528 42484 230580
rect 43812 230528 43864 230580
rect 48412 230528 48464 230580
rect 659752 230528 659804 230580
rect 48780 230460 48832 230512
rect 662604 230460 662656 230512
rect 48872 230392 48924 230444
rect 662696 230392 662748 230444
rect 42156 230324 42208 230376
rect 43720 230324 43772 230376
rect 350172 230188 350224 230240
rect 423864 230188 423916 230240
rect 348792 230120 348844 230172
rect 420460 230120 420512 230172
rect 345940 230052 345992 230104
rect 414020 230052 414072 230104
rect 351644 229984 351696 230036
rect 427176 229984 427228 230036
rect 354496 229916 354548 229968
rect 433892 229916 433944 229968
rect 353024 229848 353076 229900
rect 430580 229848 430632 229900
rect 357348 229780 357400 229832
rect 440700 229780 440752 229832
rect 359832 229712 359884 229764
rect 445668 229712 445720 229764
rect 360200 229644 360252 229696
rect 447416 229644 447468 229696
rect 364432 229576 364484 229628
rect 457444 229576 457496 229628
rect 365536 229508 365588 229560
rect 459192 229508 459244 229560
rect 364064 229440 364116 229492
rect 455788 229440 455840 229492
rect 370136 229372 370188 229424
rect 470968 229372 471020 229424
rect 371240 229304 371292 229356
rect 472624 229304 472676 229356
rect 374828 229236 374880 229288
rect 483020 229236 483072 229288
rect 388352 229168 388404 229220
rect 515496 229168 515548 229220
rect 63500 229032 63552 229084
rect 74448 229100 74500 229152
rect 396908 229100 396960 229152
rect 535460 229100 535512 229152
rect 156972 229032 157024 229084
rect 237196 229032 237248 229084
rect 256976 229032 257028 229084
rect 264612 229032 264664 229084
rect 264704 229032 264756 229084
rect 273904 229032 273956 229084
rect 296352 229032 296404 229084
rect 298468 229032 298520 229084
rect 306656 229032 306708 229084
rect 323860 229032 323912 229084
rect 338028 229032 338080 229084
rect 373908 229032 373960 229084
rect 389732 229032 389784 229084
rect 469128 229032 469180 229084
rect 152832 228964 152884 229016
rect 233976 228964 234028 229016
rect 239864 228964 239916 229016
rect 265348 228964 265400 229016
rect 290740 228964 290792 229016
rect 292396 228964 292448 229016
rect 293224 228964 293276 229016
rect 294604 228964 294656 229016
rect 297456 228964 297508 229016
rect 299388 228964 299440 229016
rect 304172 228964 304224 229016
rect 314660 228964 314712 229016
rect 321652 228964 321704 229016
rect 340696 228964 340748 229016
rect 342352 228964 342404 229016
rect 362960 228964 363012 229016
rect 363052 228964 363104 229016
rect 365904 228964 365956 229016
rect 391940 228964 391992 229016
rect 472072 228964 472124 229016
rect 156144 228896 156196 228948
rect 235356 228896 235408 228948
rect 240324 228896 240376 228948
rect 269580 228896 269632 228948
rect 304540 228896 304592 228948
rect 316132 228896 316184 228948
rect 342720 228896 342772 228948
rect 380992 228896 381044 228948
rect 398288 228896 398340 228948
rect 477500 228896 477552 228948
rect 150256 228828 150308 228880
rect 234344 228828 234396 228880
rect 239956 228828 240008 228880
rect 266728 228828 266780 228880
rect 305644 228828 305696 228880
rect 317880 228828 317932 228880
rect 340880 228828 340932 228880
rect 380900 228828 380952 228880
rect 396172 228828 396224 228880
rect 474832 228828 474884 228880
rect 121184 228760 121236 228812
rect 203340 228760 203392 228812
rect 209596 228760 209648 228812
rect 258172 228760 258224 228812
rect 258264 228760 258316 228812
rect 277492 228760 277544 228812
rect 306012 228760 306064 228812
rect 319536 228760 319588 228812
rect 337752 228760 337804 228812
rect 383752 228760 383804 228812
rect 394056 228760 394108 228812
rect 474740 228760 474792 228812
rect 151728 228692 151780 228744
rect 234712 228692 234764 228744
rect 241980 228692 242032 228744
rect 272156 228692 272208 228744
rect 298836 228692 298888 228744
rect 302700 228692 302752 228744
rect 305276 228692 305328 228744
rect 320364 228692 320416 228744
rect 322020 228692 322072 228744
rect 359096 228692 359148 228744
rect 376576 228692 376628 228744
rect 466368 228692 466420 228744
rect 146024 228624 146076 228676
rect 231124 228624 231176 228676
rect 245292 228624 245344 228676
rect 273536 228624 273588 228676
rect 308864 228624 308916 228676
rect 316224 228624 316276 228676
rect 328828 228624 328880 228676
rect 345940 228624 345992 228676
rect 375472 228624 375524 228676
rect 484400 228624 484452 228676
rect 145196 228556 145248 228608
rect 231860 228556 231912 228608
rect 238484 228556 238536 228608
rect 268200 228556 268252 228608
rect 307392 228556 307444 228608
rect 322940 228556 322992 228608
rect 336648 228556 336700 228608
rect 376668 228556 376720 228608
rect 379428 228556 379480 228608
rect 494520 228556 494572 228608
rect 138480 228488 138532 228540
rect 229008 228488 229060 228540
rect 240140 228488 240192 228540
rect 271052 228488 271104 228540
rect 307760 228488 307812 228540
rect 325700 228488 325752 228540
rect 329196 228488 329248 228540
rect 375932 228488 375984 228540
rect 384396 228488 384448 228540
rect 506296 228488 506348 228540
rect 143448 228420 143500 228472
rect 231492 228420 231544 228472
rect 235264 228420 235316 228472
rect 269304 228420 269356 228472
rect 310244 228420 310296 228472
rect 329656 228420 329708 228472
rect 362960 228420 363012 228472
rect 378232 228420 378284 228472
rect 386512 228420 386564 228472
rect 511356 228420 511408 228472
rect 136824 228352 136876 228404
rect 228640 228352 228692 228404
rect 229284 228352 229336 228404
rect 267464 228352 267516 228404
rect 298744 228352 298796 228404
rect 301044 228352 301096 228404
rect 308128 228352 308180 228404
rect 327080 228352 327132 228404
rect 333428 228352 333480 228404
rect 385960 228352 386012 228404
rect 400496 228352 400548 228404
rect 544108 228352 544160 228404
rect 130108 228284 130160 228336
rect 225788 228284 225840 228336
rect 238576 228284 238628 228336
rect 270684 228284 270736 228336
rect 309508 228284 309560 228336
rect 330484 228284 330536 228336
rect 334900 228284 334952 228336
rect 389088 228284 389140 228336
rect 401876 228284 401928 228336
rect 547788 228284 547840 228336
rect 125048 228216 125100 228268
rect 223304 228216 223356 228268
rect 227720 228216 227772 228268
rect 267096 228216 267148 228268
rect 296720 228216 296772 228268
rect 300216 228216 300268 228268
rect 302792 228216 302844 228268
rect 311164 228216 311216 228268
rect 131764 228148 131816 228200
rect 226156 228148 226208 228200
rect 231676 228148 231728 228200
rect 267832 228148 267884 228200
rect 309232 228148 309284 228200
rect 328828 228216 328880 228268
rect 337016 228216 337068 228268
rect 391940 228216 391992 228268
rect 402612 228216 402664 228268
rect 549260 228216 549312 228268
rect 316224 228148 316276 228200
rect 326252 228148 326304 228200
rect 339132 228148 339184 228200
rect 393780 228148 393832 228200
rect 403624 228148 403676 228200
rect 552020 228148 552072 228200
rect 123392 228080 123444 228132
rect 222936 228080 222988 228132
rect 223488 228080 223540 228132
rect 263876 228080 263928 228132
rect 311716 228080 311768 228132
rect 332968 228080 333020 228132
rect 336280 228080 336332 228132
rect 389916 228080 389968 228132
rect 406844 228080 406896 228132
rect 559288 228080 559340 228132
rect 108212 228012 108264 228064
rect 216128 228012 216180 228064
rect 216680 228012 216732 228064
rect 261024 228012 261076 228064
rect 311348 228012 311400 228064
rect 331312 228012 331364 228064
rect 341248 228012 341300 228064
rect 396172 228012 396224 228064
rect 406200 228012 406252 228064
rect 557632 228012 557684 228064
rect 78772 227944 78824 227996
rect 193404 227944 193456 227996
rect 72056 227876 72108 227928
rect 199752 227944 199804 227996
rect 203248 227944 203300 227996
rect 255320 227944 255372 227996
rect 257712 227944 257764 227996
rect 276020 227944 276072 227996
rect 303160 227944 303212 227996
rect 312820 227944 312872 227996
rect 193588 227876 193640 227928
rect 64512 227808 64564 227860
rect 197636 227808 197688 227860
rect 199016 227876 199068 227928
rect 254676 227876 254728 227928
rect 256608 227876 256660 227928
rect 277124 227876 277176 227928
rect 301688 227876 301740 227928
rect 309416 227876 309468 227928
rect 310612 227876 310664 227928
rect 332140 227944 332192 227996
rect 338396 227944 338448 227996
rect 395252 227944 395304 227996
rect 409052 227944 409104 227996
rect 564440 227944 564492 227996
rect 202604 227808 202656 227860
rect 204076 227808 204128 227860
rect 257160 227808 257212 227860
rect 259644 227808 259696 227860
rect 278872 227808 278924 227860
rect 65340 227740 65392 227792
rect 196900 227740 196952 227792
rect 197360 227740 197412 227792
rect 254308 227740 254360 227792
rect 256148 227740 256200 227792
rect 274272 227740 274324 227792
rect 302056 227740 302108 227792
rect 311992 227740 312044 227792
rect 312728 227740 312780 227792
rect 334716 227876 334768 227928
rect 341616 227876 341668 227928
rect 400036 227876 400088 227928
rect 407212 227876 407264 227928
rect 560392 227876 560444 227928
rect 315948 227808 316000 227860
rect 338120 227808 338172 227860
rect 340604 227808 340656 227860
rect 402796 227808 402848 227860
rect 408316 227808 408368 227860
rect 562876 227808 562928 227860
rect 318800 227740 318852 227792
rect 339592 227740 339644 227792
rect 341984 227740 342036 227792
rect 403716 227740 403768 227792
rect 410432 227740 410484 227792
rect 567936 227740 567988 227792
rect 52736 227672 52788 227724
rect 192944 227672 192996 227724
rect 193036 227672 193088 227724
rect 251824 227672 251876 227724
rect 253664 227672 253716 227724
rect 276756 227672 276808 227724
rect 320272 227672 320324 227724
rect 341524 227672 341576 227724
rect 344468 227672 344520 227724
rect 410340 227672 410392 227724
rect 411536 227672 411588 227724
rect 570236 227672 570288 227724
rect 158720 227604 158772 227656
rect 237564 227604 237616 227656
rect 243636 227604 243688 227656
rect 272432 227604 272484 227656
rect 308496 227604 308548 227656
rect 324596 227604 324648 227656
rect 339500 227604 339552 227656
rect 376852 227604 376904 227656
rect 387248 227604 387300 227656
rect 460940 227604 460992 227656
rect 165436 227536 165488 227588
rect 240416 227536 240468 227588
rect 250352 227536 250404 227588
rect 275284 227536 275336 227588
rect 307024 227536 307076 227588
rect 321192 227536 321244 227588
rect 343732 227536 343784 227588
rect 378140 227536 378192 227588
rect 385132 227536 385184 227588
rect 458180 227536 458232 227588
rect 162768 227468 162820 227520
rect 238208 227468 238260 227520
rect 248696 227468 248748 227520
rect 275008 227468 275060 227520
rect 320640 227468 320692 227520
rect 356060 227468 356112 227520
rect 383016 227468 383068 227520
rect 453856 227468 453908 227520
rect 163688 227400 163740 227452
rect 240048 227400 240100 227452
rect 252008 227400 252060 227452
rect 276388 227400 276440 227452
rect 306380 227400 306432 227452
rect 322020 227400 322072 227452
rect 323124 227400 323176 227452
rect 344008 227400 344060 227452
rect 347320 227400 347372 227452
rect 411076 227400 411128 227452
rect 167092 227332 167144 227384
rect 241428 227332 241480 227384
rect 248604 227332 248656 227384
rect 268568 227332 268620 227384
rect 300952 227332 301004 227384
rect 173624 227264 173676 227316
rect 244280 227264 244332 227316
rect 253756 227264 253808 227316
rect 272800 227264 272852 227316
rect 295248 227264 295300 227316
rect 296812 227264 296864 227316
rect 297824 227264 297876 227316
rect 301872 227264 301924 227316
rect 302424 227332 302476 227384
rect 313648 227332 313700 227384
rect 332048 227332 332100 227384
rect 364340 227332 364392 227384
rect 374460 227332 374512 227384
rect 433248 227332 433300 227384
rect 310244 227264 310296 227316
rect 325976 227264 326028 227316
rect 345112 227264 345164 227316
rect 368756 227264 368808 227316
rect 425704 227264 425756 227316
rect 169576 227196 169628 227248
rect 241060 227196 241112 227248
rect 248420 227196 248472 227248
rect 269948 227196 270000 227248
rect 303528 227196 303580 227248
rect 315304 227196 315356 227248
rect 371608 227196 371660 227248
rect 430488 227196 430540 227248
rect 172152 227128 172204 227180
rect 243268 227128 243320 227180
rect 252928 227128 252980 227180
rect 271420 227128 271472 227180
rect 376208 227128 376260 227180
rect 434628 227128 434680 227180
rect 176384 227060 176436 227112
rect 243912 227060 243964 227112
rect 255228 227060 255280 227112
rect 275652 227060 275704 227112
rect 317420 227060 317472 227112
rect 337660 227060 337712 227112
rect 366180 227060 366232 227112
rect 419540 227060 419592 227112
rect 181904 226992 181956 227044
rect 246120 226992 246172 227044
rect 248512 226992 248564 227044
rect 265716 226992 265768 227044
rect 312084 226992 312136 227044
rect 335544 226992 335596 227044
rect 361580 226992 361632 227044
rect 418896 226992 418948 227044
rect 180524 226924 180576 226976
rect 247132 226924 247184 226976
rect 255596 226924 255648 226976
rect 271788 226924 271840 226976
rect 358728 226924 358780 226976
rect 411996 226924 412048 226976
rect 185584 226856 185636 226908
rect 248972 226856 249024 226908
rect 258448 226856 258500 226908
rect 274640 226856 274692 226908
rect 300676 226856 300728 226908
rect 308588 226856 308640 226908
rect 355876 226856 355928 226908
rect 408316 226856 408368 226908
rect 408684 226856 408736 226908
rect 449716 226856 449768 226908
rect 190368 226788 190420 226840
rect 251456 226788 251508 226840
rect 255412 226788 255464 226840
rect 270316 226788 270368 226840
rect 299572 226788 299624 226840
rect 306932 226788 306984 226840
rect 323492 226788 323544 226840
rect 362408 226788 362460 226840
rect 366916 226788 366968 226840
rect 408408 226788 408460 226840
rect 409696 226788 409748 226840
rect 448796 226788 448848 226840
rect 186412 226720 186464 226772
rect 248236 226720 248288 226772
rect 299204 226720 299256 226772
rect 305276 226720 305328 226772
rect 345204 226720 345256 226772
rect 376576 226720 376628 226772
rect 379796 226720 379848 226772
rect 391756 226720 391808 226772
rect 402244 226720 402296 226772
rect 441620 226720 441672 226772
rect 42156 226652 42208 226704
rect 43996 226652 44048 226704
rect 192944 226652 192996 226704
rect 251088 226652 251140 226704
rect 259368 226652 259420 226704
rect 273168 226652 273220 226704
rect 298100 226652 298152 226704
rect 303620 226652 303672 226704
rect 361212 226652 361264 226704
rect 383660 226652 383712 226704
rect 399024 226652 399076 226704
rect 436100 226652 436152 226704
rect 234712 226584 234764 226636
rect 256792 226584 256844 226636
rect 300308 226584 300360 226636
rect 306380 226584 306432 226636
rect 371976 226584 372028 226636
rect 397552 226584 397604 226636
rect 404360 226584 404412 226636
rect 438860 226584 438912 226636
rect 247040 226516 247092 226568
rect 264704 226516 264756 226568
rect 301320 226516 301372 226568
rect 307760 226516 307812 226568
rect 374092 226516 374144 226568
rect 402980 226516 403032 226568
rect 197820 226448 197872 226500
rect 207940 226448 207992 226500
rect 245660 226448 245712 226500
rect 258540 226448 258592 226500
rect 303804 226448 303856 226500
rect 317420 226448 317472 226500
rect 330576 226448 330628 226500
rect 379244 226448 379296 226500
rect 395804 226448 395856 226500
rect 422300 226448 422352 226500
rect 304908 226380 304960 226432
rect 318708 226380 318760 226432
rect 373356 226380 373408 226432
rect 397460 226380 397512 226432
rect 254676 226312 254728 226364
rect 268936 226312 268988 226364
rect 299940 226312 299992 226364
rect 304356 226312 304408 226364
rect 309876 226312 309928 226364
rect 327908 226312 327960 226364
rect 331680 226312 331732 226364
rect 347412 226312 347464 226364
rect 368020 226312 368072 226364
rect 369952 226312 370004 226364
rect 389364 226312 389416 226364
rect 411168 226312 411220 226364
rect 411902 226356 411954 226408
rect 485552 226354 485604 226406
rect 154488 226244 154540 226296
rect 235080 226244 235132 226296
rect 354128 226244 354180 226296
rect 432236 226244 432288 226296
rect 144368 226176 144420 226228
rect 230756 226176 230808 226228
rect 353760 226176 353812 226228
rect 434812 226244 434864 226296
rect 147772 226108 147824 226160
rect 232228 226108 232280 226160
rect 352288 226108 352340 226160
rect 431408 226108 431460 226160
rect 141056 226040 141108 226092
rect 229376 226040 229428 226092
rect 355508 226040 355560 226092
rect 435640 226176 435692 226228
rect 466368 226176 466420 226228
rect 487804 226176 487856 226228
rect 433248 226108 433300 226160
rect 480996 226108 481048 226160
rect 434628 226040 434680 226092
rect 487160 226040 487212 226092
rect 137652 225972 137704 226024
rect 227904 225972 227956 226024
rect 340236 225972 340288 226024
rect 370228 225972 370280 226024
rect 397460 225972 397512 226024
rect 480352 225972 480404 226024
rect 130936 225904 130988 225956
rect 225052 225904 225104 225956
rect 356612 225904 356664 225956
rect 441712 225904 441764 225956
rect 480260 225904 480312 225956
rect 502340 225904 502392 225956
rect 134248 225836 134300 225888
rect 226524 225836 226576 225888
rect 360844 225836 360896 225888
rect 451556 225836 451608 225888
rect 472072 225836 472124 225888
rect 523960 225836 524012 225888
rect 127532 225768 127584 225820
rect 223672 225768 223724 225820
rect 362316 225768 362368 225820
rect 454960 225768 455012 225820
rect 458180 225768 458232 225820
rect 507952 225768 508004 225820
rect 119160 225700 119212 225752
rect 219716 225700 219768 225752
rect 220636 225700 220688 225752
rect 249616 225700 249668 225752
rect 362684 225700 362736 225752
rect 452660 225700 452712 225752
rect 453856 225700 453908 225752
rect 503168 225700 503220 225752
rect 124128 225632 124180 225684
rect 222200 225632 222252 225684
rect 231860 225632 231912 225684
rect 253940 225632 253992 225684
rect 363696 225632 363748 225684
rect 458456 225632 458508 225684
rect 460940 225632 460992 225684
rect 513472 225632 513524 225684
rect 42432 225564 42484 225616
rect 48688 225564 48740 225616
rect 114100 225564 114152 225616
rect 217968 225564 218020 225616
rect 228456 225564 228508 225616
rect 266452 225564 266504 225616
rect 365168 225564 365220 225616
rect 461676 225564 461728 225616
rect 474740 225564 474792 225616
rect 529020 225564 529072 225616
rect 117504 225496 117556 225548
rect 219348 225496 219400 225548
rect 105728 225428 105780 225480
rect 214012 225428 214064 225480
rect 218428 225428 218480 225480
rect 262128 225496 262180 225548
rect 343088 225496 343140 225548
rect 368204 225496 368256 225548
rect 369768 225496 369820 225548
rect 468392 225496 468444 225548
rect 469128 225496 469180 225548
rect 518900 225496 518952 225548
rect 221740 225428 221792 225480
rect 263600 225428 263652 225480
rect 366548 225428 366600 225480
rect 465080 225428 465132 225480
rect 474832 225428 474884 225480
rect 533988 225428 534040 225480
rect 107384 225360 107436 225412
rect 215116 225360 215168 225412
rect 225144 225360 225196 225412
rect 264980 225360 265032 225412
rect 339868 225360 339920 225412
rect 369584 225360 369636 225412
rect 369676 225360 369728 225412
rect 469220 225360 469272 225412
rect 477500 225360 477552 225412
rect 539048 225360 539100 225412
rect 90548 225292 90600 225344
rect 197820 225292 197872 225344
rect 198188 225292 198240 225344
rect 253572 225292 253624 225344
rect 355140 225292 355192 225344
rect 103980 225224 104032 225276
rect 213644 225224 213696 225276
rect 215024 225224 215076 225276
rect 260748 225224 260800 225276
rect 313464 225224 313516 225276
rect 338856 225224 338908 225276
rect 358360 225224 358412 225276
rect 429108 225224 429160 225276
rect 436100 225292 436152 225344
rect 541440 225292 541492 225344
rect 438124 225224 438176 225276
rect 441620 225224 441672 225276
rect 546500 225224 546552 225276
rect 100668 225156 100720 225208
rect 197452 225156 197504 225208
rect 208308 225156 208360 225208
rect 95608 225088 95660 225140
rect 209688 225088 209740 225140
rect 211712 225156 211764 225208
rect 259276 225156 259328 225208
rect 314936 225156 314988 225208
rect 342444 225156 342496 225208
rect 349804 225156 349856 225208
rect 422208 225156 422260 225208
rect 422300 225156 422352 225208
rect 532792 225156 532844 225208
rect 257896 225088 257948 225140
rect 317788 225088 317840 225140
rect 348976 225088 349028 225140
rect 356980 225088 357032 225140
rect 438768 225088 438820 225140
rect 438860 225088 438912 225140
rect 554320 225088 554372 225140
rect 88892 225020 88944 225072
rect 206744 225020 206796 225072
rect 206928 225020 206980 225072
rect 256424 225020 256476 225072
rect 316316 225020 316368 225072
rect 345572 225020 345624 225072
rect 357992 225020 358044 225072
rect 444840 225020 444892 225072
rect 449716 225020 449768 225072
rect 563704 225020 563756 225072
rect 73712 224952 73764 225004
rect 200856 224952 200908 225004
rect 60280 224884 60332 224936
rect 195152 224884 195204 224936
rect 201408 224884 201460 224936
rect 255044 224952 255096 225004
rect 319168 224952 319220 225004
rect 352380 224952 352432 225004
rect 359464 224952 359516 225004
rect 448244 224952 448296 225004
rect 448796 224952 448848 225004
rect 566004 224952 566056 225004
rect 207020 224884 207072 224936
rect 252192 224884 252244 224936
rect 335176 224884 335228 224936
rect 391020 224884 391072 224936
rect 406476 224884 406528 224936
rect 559104 224884 559156 224936
rect 151084 224816 151136 224868
rect 233608 224816 233660 224868
rect 350908 224816 350960 224868
rect 428004 224816 428056 224868
rect 430488 224816 430540 224868
rect 474280 224816 474332 224868
rect 157800 224748 157852 224800
rect 236460 224748 236512 224800
rect 349436 224748 349488 224800
rect 425060 224748 425112 224800
rect 425704 224748 425756 224800
rect 467564 224748 467616 224800
rect 161204 224680 161256 224732
rect 237932 224680 237984 224732
rect 352656 224680 352708 224732
rect 428924 224680 428976 224732
rect 429108 224680 429160 224732
rect 442356 224680 442408 224732
rect 167920 224612 167972 224664
rect 240784 224612 240836 224664
rect 380900 224612 380952 224664
rect 402796 224612 402848 224664
rect 402980 224612 403032 224664
rect 479340 224612 479392 224664
rect 164608 224544 164660 224596
rect 239312 224544 239364 224596
rect 351276 224544 351328 224596
rect 425520 224544 425572 224596
rect 170956 224476 171008 224528
rect 242164 224476 242216 224528
rect 348056 224476 348108 224528
rect 174636 224408 174688 224460
rect 243360 224408 243412 224460
rect 346584 224408 346636 224460
rect 181352 224340 181404 224392
rect 246488 224340 246540 224392
rect 348424 224340 348476 224392
rect 402612 224340 402664 224392
rect 402796 224408 402848 224460
rect 404452 224408 404504 224460
rect 419540 224476 419592 224528
rect 460940 224476 460992 224528
rect 417976 224340 418028 224392
rect 421288 224340 421340 224392
rect 178040 224272 178092 224324
rect 245016 224272 245068 224324
rect 346952 224272 347004 224324
rect 415400 224272 415452 224324
rect 418896 224272 418948 224324
rect 450728 224272 450780 224324
rect 184756 224204 184808 224256
rect 247868 224204 247920 224256
rect 344100 224204 344152 224256
rect 408684 224204 408736 224256
rect 411996 224204 412048 224256
rect 444380 224204 444432 224256
rect 188160 224136 188212 224188
rect 249340 224136 249392 224188
rect 345664 224136 345716 224188
rect 412088 224136 412140 224188
rect 191472 224068 191524 224120
rect 250720 224068 250772 224120
rect 383660 224068 383712 224120
rect 449072 224068 449124 224120
rect 155408 224000 155460 224052
rect 197452 224000 197504 224052
rect 212264 224000 212316 224052
rect 214288 224000 214340 224052
rect 245384 224000 245436 224052
rect 378232 224000 378284 224052
rect 407856 224000 407908 224052
rect 408408 224000 408460 224052
rect 462504 224000 462556 224052
rect 204260 223932 204312 223984
rect 252468 223932 252520 223984
rect 376576 223932 376628 223984
rect 414572 223932 414624 223984
rect 190276 223864 190328 223916
rect 232504 223864 232556 223916
rect 378140 223864 378192 223916
rect 411260 223864 411312 223916
rect 209412 223796 209464 223848
rect 216220 223796 216272 223848
rect 246764 223796 246816 223848
rect 380992 223796 381044 223848
rect 405740 223796 405792 223848
rect 171048 223728 171100 223780
rect 206560 223728 206612 223780
rect 209688 223728 209740 223780
rect 236828 223728 236880 223780
rect 402612 223728 402664 223780
rect 418804 223728 418856 223780
rect 194876 223660 194928 223712
rect 206928 223660 206980 223712
rect 215208 223660 215260 223712
rect 242532 223660 242584 223712
rect 57980 223592 58032 223644
rect 63500 223592 63552 223644
rect 169668 223592 169720 223644
rect 180708 223592 180760 223644
rect 182180 223592 182232 223644
rect 192300 223592 192352 223644
rect 411076 223592 411128 223644
rect 417148 223592 417200 223644
rect 488448 223592 488500 223644
rect 489736 223592 489788 223644
rect 153660 223524 153712 223576
rect 222108 223524 222160 223576
rect 224408 223524 224460 223576
rect 232872 223524 232924 223576
rect 241152 223524 241204 223576
rect 253756 223524 253808 223576
rect 278688 223524 278740 223576
rect 287796 223524 287848 223576
rect 324136 223524 324188 223576
rect 361764 223524 361816 223576
rect 364340 223524 364392 223576
rect 365904 223524 365956 223576
rect 494060 223524 494112 223576
rect 607588 223524 607640 223576
rect 87144 223456 87196 223508
rect 171048 223456 171100 223508
rect 175464 223456 175516 223508
rect 244648 223456 244700 223508
rect 322388 223456 322440 223508
rect 360752 223456 360804 223508
rect 387616 223456 387668 223508
rect 513840 223456 513892 223508
rect 535460 223456 535512 223508
rect 536104 223456 536156 223508
rect 615040 223456 615092 223508
rect 148600 223388 148652 223440
rect 223856 223388 223908 223440
rect 227444 223388 227496 223440
rect 242900 223388 242952 223440
rect 323768 223388 323820 223440
rect 364340 223388 364392 223440
rect 499488 223388 499540 223440
rect 608048 223388 608100 223440
rect 146944 223320 146996 223372
rect 224132 223320 224184 223372
rect 141884 223252 141936 223304
rect 230388 223320 230440 223372
rect 237748 223320 237800 223372
rect 252928 223320 252980 223372
rect 273076 223320 273128 223372
rect 286048 223320 286100 223372
rect 324504 223320 324556 223372
rect 363236 223320 363288 223372
rect 388720 223320 388772 223372
rect 516416 223320 516468 223372
rect 541440 223320 541492 223372
rect 615960 223320 616012 223372
rect 227628 223252 227680 223304
rect 249984 223252 250036 223304
rect 325608 223252 325660 223304
rect 364984 223252 365036 223304
rect 390836 223252 390888 223304
rect 521660 223252 521712 223304
rect 538864 223252 538916 223304
rect 539324 223252 539376 223304
rect 615500 223252 615552 223304
rect 140136 223184 140188 223236
rect 230020 223184 230072 223236
rect 239404 223184 239456 223236
rect 255596 223184 255648 223236
rect 326988 223184 327040 223236
rect 368296 223184 368348 223236
rect 392952 223184 393004 223236
rect 526444 223184 526496 223236
rect 546500 223184 546552 223236
rect 548616 223184 548668 223236
rect 617340 223184 617392 223236
rect 135168 223116 135220 223168
rect 227536 223116 227588 223168
rect 227812 223116 227864 223168
rect 235724 223116 235776 223168
rect 242808 223116 242860 223168
rect 259368 223116 259420 223168
rect 274732 223116 274784 223168
rect 287060 223116 287112 223168
rect 328460 223116 328512 223168
rect 371700 223116 371752 223168
rect 395068 223116 395120 223168
rect 531504 223116 531556 223168
rect 557448 223116 557500 223168
rect 618720 223116 618772 223168
rect 133420 223048 133472 223100
rect 227168 223048 227220 223100
rect 231032 223048 231084 223100
rect 248604 223048 248656 223100
rect 271420 223048 271472 223100
rect 128360 222980 128412 223032
rect 224684 222980 224736 223032
rect 77944 222912 77996 222964
rect 121184 222912 121236 222964
rect 126704 222912 126756 222964
rect 224040 222912 224092 222964
rect 233240 222980 233292 223032
rect 236092 222980 236144 223032
rect 255412 222980 255464 223032
rect 116584 222844 116636 222896
rect 220084 222844 220136 222896
rect 223856 222844 223908 222896
rect 232688 222912 232740 222964
rect 254676 222912 254728 222964
rect 263784 222912 263836 222964
rect 280988 222912 281040 222964
rect 224316 222844 224368 222896
rect 248512 222844 248564 222896
rect 257068 222844 257120 222896
rect 278136 222844 278188 222896
rect 326344 223048 326396 223100
rect 369124 223048 369176 223100
rect 395436 223048 395488 223100
rect 532700 223048 532752 223100
rect 566004 223048 566056 223100
rect 620560 223048 620612 223100
rect 324872 222980 324924 223032
rect 365812 222980 365864 223032
rect 365904 222980 365956 223032
rect 382648 222980 382700 223032
rect 397276 222980 397328 223032
rect 536564 222980 536616 223032
rect 326620 222912 326672 222964
rect 370872 222912 370924 222964
rect 399392 222912 399444 222964
rect 541624 222912 541676 222964
rect 285680 222844 285732 222896
rect 327356 222844 327408 222896
rect 370044 222844 370096 222896
rect 370228 222844 370280 222896
rect 400404 222844 400456 222896
rect 400772 222844 400824 222896
rect 545120 222844 545172 222896
rect 568580 222844 568632 222896
rect 621020 222844 621072 222896
rect 119988 222776 120040 222828
rect 221464 222776 221516 222828
rect 222568 222776 222620 222828
rect 256976 222776 257028 222828
rect 261300 222776 261352 222828
rect 281356 222776 281408 222828
rect 325240 222776 325292 222828
rect 367468 222776 367520 222828
rect 369584 222776 369636 222828
rect 398564 222776 398616 222828
rect 400128 222776 400180 222828
rect 543648 222776 543700 222828
rect 545764 222776 545816 222828
rect 616880 222776 616932 222828
rect 91376 222708 91428 222760
rect 197268 222708 197320 222760
rect 207480 222708 207532 222760
rect 245660 222708 245712 222760
rect 266360 222708 266412 222760
rect 283196 222708 283248 222760
rect 328092 222708 328144 222760
rect 374184 222708 374236 222760
rect 401508 222708 401560 222760
rect 546684 222708 546736 222760
rect 85488 222640 85540 222692
rect 192852 222640 192904 222692
rect 82176 222572 82228 222624
rect 203984 222640 204036 222692
rect 215852 222640 215904 222692
rect 256700 222640 256752 222692
rect 260472 222640 260524 222692
rect 279608 222640 279660 222692
rect 329472 222640 329524 222692
rect 377588 222640 377640 222692
rect 403348 222640 403400 222692
rect 549352 222640 549404 222692
rect 563704 222640 563756 222692
rect 620100 222640 620152 222692
rect 193128 222572 193180 222624
rect 201316 222572 201368 222624
rect 209136 222572 209188 222624
rect 258908 222572 258960 222624
rect 262956 222572 263008 222624
rect 281724 222572 281776 222624
rect 75368 222504 75420 222556
rect 201132 222504 201184 222556
rect 205824 222504 205876 222556
rect 257528 222504 257580 222556
rect 262128 222504 262180 222556
rect 280712 222504 280764 222556
rect 72884 222436 72936 222488
rect 193128 222436 193180 222488
rect 193220 222436 193272 222488
rect 195796 222436 195848 222488
rect 202420 222436 202472 222488
rect 256056 222436 256108 222488
rect 257896 222436 257948 222488
rect 279976 222436 280028 222488
rect 68652 222368 68704 222420
rect 198280 222368 198332 222420
rect 200764 222368 200816 222420
rect 255688 222368 255740 222420
rect 272248 222368 272300 222420
rect 284944 222572 284996 222624
rect 329840 222572 329892 222624
rect 375380 222572 375432 222624
rect 376668 222572 376720 222624
rect 394700 222572 394752 222624
rect 403256 222572 403308 222624
rect 549996 222572 550048 222624
rect 553768 222572 553820 222624
rect 561220 222572 561272 222624
rect 619640 222572 619692 222624
rect 283196 222504 283248 222556
rect 290280 222504 290332 222556
rect 331588 222504 331640 222556
rect 378416 222504 378468 222556
rect 404728 222504 404780 222556
rect 554228 222504 554280 222556
rect 554320 222504 554372 222556
rect 618260 222504 618312 222556
rect 327724 222436 327776 222488
rect 372620 222436 372672 222488
rect 373908 222436 373960 222488
rect 397736 222436 397788 222488
rect 405832 222436 405884 222488
rect 556712 222436 556764 222488
rect 559104 222436 559156 222488
rect 619180 222436 619232 222488
rect 332692 222368 332744 222420
rect 351920 222368 351972 222420
rect 352012 222368 352064 222420
rect 376760 222368 376812 222420
rect 376852 222368 376904 222420
rect 401140 222368 401192 222420
rect 405096 222368 405148 222420
rect 555056 222368 555108 222420
rect 562876 222368 562928 222420
rect 634544 222368 634596 222420
rect 53564 222300 53616 222352
rect 182180 222300 182232 222352
rect 187240 222300 187292 222352
rect 227628 222300 227680 222352
rect 259368 222300 259420 222352
rect 280344 222300 280396 222352
rect 310980 222300 311032 222352
rect 333980 222300 334032 222352
rect 334164 222300 334216 222352
rect 385132 222300 385184 222352
rect 405464 222300 405516 222352
rect 556252 222300 556304 222352
rect 557448 222300 557500 222352
rect 557632 222300 557684 222352
rect 633624 222300 633676 222352
rect 61936 222232 61988 222284
rect 195428 222232 195480 222284
rect 195704 222232 195756 222284
rect 253204 222232 253256 222284
rect 254584 222232 254636 222284
rect 278504 222232 278556 222284
rect 337384 222232 337436 222284
rect 59452 222164 59504 222216
rect 193220 222164 193272 222216
rect 194048 222164 194100 222216
rect 252836 222164 252888 222216
rect 255412 222164 255464 222216
rect 277860 222164 277912 222216
rect 314200 222164 314252 222216
rect 338028 222164 338080 222216
rect 338120 222164 338172 222216
rect 343088 222164 343140 222216
rect 351920 222232 351972 222284
rect 381820 222232 381872 222284
rect 396172 222232 396224 222284
rect 401968 222232 402020 222284
rect 409328 222232 409380 222284
rect 565176 222232 565228 222284
rect 393596 222164 393648 222216
rect 400036 222164 400088 222216
rect 403624 222164 403676 222216
rect 543648 222164 543700 222216
rect 616420 222164 616472 222216
rect 155316 222096 155368 222148
rect 219992 222096 220044 222148
rect 220084 222096 220136 222148
rect 234620 222096 234672 222148
rect 269672 222096 269724 222148
rect 284576 222096 284628 222148
rect 320916 222096 320968 222148
rect 357348 222096 357400 222148
rect 384028 222096 384080 222148
rect 505744 222096 505796 222148
rect 532792 222096 532844 222148
rect 533436 222096 533488 222148
rect 614580 222096 614632 222148
rect 93768 222028 93820 222080
rect 155408 222028 155460 222080
rect 160376 222028 160428 222080
rect 238300 222028 238352 222080
rect 244464 222028 244516 222080
rect 256148 222028 256200 222080
rect 319812 222028 319864 222080
rect 354036 222028 354088 222080
rect 383384 222028 383436 222080
rect 503720 222028 503772 222080
rect 552572 222028 552624 222080
rect 553216 222028 553268 222080
rect 632704 222028 632756 222080
rect 162032 221960 162084 222012
rect 238944 221960 238996 222012
rect 322756 221960 322808 222012
rect 358268 221960 358320 222012
rect 381912 221960 381964 222012
rect 501052 221960 501104 222012
rect 547788 221960 547840 222012
rect 631784 221960 631836 222012
rect 170496 221892 170548 221944
rect 227444 221892 227496 221944
rect 168748 221824 168800 221876
rect 241796 221892 241848 221944
rect 275560 221892 275612 221944
rect 286416 221892 286468 221944
rect 316684 221892 316736 221944
rect 347320 221892 347372 221944
rect 347412 221892 347464 221944
rect 380072 221892 380124 221944
rect 382280 221892 382332 221944
rect 501236 221892 501288 221944
rect 530676 221892 530728 221944
rect 614028 221892 614080 221944
rect 166264 221756 166316 221808
rect 239680 221824 239732 221876
rect 321284 221824 321336 221876
rect 354864 221824 354916 221876
rect 380532 221824 380584 221876
rect 497372 221824 497424 221876
rect 499488 221824 499540 221876
rect 528100 221824 528152 221876
rect 613568 221824 613620 221876
rect 234344 221756 234396 221808
rect 248420 221756 248472 221808
rect 278136 221756 278188 221808
rect 288532 221756 288584 221808
rect 319904 221756 319956 221808
rect 351460 221756 351512 221808
rect 377956 221756 378008 221808
rect 491300 221756 491352 221808
rect 542728 221756 542780 221808
rect 630864 221756 630916 221808
rect 177212 221688 177264 221740
rect 245752 221688 245804 221740
rect 281448 221688 281500 221740
rect 289912 221688 289964 221740
rect 318064 221688 318116 221740
rect 350632 221688 350684 221740
rect 380808 221688 380860 221740
rect 497832 221688 497884 221740
rect 538312 221688 538364 221740
rect 540152 221688 540204 221740
rect 630404 221688 630456 221740
rect 183928 221620 183980 221672
rect 248328 221620 248380 221672
rect 264612 221620 264664 221672
rect 282828 221620 282880 221672
rect 317052 221620 317104 221672
rect 345020 221620 345072 221672
rect 345940 221620 345992 221672
rect 373356 221620 373408 221672
rect 377680 221620 377732 221672
rect 490288 221620 490340 221672
rect 534908 221620 534960 221672
rect 629484 221620 629536 221672
rect 182088 221552 182140 221604
rect 188988 221484 189040 221536
rect 159548 221416 159600 221468
rect 209688 221416 209740 221468
rect 178868 221348 178920 221400
rect 181904 221348 181956 221400
rect 181996 221348 182048 221400
rect 215208 221348 215260 221400
rect 219992 221484 220044 221536
rect 235816 221484 235868 221536
rect 258816 221552 258868 221604
rect 279240 221552 279292 221604
rect 283932 221552 283984 221604
rect 289544 221552 289596 221604
rect 318432 221552 318484 221604
rect 348148 221552 348200 221604
rect 379060 221552 379112 221604
rect 494060 221552 494112 221604
rect 530124 221552 530176 221604
rect 628472 221552 628524 221604
rect 247500 221484 247552 221536
rect 273904 221484 273956 221536
rect 285312 221484 285364 221536
rect 286508 221484 286560 221536
rect 291752 221484 291804 221536
rect 314568 221484 314620 221536
rect 339684 221484 339736 221536
rect 345112 221484 345164 221536
rect 366640 221484 366692 221536
rect 375104 221484 375156 221536
rect 483572 221484 483624 221536
rect 510620 221484 510672 221536
rect 610348 221484 610400 221536
rect 219900 221416 219952 221468
rect 245844 221416 245896 221468
rect 249524 221416 249576 221468
rect 257712 221416 257764 221468
rect 268844 221416 268896 221468
rect 283564 221416 283616 221468
rect 288256 221416 288308 221468
rect 292764 221416 292816 221468
rect 315212 221416 315264 221468
rect 343916 221416 343968 221468
rect 344008 221416 344060 221468
rect 359924 221416 359976 221468
rect 372988 221416 373040 221468
rect 477776 221416 477828 221468
rect 525064 221416 525116 221468
rect 627552 221416 627604 221468
rect 250076 221348 250128 221400
rect 251088 221348 251140 221400
rect 256608 221348 256660 221400
rect 267188 221348 267240 221400
rect 282460 221348 282512 221400
rect 289084 221348 289136 221400
rect 292120 221348 292172 221400
rect 292396 221348 292448 221400
rect 293500 221348 293552 221400
rect 313832 221348 313884 221400
rect 340604 221348 340656 221400
rect 340696 221348 340748 221400
rect 356520 221348 356572 221400
rect 367284 221348 367336 221400
rect 464252 221348 464304 221400
rect 505744 221348 505796 221400
rect 609428 221348 609480 221400
rect 149428 221280 149480 221332
rect 190276 221280 190328 221332
rect 199936 221280 199988 221332
rect 231860 221280 231912 221332
rect 236920 221280 236972 221332
rect 240324 221280 240376 221332
rect 247868 221280 247920 221332
rect 255228 221280 255280 221332
rect 256240 221280 256292 221332
rect 259644 221280 259696 221332
rect 280620 221280 280672 221332
rect 288164 221280 288216 221332
rect 289728 221280 289780 221332
rect 293132 221280 293184 221332
rect 294972 221280 295024 221332
rect 295616 221280 295668 221332
rect 315580 221280 315632 221332
rect 341432 221280 341484 221332
rect 341524 221280 341576 221332
rect 353300 221280 353352 221332
rect 365996 221280 366048 221332
rect 454132 221280 454184 221332
rect 501052 221280 501104 221332
rect 608508 221280 608560 221332
rect 179696 221212 179748 221264
rect 214288 221212 214340 221264
rect 226800 221212 226852 221264
rect 239864 221212 239916 221264
rect 252928 221212 252980 221264
rect 258264 221212 258316 221264
rect 270408 221212 270460 221264
rect 283840 221212 283892 221264
rect 284852 221212 284904 221264
rect 291384 221212 291436 221264
rect 291568 221212 291620 221264
rect 294236 221212 294288 221264
rect 312360 221212 312412 221264
rect 337200 221212 337252 221264
rect 337660 221212 337712 221264
rect 346492 221212 346544 221264
rect 389916 221212 389968 221264
rect 392676 221212 392728 221264
rect 397552 221212 397604 221264
rect 476856 221212 476908 221264
rect 518992 221212 519044 221264
rect 520004 221212 520056 221264
rect 626632 221212 626684 221264
rect 172980 221144 173032 221196
rect 181996 221144 182048 221196
rect 183100 221144 183152 221196
rect 216220 221144 216272 221196
rect 246120 221144 246172 221196
rect 258448 221144 258500 221196
rect 276480 221144 276532 221196
rect 287428 221144 287480 221196
rect 330208 221144 330260 221196
rect 189816 221076 189868 221128
rect 220636 221076 220688 221128
rect 192300 221008 192352 221060
rect 193036 221008 193088 221060
rect 192852 220940 192904 220992
rect 205456 221008 205508 221060
rect 206652 221008 206704 221060
rect 234712 221076 234764 221128
rect 277308 221076 277360 221128
rect 286692 221076 286744 221128
rect 230204 221008 230256 221060
rect 239956 221008 240008 221060
rect 265532 221008 265584 221060
rect 282092 221008 282144 221060
rect 282368 221008 282420 221060
rect 289268 221076 289320 221128
rect 313096 221076 313148 221128
rect 336740 221076 336792 221128
rect 339592 221144 339644 221196
rect 349804 221144 349856 221196
rect 368204 221144 368256 221196
rect 352012 221076 352064 221128
rect 383752 221076 383804 221128
rect 396080 221076 396132 221128
rect 403716 221144 403768 221196
rect 406200 221144 406252 221196
rect 408316 221144 408368 221196
rect 437296 221144 437348 221196
rect 513380 221144 513432 221196
rect 514944 221144 514996 221196
rect 625712 221144 625764 221196
rect 655796 221144 655848 221196
rect 675944 221144 675996 221196
rect 407028 221076 407080 221128
rect 407948 221076 408000 221128
rect 561772 221076 561824 221128
rect 287336 221008 287388 221060
rect 291016 221008 291068 221060
rect 386236 221008 386288 221060
rect 510620 221008 510672 221060
rect 549352 221008 549404 221060
rect 551100 221008 551152 221060
rect 617800 221008 617852 221060
rect 655612 221008 655664 221060
rect 676036 221008 676088 221060
rect 197268 220940 197320 220992
rect 209044 220940 209096 220992
rect 213368 220940 213420 220992
rect 234804 220940 234856 220992
rect 268016 220940 268068 220992
rect 284208 220940 284260 220992
rect 285680 220940 285732 220992
rect 290648 220940 290700 220992
rect 385500 220940 385552 220992
rect 508780 220940 508832 220992
rect 509608 220940 509660 220992
rect 624792 220940 624844 220992
rect 279792 220872 279844 220924
rect 288900 220872 288952 220924
rect 393780 220872 393832 220924
rect 399484 220872 399536 220924
rect 504824 220872 504876 220924
rect 623872 220872 623924 220924
rect 196532 220804 196584 220856
rect 204260 220804 204312 220856
rect 204904 220804 204956 220856
rect 206836 220804 206888 220856
rect 233516 220804 233568 220856
rect 238484 220804 238536 220856
rect 499304 220804 499356 220856
rect 622952 220804 623004 220856
rect 655520 220804 655572 220856
rect 675852 220804 675904 220856
rect 350540 220736 350592 220788
rect 426348 220736 426400 220788
rect 675208 220736 675260 220788
rect 676036 220736 676088 220788
rect 352104 220668 352156 220720
rect 429752 220668 429804 220720
rect 353392 220600 353444 220652
rect 433340 220600 433392 220652
rect 355048 220532 355100 220584
rect 436468 220532 436520 220584
rect 356244 220464 356296 220516
rect 439780 220464 439832 220516
rect 359372 220396 359424 220448
rect 446588 220396 446640 220448
rect 357716 220328 357768 220380
rect 443184 220328 443236 220380
rect 361948 220260 362000 220312
rect 453304 220260 453356 220312
rect 142712 220192 142764 220244
rect 229652 220192 229704 220244
rect 360568 220192 360620 220244
rect 449900 220192 449952 220244
rect 139308 220124 139360 220176
rect 228272 220124 228324 220176
rect 364800 220124 364852 220176
rect 460020 220124 460072 220176
rect 135996 220056 136048 220108
rect 226616 220056 226668 220108
rect 363420 220056 363472 220108
rect 456616 220056 456668 220108
rect 132408 219988 132460 220040
rect 225420 219988 225472 220040
rect 368388 219988 368440 220040
rect 465908 219988 465960 220040
rect 129280 219920 129332 219972
rect 223764 219920 223816 219972
rect 367652 219920 367704 219972
rect 466736 219920 466788 219972
rect 125876 219852 125928 219904
rect 222292 219852 222344 219904
rect 366272 219852 366324 219904
rect 463700 219852 463752 219904
rect 122472 219784 122524 219836
rect 221096 219784 221148 219836
rect 370504 219784 370556 219836
rect 473452 219784 473504 219836
rect 58624 219716 58676 219768
rect 193772 219716 193824 219768
rect 369308 219716 369360 219768
rect 470140 219716 470192 219768
rect 45468 219648 45520 219700
rect 648528 219648 648580 219700
rect 45560 219580 45612 219632
rect 649908 219580 649960 219632
rect 45744 219512 45796 219564
rect 651288 219512 651340 219564
rect 45836 219444 45888 219496
rect 652760 219444 652812 219496
rect 45928 219376 45980 219428
rect 654140 219376 654192 219428
rect 347688 219308 347740 219360
rect 419724 219308 419776 219360
rect 349160 219240 349212 219292
rect 423036 219240 423088 219292
rect 346308 219172 346360 219224
rect 416228 219172 416280 219224
rect 344836 219104 344888 219156
rect 412916 219104 412968 219156
rect 343456 219036 343508 219088
rect 409512 219036 409564 219088
rect 666560 218560 666612 218612
rect 666836 218560 666888 218612
rect 525800 218424 525852 218476
rect 613108 218424 613160 218476
rect 523408 218356 523460 218408
rect 612648 218356 612700 218408
rect 520832 218288 520884 218340
rect 612188 218288 612240 218340
rect 674564 218288 674616 218340
rect 676036 218288 676088 218340
rect 518624 218220 518676 218272
rect 611728 218220 611780 218272
rect 515496 218152 515548 218204
rect 611268 218152 611320 218204
rect 490288 218084 490340 218136
rect 607128 218084 607180 218136
rect 487160 218016 487212 218068
rect 606668 218016 606720 218068
rect 674840 218016 674892 218068
rect 676036 218016 676088 218068
rect 418160 217948 418212 218000
rect 418620 217948 418672 218000
rect 213874 217608 213926 217660
rect 219900 217608 219952 217660
rect 492266 217540 492318 217592
rect 622032 217540 622084 217592
rect 24952 217472 25004 217524
rect 665732 217472 665784 217524
rect 570880 217404 570932 217456
rect 635924 217404 635976 217456
rect 568304 217336 568356 217388
rect 635464 217336 635516 217388
rect 565636 217268 565688 217320
rect 635004 217268 635056 217320
rect 560760 217200 560812 217252
rect 634084 217200 634136 217252
rect 555700 217132 555752 217184
rect 633164 217132 633216 217184
rect 508596 217064 508648 217116
rect 533068 217064 533120 217116
rect 550456 217064 550508 217116
rect 632244 217064 632296 217116
rect 418528 216996 418580 217048
rect 639696 216996 639748 217048
rect 418620 216928 418672 216980
rect 640156 216928 640208 216980
rect 418436 216860 418488 216912
rect 640616 216860 640668 216912
rect 52184 216792 52236 216844
rect 57980 216792 58032 216844
rect 417884 216792 417936 216844
rect 641076 216792 641128 216844
rect 52276 216724 52328 216776
rect 169668 216724 169720 216776
rect 187608 216724 187660 216776
rect 603448 216724 603500 216776
rect 46296 216656 46348 216708
rect 664812 216656 664864 216708
rect 673828 216656 673880 216708
rect 676036 216656 676088 216708
rect 45652 216588 45704 216640
rect 664352 216588 664404 216640
rect 503536 216520 503588 216572
rect 524052 216520 524104 216572
rect 532976 216520 533028 216572
rect 502708 216452 502760 216504
rect 486700 216384 486752 216436
rect 490104 216384 490156 216436
rect 493232 216384 493284 216436
rect 507768 216384 507820 216436
rect 512828 216384 512880 216436
rect 513656 216384 513708 216436
rect 517888 216384 517940 216436
rect 522856 216384 522908 216436
rect 524052 216384 524104 216436
rect 527916 216384 527968 216436
rect 533068 216384 533120 216436
rect 545580 216520 545632 216572
rect 631324 216520 631376 216572
rect 538036 216452 538088 216504
rect 629944 216452 629996 216504
rect 628932 216384 628984 216436
rect 610808 216316 610860 216368
rect 609888 216248 609940 216300
rect 673552 216248 673604 216300
rect 675944 216248 675996 216300
rect 628012 216180 628064 216232
rect 608968 216112 609020 216164
rect 627092 216044 627144 216096
rect 626172 215976 626224 216028
rect 625252 215908 625304 215960
rect 623412 215840 623464 215892
rect 624332 215772 624384 215824
rect 580908 215704 580960 215756
rect 638776 215704 638828 215756
rect 636936 215636 636988 215688
rect 636384 215568 636436 215620
rect 638316 215500 638368 215552
rect 673460 215500 673512 215552
rect 675576 215500 675628 215552
rect 25136 215432 25188 215484
rect 666192 215432 666244 215484
rect 674472 215432 674524 215484
rect 675852 215432 675904 215484
rect 24860 215364 24912 215416
rect 665272 215364 665324 215416
rect 674656 215364 674708 215416
rect 675944 215364 675996 215416
rect 582288 215296 582340 215348
rect 599860 215296 599912 215348
rect 603448 215296 603500 215348
rect 604368 215296 604420 215348
rect 639236 215296 639288 215348
rect 674932 215296 674984 215348
rect 676036 215296 676088 215348
rect 41512 215092 41564 215144
rect 46204 215092 46256 215144
rect 41512 214684 41564 214736
rect 46112 214684 46164 214736
rect 41512 214276 41564 214328
rect 50988 214276 51040 214328
rect 41512 214072 41564 214124
rect 43536 214072 43588 214124
rect 33048 213596 33100 213648
rect 32956 213528 33008 213580
rect 32864 213460 32916 213512
rect 41512 213392 41564 213444
rect 659660 215092 659712 215144
rect 660764 215092 660816 215144
rect 673736 214616 673788 214668
rect 676036 214616 676088 214668
rect 673644 213800 673696 213852
rect 675944 213800 675996 213852
rect 670884 213596 670936 213648
rect 671804 213528 671856 213580
rect 673092 213460 673144 213512
rect 671896 213392 671948 213444
rect 580172 212576 580224 212628
rect 598940 212576 598992 212628
rect 674288 212576 674340 212628
rect 675944 212576 675996 212628
rect 580448 212508 580500 212560
rect 599952 212508 600004 212560
rect 674748 212508 674800 212560
rect 676036 212508 676088 212560
rect 655428 212440 655480 212492
rect 669688 212440 669740 212492
rect 41512 212236 41564 212288
rect 43168 212236 43220 212288
rect 41512 212100 41564 212152
rect 43628 212100 43680 212152
rect 673000 212032 673052 212084
rect 676036 212032 676088 212084
rect 662696 210060 662748 210112
rect 663524 210060 663576 210112
rect 582288 209856 582340 209908
rect 599124 209856 599176 209908
rect 580080 209788 580132 209840
rect 601148 209788 601200 209840
rect 641812 209788 641864 209840
rect 642088 209788 642140 209840
rect 644664 209788 644716 209840
rect 644940 209788 644992 209840
rect 647424 209788 647476 209840
rect 647700 209788 647752 209840
rect 675024 208360 675076 208412
rect 675300 208360 675352 208412
rect 675116 208292 675168 208344
rect 675392 208292 675444 208344
rect 41512 208224 41564 208276
rect 43352 208224 43404 208276
rect 674840 208224 674892 208276
rect 675300 208224 675352 208276
rect 41512 207272 41564 207324
rect 43444 207272 43496 207324
rect 41788 207136 41840 207188
rect 43720 207136 43772 207188
rect 582288 207068 582340 207120
rect 601516 207068 601568 207120
rect 579804 207000 579856 207052
rect 600964 207000 601016 207052
rect 666928 206932 666980 206984
rect 675392 206932 675444 206984
rect 674840 206252 674892 206304
rect 675760 206252 675812 206304
rect 673368 206184 673420 206236
rect 675484 206184 675536 206236
rect 675668 206184 675720 206236
rect 674564 205164 674616 205216
rect 675300 205164 675352 205216
rect 674564 205028 674616 205080
rect 674932 204960 674984 205012
rect 675392 204960 675444 205012
rect 581460 204280 581512 204332
rect 599952 204280 600004 204332
rect 675116 203872 675168 203924
rect 675300 203872 675352 203924
rect 674840 203804 674892 203856
rect 675116 203736 675168 203788
rect 674288 203668 674340 203720
rect 674840 203668 674892 203720
rect 673828 202716 673880 202768
rect 675392 202716 675444 202768
rect 674656 202036 674708 202088
rect 675392 202036 675444 202088
rect 582288 201560 582340 201612
rect 599952 201560 600004 201612
rect 580632 201492 580684 201544
rect 598940 201492 598992 201544
rect 674472 201492 674524 201544
rect 675392 201492 675444 201544
rect 38016 201424 38068 201476
rect 43536 201424 43588 201476
rect 41420 201356 41472 201408
rect 43076 201356 43128 201408
rect 674748 200880 674800 200932
rect 675392 200880 675444 200932
rect 673552 200744 673604 200796
rect 674748 200744 674800 200796
rect 30196 200608 30248 200660
rect 42708 200608 42760 200660
rect 30288 200472 30340 200524
rect 42248 200472 42300 200524
rect 582288 200064 582340 200116
rect 599952 200064 600004 200116
rect 41604 199112 41656 199164
rect 43168 199112 43220 199164
rect 41696 198976 41748 199028
rect 43260 198976 43312 199028
rect 41788 198908 41840 198960
rect 43628 198908 43680 198960
rect 41512 198772 41564 198824
rect 42340 198772 42392 198824
rect 581092 198704 581144 198756
rect 599124 198704 599176 198756
rect 673460 198364 673512 198416
rect 675392 198364 675444 198416
rect 673644 197752 673696 197804
rect 675484 197752 675536 197804
rect 582288 197344 582340 197396
rect 599308 197344 599360 197396
rect 580724 197276 580776 197328
rect 599952 197276 600004 197328
rect 673736 197004 673788 197056
rect 675392 197004 675444 197056
rect 42248 196528 42300 196580
rect 42708 196528 42760 196580
rect 674840 196528 674892 196580
rect 675392 196528 675444 196580
rect 673552 195304 673604 195356
rect 675392 195304 675444 195356
rect 582196 194624 582248 194676
rect 599124 194624 599176 194676
rect 582288 194556 582340 194608
rect 599952 194556 600004 194608
rect 42064 193468 42116 193520
rect 43076 193468 43128 193520
rect 674472 192788 674524 192840
rect 675300 192788 675352 192840
rect 582196 191836 582248 191888
rect 599124 191836 599176 191888
rect 582288 191768 582340 191820
rect 599952 191768 600004 191820
rect 42340 191632 42392 191684
rect 43168 191632 43220 191684
rect 674748 191632 674800 191684
rect 675392 191632 675444 191684
rect 42064 191428 42116 191480
rect 43260 191428 43312 191480
rect 581368 190408 581420 190460
rect 599860 190408 599912 190460
rect 42248 190136 42300 190188
rect 43444 190136 43496 190188
rect 42156 190068 42208 190120
rect 43536 190068 43588 190120
rect 42432 189116 42484 189168
rect 43352 189116 43404 189168
rect 42156 187824 42208 187876
rect 43628 187824 43680 187876
rect 582196 187620 582248 187672
rect 601608 187620 601660 187672
rect 582288 187552 582340 187604
rect 600964 187552 601016 187604
rect 42156 187144 42208 187196
rect 43720 187144 43772 187196
rect 579804 184832 579856 184884
rect 599952 184832 600004 184884
rect 582288 184764 582340 184816
rect 601516 184764 601568 184816
rect 42156 182112 42208 182164
rect 48504 182112 48556 182164
rect 580172 182112 580224 182164
rect 599860 182112 599912 182164
rect 582288 182044 582340 182096
rect 600044 182044 600096 182096
rect 580540 179324 580592 179376
rect 599768 179324 599820 179376
rect 580264 179256 580316 179308
rect 599952 179256 600004 179308
rect 669412 178780 669464 178832
rect 676220 178780 676272 178832
rect 675208 178576 675260 178628
rect 676036 178576 676088 178628
rect 669504 178100 669556 178152
rect 675944 178100 675996 178152
rect 669596 177692 669648 177744
rect 675944 177692 675996 177744
rect 671712 176808 671764 176860
rect 676036 176808 676088 176860
rect 581276 176672 581328 176724
rect 598940 176672 598992 176724
rect 580540 176604 580592 176656
rect 599860 176604 599912 176656
rect 675116 176604 675168 176656
rect 676036 176604 676088 176656
rect 580816 176536 580868 176588
rect 600136 176536 600188 176588
rect 675024 176332 675076 176384
rect 676036 176332 676088 176384
rect 673184 175992 673236 176044
rect 675944 175992 675996 176044
rect 673276 175176 673328 175228
rect 675944 175176 675996 175228
rect 673368 174360 673420 174412
rect 676036 174360 676088 174412
rect 581000 173884 581052 173936
rect 599952 173884 600004 173936
rect 674564 173884 674616 173936
rect 676036 173884 676088 173936
rect 582288 173816 582340 173868
rect 599676 173816 599728 173868
rect 582196 173748 582248 173800
rect 600044 173748 600096 173800
rect 673552 172864 673604 172916
rect 676036 172864 676088 172916
rect 673736 172048 673788 172100
rect 675944 172048 675996 172100
rect 674748 171640 674800 171692
rect 675944 171640 675996 171692
rect 582012 171164 582064 171216
rect 599952 171164 600004 171216
rect 674932 171164 674984 171216
rect 675944 171164 675996 171216
rect 579896 171096 579948 171148
rect 599860 171096 599912 171148
rect 675024 171096 675076 171148
rect 676036 171096 676088 171148
rect 582288 171028 582340 171080
rect 599768 171028 599820 171080
rect 674288 169600 674340 169652
rect 675944 169600 675996 169652
rect 673644 169192 673696 169244
rect 675852 169192 675904 169244
rect 673828 168580 673880 168632
rect 675760 168580 675812 168632
rect 579804 168512 579856 168564
rect 599952 168512 600004 168564
rect 674472 168512 674524 168564
rect 675852 168512 675904 168564
rect 581736 168444 581788 168496
rect 599032 168444 599084 168496
rect 674840 168444 674892 168496
rect 675944 168444 675996 168496
rect 579712 168376 579764 168428
rect 599860 168376 599912 168428
rect 675208 168376 675260 168428
rect 676036 168376 676088 168428
rect 581460 168308 581512 168360
rect 600320 168308 600372 168360
rect 671988 167016 672040 167068
rect 676036 167016 676088 167068
rect 666560 165928 666612 165980
rect 666928 165928 666980 165980
rect 582288 165724 582340 165776
rect 599860 165724 599912 165776
rect 581920 165656 581972 165708
rect 600044 165656 600096 165708
rect 581828 165588 581880 165640
rect 599952 165588 600004 165640
rect 580264 165520 580316 165572
rect 600136 165520 600188 165572
rect 582104 162936 582156 162988
rect 599860 162936 599912 162988
rect 581460 162868 581512 162920
rect 599952 162868 600004 162920
rect 675116 160488 675168 160540
rect 675392 160488 675444 160540
rect 675024 160352 675076 160404
rect 581276 160216 581328 160268
rect 599860 160216 599912 160268
rect 581000 160148 581052 160200
rect 599952 160148 600004 160200
rect 674748 160148 674800 160200
rect 675300 160148 675352 160200
rect 581368 160080 581420 160132
rect 599308 160080 599360 160132
rect 674932 160080 674984 160132
rect 675024 160012 675076 160064
rect 675392 160012 675444 160064
rect 674932 159944 674984 159996
rect 674840 159740 674892 159792
rect 674564 159536 674616 159588
rect 675484 159536 675536 159588
rect 581552 157496 581604 157548
rect 599952 157496 600004 157548
rect 581092 157428 581144 157480
rect 600044 157428 600096 157480
rect 580724 157360 580776 157412
rect 599860 157360 599912 157412
rect 666836 157292 666888 157344
rect 675116 157292 675168 157344
rect 674472 155252 674524 155304
rect 675116 155252 675168 155304
rect 673736 155184 673788 155236
rect 675208 155184 675260 155236
rect 581184 154640 581236 154692
rect 599952 154640 600004 154692
rect 580448 154572 580500 154624
rect 599860 154572 599912 154624
rect 674288 152192 674340 152244
rect 675116 152192 675168 152244
rect 673828 152124 673880 152176
rect 675208 152124 675260 152176
rect 673644 152056 673696 152108
rect 675300 152056 675352 152108
rect 582196 151920 582248 151972
rect 599308 151920 599360 151972
rect 580816 151852 580868 151904
rect 599952 151852 600004 151904
rect 580632 151784 580684 151836
rect 599860 151784 599912 151836
rect 582012 149200 582064 149252
rect 599768 149200 599820 149252
rect 582288 149132 582340 149184
rect 598940 149132 598992 149184
rect 581828 149064 581880 149116
rect 599952 149064 600004 149116
rect 673552 148452 673604 148504
rect 675392 148452 675444 148504
rect 581644 146344 581696 146396
rect 599952 146344 600004 146396
rect 580540 146276 580592 146328
rect 599860 146276 599912 146328
rect 582104 143692 582156 143744
rect 600044 143692 600096 143744
rect 581736 143624 581788 143676
rect 599860 143624 599912 143676
rect 581460 143556 581512 143608
rect 599952 143556 600004 143608
rect 581920 140904 581972 140956
rect 599860 140904 599912 140956
rect 581276 140836 581328 140888
rect 599952 140836 600004 140888
rect 581000 140768 581052 140820
rect 599308 140768 599360 140820
rect 581552 138116 581604 138168
rect 599860 138116 599912 138168
rect 581092 138048 581144 138100
rect 599952 138048 600004 138100
rect 579896 137980 579948 138032
rect 600044 137980 600096 138032
rect 581368 135328 581420 135380
rect 599860 135328 599912 135380
rect 579988 135260 580040 135312
rect 599952 135260 600004 135312
rect 669688 132880 669740 132932
rect 676036 132880 676088 132932
rect 669320 132744 669372 132796
rect 676220 132744 676272 132796
rect 580908 132608 580960 132660
rect 599860 132608 599912 132660
rect 669228 132608 669280 132660
rect 676128 132608 676180 132660
rect 580448 132540 580500 132592
rect 599952 132540 600004 132592
rect 579804 132472 579856 132524
rect 600044 132472 600096 132524
rect 671712 132268 671764 132320
rect 676220 132268 676272 132320
rect 671896 131656 671948 131708
rect 672172 131656 672224 131708
rect 676036 131656 676088 131708
rect 673184 131452 673236 131504
rect 676220 131452 676272 131504
rect 672264 130840 672316 130892
rect 676036 130840 676088 130892
rect 673276 130636 673328 130688
rect 676220 130636 676272 130688
rect 671804 130024 671856 130076
rect 672080 130024 672132 130076
rect 676036 130024 676088 130076
rect 581184 129888 581236 129940
rect 599952 129888 600004 129940
rect 580632 129820 580684 129872
rect 599768 129820 599820 129872
rect 580080 129752 580132 129804
rect 598940 129752 598992 129804
rect 673368 129684 673420 129736
rect 676036 129684 676088 129736
rect 672356 129412 672408 129464
rect 673092 129412 673144 129464
rect 676220 129412 676272 129464
rect 674656 127712 674708 127764
rect 676036 127712 676088 127764
rect 673552 127304 673604 127356
rect 675944 127304 675996 127356
rect 582196 127032 582248 127084
rect 599860 127032 599912 127084
rect 673828 127032 673880 127084
rect 675944 127032 675996 127084
rect 580264 126964 580316 127016
rect 599952 126964 600004 127016
rect 674748 126964 674800 127016
rect 676036 126964 676088 127016
rect 674564 126080 674616 126132
rect 676036 126080 676088 126132
rect 673644 124584 673696 124636
rect 676128 124584 676180 124636
rect 674932 124448 674984 124500
rect 676036 124448 676088 124500
rect 580724 124312 580776 124364
rect 599952 124312 600004 124364
rect 673736 124312 673788 124364
rect 676128 124312 676180 124364
rect 580356 124244 580408 124296
rect 599860 124244 599912 124296
rect 674840 124244 674892 124296
rect 675944 124244 675996 124296
rect 580172 124176 580224 124228
rect 600044 124176 600096 124228
rect 675208 124176 675260 124228
rect 676036 124176 676088 124228
rect 674288 123632 674340 123684
rect 676036 123632 676088 123684
rect 582012 121592 582064 121644
rect 599584 121592 599636 121644
rect 672448 121592 672500 121644
rect 676220 121592 676272 121644
rect 580816 121524 580868 121576
rect 599952 121524 600004 121576
rect 580540 121456 580592 121508
rect 599860 121456 599912 121508
rect 675024 121456 675076 121508
rect 676036 121456 676088 121508
rect 586428 118804 586480 118856
rect 599860 118804 599912 118856
rect 583668 118736 583720 118788
rect 599952 118736 600004 118788
rect 582288 118668 582340 118720
rect 600044 118668 600096 118720
rect 582104 116016 582156 116068
rect 599860 116016 599912 116068
rect 581828 115948 581880 116000
rect 599952 115948 600004 116000
rect 666744 115880 666796 115932
rect 675392 115880 675444 115932
rect 674656 114316 674708 114368
rect 675208 114316 675260 114368
rect 674748 113704 674800 113756
rect 675208 113704 675260 113756
rect 581920 113296 581972 113348
rect 600044 113296 600096 113348
rect 581644 113228 581696 113280
rect 599952 113228 600004 113280
rect 581736 113160 581788 113212
rect 599860 113160 599912 113212
rect 674932 111868 674984 111920
rect 675208 111868 675260 111920
rect 674840 111120 674892 111172
rect 675392 111120 675444 111172
rect 581276 110508 581328 110560
rect 599952 110508 600004 110560
rect 581460 110440 581512 110492
rect 598940 110440 598992 110492
rect 673736 110032 673788 110084
rect 675116 110032 675168 110084
rect 673828 108196 673880 108248
rect 675392 108196 675444 108248
rect 581552 107720 581604 107772
rect 599860 107720 599912 107772
rect 581000 107652 581052 107704
rect 599952 107652 600004 107704
rect 674288 107516 674340 107568
rect 675392 107516 675444 107568
rect 673644 105680 673696 105732
rect 675116 105680 675168 105732
rect 581368 104932 581420 104984
rect 599860 104932 599912 104984
rect 581092 104864 581144 104916
rect 599952 104864 600004 104916
rect 673552 104524 673604 104576
rect 675116 104524 675168 104576
rect 657728 99764 657780 99816
rect 660902 99764 660954 99816
rect 580908 99356 580960 99408
rect 599952 99356 600004 99408
rect 633808 96568 633860 96620
rect 636384 96568 636436 96620
rect 637028 96568 637080 96620
rect 642180 96568 642232 96620
rect 655980 96568 656032 96620
rect 659568 96568 659620 96620
rect 661868 96568 661920 96620
rect 663064 96568 663116 96620
rect 634452 96500 634504 96552
rect 637580 96500 637632 96552
rect 654692 96500 654744 96552
rect 658280 96500 658332 96552
rect 659108 96500 659160 96552
rect 662512 96500 662564 96552
rect 635740 96432 635792 96484
rect 639880 96432 639932 96484
rect 652024 96432 652076 96484
rect 661960 96432 662012 96484
rect 636292 96364 636344 96416
rect 640984 96364 641036 96416
rect 633072 96296 633124 96348
rect 635280 96296 635332 96348
rect 640340 96228 640392 96280
rect 641720 96228 641772 96280
rect 638960 96160 639012 96212
rect 646228 96160 646280 96212
rect 622032 96092 622084 96144
rect 642824 96092 642876 96144
rect 631140 96024 631192 96076
rect 632106 96024 632158 96076
rect 632428 96024 632480 96076
rect 634406 96024 634458 96076
rect 635096 96024 635148 96076
rect 639006 96024 639058 96076
rect 640064 95956 640116 96008
rect 646044 95956 646096 96008
rect 631784 95888 631836 95940
rect 632980 95888 633032 95940
rect 639604 95888 639656 95940
rect 645952 95888 646004 95940
rect 623688 95820 623740 95872
rect 642916 95820 642968 95872
rect 647516 95820 647568 95872
rect 651564 95820 651616 95872
rect 621388 95752 621440 95804
rect 643008 95752 643060 95804
rect 626540 95684 626592 95736
rect 640340 95684 640392 95736
rect 640892 95684 640944 95736
rect 645860 95684 645912 95736
rect 596180 95616 596232 95668
rect 607680 95616 607732 95668
rect 638316 95616 638368 95668
rect 642640 95616 642692 95668
rect 652668 95616 652720 95668
rect 663800 95616 663852 95668
rect 607496 95548 607548 95600
rect 608968 95548 609020 95600
rect 610348 95548 610400 95600
rect 611544 95548 611596 95600
rect 616144 95548 616196 95600
rect 623228 95548 623280 95600
rect 623780 95548 623832 95600
rect 624608 95548 624660 95600
rect 637488 95548 637540 95600
rect 641628 95548 641680 95600
rect 643100 95548 643152 95600
rect 656992 95548 657044 95600
rect 659200 95548 659252 95600
rect 619364 95480 619416 95532
rect 621204 95480 621256 95532
rect 642732 95480 642784 95532
rect 660580 95480 660632 95532
rect 661408 95480 661460 95532
rect 620008 95412 620060 95464
rect 623504 95412 623556 95464
rect 642824 95412 642876 95464
rect 588084 95344 588136 95396
rect 610900 95344 610952 95396
rect 581184 95276 581236 95328
rect 612188 95276 612240 95328
rect 620744 95276 620796 95328
rect 642824 95276 642876 95328
rect 575664 95208 575716 95260
rect 606392 95208 606444 95260
rect 622676 95208 622728 95260
rect 623688 95208 623740 95260
rect 617432 95072 617484 95124
rect 621940 95072 621992 95124
rect 614856 94936 614908 94988
rect 615408 94936 615460 94988
rect 618720 94936 618772 94988
rect 623320 94936 623372 94988
rect 616788 94868 616840 94920
rect 622492 94868 622544 94920
rect 646780 95276 646832 95328
rect 663340 95276 663392 95328
rect 657084 95208 657136 95260
rect 657912 95208 657964 95260
rect 646136 95140 646188 95192
rect 663432 95140 663484 95192
rect 643468 95072 643520 95124
rect 644848 95072 644900 95124
rect 648620 94936 648672 94988
rect 650736 94936 650788 94988
rect 646044 94868 646096 94920
rect 646228 94868 646280 94920
rect 648712 94800 648764 94852
rect 649448 94800 649500 94852
rect 642916 94732 642968 94784
rect 653312 94732 653364 94784
rect 663708 94732 663760 94784
rect 647516 94664 647568 94716
rect 648160 94664 648212 94716
rect 651840 94664 651892 94716
rect 653404 94664 653456 94716
rect 656624 94664 656676 94716
rect 663892 94664 663944 94716
rect 657268 94596 657320 94648
rect 663524 94596 663576 94648
rect 618076 94528 618128 94580
rect 623136 94528 623188 94580
rect 648804 94528 648856 94580
rect 650092 94528 650144 94580
rect 656900 94528 656952 94580
rect 658556 94528 658608 94580
rect 648068 94460 648120 94512
rect 659844 94460 659896 94512
rect 660396 94460 660448 94512
rect 643560 94188 643612 94240
rect 644756 94120 644808 94172
rect 652760 94120 652812 94172
rect 644204 94052 644256 94104
rect 654048 94052 654100 94104
rect 607220 93848 607272 93900
rect 613568 93848 613620 93900
rect 649356 93848 649408 93900
rect 656900 93848 656952 93900
rect 585140 89632 585192 89684
rect 607220 89632 607272 89684
rect 657084 88816 657136 88868
rect 658004 88816 658056 88868
rect 659476 88816 659528 88868
rect 663616 88816 663668 88868
rect 582196 88340 582248 88392
rect 588084 88340 588136 88392
rect 591948 85960 592000 86012
rect 596180 85960 596232 86012
rect 648804 85484 648856 85536
rect 657728 85484 657780 85536
rect 651840 85416 651892 85468
rect 658832 85416 658884 85468
rect 648712 85348 648764 85400
rect 660672 85348 660724 85400
rect 648620 85280 648672 85332
rect 657176 85280 657228 85332
rect 643468 85212 643520 85264
rect 660120 85212 660172 85264
rect 647516 85144 647568 85196
rect 661408 85144 661460 85196
rect 583760 84396 583812 84448
rect 600504 84396 600556 84448
rect 583852 84328 583904 84380
rect 600688 84328 600740 84380
rect 580816 84260 580868 84312
rect 600320 84260 600372 84312
rect 580724 84192 580776 84244
rect 600228 84192 600280 84244
rect 580632 84124 580684 84176
rect 600412 84124 600464 84176
rect 602988 82832 603040 82884
rect 610164 82832 610216 82884
rect 579988 82764 580040 82816
rect 586428 82764 586480 82816
rect 579620 82288 579672 82340
rect 583668 82288 583720 82340
rect 604368 81268 604420 81320
rect 631324 81268 631376 81320
rect 628564 81200 628616 81252
rect 637028 81200 637080 81252
rect 575756 80112 575808 80164
rect 585140 80112 585192 80164
rect 629208 80044 629260 80096
rect 639880 80044 639932 80096
rect 615316 77188 615368 77240
rect 640340 77188 640392 77240
rect 623688 75964 623740 76016
rect 641076 75964 641128 76016
rect 623596 75828 623648 75880
rect 640984 75828 641036 75880
rect 612740 75760 612792 75812
rect 623090 75760 623142 75812
rect 631508 75760 631560 75812
rect 578148 74740 578200 74792
rect 625620 74944 625672 74996
rect 638960 74944 639012 74996
rect 598940 66444 598992 66496
rect 612740 66444 612792 66496
rect 579620 60392 579672 60444
rect 583760 60392 583812 60444
rect 597468 58352 597520 58404
rect 602988 58352 603040 58404
rect 579620 58284 579672 58336
rect 583852 58284 583904 58336
rect 594800 57944 594852 57996
rect 598940 57944 598992 57996
rect 52184 53864 52236 53916
rect 145380 53580 145432 53632
rect 339408 53560 339460 53612
rect 582196 53864 582248 53916
rect 594800 53796 594852 53848
rect 543648 53560 543700 53612
rect 600044 52436 600096 52488
rect 613016 52436 613068 52488
rect 52276 52368 52328 52420
rect 149980 52368 150032 52420
rect 568580 51008 568632 51060
rect 581184 51008 581236 51060
rect 150348 49648 150400 49700
rect 184940 49648 184992 49700
rect 615408 49512 615460 49564
rect 650000 49580 650052 49632
rect 478144 48424 478196 48476
rect 526168 48424 526220 48476
rect 412640 48356 412692 48408
rect 506388 48356 506440 48408
rect 281448 48288 281500 48340
rect 507860 48288 507912 48340
rect 661040 47336 661092 47388
rect 650000 46928 650052 46980
rect 460664 45772 460716 45824
rect 610348 45772 610400 45824
rect 367100 45704 367152 45756
rect 607404 45704 607456 45756
rect 312820 45636 312872 45688
rect 607588 45636 607640 45688
rect 85120 45568 85172 45620
rect 475568 45568 475620 45620
rect 187332 45500 187384 45552
rect 578148 45500 578200 45552
rect 312820 44140 312872 44192
rect 367100 44140 367152 44192
rect 310428 44072 310480 44124
rect 365168 44072 365220 44124
rect 390192 43120 390244 43172
rect 575664 43120 575716 43172
rect 223580 43052 223632 43104
rect 661460 43052 661512 43104
rect 475476 42576 475528 42628
rect 513288 41964 513340 42016
rect 518532 41964 518584 42016
rect 405832 41896 405884 41948
rect 420644 41896 420696 41948
rect 514024 41896 514076 41948
rect 514852 41896 514904 41948
rect 529664 41896 529716 41948
rect 530492 41896 530544 41948
rect 420644 41692 420696 41744
rect 607496 41420 607548 41472
rect 506388 41352 506440 41404
rect 513288 41352 513340 41404
rect 530308 41352 530360 41404
rect 610256 41352 610308 41404
rect 507860 41284 507912 41336
rect 513196 41284 513248 41336
rect 530400 41284 530452 41336
rect 575756 41284 575808 41336
rect 475568 38564 475620 38616
rect 514024 38564 514076 38616
rect 530492 38564 530544 38616
rect 543004 38564 543056 38616
<< metal2 >>
rect 703694 897668 703722 897804
rect 704154 897668 704182 897804
rect 704614 897668 704642 897804
rect 705074 897668 705102 897804
rect 705534 897668 705562 897804
rect 705994 897668 706022 897804
rect 706454 897668 706482 897804
rect 706914 897668 706942 897804
rect 707374 897668 707402 897804
rect 707834 897668 707862 897804
rect 708294 897668 708322 897804
rect 708754 897668 708782 897804
rect 709214 897668 709242 897804
rect 676034 897152 676090 897161
rect 676034 897087 676090 897096
rect 676048 897054 676076 897087
rect 655428 897048 655480 897054
rect 655428 896990 655480 896996
rect 676036 897048 676088 897054
rect 676036 896990 676088 896996
rect 655440 867649 655468 896990
rect 676034 896744 676090 896753
rect 676034 896679 676090 896688
rect 675942 894704 675998 894713
rect 673368 894668 673420 894674
rect 675942 894639 675944 894648
rect 673368 894610 673420 894616
rect 675996 894639 675998 894648
rect 675944 894610 675996 894616
rect 655612 894396 655664 894402
rect 655612 894338 655664 894344
rect 655520 894328 655572 894334
rect 655520 894270 655572 894276
rect 655426 867640 655482 867649
rect 655426 867575 655482 867584
rect 655532 866561 655560 894270
rect 655624 868873 655652 894338
rect 673276 893036 673328 893042
rect 673276 892978 673328 892984
rect 671988 885012 672040 885018
rect 671988 884954 672040 884960
rect 655704 883312 655756 883318
rect 655704 883254 655756 883260
rect 655610 868864 655666 868873
rect 655610 868799 655666 868808
rect 655518 866552 655574 866561
rect 655518 866487 655574 866496
rect 655716 865337 655744 883254
rect 655796 872228 655848 872234
rect 655796 872170 655848 872176
rect 655702 865328 655758 865337
rect 655702 865263 655758 865272
rect 655808 863841 655836 872170
rect 656808 863864 656860 863870
rect 655794 863832 655850 863841
rect 656808 863806 656860 863812
rect 655794 863767 655850 863776
rect 656820 862617 656848 863806
rect 656806 862608 656862 862617
rect 656806 862543 656862 862552
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 41786 817728 41842 817737
rect 41786 817663 41788 817672
rect 41840 817663 41842 817672
rect 50988 817692 51040 817698
rect 41788 817634 41840 817640
rect 50988 817634 51040 817640
rect 41786 817320 41842 817329
rect 41786 817255 41788 817264
rect 41840 817255 41842 817264
rect 48228 817284 48280 817290
rect 41788 817226 41840 817232
rect 48228 817226 48280 817232
rect 41786 816912 41842 816921
rect 41786 816847 41788 816856
rect 41840 816847 41842 816856
rect 45560 816876 45612 816882
rect 41788 816818 41840 816824
rect 45560 816818 45612 816824
rect 41786 816096 41842 816105
rect 41786 816031 41842 816040
rect 41800 815726 41828 816031
rect 41788 815720 41840 815726
rect 41788 815662 41840 815668
rect 43812 815720 43864 815726
rect 43812 815662 43864 815668
rect 41786 815280 41842 815289
rect 41786 815215 41842 815224
rect 41800 814570 41828 815215
rect 41788 814564 41840 814570
rect 41788 814506 41840 814512
rect 43628 814564 43680 814570
rect 43628 814506 43680 814512
rect 41786 814464 41842 814473
rect 41786 814399 41788 814408
rect 41840 814399 41842 814408
rect 43536 814428 43588 814434
rect 41788 814370 41840 814376
rect 43536 814370 43588 814376
rect 41786 813648 41842 813657
rect 41786 813583 41842 813592
rect 41800 813346 41828 813583
rect 41788 813340 41840 813346
rect 41788 813282 41840 813288
rect 43352 813340 43404 813346
rect 43352 813282 43404 813288
rect 41786 813240 41842 813249
rect 41786 813175 41842 813184
rect 41800 812938 41828 813175
rect 41788 812932 41840 812938
rect 41788 812874 41840 812880
rect 42800 812932 42852 812938
rect 42800 812874 42852 812880
rect 41786 812832 41842 812841
rect 41786 812767 41788 812776
rect 41840 812767 41842 812776
rect 42708 812796 42760 812802
rect 41788 812738 41840 812744
rect 42708 812738 42760 812744
rect 41786 812424 41842 812433
rect 41786 812359 41842 812368
rect 41800 811510 41828 812359
rect 41970 811608 42026 811617
rect 41970 811543 42026 811552
rect 41788 811504 41840 811510
rect 41788 811446 41840 811452
rect 41786 810792 41842 810801
rect 41786 810727 41842 810736
rect 41800 810150 41828 810727
rect 41878 810384 41934 810393
rect 41878 810319 41934 810328
rect 41788 810144 41840 810150
rect 41788 810086 41840 810092
rect 41786 809568 41842 809577
rect 41786 809503 41842 809512
rect 41800 808722 41828 809503
rect 41892 808858 41920 810319
rect 41880 808852 41932 808858
rect 41880 808794 41932 808800
rect 41878 808752 41934 808761
rect 41788 808716 41840 808722
rect 41878 808687 41934 808696
rect 41788 808658 41840 808664
rect 41786 808344 41842 808353
rect 41786 808279 41842 808288
rect 41800 808042 41828 808279
rect 41788 808036 41840 808042
rect 41788 807978 41840 807984
rect 41786 807936 41842 807945
rect 41786 807871 41842 807880
rect 41800 806070 41828 807871
rect 41788 806064 41840 806070
rect 41788 806006 41840 806012
rect 41892 803146 41920 808687
rect 41880 803140 41932 803146
rect 41880 803082 41932 803088
rect 41984 803078 42012 811543
rect 42246 811200 42302 811209
rect 42246 811135 42302 811144
rect 42062 807528 42118 807537
rect 42062 807463 42118 807472
rect 42076 806313 42104 807463
rect 42062 806304 42118 806313
rect 42062 806239 42118 806248
rect 42076 806002 42104 806239
rect 42064 805996 42116 806002
rect 42064 805938 42116 805944
rect 41972 803072 42024 803078
rect 41972 803014 42024 803020
rect 42260 799459 42288 811135
rect 42614 809976 42670 809985
rect 42614 809911 42670 809920
rect 42340 800488 42392 800494
rect 42340 800430 42392 800436
rect 42182 799431 42288 799459
rect 42352 799082 42380 800430
rect 42260 799054 42380 799082
rect 42156 798176 42208 798182
rect 42156 798118 42208 798124
rect 42168 797605 42196 798118
rect 42260 796974 42288 799054
rect 42340 798992 42392 798998
rect 42340 798934 42392 798940
rect 42182 796946 42288 796974
rect 42352 796906 42380 798934
rect 42260 796878 42380 796906
rect 42260 795938 42288 796878
rect 42340 796748 42392 796754
rect 42340 796690 42392 796696
rect 42248 795932 42300 795938
rect 42248 795874 42300 795880
rect 42352 795779 42380 796690
rect 42182 795751 42380 795779
rect 42182 795110 42380 795138
rect 42248 795048 42300 795054
rect 42248 794990 42300 794996
rect 42260 794594 42288 794990
rect 42182 794566 42288 794594
rect 42248 794504 42300 794510
rect 41878 794472 41934 794481
rect 42248 794446 42300 794452
rect 41878 794407 41934 794416
rect 41892 793900 41920 794407
rect 42156 793824 42208 793830
rect 42156 793766 42208 793772
rect 42168 793288 42196 793766
rect 42260 792758 42288 794446
rect 42182 792730 42288 792758
rect 42352 792266 42380 795110
rect 42340 792260 42392 792266
rect 42340 792202 42392 792208
rect 42628 792010 42656 809911
rect 42720 798182 42748 812738
rect 42812 798998 42840 812874
rect 43260 808716 43312 808722
rect 43260 808658 43312 808664
rect 43076 808036 43128 808042
rect 43076 807978 43128 807984
rect 42984 806064 43036 806070
rect 42984 806006 43036 806012
rect 42892 803140 42944 803146
rect 42892 803082 42944 803088
rect 42800 798992 42852 798998
rect 42800 798934 42852 798940
rect 42708 798176 42760 798182
rect 42708 798118 42760 798124
rect 42708 798040 42760 798046
rect 42708 797982 42760 797988
rect 42720 794510 42748 797982
rect 42708 794504 42760 794510
rect 42708 794446 42760 794452
rect 42708 792260 42760 792266
rect 42708 792202 42760 792208
rect 42444 791982 42656 792010
rect 42156 790696 42208 790702
rect 42156 790638 42208 790644
rect 42168 790228 42196 790638
rect 42444 789630 42472 791982
rect 42182 789602 42472 789630
rect 42248 789540 42300 789546
rect 42248 789482 42300 789488
rect 42156 789268 42208 789274
rect 42156 789210 42208 789216
rect 42168 788936 42196 789210
rect 42260 788406 42288 789482
rect 42432 789404 42484 789410
rect 42432 789346 42484 789352
rect 42340 789200 42392 789206
rect 42340 789142 42392 789148
rect 42182 788378 42288 788406
rect 42352 786570 42380 789142
rect 42182 786542 42380 786570
rect 42340 786480 42392 786486
rect 42340 786422 42392 786428
rect 42064 786276 42116 786282
rect 42064 786218 42116 786224
rect 42076 785944 42104 786218
rect 42352 785278 42380 786422
rect 42182 785250 42380 785278
rect 42444 784734 42472 789346
rect 42720 789342 42748 792202
rect 42904 790702 42932 803082
rect 42996 795054 43024 806006
rect 42984 795048 43036 795054
rect 42984 794990 43036 794996
rect 43088 793830 43116 807978
rect 43168 803072 43220 803078
rect 43168 803014 43220 803020
rect 43180 798046 43208 803014
rect 43168 798040 43220 798046
rect 43168 797982 43220 797988
rect 43168 797904 43220 797910
rect 43168 797846 43220 797852
rect 43076 793824 43128 793830
rect 43076 793766 43128 793772
rect 42892 790696 42944 790702
rect 42892 790638 42944 790644
rect 42708 789336 42760 789342
rect 42708 789278 42760 789284
rect 42182 784706 42472 784734
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 41786 774480 41842 774489
rect 41786 774415 41788 774424
rect 41840 774415 41842 774424
rect 41788 774386 41840 774392
rect 41512 774308 41564 774314
rect 41512 774250 41564 774256
rect 41418 773936 41474 773945
rect 41418 773871 41420 773880
rect 41472 773871 41474 773880
rect 41420 773842 41472 773848
rect 41524 773537 41552 774250
rect 41786 773664 41842 773673
rect 41786 773599 41788 773608
rect 41840 773599 41842 773608
rect 41788 773570 41840 773576
rect 41510 773528 41566 773537
rect 41510 773463 41566 773472
rect 41880 772880 41932 772886
rect 41878 772848 41880 772857
rect 41932 772848 41934 772857
rect 41788 772812 41840 772818
rect 41878 772783 41934 772792
rect 41788 772754 41840 772760
rect 41512 772744 41564 772750
rect 41510 772712 41512 772721
rect 41564 772712 41566 772721
rect 41510 772647 41566 772656
rect 41510 771896 41566 771905
rect 41510 771831 41566 771840
rect 41418 771080 41474 771089
rect 41418 771015 41420 771024
rect 41472 771015 41474 771024
rect 41420 770986 41472 770992
rect 41524 770370 41552 771831
rect 41800 771633 41828 772754
rect 41786 771624 41842 771633
rect 41786 771559 41842 771568
rect 43180 771526 43208 797846
rect 43272 796754 43300 808658
rect 43364 797910 43392 813282
rect 43444 811504 43496 811510
rect 43444 811446 43496 811452
rect 43352 797904 43404 797910
rect 43352 797846 43404 797852
rect 43352 797768 43404 797774
rect 43352 797710 43404 797716
rect 43260 796748 43312 796754
rect 43260 796690 43312 796696
rect 43260 795932 43312 795938
rect 43260 795874 43312 795880
rect 43272 789206 43300 795874
rect 43260 789200 43312 789206
rect 43260 789142 43312 789148
rect 43364 772818 43392 797710
rect 43456 786486 43484 811446
rect 43548 797978 43576 814370
rect 43536 797972 43588 797978
rect 43536 797914 43588 797920
rect 43640 797858 43668 814506
rect 43718 811880 43774 811889
rect 43718 811815 43774 811824
rect 43548 797830 43668 797858
rect 43732 797842 43760 811815
rect 43720 797836 43772 797842
rect 43444 786480 43496 786486
rect 43444 786422 43496 786428
rect 43352 772812 43404 772818
rect 43352 772754 43404 772760
rect 43548 772750 43576 797830
rect 43720 797778 43772 797784
rect 43720 797700 43772 797706
rect 43720 797642 43772 797648
rect 43628 794096 43680 794102
rect 43628 794038 43680 794044
rect 43640 774314 43668 794038
rect 43732 789546 43760 797642
rect 43824 794102 43852 815662
rect 43904 810144 43956 810150
rect 43904 810086 43956 810092
rect 43812 794096 43864 794102
rect 43812 794038 43864 794044
rect 43720 789540 43772 789546
rect 43720 789482 43772 789488
rect 43916 786282 43944 810086
rect 44088 808852 44140 808858
rect 44088 808794 44140 808800
rect 44100 789274 44128 808794
rect 45468 805996 45520 806002
rect 45468 805938 45520 805944
rect 44088 789268 44140 789274
rect 44088 789210 44140 789216
rect 43904 786276 43956 786282
rect 43904 786218 43956 786224
rect 43628 774308 43680 774314
rect 43628 774250 43680 774256
rect 44088 772880 44140 772886
rect 44088 772822 44140 772828
rect 43536 772744 43588 772750
rect 43536 772686 43588 772692
rect 41788 771520 41840 771526
rect 41788 771462 41840 771468
rect 43168 771520 43220 771526
rect 43168 771462 43220 771468
rect 41800 770817 41828 771462
rect 43168 771044 43220 771050
rect 43168 770986 43220 770992
rect 41786 770808 41842 770817
rect 41786 770743 41842 770752
rect 42154 770400 42210 770409
rect 41512 770364 41564 770370
rect 42154 770335 42210 770344
rect 42432 770364 42484 770370
rect 41512 770306 41564 770312
rect 41510 769856 41566 769865
rect 41510 769791 41566 769800
rect 41524 769554 41552 769791
rect 41512 769548 41564 769554
rect 41512 769490 41564 769496
rect 41510 769448 41566 769457
rect 41510 769383 41512 769392
rect 41564 769383 41566 769392
rect 41512 769354 41564 769360
rect 41510 769040 41566 769049
rect 41510 768975 41512 768984
rect 41564 768975 41566 768984
rect 41512 768946 41564 768952
rect 41510 768632 41566 768641
rect 41510 768567 41566 768576
rect 41524 768330 41552 768567
rect 41512 768324 41564 768330
rect 41512 768266 41564 768272
rect 41510 768224 41566 768233
rect 41510 768159 41512 768168
rect 41564 768159 41566 768168
rect 41512 768130 41564 768136
rect 41786 767952 41842 767961
rect 41786 767887 41842 767896
rect 41512 767440 41564 767446
rect 41510 767408 41512 767417
rect 41564 767408 41566 767417
rect 41510 767343 41566 767352
rect 41694 767000 41750 767009
rect 41694 766935 41750 766944
rect 41418 766592 41474 766601
rect 41418 766527 41474 766536
rect 41432 759082 41460 766527
rect 41510 766184 41566 766193
rect 41510 766119 41512 766128
rect 41564 766119 41566 766128
rect 41512 766090 41564 766096
rect 41510 765776 41566 765785
rect 41510 765711 41512 765720
rect 41564 765711 41566 765720
rect 41512 765682 41564 765688
rect 41602 765368 41658 765377
rect 41602 765303 41658 765312
rect 41510 764960 41566 764969
rect 41510 764895 41512 764904
rect 41564 764895 41566 764904
rect 41512 764866 41564 764872
rect 41512 764584 41564 764590
rect 41510 764552 41512 764561
rect 41564 764552 41566 764561
rect 41510 764487 41566 764496
rect 41510 764144 41566 764153
rect 41510 764079 41566 764088
rect 41524 762929 41552 764079
rect 41510 762920 41566 762929
rect 41510 762855 41512 762864
rect 41564 762855 41566 762864
rect 41512 762826 41564 762832
rect 41616 759354 41644 765303
rect 41708 761682 41736 766935
rect 41800 761802 41828 767887
rect 41788 761796 41840 761802
rect 41788 761738 41840 761744
rect 41708 761654 41828 761682
rect 41604 759348 41656 759354
rect 41604 759290 41656 759296
rect 41420 759076 41472 759082
rect 41420 759018 41472 759024
rect 41800 757081 41828 761654
rect 42168 757081 42196 770335
rect 42432 770306 42484 770312
rect 42444 767294 42472 770306
rect 43076 769412 43128 769418
rect 43076 769354 43128 769360
rect 42605 767378 42748 767394
rect 42605 767372 42760 767378
rect 42605 767366 42708 767372
rect 42708 767314 42760 767320
rect 42352 767266 42472 767294
rect 42248 761796 42300 761802
rect 42248 761738 42300 761744
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 42154 757072 42210 757081
rect 42154 757007 42210 757016
rect 42260 756786 42288 761738
rect 42352 760986 42380 767266
rect 42432 766148 42484 766154
rect 42432 766090 42484 766096
rect 42340 760980 42392 760986
rect 42340 760922 42392 760928
rect 42340 760844 42392 760850
rect 42340 760786 42392 760792
rect 42168 756758 42288 756786
rect 42168 756228 42196 756758
rect 42248 756288 42300 756294
rect 42248 756230 42300 756236
rect 42156 754928 42208 754934
rect 42156 754870 42208 754876
rect 42168 754392 42196 754870
rect 42168 753370 42196 753780
rect 42156 753364 42208 753370
rect 42156 753306 42208 753312
rect 42156 753092 42208 753098
rect 42156 753034 42208 753040
rect 42168 752556 42196 753034
rect 42168 751890 42196 751944
rect 42260 751890 42288 756230
rect 42352 754934 42380 760786
rect 42444 760714 42472 766090
rect 42708 764584 42760 764590
rect 42708 764526 42760 764532
rect 42432 760708 42484 760714
rect 42432 760650 42484 760656
rect 42340 754928 42392 754934
rect 42340 754870 42392 754876
rect 42720 754322 42748 764526
rect 43088 760850 43116 769354
rect 43076 760844 43128 760850
rect 43076 760786 43128 760792
rect 43076 760708 43128 760714
rect 43076 760650 43128 760656
rect 42340 754316 42392 754322
rect 42340 754258 42392 754264
rect 42708 754316 42760 754322
rect 42708 754258 42760 754264
rect 42168 751862 42288 751890
rect 42352 751383 42380 754258
rect 42708 753364 42760 753370
rect 42708 753306 42760 753312
rect 42182 751355 42380 751383
rect 42340 751256 42392 751262
rect 42340 751198 42392 751204
rect 42352 750734 42380 751198
rect 42182 750706 42380 750734
rect 42064 750644 42116 750650
rect 42064 750586 42116 750592
rect 42076 750108 42104 750586
rect 42340 750576 42392 750582
rect 42340 750518 42392 750524
rect 42248 750508 42300 750514
rect 42248 750450 42300 750456
rect 42260 749543 42288 750450
rect 42182 749515 42288 749543
rect 42352 747062 42380 750518
rect 42720 750446 42748 753306
rect 43088 753098 43116 760650
rect 43180 757602 43208 770986
rect 43260 769548 43312 769554
rect 43260 769490 43312 769496
rect 43272 757738 43300 769490
rect 43720 769004 43772 769010
rect 43720 768946 43772 768952
rect 43444 768324 43496 768330
rect 43444 768266 43496 768272
rect 43352 768188 43404 768194
rect 43352 768130 43404 768136
rect 43364 765882 43392 768130
rect 43352 765876 43404 765882
rect 43352 765818 43404 765824
rect 43352 765740 43404 765746
rect 43352 765682 43404 765688
rect 43364 757858 43392 765682
rect 43352 757852 43404 757858
rect 43352 757794 43404 757800
rect 43272 757710 43392 757738
rect 43180 757574 43300 757602
rect 43168 757512 43220 757518
rect 43168 757454 43220 757460
rect 43076 753092 43128 753098
rect 43076 753034 43128 753040
rect 43074 752992 43130 753001
rect 43074 752927 43130 752936
rect 42708 750440 42760 750446
rect 42708 750382 42760 750388
rect 43088 750378 43116 752927
rect 43076 750372 43128 750378
rect 43076 750314 43128 750320
rect 42430 748776 42486 748785
rect 42430 748711 42486 748720
rect 42182 747034 42380 747062
rect 42340 746972 42392 746978
rect 42340 746914 42392 746920
rect 42352 746415 42380 746914
rect 42182 746387 42380 746415
rect 42444 745770 42472 748711
rect 42182 745742 42472 745770
rect 42248 745612 42300 745618
rect 42248 745554 42300 745560
rect 42260 745226 42288 745554
rect 42182 745198 42288 745226
rect 42340 745272 42392 745278
rect 42340 745214 42392 745220
rect 42248 745136 42300 745142
rect 42248 745078 42300 745084
rect 42260 743390 42288 745078
rect 42182 743362 42288 743390
rect 42248 743300 42300 743306
rect 42248 743242 42300 743248
rect 42156 743096 42208 743102
rect 42156 743038 42208 743044
rect 42168 742696 42196 743038
rect 42260 742098 42288 743242
rect 42182 742070 42288 742098
rect 42352 741554 42380 745214
rect 43180 745142 43208 757454
rect 43168 745136 43220 745142
rect 43168 745078 43220 745084
rect 42182 741526 42380 741554
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 41510 731096 41566 731105
rect 41510 731031 41512 731040
rect 41564 731031 41566 731040
rect 41512 731002 41564 731008
rect 41788 730788 41840 730794
rect 41788 730730 41840 730736
rect 41510 730688 41566 730697
rect 41510 730623 41512 730632
rect 41564 730623 41566 730632
rect 41512 730594 41564 730600
rect 41510 730280 41566 730289
rect 41510 730215 41512 730224
rect 41564 730215 41566 730224
rect 41512 730186 41564 730192
rect 41510 729464 41566 729473
rect 41510 729399 41566 729408
rect 41524 729162 41552 729399
rect 41800 729337 41828 730730
rect 41880 730516 41932 730522
rect 41880 730458 41932 730464
rect 41892 730153 41920 730458
rect 41878 730144 41934 730153
rect 41878 730079 41934 730088
rect 41786 729328 41842 729337
rect 41786 729263 41842 729272
rect 41512 729156 41564 729162
rect 41512 729098 41564 729104
rect 42430 728920 42486 728929
rect 42430 728855 42486 728864
rect 41510 728648 41566 728657
rect 41510 728583 41512 728592
rect 41564 728583 41566 728592
rect 41512 728554 41564 728560
rect 41786 728104 41842 728113
rect 41786 728039 41842 728048
rect 41512 727932 41564 727938
rect 41512 727874 41564 727880
rect 41524 727841 41552 727874
rect 41510 727832 41566 727841
rect 41510 727767 41566 727776
rect 41510 726608 41566 726617
rect 41510 726543 41512 726552
rect 41564 726543 41566 726552
rect 41512 726514 41564 726520
rect 41800 726238 41828 728039
rect 41970 727288 42026 727297
rect 41970 727223 42026 727232
rect 41788 726232 41840 726238
rect 41510 726200 41566 726209
rect 41788 726174 41840 726180
rect 41510 726135 41512 726144
rect 41564 726135 41566 726144
rect 41512 726106 41564 726112
rect 41786 726064 41842 726073
rect 41786 725999 41788 726008
rect 41840 725999 41842 726008
rect 41788 725970 41840 725976
rect 41510 725384 41566 725393
rect 41510 725319 41566 725328
rect 41524 724266 41552 725319
rect 41786 725248 41842 725257
rect 41786 725183 41842 725192
rect 41512 724260 41564 724266
rect 41512 724202 41564 724208
rect 41510 724160 41566 724169
rect 41510 724095 41566 724104
rect 30286 723752 30342 723761
rect 30286 723687 30342 723696
rect 30300 716310 30328 723687
rect 41524 723314 41552 724095
rect 41800 723450 41828 725183
rect 41788 723444 41840 723450
rect 41788 723386 41840 723392
rect 41694 723344 41750 723353
rect 41512 723308 41564 723314
rect 41694 723279 41750 723288
rect 41512 723250 41564 723256
rect 41510 722120 41566 722129
rect 41510 722055 41512 722064
rect 41564 722055 41566 722064
rect 41512 722026 41564 722032
rect 41510 721712 41566 721721
rect 41510 721647 41566 721656
rect 41418 720896 41474 720905
rect 41418 720831 41474 720840
rect 41432 719658 41460 720831
rect 41524 720458 41552 721647
rect 41602 721304 41658 721313
rect 41602 721239 41658 721248
rect 41616 720730 41644 721239
rect 41604 720724 41656 720730
rect 41604 720666 41656 720672
rect 41512 720452 41564 720458
rect 41512 720394 41564 720400
rect 41510 719672 41566 719681
rect 41432 719630 41510 719658
rect 41510 719607 41512 719616
rect 41564 719607 41566 719616
rect 41512 719578 41564 719584
rect 30288 716304 30340 716310
rect 30288 716246 30340 716252
rect 41708 714950 41736 723279
rect 41786 723208 41842 723217
rect 41786 723143 41788 723152
rect 41840 723143 41842 723152
rect 41788 723114 41840 723120
rect 41878 722800 41934 722809
rect 41878 722735 41934 722744
rect 41696 714944 41748 714950
rect 41696 714886 41748 714892
rect 41892 713862 41920 722735
rect 41984 713930 42012 727223
rect 42246 724840 42302 724849
rect 42246 724775 42302 724784
rect 41972 713924 42024 713930
rect 41972 713866 42024 713872
rect 41880 713856 41932 713862
rect 41880 713798 41932 713804
rect 42260 713062 42288 724775
rect 42340 714876 42392 714882
rect 42340 714818 42392 714824
rect 42182 713034 42288 713062
rect 42248 712972 42300 712978
rect 42248 712914 42300 712920
rect 42156 711748 42208 711754
rect 42156 711690 42208 711696
rect 42168 711212 42196 711690
rect 42156 710932 42208 710938
rect 42156 710874 42208 710880
rect 42168 710561 42196 710874
rect 42260 709986 42288 712914
rect 42352 710938 42380 714818
rect 42340 710932 42392 710938
rect 42340 710874 42392 710880
rect 42340 710456 42392 710462
rect 42340 710398 42392 710404
rect 42248 709980 42300 709986
rect 42248 709922 42300 709928
rect 42352 709866 42380 710398
rect 42076 709838 42380 709866
rect 42076 709376 42104 709838
rect 42340 709776 42392 709782
rect 42340 709718 42392 709724
rect 42248 709436 42300 709442
rect 42248 709378 42300 709384
rect 42260 709050 42288 709378
rect 42168 709022 42288 709050
rect 42168 708696 42196 709022
rect 42246 708928 42302 708937
rect 42246 708863 42302 708872
rect 42156 708620 42208 708626
rect 42156 708562 42208 708568
rect 42168 708152 42196 708562
rect 42156 708076 42208 708082
rect 42156 708018 42208 708024
rect 42168 707540 42196 708018
rect 42156 707260 42208 707266
rect 42156 707202 42208 707208
rect 42168 706860 42196 707202
rect 42156 706784 42208 706790
rect 42156 706726 42208 706732
rect 42168 706316 42196 706726
rect 42064 704268 42116 704274
rect 42064 704210 42116 704216
rect 42076 703868 42104 704210
rect 42156 703588 42208 703594
rect 42156 703530 42208 703536
rect 42168 703188 42196 703530
rect 42064 703112 42116 703118
rect 42064 703054 42116 703060
rect 42076 702576 42104 703054
rect 42064 702432 42116 702438
rect 42064 702374 42116 702380
rect 42076 702032 42104 702374
rect 42156 700596 42208 700602
rect 42156 700538 42208 700544
rect 42168 700165 42196 700538
rect 42156 700052 42208 700058
rect 42156 699994 42208 700000
rect 42168 699516 42196 699994
rect 42168 698850 42196 698904
rect 42260 698850 42288 708863
rect 42352 708082 42380 709718
rect 42340 708076 42392 708082
rect 42340 708018 42392 708024
rect 42340 703860 42392 703866
rect 42340 703802 42392 703808
rect 42168 698822 42288 698850
rect 42352 698339 42380 703802
rect 42182 698311 42380 698339
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 41786 688120 41842 688129
rect 41786 688055 41788 688064
rect 41840 688055 41842 688064
rect 41788 688026 41840 688032
rect 41786 687712 41842 687721
rect 41786 687647 41788 687656
rect 41840 687647 41842 687656
rect 41788 687618 41840 687624
rect 41788 687336 41840 687342
rect 41786 687304 41788 687313
rect 41840 687304 41842 687313
rect 41786 687239 41842 687248
rect 41788 687200 41840 687206
rect 41788 687142 41840 687148
rect 41800 686905 41828 687142
rect 41786 686896 41842 686905
rect 41786 686831 41842 686840
rect 41786 686488 41842 686497
rect 41786 686423 41842 686432
rect 41800 686186 41828 686423
rect 41788 686180 41840 686186
rect 41788 686122 41840 686128
rect 42444 686089 42472 728855
rect 43272 728618 43300 757574
rect 43364 757518 43392 757710
rect 43456 757602 43484 768266
rect 43536 767440 43588 767446
rect 43536 767382 43588 767388
rect 43548 766358 43576 767382
rect 43536 766352 43588 766358
rect 43536 766294 43588 766300
rect 43628 765876 43680 765882
rect 43628 765818 43680 765824
rect 43640 761138 43668 765818
rect 43548 761110 43668 761138
rect 43548 757722 43576 761110
rect 43628 760980 43680 760986
rect 43628 760922 43680 760928
rect 43536 757716 43588 757722
rect 43536 757658 43588 757664
rect 43456 757574 43576 757602
rect 43352 757512 43404 757518
rect 43352 757454 43404 757460
rect 43444 757512 43496 757518
rect 43444 757454 43496 757460
rect 43352 757376 43404 757382
rect 43352 757318 43404 757324
rect 43364 743306 43392 757318
rect 43456 751262 43484 757454
rect 43444 751256 43496 751262
rect 43444 751198 43496 751204
rect 43548 751194 43576 757574
rect 43536 751188 43588 751194
rect 43536 751130 43588 751136
rect 43640 751074 43668 760922
rect 43732 757382 43760 768946
rect 43996 766352 44048 766358
rect 43996 766294 44048 766300
rect 43812 764924 43864 764930
rect 43812 764866 43864 764872
rect 43720 757376 43772 757382
rect 43720 757318 43772 757324
rect 43720 757240 43772 757246
rect 43720 757182 43772 757188
rect 43456 751046 43668 751074
rect 43352 743300 43404 743306
rect 43352 743242 43404 743248
rect 43456 730794 43484 751046
rect 43536 750984 43588 750990
rect 43536 750926 43588 750932
rect 43548 745618 43576 750926
rect 43732 750514 43760 757182
rect 43824 750650 43852 764866
rect 43904 759348 43956 759354
rect 43904 759290 43956 759296
rect 43812 750644 43864 750650
rect 43812 750586 43864 750592
rect 43916 750582 43944 759290
rect 43904 750576 43956 750582
rect 43904 750518 43956 750524
rect 43720 750508 43772 750514
rect 43720 750450 43772 750456
rect 43812 750508 43864 750514
rect 43812 750450 43864 750456
rect 43720 750372 43772 750378
rect 43720 750314 43772 750320
rect 43536 745612 43588 745618
rect 43536 745554 43588 745560
rect 43444 730788 43496 730794
rect 43444 730730 43496 730736
rect 43260 728612 43312 728618
rect 43260 728554 43312 728560
rect 43732 727938 43760 750314
rect 43824 746978 43852 750450
rect 43904 750440 43956 750446
rect 43904 750382 43956 750388
rect 43916 747930 43944 750382
rect 43904 747924 43956 747930
rect 43904 747866 43956 747872
rect 43812 746972 43864 746978
rect 43812 746914 43864 746920
rect 44008 743102 44036 766294
rect 43996 743096 44048 743102
rect 43996 743038 44048 743044
rect 44100 730522 44128 772822
rect 44180 759076 44232 759082
rect 44180 759018 44232 759024
rect 44192 750514 44220 759018
rect 44180 750508 44232 750514
rect 44180 750450 44232 750456
rect 44088 730516 44140 730522
rect 44088 730458 44140 730464
rect 43996 729156 44048 729162
rect 43996 729098 44048 729104
rect 43720 727932 43772 727938
rect 43720 727874 43772 727880
rect 43168 726572 43220 726578
rect 43168 726514 43220 726520
rect 43076 726232 43128 726238
rect 43076 726174 43128 726180
rect 42708 723172 42760 723178
rect 42708 723114 42760 723120
rect 42720 710462 42748 723114
rect 43088 714377 43116 726174
rect 43074 714368 43130 714377
rect 43074 714303 43130 714312
rect 43180 714241 43208 726514
rect 43352 726164 43404 726170
rect 43352 726106 43404 726112
rect 43260 720452 43312 720458
rect 43260 720394 43312 720400
rect 43166 714232 43222 714241
rect 43166 714167 43222 714176
rect 42708 710456 42760 710462
rect 42708 710398 42760 710404
rect 43272 710326 43300 720394
rect 43364 711754 43392 726106
rect 43720 726028 43772 726034
rect 43720 725970 43772 725976
rect 43536 723308 43588 723314
rect 43536 723250 43588 723256
rect 43444 722084 43496 722090
rect 43444 722026 43496 722032
rect 43352 711748 43404 711754
rect 43352 711690 43404 711696
rect 43456 711634 43484 722026
rect 43364 711606 43484 711634
rect 42708 710320 42760 710326
rect 42708 710262 42760 710268
rect 43260 710320 43312 710326
rect 43260 710262 43312 710268
rect 42720 707266 42748 710262
rect 43260 710184 43312 710190
rect 43260 710126 43312 710132
rect 42708 707260 42760 707266
rect 42708 707202 42760 707208
rect 43272 702438 43300 710126
rect 43364 704274 43392 711606
rect 43442 711512 43498 711521
rect 43442 711447 43498 711456
rect 43352 704268 43404 704274
rect 43352 704210 43404 704216
rect 43260 702432 43312 702438
rect 43260 702374 43312 702380
rect 42430 686080 42486 686089
rect 41788 686044 41840 686050
rect 43456 686050 43484 711447
rect 43548 700058 43576 723250
rect 43628 716304 43680 716310
rect 43628 716246 43680 716252
rect 43640 703118 43668 716246
rect 43732 709481 43760 725970
rect 43904 724260 43956 724266
rect 43904 724202 43956 724208
rect 43812 720724 43864 720730
rect 43812 720666 43864 720672
rect 43718 709472 43774 709481
rect 43718 709407 43774 709416
rect 43720 709368 43772 709374
rect 43720 709310 43772 709316
rect 43732 706790 43760 709310
rect 43824 708626 43852 720666
rect 43916 710190 43944 724202
rect 43904 710184 43956 710190
rect 43904 710126 43956 710132
rect 43904 710048 43956 710054
rect 43904 709990 43956 709996
rect 43812 708620 43864 708626
rect 43812 708562 43864 708568
rect 43810 708520 43866 708529
rect 43810 708455 43866 708464
rect 43720 706784 43772 706790
rect 43720 706726 43772 706732
rect 43628 703112 43680 703118
rect 43628 703054 43680 703060
rect 43824 700602 43852 708455
rect 43812 700596 43864 700602
rect 43812 700538 43864 700544
rect 43536 700052 43588 700058
rect 43536 699994 43588 700000
rect 42430 686015 42486 686024
rect 43444 686044 43496 686050
rect 41788 685986 41840 685992
rect 43444 685986 43496 685992
rect 41800 685273 41828 685986
rect 42062 685672 42118 685681
rect 42062 685607 42118 685616
rect 41786 685264 41842 685273
rect 41786 685199 41842 685208
rect 41788 684480 41840 684486
rect 41786 684448 41788 684457
rect 41840 684448 41842 684457
rect 41786 684383 41842 684392
rect 41786 684040 41842 684049
rect 41786 683975 41842 683984
rect 41800 683738 41828 683975
rect 41788 683732 41840 683738
rect 41788 683674 41840 683680
rect 41786 683632 41842 683641
rect 41786 683567 41842 683576
rect 41694 682680 41750 682689
rect 41694 682615 41750 682624
rect 41708 682514 41736 682615
rect 41696 682508 41748 682514
rect 41696 682450 41748 682456
rect 41694 682272 41750 682281
rect 41694 682207 41696 682216
rect 41748 682207 41750 682216
rect 41696 682178 41748 682184
rect 30286 682000 30342 682009
rect 30286 681935 30342 681944
rect 27434 680368 27490 680377
rect 27434 680303 27490 680312
rect 27448 672110 27476 680303
rect 27526 679144 27582 679153
rect 27526 679079 27582 679088
rect 27540 672178 27568 679079
rect 30300 672246 30328 681935
rect 41800 681766 41828 683567
rect 41788 681760 41840 681766
rect 41788 681702 41840 681708
rect 41786 681184 41842 681193
rect 41786 681119 41842 681128
rect 41800 680066 41828 681119
rect 41970 680776 42026 680785
rect 41970 680711 42026 680720
rect 41788 680060 41840 680066
rect 41788 680002 41840 680008
rect 41786 679960 41842 679969
rect 41786 679895 41788 679904
rect 41840 679895 41842 679904
rect 41788 679866 41840 679872
rect 41694 679416 41750 679425
rect 41694 679351 41696 679360
rect 41748 679351 41750 679360
rect 41696 679322 41748 679328
rect 41786 678736 41842 678745
rect 41786 678671 41842 678680
rect 41694 678192 41750 678201
rect 41694 678127 41750 678136
rect 41708 676666 41736 678127
rect 41696 676660 41748 676666
rect 41696 676602 41748 676608
rect 41694 676560 41750 676569
rect 41694 676495 41696 676504
rect 41748 676495 41750 676504
rect 41696 676466 41748 676472
rect 41800 676258 41828 678671
rect 41788 676252 41840 676258
rect 41788 676194 41840 676200
rect 30288 672240 30340 672246
rect 30288 672182 30340 672188
rect 27528 672172 27580 672178
rect 27528 672114 27580 672120
rect 27436 672104 27488 672110
rect 27436 672046 27488 672052
rect 41984 670721 42012 680711
rect 42076 670750 42104 685607
rect 42430 684856 42486 684865
rect 42430 684791 42486 684800
rect 42246 683224 42302 683233
rect 42246 683159 42302 683168
rect 42064 670744 42116 670750
rect 41970 670712 42026 670721
rect 42064 670686 42116 670692
rect 41970 670647 42026 670656
rect 42260 670002 42288 683159
rect 42338 681592 42394 681601
rect 42338 681527 42394 681536
rect 42248 669996 42300 670002
rect 42248 669938 42300 669944
rect 42352 669882 42380 681527
rect 42444 670993 42472 684791
rect 43916 684486 43944 709990
rect 44008 687206 44036 729098
rect 44088 723444 44140 723450
rect 44088 723386 44140 723392
rect 44100 712314 44128 723386
rect 44272 714944 44324 714950
rect 44272 714886 44324 714892
rect 44100 712286 44220 712314
rect 44088 712156 44140 712162
rect 44088 712098 44140 712104
rect 44100 709714 44128 712098
rect 44088 709708 44140 709714
rect 44088 709650 44140 709656
rect 44192 709594 44220 712286
rect 44100 709566 44220 709594
rect 44100 709442 44128 709566
rect 44088 709436 44140 709442
rect 44088 709378 44140 709384
rect 44284 709334 44312 714886
rect 44364 713924 44416 713930
rect 44364 713866 44416 713872
rect 44376 710054 44404 713866
rect 44364 710048 44416 710054
rect 44364 709990 44416 709996
rect 44100 709306 44312 709334
rect 44100 703594 44128 709306
rect 44088 703588 44140 703594
rect 44088 703530 44140 703536
rect 43996 687200 44048 687206
rect 43996 687142 44048 687148
rect 43996 686180 44048 686186
rect 43996 686122 44048 686128
rect 43904 684480 43956 684486
rect 43904 684422 43956 684428
rect 43536 683732 43588 683738
rect 43536 683674 43588 683680
rect 43444 681760 43496 681766
rect 43444 681702 43496 681708
rect 43352 676660 43404 676666
rect 43352 676602 43404 676608
rect 42708 676252 42760 676258
rect 42708 676194 42760 676200
rect 42430 670984 42486 670993
rect 42430 670919 42486 670928
rect 42432 670880 42484 670886
rect 42432 670822 42484 670828
rect 42444 670274 42472 670822
rect 42720 670410 42748 676194
rect 43076 672240 43128 672246
rect 43076 672182 43128 672188
rect 43088 670562 43116 672182
rect 43168 672172 43220 672178
rect 43168 672114 43220 672120
rect 43180 670682 43208 672114
rect 43260 672104 43312 672110
rect 43260 672046 43312 672052
rect 43272 670721 43300 672046
rect 43258 670712 43314 670721
rect 43168 670676 43220 670682
rect 43258 670647 43314 670656
rect 43168 670618 43220 670624
rect 43258 670576 43314 670585
rect 43088 670534 43208 670562
rect 42708 670404 42760 670410
rect 42708 670346 42760 670352
rect 43076 670404 43128 670410
rect 43076 670346 43128 670352
rect 42432 670268 42484 670274
rect 42432 670210 42484 670216
rect 42708 670268 42760 670274
rect 42708 670210 42760 670216
rect 42168 669746 42196 669868
rect 42260 669854 42380 669882
rect 42260 669746 42288 669854
rect 42168 669718 42288 669746
rect 42340 669792 42392 669798
rect 42340 669734 42392 669740
rect 42352 668046 42380 669734
rect 42168 667978 42196 668032
rect 42260 668018 42380 668046
rect 42260 667978 42288 668018
rect 42168 667950 42288 667978
rect 42720 667962 42748 670210
rect 42340 667956 42392 667962
rect 42340 667898 42392 667904
rect 42708 667956 42760 667962
rect 42708 667898 42760 667904
rect 42352 667366 42380 667898
rect 42708 667820 42760 667826
rect 42708 667762 42760 667768
rect 42182 667338 42380 667366
rect 42340 667276 42392 667282
rect 42340 667218 42392 667224
rect 42352 666179 42380 667218
rect 42182 666151 42380 666179
rect 42182 665502 42380 665530
rect 42248 665440 42300 665446
rect 42248 665382 42300 665388
rect 42156 665236 42208 665242
rect 42156 665178 42208 665184
rect 42168 664972 42196 665178
rect 42156 664692 42208 664698
rect 42156 664634 42208 664640
rect 42168 664325 42196 664634
rect 42260 663694 42288 665382
rect 42182 663666 42288 663694
rect 42248 663604 42300 663610
rect 42248 663546 42300 663552
rect 42260 663150 42288 663546
rect 42182 663122 42288 663150
rect 42248 663060 42300 663066
rect 42248 663002 42300 663008
rect 42156 661088 42208 661094
rect 42156 661030 42208 661036
rect 42168 660620 42196 661030
rect 42260 660022 42288 663002
rect 42182 659994 42288 660022
rect 42352 659666 42380 665502
rect 42720 664698 42748 667762
rect 43088 665446 43116 670346
rect 43076 665440 43128 665446
rect 43076 665382 43128 665388
rect 43074 665272 43130 665281
rect 43074 665207 43130 665216
rect 42708 664692 42760 664698
rect 42708 664634 42760 664640
rect 42432 659728 42484 659734
rect 42432 659670 42484 659676
rect 42340 659660 42392 659666
rect 42340 659602 42392 659608
rect 42340 659524 42392 659530
rect 42340 659466 42392 659472
rect 42352 659371 42380 659466
rect 42182 659343 42380 659371
rect 42340 659252 42392 659258
rect 42340 659194 42392 659200
rect 42156 659048 42208 659054
rect 42156 658990 42208 658996
rect 42168 658784 42196 658990
rect 42156 657416 42208 657422
rect 42156 657358 42208 657364
rect 42168 656948 42196 657358
rect 42352 656350 42380 659194
rect 42182 656322 42380 656350
rect 42156 656192 42208 656198
rect 42156 656134 42208 656140
rect 42168 655656 42196 656134
rect 42444 655126 42472 659670
rect 43088 656198 43116 665207
rect 43180 663610 43208 670534
rect 43258 670511 43314 670520
rect 43168 663604 43220 663610
rect 43168 663546 43220 663552
rect 43272 659530 43300 670511
rect 43364 665242 43392 676602
rect 43456 671129 43484 681702
rect 43442 671120 43498 671129
rect 43442 671055 43498 671064
rect 43548 670834 43576 683674
rect 43628 682508 43680 682514
rect 43628 682450 43680 682456
rect 43640 670857 43668 682450
rect 43720 682236 43772 682242
rect 43720 682178 43772 682184
rect 43456 670806 43576 670834
rect 43626 670848 43682 670857
rect 43352 665236 43404 665242
rect 43352 665178 43404 665184
rect 43352 665100 43404 665106
rect 43352 665042 43404 665048
rect 43260 659524 43312 659530
rect 43260 659466 43312 659472
rect 43364 659258 43392 665042
rect 43352 659252 43404 659258
rect 43352 659194 43404 659200
rect 43076 656192 43128 656198
rect 43076 656134 43128 656140
rect 42182 655098 42472 655126
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 41510 644736 41566 644745
rect 41510 644671 41512 644680
rect 41564 644671 41566 644680
rect 41512 644642 41564 644648
rect 41510 644328 41566 644337
rect 41510 644263 41512 644272
rect 41564 644263 41566 644272
rect 41512 644234 41564 644240
rect 41786 644124 41842 644133
rect 41786 644059 41788 644068
rect 41840 644059 41842 644068
rect 41788 644030 41840 644036
rect 41512 644020 41564 644026
rect 41512 643962 41564 643968
rect 41524 643929 41552 643962
rect 41510 643920 41566 643929
rect 41510 643855 41566 643864
rect 41786 643308 41842 643317
rect 41786 643243 41788 643252
rect 41840 643243 41842 643252
rect 41788 643214 41840 643220
rect 41510 643104 41566 643113
rect 41510 643039 41512 643048
rect 41564 643039 41566 643048
rect 41512 643010 41564 643016
rect 43456 642870 43484 670806
rect 43626 670783 43682 670792
rect 43536 670744 43588 670750
rect 43536 670686 43588 670692
rect 43548 643074 43576 670686
rect 43732 670682 43760 682178
rect 43904 680060 43956 680066
rect 43904 680002 43956 680008
rect 43812 679924 43864 679930
rect 43812 679866 43864 679872
rect 43720 670676 43772 670682
rect 43720 670618 43772 670624
rect 43628 670608 43680 670614
rect 43628 670550 43680 670556
rect 43718 670576 43774 670585
rect 43640 661094 43668 670550
rect 43718 670511 43774 670520
rect 43732 663066 43760 670511
rect 43824 667282 43852 679866
rect 43916 670546 43944 680002
rect 43904 670540 43956 670546
rect 43904 670482 43956 670488
rect 43902 670440 43958 670449
rect 43902 670375 43958 670384
rect 43812 667276 43864 667282
rect 43812 667218 43864 667224
rect 43812 667140 43864 667146
rect 43812 667082 43864 667088
rect 43720 663060 43772 663066
rect 43720 663002 43772 663008
rect 43628 661088 43680 661094
rect 43628 661030 43680 661036
rect 43824 659054 43852 667082
rect 43812 659048 43864 659054
rect 43812 658990 43864 658996
rect 43916 657422 43944 670375
rect 43904 657416 43956 657422
rect 43904 657358 43956 657364
rect 44008 644026 44036 686122
rect 44088 679380 44140 679386
rect 44088 679322 44140 679328
rect 44100 670834 44128 679322
rect 44100 670806 44220 670834
rect 44086 670712 44142 670721
rect 44086 670647 44142 670656
rect 43996 644020 44048 644026
rect 43996 643962 44048 643968
rect 43812 643272 43864 643278
rect 43812 643214 43864 643220
rect 43536 643068 43588 643074
rect 43536 643010 43588 643016
rect 41512 642864 41564 642870
rect 41512 642806 41564 642812
rect 43444 642864 43496 642870
rect 43444 642806 43496 642812
rect 41524 641481 41552 642806
rect 41788 642728 41840 642734
rect 41788 642670 41840 642676
rect 41602 642288 41658 642297
rect 41602 642223 41658 642232
rect 41510 641472 41566 641481
rect 41510 641407 41566 641416
rect 41510 640656 41566 640665
rect 41510 640591 41512 640600
rect 41564 640591 41566 640600
rect 41512 640562 41564 640568
rect 41616 640354 41644 642223
rect 41800 642093 41828 642670
rect 41786 642084 41842 642093
rect 41786 642019 41842 642028
rect 41786 641676 41842 641685
rect 41786 641611 41842 641620
rect 41800 640558 41828 641611
rect 43720 640620 43772 640626
rect 43720 640562 43772 640568
rect 41788 640552 41840 640558
rect 41788 640494 41840 640500
rect 43260 640552 43312 640558
rect 43260 640494 43312 640500
rect 41786 640452 41842 640461
rect 41786 640387 41788 640396
rect 41840 640387 41842 640396
rect 42708 640416 42760 640422
rect 41788 640358 41840 640364
rect 42708 640358 42760 640364
rect 41604 640348 41656 640354
rect 41604 640290 41656 640296
rect 42338 639976 42394 639985
rect 42338 639911 42394 639920
rect 41510 639432 41566 639441
rect 41510 639367 41566 639376
rect 41524 639130 41552 639367
rect 41512 639124 41564 639130
rect 41512 639066 41564 639072
rect 41510 639024 41566 639033
rect 41510 638959 41566 638968
rect 41524 638042 41552 638959
rect 41786 638820 41842 638829
rect 41786 638755 41842 638764
rect 41800 638518 41828 638755
rect 41788 638512 41840 638518
rect 41788 638454 41840 638460
rect 41786 638412 41842 638421
rect 41786 638347 41842 638356
rect 41512 638036 41564 638042
rect 41512 637978 41564 637984
rect 41510 637800 41566 637809
rect 41510 637735 41512 637744
rect 41564 637735 41566 637744
rect 41512 637706 41564 637712
rect 38106 636984 38162 636993
rect 38106 636919 38162 636928
rect 38120 631922 38148 636919
rect 41510 636576 41566 636585
rect 41510 636511 41566 636520
rect 38198 635760 38254 635769
rect 38198 635695 38254 635704
rect 38108 631916 38160 631922
rect 38108 631858 38160 631864
rect 38212 631854 38240 635695
rect 41524 634914 41552 636511
rect 41602 636168 41658 636177
rect 41602 636103 41658 636112
rect 41616 635458 41644 636103
rect 41604 635452 41656 635458
rect 41604 635394 41656 635400
rect 41602 635352 41658 635361
rect 41602 635287 41658 635296
rect 41616 635186 41644 635287
rect 41604 635180 41656 635186
rect 41604 635122 41656 635128
rect 41602 634944 41658 634953
rect 41512 634908 41564 634914
rect 41602 634879 41658 634888
rect 41512 634850 41564 634856
rect 41616 634846 41644 634879
rect 41604 634840 41656 634846
rect 41604 634782 41656 634788
rect 41510 634536 41566 634545
rect 41510 634471 41566 634480
rect 41524 633321 41552 634471
rect 41510 633312 41566 633321
rect 41510 633247 41512 633256
rect 41564 633247 41566 633256
rect 41512 633218 41564 633224
rect 41694 631952 41750 631961
rect 41694 631887 41750 631896
rect 38200 631848 38252 631854
rect 38200 631790 38252 631796
rect 41708 627722 41736 631887
rect 41800 629354 41828 638347
rect 41878 637596 41934 637605
rect 41878 637531 41934 637540
rect 41892 629474 41920 637531
rect 41880 629468 41932 629474
rect 41880 629410 41932 629416
rect 41800 629326 42288 629354
rect 41708 627694 41828 627722
rect 41800 627473 41828 627694
rect 41786 627464 41842 627473
rect 41786 627399 41842 627408
rect 42260 627178 42288 629326
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42248 626748 42300 626754
rect 42248 626690 42300 626696
rect 42156 625320 42208 625326
rect 42156 625262 42208 625268
rect 42168 624784 42196 625262
rect 42260 624306 42288 626690
rect 42352 625326 42380 639911
rect 42432 629740 42484 629746
rect 42432 629682 42484 629688
rect 42444 627473 42472 629682
rect 42430 627464 42486 627473
rect 42430 627399 42486 627408
rect 42720 626754 42748 640358
rect 43168 638036 43220 638042
rect 43168 637978 43220 637984
rect 43076 637764 43128 637770
rect 43076 637706 43128 637712
rect 43088 631990 43116 637706
rect 43180 632058 43208 637978
rect 43168 632052 43220 632058
rect 43168 631994 43220 632000
rect 43076 631984 43128 631990
rect 43076 631926 43128 631932
rect 43168 631916 43220 631922
rect 43168 631858 43220 631864
rect 43076 631848 43128 631854
rect 43076 631790 43128 631796
rect 42708 626748 42760 626754
rect 42708 626690 42760 626696
rect 42708 626612 42760 626618
rect 42708 626554 42760 626560
rect 42340 625320 42392 625326
rect 42340 625262 42392 625268
rect 42720 624510 42748 626554
rect 42340 624504 42392 624510
rect 42340 624446 42392 624452
rect 42708 624504 42760 624510
rect 42708 624446 42760 624452
rect 42248 624300 42300 624306
rect 42248 624242 42300 624248
rect 42182 624158 42288 624186
rect 42156 623484 42208 623490
rect 42156 623426 42208 623432
rect 42168 622948 42196 623426
rect 42156 622872 42208 622878
rect 42156 622814 42208 622820
rect 42168 622336 42196 622814
rect 42260 622690 42288 624158
rect 42352 622878 42380 624446
rect 42708 624300 42760 624306
rect 42708 624242 42760 624248
rect 42340 622872 42392 622878
rect 42340 622814 42392 622820
rect 42260 622662 42380 622690
rect 42062 622024 42118 622033
rect 42062 621959 42118 621968
rect 42076 621792 42104 621959
rect 41878 621480 41934 621489
rect 41878 621415 41934 621424
rect 41892 621112 41920 621415
rect 42064 620832 42116 620838
rect 42064 620774 42116 620780
rect 42076 620500 42104 620774
rect 42064 620356 42116 620362
rect 42064 620298 42116 620304
rect 42076 619956 42104 620298
rect 42352 618254 42380 622662
rect 42432 619200 42484 619206
rect 42432 619142 42484 619148
rect 42340 618248 42392 618254
rect 42340 618190 42392 618196
rect 42444 617454 42472 619142
rect 42182 617426 42472 617454
rect 42432 617364 42484 617370
rect 42432 617306 42484 617312
rect 42444 616842 42472 617306
rect 42168 616706 42196 616828
rect 42260 616814 42472 616842
rect 42260 616706 42288 616814
rect 42168 616678 42288 616706
rect 42432 616752 42484 616758
rect 42432 616694 42484 616700
rect 42444 616162 42472 616694
rect 42182 616134 42472 616162
rect 42432 616072 42484 616078
rect 42432 616014 42484 616020
rect 42444 615618 42472 616014
rect 42182 615590 42472 615618
rect 42340 615528 42392 615534
rect 42340 615470 42392 615476
rect 42156 614236 42208 614242
rect 42156 614178 42208 614184
rect 42168 613768 42196 614178
rect 42248 614100 42300 614106
rect 42248 614042 42300 614048
rect 42156 613488 42208 613494
rect 42156 613430 42208 613436
rect 42168 613121 42196 613430
rect 42260 612490 42288 614042
rect 42182 612462 42288 612490
rect 42352 611946 42380 615470
rect 42720 614242 42748 624242
rect 43088 619206 43116 631790
rect 43076 619200 43128 619206
rect 43076 619142 43128 619148
rect 43180 617370 43208 631858
rect 43168 617364 43220 617370
rect 43168 617306 43220 617312
rect 42708 614236 42760 614242
rect 42708 614178 42760 614184
rect 42182 611918 42380 611946
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 41786 601760 41842 601769
rect 41786 601695 41788 601704
rect 41840 601695 41842 601704
rect 41788 601666 41840 601672
rect 41786 601352 41842 601361
rect 41786 601287 41788 601296
rect 41840 601287 41842 601296
rect 41788 601258 41840 601264
rect 41512 601044 41564 601050
rect 41512 600986 41564 600992
rect 41524 600681 41552 600986
rect 41786 600944 41842 600953
rect 41786 600879 41788 600888
rect 41840 600879 41842 600888
rect 41788 600850 41840 600856
rect 41510 600672 41566 600681
rect 41510 600607 41566 600616
rect 41512 600364 41564 600370
rect 41512 600306 41564 600312
rect 41524 599865 41552 600306
rect 41786 600128 41842 600137
rect 41786 600063 41842 600072
rect 41510 599856 41566 599865
rect 41510 599791 41566 599800
rect 41800 599078 41828 600063
rect 41788 599072 41840 599078
rect 41510 599040 41566 599049
rect 41788 599014 41840 599020
rect 41510 598975 41512 598984
rect 41564 598975 41566 598984
rect 41512 598946 41564 598952
rect 43272 598942 43300 640494
rect 43352 640348 43404 640354
rect 43352 640290 43404 640296
rect 43364 600370 43392 640290
rect 43628 639124 43680 639130
rect 43628 639066 43680 639072
rect 43444 638512 43496 638518
rect 43444 638454 43496 638460
rect 43456 629610 43484 638454
rect 43536 634908 43588 634914
rect 43536 634850 43588 634856
rect 43444 629604 43496 629610
rect 43444 629546 43496 629552
rect 43444 629468 43496 629474
rect 43444 629410 43496 629416
rect 43456 616758 43484 629410
rect 43548 623490 43576 634850
rect 43536 623484 43588 623490
rect 43536 623426 43588 623432
rect 43536 623348 43588 623354
rect 43536 623290 43588 623296
rect 43548 620838 43576 623290
rect 43536 620832 43588 620838
rect 43536 620774 43588 620780
rect 43444 616752 43496 616758
rect 43444 616694 43496 616700
rect 43640 614106 43668 639066
rect 43628 614100 43680 614106
rect 43628 614042 43680 614048
rect 43352 600364 43404 600370
rect 43352 600306 43404 600312
rect 43352 599004 43404 599010
rect 43352 598946 43404 598952
rect 41788 598936 41840 598942
rect 41786 598904 41788 598913
rect 43260 598936 43312 598942
rect 41840 598904 41842 598913
rect 43260 598878 43312 598884
rect 41786 598839 41842 598848
rect 41512 598528 41564 598534
rect 41512 598470 41564 598476
rect 42430 598496 42486 598505
rect 41524 598233 41552 598470
rect 42430 598431 42486 598440
rect 41510 598224 41566 598233
rect 41510 598159 41566 598168
rect 41510 597408 41566 597417
rect 41510 597343 41566 597352
rect 41524 597106 41552 597343
rect 41512 597100 41564 597106
rect 41512 597042 41564 597048
rect 41510 597000 41566 597009
rect 41510 596935 41566 596944
rect 41524 596698 41552 596935
rect 41512 596692 41564 596698
rect 41512 596634 41564 596640
rect 41510 596592 41566 596601
rect 41510 596527 41566 596536
rect 41524 596426 41552 596527
rect 42154 596456 42210 596465
rect 41512 596420 41564 596426
rect 42154 596391 42210 596400
rect 41512 596362 41564 596368
rect 41510 595776 41566 595785
rect 41510 595711 41566 595720
rect 41524 595474 41552 595711
rect 41512 595468 41564 595474
rect 41512 595410 41564 595416
rect 41510 595368 41566 595377
rect 41510 595303 41566 595312
rect 41524 594658 41552 595303
rect 41878 595232 41934 595241
rect 41878 595167 41934 595176
rect 41512 594652 41564 594658
rect 41512 594594 41564 594600
rect 41510 594552 41566 594561
rect 41510 594487 41566 594496
rect 38014 594144 38070 594153
rect 41524 594114 41552 594487
rect 38014 594079 38070 594088
rect 41512 594108 41564 594114
rect 38028 587858 38056 594079
rect 41512 594050 41564 594056
rect 38106 593736 38162 593745
rect 38106 593671 38162 593680
rect 38016 587852 38068 587858
rect 38016 587794 38068 587800
rect 38120 587790 38148 593671
rect 41786 593600 41842 593609
rect 41786 593535 41788 593544
rect 41840 593535 41842 593544
rect 41788 593506 41840 593512
rect 41892 593414 41920 595167
rect 41800 593386 41920 593414
rect 41510 592920 41566 592929
rect 41510 592855 41566 592864
rect 41524 592210 41552 592855
rect 41694 592512 41750 592521
rect 41694 592447 41750 592456
rect 41512 592204 41564 592210
rect 41512 592146 41564 592152
rect 41510 592104 41566 592113
rect 41510 592039 41566 592048
rect 41524 591802 41552 592039
rect 41512 591796 41564 591802
rect 41512 591738 41564 591744
rect 41510 591696 41566 591705
rect 41510 591631 41566 591640
rect 41418 591288 41474 591297
rect 41524 591258 41552 591631
rect 41418 591223 41474 591232
rect 41512 591252 41564 591258
rect 41432 590050 41460 591223
rect 41512 591194 41564 591200
rect 41510 590064 41566 590073
rect 41432 590022 41510 590050
rect 41510 589999 41512 590008
rect 41564 589999 41566 590008
rect 41512 589970 41564 589976
rect 41708 588282 41736 592447
rect 41800 588418 41828 593386
rect 42168 588538 42196 596391
rect 42340 591932 42392 591938
rect 42340 591874 42392 591880
rect 42156 588532 42208 588538
rect 42156 588474 42208 588480
rect 41800 588390 42288 588418
rect 41708 588254 41828 588282
rect 38108 587784 38160 587790
rect 38108 587726 38160 587732
rect 41420 587784 41472 587790
rect 41420 587726 41472 587732
rect 41432 585274 41460 587726
rect 41420 585268 41472 585274
rect 41420 585210 41472 585216
rect 41800 584225 41828 588254
rect 41786 584216 41842 584225
rect 41786 584151 41842 584160
rect 42260 583454 42288 588390
rect 42352 585313 42380 591874
rect 42338 585304 42394 585313
rect 42338 585239 42394 585248
rect 42340 585200 42392 585206
rect 42340 585142 42392 585148
rect 42182 583426 42288 583454
rect 42248 582616 42300 582622
rect 42248 582558 42300 582564
rect 42156 582140 42208 582146
rect 42156 582082 42208 582088
rect 42168 581604 42196 582082
rect 42260 581330 42288 582558
rect 42248 581324 42300 581330
rect 42248 581266 42300 581272
rect 42352 581210 42380 585142
rect 42444 584254 42472 598431
rect 43168 594108 43220 594114
rect 43168 594050 43220 594056
rect 43076 593564 43128 593570
rect 43076 593506 43128 593512
rect 42708 587852 42760 587858
rect 42708 587794 42760 587800
rect 42432 584248 42484 584254
rect 42432 584190 42484 584196
rect 42720 583953 42748 587794
rect 42706 583944 42762 583953
rect 42706 583879 42762 583888
rect 42708 583772 42760 583778
rect 42708 583714 42760 583720
rect 42168 581182 42380 581210
rect 42168 580961 42196 581182
rect 42248 581120 42300 581126
rect 42300 581068 42380 581074
rect 42248 581062 42380 581068
rect 42260 581046 42380 581062
rect 42352 580802 42380 581046
rect 42168 580774 42380 580802
rect 42168 580530 42196 580774
rect 42246 580680 42302 580689
rect 42302 580638 42380 580666
rect 42246 580615 42302 580624
rect 42168 580502 42288 580530
rect 42156 580304 42208 580310
rect 42156 580246 42208 580252
rect 42168 579768 42196 580246
rect 42260 579135 42288 580502
rect 42182 579107 42288 579135
rect 42248 579012 42300 579018
rect 42248 578954 42300 578960
rect 42156 578808 42208 578814
rect 42156 578750 42208 578756
rect 42168 578544 42196 578750
rect 42156 578468 42208 578474
rect 42156 578410 42208 578416
rect 42168 577932 42196 578410
rect 42260 577295 42288 578954
rect 42182 577267 42288 577295
rect 42154 577008 42210 577017
rect 42154 576943 42210 576952
rect 42168 576708 42196 576943
rect 42352 574274 42380 580638
rect 42182 574246 42380 574274
rect 42340 574184 42392 574190
rect 42340 574126 42392 574132
rect 42352 574094 42380 574126
rect 42260 574066 42380 574094
rect 42432 574116 42484 574122
rect 42156 573844 42208 573850
rect 42156 573786 42208 573792
rect 42168 573580 42196 573786
rect 42260 573458 42288 574066
rect 42432 574058 42484 574064
rect 42168 573430 42288 573458
rect 42168 572968 42196 573430
rect 42064 572688 42116 572694
rect 42064 572630 42116 572636
rect 42076 572424 42104 572630
rect 42248 572008 42300 572014
rect 42248 571950 42300 571956
rect 42064 570988 42116 570994
rect 42064 570930 42116 570936
rect 42076 570588 42104 570930
rect 42260 569922 42288 571950
rect 42182 569894 42288 569922
rect 42064 569628 42116 569634
rect 42064 569570 42116 569576
rect 42076 569296 42104 569570
rect 42444 568766 42472 574058
rect 42720 572014 42748 583714
rect 43088 580310 43116 593506
rect 43180 583778 43208 594050
rect 43260 591252 43312 591258
rect 43260 591194 43312 591200
rect 43168 583772 43220 583778
rect 43168 583714 43220 583720
rect 43168 583636 43220 583642
rect 43168 583578 43220 583584
rect 43180 582010 43208 583578
rect 43168 582004 43220 582010
rect 43168 581946 43220 581952
rect 43166 581904 43222 581913
rect 43166 581839 43222 581848
rect 43076 580304 43128 580310
rect 43076 580246 43128 580252
rect 43076 580168 43128 580174
rect 43076 580110 43128 580116
rect 42708 572008 42760 572014
rect 42708 571950 42760 571956
rect 43088 570994 43116 580110
rect 43180 574190 43208 581839
rect 43272 578814 43300 591194
rect 43260 578808 43312 578814
rect 43260 578750 43312 578756
rect 43168 574184 43220 574190
rect 43168 574126 43220 574132
rect 43076 570988 43128 570994
rect 43076 570930 43128 570936
rect 42168 568698 42196 568752
rect 42260 568738 42472 568766
rect 42260 568698 42288 568738
rect 42168 568670 42288 568698
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 41510 558376 41566 558385
rect 41510 558311 41512 558320
rect 41564 558311 41566 558320
rect 41512 558282 41564 558288
rect 41510 557968 41566 557977
rect 41510 557903 41512 557912
rect 41564 557903 41566 557912
rect 41512 557874 41564 557880
rect 41512 557592 41564 557598
rect 41510 557560 41512 557569
rect 41564 557560 41566 557569
rect 41510 557495 41566 557504
rect 41788 557320 41840 557326
rect 41786 557288 41788 557297
rect 41840 557288 41842 557297
rect 41786 557223 41842 557232
rect 43364 556850 43392 598946
rect 43732 598534 43760 640562
rect 43824 601050 43852 643214
rect 44100 642734 44128 670647
rect 44192 667826 44220 670806
rect 44272 670676 44324 670682
rect 44272 670618 44324 670624
rect 44180 667820 44232 667826
rect 44180 667762 44232 667768
rect 44284 667146 44312 670618
rect 44364 670540 44416 670546
rect 44364 670482 44416 670488
rect 44272 667140 44324 667146
rect 44272 667082 44324 667088
rect 44376 665106 44404 670482
rect 44364 665100 44416 665106
rect 44364 665042 44416 665048
rect 44088 642728 44140 642734
rect 44088 642670 44140 642676
rect 43904 635452 43956 635458
rect 43904 635394 43956 635400
rect 43916 632097 43944 635394
rect 44088 635180 44140 635186
rect 44088 635122 44140 635128
rect 43996 634840 44048 634846
rect 43996 634782 44048 634788
rect 43902 632088 43958 632097
rect 43902 632023 43958 632032
rect 44008 631938 44036 634782
rect 43916 631910 44036 631938
rect 44100 631938 44128 635122
rect 44100 631910 44220 631938
rect 43916 629746 43944 631910
rect 43996 631848 44048 631854
rect 43996 631790 44048 631796
rect 43904 629740 43956 629746
rect 43904 629682 43956 629688
rect 43904 629604 43956 629610
rect 43904 629546 43956 629552
rect 43916 620362 43944 629546
rect 43904 620356 43956 620362
rect 43904 620298 43956 620304
rect 44008 616078 44036 631790
rect 44088 631780 44140 631786
rect 44088 631722 44140 631728
rect 43996 616072 44048 616078
rect 43996 616014 44048 616020
rect 44100 613494 44128 631722
rect 44192 623354 44220 631910
rect 44180 623348 44232 623354
rect 44180 623290 44232 623296
rect 44088 613488 44140 613494
rect 44088 613430 44140 613436
rect 43812 601044 43864 601050
rect 43812 600986 43864 600992
rect 43996 599072 44048 599078
rect 43996 599014 44048 599020
rect 43720 598528 43772 598534
rect 43720 598470 43772 598476
rect 43812 596692 43864 596698
rect 43812 596634 43864 596640
rect 43628 596420 43680 596426
rect 43628 596362 43680 596368
rect 43444 595468 43496 595474
rect 43444 595410 43496 595416
rect 43456 572694 43484 595410
rect 43536 594652 43588 594658
rect 43536 594594 43588 594600
rect 43548 591938 43576 594594
rect 43536 591932 43588 591938
rect 43536 591874 43588 591880
rect 43536 591796 43588 591802
rect 43536 591738 43588 591744
rect 43548 579018 43576 591738
rect 43640 582146 43668 596362
rect 43720 592204 43772 592210
rect 43720 592146 43772 592152
rect 43628 582140 43680 582146
rect 43628 582082 43680 582088
rect 43628 582004 43680 582010
rect 43628 581946 43680 581952
rect 43536 579012 43588 579018
rect 43536 578954 43588 578960
rect 43536 578876 43588 578882
rect 43536 578818 43588 578824
rect 43444 572688 43496 572694
rect 43444 572630 43496 572636
rect 43548 569634 43576 578818
rect 43536 569628 43588 569634
rect 43536 569570 43588 569576
rect 41788 556844 41840 556850
rect 41788 556786 41840 556792
rect 43352 556844 43404 556850
rect 43352 556786 43404 556792
rect 41512 556708 41564 556714
rect 41512 556650 41564 556656
rect 41524 555937 41552 556650
rect 41800 556481 41828 556786
rect 43640 556714 43668 581946
rect 43732 578474 43760 592146
rect 43824 580174 43852 596634
rect 43904 588532 43956 588538
rect 43904 588474 43956 588480
rect 43916 583914 43944 588474
rect 43904 583908 43956 583914
rect 43904 583850 43956 583856
rect 43902 583808 43958 583817
rect 43902 583743 43958 583752
rect 43812 580168 43864 580174
rect 43812 580110 43864 580116
rect 43720 578468 43772 578474
rect 43720 578410 43772 578416
rect 43628 556708 43680 556714
rect 43628 556650 43680 556656
rect 41786 556472 41842 556481
rect 41786 556407 41842 556416
rect 41510 555928 41566 555937
rect 41510 555863 41566 555872
rect 43916 554810 43944 583743
rect 44008 557326 44036 599014
rect 44088 597100 44140 597106
rect 44088 597042 44140 597048
rect 44100 583817 44128 597042
rect 44180 585268 44232 585274
rect 44180 585210 44232 585216
rect 44086 583808 44142 583817
rect 44086 583743 44142 583752
rect 44088 583704 44140 583710
rect 44088 583646 44140 583652
rect 44100 578882 44128 583646
rect 44088 578876 44140 578882
rect 44088 578818 44140 578824
rect 44192 578762 44220 585210
rect 44100 578734 44220 578762
rect 44100 573850 44128 578734
rect 44088 573844 44140 573850
rect 44088 573786 44140 573792
rect 43996 557320 44048 557326
rect 43996 557262 44048 557268
rect 38568 554804 38620 554810
rect 38568 554746 38620 554752
rect 43904 554804 43956 554810
rect 43904 554746 43956 554752
rect 38580 554713 38608 554746
rect 38566 554704 38622 554713
rect 38566 554639 38622 554648
rect 41510 553480 41566 553489
rect 41510 553415 41566 553424
rect 41524 552362 41552 553415
rect 41512 552356 41564 552362
rect 41512 552298 41564 552304
rect 43260 552356 43312 552362
rect 43260 552298 43312 552304
rect 41786 551984 41842 551993
rect 41786 551919 41842 551928
rect 41510 550216 41566 550225
rect 41510 550151 41566 550160
rect 41418 549808 41474 549817
rect 41418 549743 41420 549752
rect 41472 549743 41474 549752
rect 41420 549714 41472 549720
rect 41524 549642 41552 550151
rect 41512 549636 41564 549642
rect 41512 549578 41564 549584
rect 41510 549400 41566 549409
rect 41510 549335 41512 549344
rect 41564 549335 41566 549344
rect 41512 549306 41564 549312
rect 41510 548992 41566 549001
rect 41510 548927 41566 548936
rect 41524 548690 41552 548927
rect 41512 548684 41564 548690
rect 41512 548626 41564 548632
rect 41510 548584 41566 548593
rect 41510 548519 41566 548528
rect 41418 548176 41474 548185
rect 41418 548111 41474 548120
rect 41432 546938 41460 548111
rect 41524 547058 41552 548519
rect 41512 547052 41564 547058
rect 41512 546994 41564 547000
rect 41510 546952 41566 546961
rect 41432 546910 41510 546938
rect 41510 546887 41512 546896
rect 41564 546887 41566 546896
rect 41512 546858 41564 546864
rect 41800 546494 41828 551919
rect 43076 549636 43128 549642
rect 43076 549578 43128 549584
rect 41800 546466 42288 546494
rect 42260 540274 42288 546466
rect 43088 541226 43116 549578
rect 43168 547052 43220 547058
rect 43168 546994 43220 547000
rect 43180 541346 43208 546994
rect 43168 541340 43220 541346
rect 43168 541282 43220 541288
rect 43088 541198 43208 541226
rect 43076 541068 43128 541074
rect 43076 541010 43128 541016
rect 42708 541000 42760 541006
rect 42708 540942 42760 540948
rect 42182 540246 42288 540274
rect 42064 538960 42116 538966
rect 42064 538902 42116 538908
rect 42076 538424 42104 538902
rect 42248 538484 42300 538490
rect 42248 538426 42300 538432
rect 42156 538280 42208 538286
rect 42156 538222 42208 538228
rect 42168 537744 42196 538222
rect 42064 537124 42116 537130
rect 42064 537066 42116 537072
rect 42076 536588 42104 537066
rect 42260 535922 42288 538426
rect 42720 538286 42748 540942
rect 43088 538490 43116 541010
rect 43076 538484 43128 538490
rect 43076 538426 43128 538432
rect 43074 538384 43130 538393
rect 43074 538319 43130 538328
rect 42708 538280 42760 538286
rect 42708 538222 42760 538228
rect 42706 538112 42762 538121
rect 42706 538047 42762 538056
rect 42182 535894 42288 535922
rect 42156 535628 42208 535634
rect 42156 535570 42208 535576
rect 42168 535364 42196 535570
rect 42246 535392 42302 535401
rect 42246 535327 42302 535336
rect 42064 535084 42116 535090
rect 42064 535026 42116 535032
rect 42076 534752 42104 535026
rect 42156 534472 42208 534478
rect 42156 534414 42208 534420
rect 42168 534072 42196 534414
rect 42156 533996 42208 534002
rect 42156 533938 42208 533944
rect 42168 533528 42196 533938
rect 42156 531480 42208 531486
rect 42156 531422 42208 531428
rect 42168 531045 42196 531422
rect 42156 530936 42208 530942
rect 42156 530878 42208 530884
rect 42168 530400 42196 530878
rect 42260 529771 42288 535327
rect 42430 532808 42486 532817
rect 42430 532743 42486 532752
rect 42338 532672 42394 532681
rect 42338 532607 42394 532616
rect 42182 529743 42288 529771
rect 42248 529644 42300 529650
rect 42248 529586 42300 529592
rect 42260 529219 42288 529586
rect 42182 529191 42288 529219
rect 42156 527808 42208 527814
rect 42156 527750 42208 527756
rect 42168 527340 42196 527750
rect 42352 526742 42380 532607
rect 42444 530126 42472 532743
rect 42720 530942 42748 538047
rect 43088 534002 43116 538319
rect 43180 537130 43208 541198
rect 43272 538966 43300 552298
rect 43352 549772 43404 549778
rect 43352 549714 43404 549720
rect 43364 541498 43392 549714
rect 43444 549364 43496 549370
rect 43444 549306 43496 549312
rect 43456 546494 43484 549306
rect 43904 548684 43956 548690
rect 43904 548626 43956 548632
rect 43456 546466 43576 546494
rect 43364 541470 43484 541498
rect 43352 541340 43404 541346
rect 43352 541282 43404 541288
rect 43260 538960 43312 538966
rect 43260 538902 43312 538908
rect 43168 537124 43220 537130
rect 43168 537066 43220 537072
rect 43364 535634 43392 541282
rect 43352 535628 43404 535634
rect 43352 535570 43404 535576
rect 43166 535392 43222 535401
rect 43166 535327 43222 535336
rect 43076 533996 43128 534002
rect 43076 533938 43128 533944
rect 43074 532672 43130 532681
rect 43074 532607 43130 532616
rect 42708 530936 42760 530942
rect 42708 530878 42760 530884
rect 42432 530120 42484 530126
rect 42432 530062 42484 530068
rect 42432 529984 42484 529990
rect 42432 529926 42484 529932
rect 42182 526714 42380 526742
rect 42340 526652 42392 526658
rect 42340 526594 42392 526600
rect 42352 526091 42380 526594
rect 42182 526063 42380 526091
rect 42168 525558 42288 525586
rect 42168 525504 42196 525558
rect 42260 525518 42288 525558
rect 42444 525518 42472 529926
rect 43088 526658 43116 532607
rect 43180 527814 43208 535327
rect 43456 535090 43484 541470
rect 43444 535084 43496 535090
rect 43444 535026 43496 535032
rect 43548 531486 43576 546466
rect 43626 538520 43682 538529
rect 43626 538455 43682 538464
rect 43536 531480 43588 531486
rect 43536 531422 43588 531428
rect 43168 527808 43220 527814
rect 43168 527750 43220 527756
rect 43640 527174 43668 538455
rect 43718 538248 43774 538257
rect 43718 538183 43774 538192
rect 43548 527146 43668 527174
rect 43076 526652 43128 526658
rect 43076 526594 43128 526600
rect 42260 525490 42472 525518
rect 43548 516134 43576 527146
rect 43364 516106 43576 516134
rect 41878 435976 41934 435985
rect 41878 435911 41934 435920
rect 8588 431596 8616 431732
rect 9048 431596 9076 431732
rect 9508 431596 9536 431732
rect 9968 431596 9996 431732
rect 10428 431596 10456 431732
rect 10888 431596 10916 431732
rect 11348 431596 11376 431732
rect 11808 431596 11836 431732
rect 12268 431596 12296 431732
rect 12728 431596 12756 431732
rect 13188 431596 13216 431732
rect 13648 431596 13676 431732
rect 14108 431596 14136 431732
rect 41786 430944 41842 430953
rect 41786 430879 41788 430888
rect 41840 430879 41842 430888
rect 41788 430850 41840 430856
rect 41786 430536 41842 430545
rect 41786 430471 41788 430480
rect 41840 430471 41842 430480
rect 41788 430442 41840 430448
rect 41786 430128 41842 430137
rect 41786 430063 41788 430072
rect 41840 430063 41842 430072
rect 41788 430034 41840 430040
rect 41788 429956 41840 429962
rect 41788 429898 41840 429904
rect 41800 429729 41828 429898
rect 41786 429720 41842 429729
rect 41786 429655 41842 429664
rect 41786 429312 41842 429321
rect 41786 429247 41842 429256
rect 41800 429078 41828 429247
rect 41788 429072 41840 429078
rect 41788 429014 41840 429020
rect 41788 428936 41840 428942
rect 41786 428904 41788 428913
rect 41840 428904 41842 428913
rect 41786 428839 41842 428848
rect 41892 427281 41920 435911
rect 43364 429962 43392 516106
rect 43352 429956 43404 429962
rect 43352 429898 43404 429904
rect 43732 428942 43760 538183
rect 43916 534478 43944 548626
rect 43904 534472 43956 534478
rect 43904 534414 43956 534420
rect 43904 429072 43956 429078
rect 43904 429014 43956 429020
rect 43720 428936 43772 428942
rect 43720 428878 43772 428884
rect 42430 428496 42486 428505
rect 42430 428431 42486 428440
rect 42062 427680 42118 427689
rect 42062 427615 42118 427624
rect 41878 427272 41934 427281
rect 41878 427207 41934 427216
rect 41786 426864 41842 426873
rect 41786 426799 41842 426808
rect 41800 426562 41828 426799
rect 41788 426556 41840 426562
rect 41788 426498 41840 426504
rect 41786 426456 41842 426465
rect 41786 426391 41788 426400
rect 41840 426391 41842 426400
rect 41788 426362 41840 426368
rect 41970 426048 42026 426057
rect 41970 425983 42026 425992
rect 41786 425640 41842 425649
rect 41786 425575 41842 425584
rect 41800 425474 41828 425575
rect 41788 425468 41840 425474
rect 41788 425410 41840 425416
rect 41786 425232 41842 425241
rect 41786 425167 41788 425176
rect 41840 425167 41842 425176
rect 41788 425138 41840 425144
rect 41786 424824 41842 424833
rect 41786 424759 41842 424768
rect 41800 422482 41828 424759
rect 41878 424008 41934 424017
rect 41878 423943 41934 423952
rect 41892 423706 41920 423943
rect 41880 423700 41932 423706
rect 41880 423642 41932 423648
rect 41878 423600 41934 423609
rect 41878 423535 41880 423544
rect 41932 423535 41934 423544
rect 41880 423506 41932 423512
rect 41878 423192 41934 423201
rect 41878 423127 41934 423136
rect 41892 422958 41920 423127
rect 41880 422952 41932 422958
rect 41880 422894 41932 422900
rect 41878 422784 41934 422793
rect 41878 422719 41934 422728
rect 41892 422686 41920 422719
rect 41880 422680 41932 422686
rect 41880 422622 41932 422628
rect 41788 422476 41840 422482
rect 41788 422418 41840 422424
rect 41786 422376 41842 422385
rect 41786 422311 41788 422320
rect 41840 422311 41842 422320
rect 41788 422282 41840 422288
rect 41786 421968 41842 421977
rect 41786 421903 41842 421912
rect 41800 421598 41828 421903
rect 41788 421592 41840 421598
rect 41788 421534 41840 421540
rect 41878 421560 41934 421569
rect 41878 421495 41934 421504
rect 41786 420744 41842 420753
rect 41786 420679 41842 420688
rect 41800 419529 41828 420679
rect 41786 419520 41842 419529
rect 41786 419455 41788 419464
rect 41840 419455 41842 419464
rect 41788 419426 41840 419432
rect 41892 416362 41920 421495
rect 41880 416356 41932 416362
rect 41880 416298 41932 416304
rect 41984 413438 42012 425983
rect 42076 413846 42104 427615
rect 42246 424416 42302 424425
rect 42246 424351 42302 424360
rect 42064 413840 42116 413846
rect 42064 413782 42116 413788
rect 41972 413432 42024 413438
rect 41972 413374 42024 413380
rect 42260 413114 42288 424351
rect 42338 421152 42394 421161
rect 42338 421087 42394 421096
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42248 413024 42300 413030
rect 42248 412966 42300 412972
rect 42260 411254 42288 412966
rect 42168 411226 42288 411254
rect 42168 410788 42196 411226
rect 42168 409766 42196 410176
rect 42352 410122 42380 421087
rect 42444 413778 42472 428431
rect 43720 426556 43772 426562
rect 43720 426498 43772 426504
rect 42708 425468 42760 425474
rect 42708 425410 42760 425416
rect 42432 413772 42484 413778
rect 42432 413714 42484 413720
rect 42260 410094 42380 410122
rect 42156 409760 42208 409766
rect 42156 409702 42208 409708
rect 42156 409488 42208 409494
rect 42156 409430 42208 409436
rect 42168 408952 42196 409430
rect 42168 407930 42196 408340
rect 42156 407924 42208 407930
rect 42156 407866 42208 407872
rect 42168 407674 42196 407796
rect 42260 407674 42288 410094
rect 42340 409760 42392 409766
rect 42340 409702 42392 409708
rect 42168 407646 42288 407674
rect 42248 407584 42300 407590
rect 42248 407526 42300 407532
rect 42260 407130 42288 407526
rect 42182 407102 42288 407130
rect 42064 407040 42116 407046
rect 42064 406982 42116 406988
rect 42076 406504 42104 406982
rect 42248 406972 42300 406978
rect 42248 406914 42300 406920
rect 42260 405943 42288 406914
rect 42182 405915 42288 405943
rect 42352 405686 42380 409702
rect 42340 405680 42392 405686
rect 42340 405622 42392 405628
rect 42340 405544 42392 405550
rect 42340 405486 42392 405492
rect 42352 403458 42380 405486
rect 42720 405210 42748 425410
rect 43260 425196 43312 425202
rect 43260 425138 43312 425144
rect 43076 423564 43128 423570
rect 43076 423506 43128 423512
rect 43088 409358 43116 423506
rect 43168 416356 43220 416362
rect 43168 416298 43220 416304
rect 43076 409352 43128 409358
rect 43076 409294 43128 409300
rect 43076 407924 43128 407930
rect 43076 407866 43128 407872
rect 42432 405204 42484 405210
rect 42432 405146 42484 405152
rect 42708 405204 42760 405210
rect 42708 405146 42760 405152
rect 42182 403430 42380 403458
rect 42340 403368 42392 403374
rect 42340 403310 42392 403316
rect 42352 402815 42380 403310
rect 42182 402787 42380 402815
rect 42248 402620 42300 402626
rect 42248 402562 42300 402568
rect 42156 402552 42208 402558
rect 42156 402494 42208 402500
rect 42168 402152 42196 402494
rect 42156 401872 42208 401878
rect 42156 401814 42208 401820
rect 42168 401608 42196 401814
rect 42156 400240 42208 400246
rect 42156 400182 42208 400188
rect 42168 399772 42196 400182
rect 42260 399135 42288 402562
rect 42182 399107 42288 399135
rect 42444 398494 42472 405146
rect 43088 402966 43116 407866
rect 43180 407046 43208 416298
rect 43272 411505 43300 425138
rect 43536 423700 43588 423706
rect 43536 423642 43588 423648
rect 43444 422680 43496 422686
rect 43444 422622 43496 422628
rect 43352 421592 43404 421598
rect 43352 421534 43404 421540
rect 43258 411496 43314 411505
rect 43258 411431 43314 411440
rect 43260 411324 43312 411330
rect 43260 411266 43312 411272
rect 43168 407040 43220 407046
rect 43168 406982 43220 406988
rect 43166 406872 43222 406881
rect 43166 406807 43222 406816
rect 43076 402960 43128 402966
rect 43076 402902 43128 402908
rect 43180 401878 43208 406807
rect 43168 401872 43220 401878
rect 43168 401814 43220 401820
rect 42182 398466 42472 398494
rect 42168 394670 42196 397936
rect 42156 394664 42208 394670
rect 42156 394606 42208 394612
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 43272 388074 43300 411266
rect 43364 405550 43392 421534
rect 43456 409494 43484 422622
rect 43444 409488 43496 409494
rect 43444 409430 43496 409436
rect 43444 409352 43496 409358
rect 43444 409294 43496 409300
rect 43352 405544 43404 405550
rect 43352 405486 43404 405492
rect 43456 402558 43484 409294
rect 43548 402626 43576 423642
rect 43628 422952 43680 422958
rect 43628 422894 43680 422900
rect 43640 403374 43668 422894
rect 43628 403368 43680 403374
rect 43628 403310 43680 403316
rect 43536 402620 43588 402626
rect 43536 402562 43588 402568
rect 43444 402552 43496 402558
rect 43444 402494 43496 402500
rect 41512 388068 41564 388074
rect 41512 388010 41564 388016
rect 43260 388068 43312 388074
rect 43260 388010 43312 388016
rect 41418 387560 41474 387569
rect 41418 387495 41420 387504
rect 41472 387495 41474 387504
rect 41420 387466 41472 387472
rect 41418 387152 41474 387161
rect 41418 387087 41420 387096
rect 41472 387087 41474 387096
rect 41420 387058 41472 387064
rect 41524 386753 41552 388010
rect 41786 386880 41842 386889
rect 41786 386815 41788 386824
rect 41840 386815 41842 386824
rect 41788 386786 41840 386792
rect 41510 386744 41566 386753
rect 41510 386679 41566 386688
rect 43732 386374 43760 426498
rect 43812 426420 43864 426426
rect 43812 426362 43864 426368
rect 43824 400246 43852 426362
rect 43916 411330 43944 429014
rect 43996 422476 44048 422482
rect 43996 422418 44048 422424
rect 44008 413982 44036 422418
rect 44088 422340 44140 422346
rect 44088 422282 44140 422288
rect 43996 413976 44048 413982
rect 43996 413918 44048 413924
rect 44100 413914 44128 422282
rect 44272 413976 44324 413982
rect 44272 413918 44324 413924
rect 44088 413908 44140 413914
rect 44088 413850 44140 413856
rect 44180 413908 44232 413914
rect 44180 413850 44232 413856
rect 43996 413840 44048 413846
rect 43996 413782 44048 413788
rect 43904 411324 43956 411330
rect 43904 411266 43956 411272
rect 43904 411188 43956 411194
rect 43904 411130 43956 411136
rect 43916 407590 43944 411130
rect 43904 407584 43956 407590
rect 43904 407526 43956 407532
rect 43812 400240 43864 400246
rect 43812 400182 43864 400188
rect 41788 386368 41840 386374
rect 41788 386310 41840 386316
rect 43720 386368 43772 386374
rect 43720 386310 43772 386316
rect 41512 386096 41564 386102
rect 41512 386038 41564 386044
rect 41524 385937 41552 386038
rect 41510 385928 41566 385937
rect 41510 385863 41566 385872
rect 41512 385824 41564 385830
rect 41512 385766 41564 385772
rect 41524 385121 41552 385766
rect 41510 385112 41566 385121
rect 41510 385047 41566 385056
rect 41510 384296 41566 384305
rect 41510 384231 41566 384240
rect 41524 383722 41552 384231
rect 41800 384033 41828 386310
rect 42430 386064 42486 386073
rect 42430 385999 42486 386008
rect 41878 385248 41934 385257
rect 41878 385183 41934 385192
rect 41786 384024 41842 384033
rect 41786 383959 41842 383968
rect 41892 383790 41920 385183
rect 41880 383784 41932 383790
rect 41880 383726 41932 383732
rect 41512 383716 41564 383722
rect 41512 383658 41564 383664
rect 41510 383480 41566 383489
rect 41510 383415 41566 383424
rect 41524 382770 41552 383415
rect 41512 382764 41564 382770
rect 41512 382706 41564 382712
rect 41510 382664 41566 382673
rect 41510 382599 41566 382608
rect 41524 381954 41552 382599
rect 41512 381948 41564 381954
rect 41512 381890 41564 381896
rect 41510 381848 41566 381857
rect 41510 381783 41512 381792
rect 41564 381783 41566 381792
rect 41512 381754 41564 381760
rect 41510 381440 41566 381449
rect 41510 381375 41566 381384
rect 41524 381274 41552 381375
rect 41512 381268 41564 381274
rect 41512 381210 41564 381216
rect 42338 381168 42394 381177
rect 42338 381103 42394 381112
rect 41970 380760 42026 380769
rect 41970 380695 42026 380704
rect 41510 380216 41566 380225
rect 41510 380151 41512 380160
rect 41564 380151 41566 380160
rect 41512 380122 41564 380128
rect 41510 379808 41566 379817
rect 41510 379743 41566 379752
rect 41524 379506 41552 379743
rect 41512 379500 41564 379506
rect 41512 379442 41564 379448
rect 41510 379400 41566 379409
rect 41510 379335 41566 379344
rect 41418 378992 41474 379001
rect 41418 378927 41420 378936
rect 41472 378927 41474 378936
rect 41420 378898 41472 378904
rect 41524 378554 41552 379335
rect 41602 378584 41658 378593
rect 41512 378548 41564 378554
rect 41602 378519 41658 378528
rect 41512 378490 41564 378496
rect 41616 378282 41644 378519
rect 41604 378276 41656 378282
rect 41604 378218 41656 378224
rect 41510 378176 41566 378185
rect 41510 378111 41566 378120
rect 41326 377768 41382 377777
rect 41326 377703 41382 377712
rect 41340 370598 41368 377703
rect 41418 377360 41474 377369
rect 41418 377295 41474 377304
rect 41432 376145 41460 377295
rect 41418 376136 41474 376145
rect 41418 376071 41420 376080
rect 41472 376071 41474 376080
rect 41420 376042 41472 376048
rect 41524 372026 41552 378111
rect 41512 372020 41564 372026
rect 41512 371962 41564 371968
rect 41328 370592 41380 370598
rect 41328 370534 41380 370540
rect 41984 370258 42012 380695
rect 41972 370252 42024 370258
rect 41972 370194 42024 370200
rect 42352 370002 42380 381103
rect 42444 374950 42472 385999
rect 44008 385830 44036 413782
rect 44088 413772 44140 413778
rect 44088 413714 44140 413720
rect 44100 386102 44128 413714
rect 44192 411194 44220 413850
rect 44180 411188 44232 411194
rect 44180 411130 44232 411136
rect 44284 406978 44312 413918
rect 44272 406972 44324 406978
rect 44272 406914 44324 406920
rect 44088 386096 44140 386102
rect 44088 386038 44140 386044
rect 43996 385824 44048 385830
rect 43996 385766 44048 385772
rect 44088 383784 44140 383790
rect 44088 383726 44140 383732
rect 43812 383716 43864 383722
rect 43812 383658 43864 383664
rect 43720 382764 43772 382770
rect 43720 382706 43772 382712
rect 42708 381948 42760 381954
rect 42708 381890 42760 381896
rect 42432 374944 42484 374950
rect 42432 374886 42484 374892
rect 42168 369974 42380 370002
rect 42168 369444 42196 369974
rect 42340 369912 42392 369918
rect 42340 369854 42392 369860
rect 42352 369458 42380 369854
rect 42260 369430 42380 369458
rect 42156 368144 42208 368150
rect 42156 368086 42208 368092
rect 42168 367608 42196 368086
rect 42260 367962 42288 369430
rect 42720 369374 42748 381890
rect 43076 381812 43128 381818
rect 43076 381754 43128 381760
rect 42340 369368 42392 369374
rect 42340 369310 42392 369316
rect 42708 369368 42760 369374
rect 42708 369310 42760 369316
rect 42352 368150 42380 369310
rect 42708 369232 42760 369238
rect 42708 369174 42760 369180
rect 42340 368144 42392 368150
rect 42340 368086 42392 368092
rect 42260 367934 42380 367962
rect 42168 366586 42196 366961
rect 42156 366580 42208 366586
rect 42156 366522 42208 366528
rect 42156 366308 42208 366314
rect 42156 366250 42208 366256
rect 42168 365772 42196 366250
rect 42168 364970 42196 365121
rect 42352 365090 42380 367934
rect 42720 366722 42748 369174
rect 42708 366716 42760 366722
rect 42708 366658 42760 366664
rect 42708 366580 42760 366586
rect 42708 366522 42760 366528
rect 42340 365084 42392 365090
rect 42340 365026 42392 365032
rect 42168 364942 42380 364970
rect 42248 364880 42300 364886
rect 42168 364828 42248 364834
rect 42168 364822 42300 364828
rect 42168 364806 42288 364822
rect 42168 364548 42196 364806
rect 42248 364744 42300 364750
rect 42248 364686 42300 364692
rect 42260 363950 42288 364686
rect 42182 363922 42288 363950
rect 42156 363860 42208 363866
rect 42156 363802 42208 363808
rect 42168 363256 42196 363802
rect 42156 363180 42208 363186
rect 42156 363122 42208 363128
rect 42168 362712 42196 363122
rect 42352 361350 42380 364942
rect 42432 361956 42484 361962
rect 42432 361898 42484 361904
rect 42340 361344 42392 361350
rect 42340 361286 42392 361292
rect 42340 360936 42392 360942
rect 42340 360878 42392 360884
rect 42352 360278 42380 360878
rect 42168 360210 42196 360264
rect 42260 360250 42380 360278
rect 42260 360210 42288 360250
rect 42168 360182 42288 360210
rect 42340 360188 42392 360194
rect 42340 360130 42392 360136
rect 42156 359984 42208 359990
rect 42156 359926 42208 359932
rect 42168 359584 42196 359926
rect 42352 358986 42380 360130
rect 42182 358958 42380 358986
rect 42444 358442 42472 361898
rect 42720 361554 42748 366522
rect 43088 361962 43116 381754
rect 43628 381268 43680 381274
rect 43628 381210 43680 381216
rect 43640 380894 43668 381210
rect 43548 380866 43668 380894
rect 43352 378956 43404 378962
rect 43352 378898 43404 378904
rect 43168 378548 43220 378554
rect 43168 378490 43220 378496
rect 43180 366314 43208 378490
rect 43260 372020 43312 372026
rect 43260 371962 43312 371968
rect 43168 366308 43220 366314
rect 43168 366250 43220 366256
rect 43168 366172 43220 366178
rect 43168 366114 43220 366120
rect 43180 364342 43208 366114
rect 43168 364336 43220 364342
rect 43168 364278 43220 364284
rect 43272 363866 43300 371962
rect 43364 364750 43392 378898
rect 43444 378276 43496 378282
rect 43444 378218 43496 378224
rect 43352 364744 43404 364750
rect 43352 364686 43404 364692
rect 43352 364608 43404 364614
rect 43352 364550 43404 364556
rect 43260 363860 43312 363866
rect 43260 363802 43312 363808
rect 43076 361956 43128 361962
rect 43076 361898 43128 361904
rect 42708 361548 42760 361554
rect 42708 361490 42760 361496
rect 43364 359990 43392 364550
rect 43456 361574 43484 378218
rect 43548 363186 43576 380866
rect 43628 380180 43680 380186
rect 43628 380122 43680 380128
rect 43640 371414 43668 380122
rect 43628 371408 43680 371414
rect 43628 371350 43680 371356
rect 43628 371272 43680 371278
rect 43628 371214 43680 371220
rect 43536 363180 43588 363186
rect 43536 363122 43588 363128
rect 43456 361546 43576 361574
rect 43548 360942 43576 361546
rect 43536 360936 43588 360942
rect 43536 360878 43588 360884
rect 43352 359984 43404 359990
rect 43352 359926 43404 359932
rect 42168 358306 42196 358428
rect 42260 358414 42472 358442
rect 42260 358306 42288 358414
rect 42168 358278 42288 358306
rect 42432 358352 42484 358358
rect 42432 358294 42484 358300
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42444 355926 42472 358294
rect 42182 355898 42472 355926
rect 41786 355736 41842 355745
rect 41786 355671 41842 355680
rect 41800 355300 41828 355671
rect 42168 350538 42196 354725
rect 42156 350532 42208 350538
rect 42156 350474 42208 350480
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 41880 345024 41932 345030
rect 41880 344966 41932 344972
rect 41510 344312 41566 344321
rect 41510 344247 41512 344256
rect 41564 344247 41566 344256
rect 41512 344218 41564 344224
rect 41788 344140 41840 344146
rect 41788 344082 41840 344088
rect 41510 343904 41566 343913
rect 41510 343839 41512 343848
rect 41564 343839 41566 343848
rect 41512 343810 41564 343816
rect 41510 343496 41566 343505
rect 41510 343431 41512 343440
rect 41564 343431 41566 343440
rect 41512 343402 41564 343408
rect 41510 342680 41566 342689
rect 41510 342615 41512 342624
rect 41564 342615 41566 342624
rect 41512 342586 41564 342592
rect 41800 342553 41828 344082
rect 41892 343369 41920 344966
rect 41878 343360 41934 343369
rect 41878 343295 41934 343304
rect 41786 342544 41842 342553
rect 41786 342479 41842 342488
rect 41786 342136 41842 342145
rect 41786 342071 41842 342080
rect 41512 341896 41564 341902
rect 41510 341864 41512 341873
rect 41564 341864 41566 341873
rect 41510 341799 41566 341808
rect 41512 341488 41564 341494
rect 41512 341430 41564 341436
rect 41524 341057 41552 341430
rect 41800 341426 41828 342071
rect 43640 341902 43668 371214
rect 43628 341896 43680 341902
rect 43628 341838 43680 341844
rect 43732 341494 43760 382706
rect 43824 371278 43852 383658
rect 44100 380894 44128 383726
rect 43916 380866 44128 380894
rect 43812 371272 43864 371278
rect 43812 371214 43864 371220
rect 43916 371090 43944 380866
rect 43996 379500 44048 379506
rect 43996 379442 44048 379448
rect 43824 371062 43944 371090
rect 43824 344146 43852 371062
rect 43904 371000 43956 371006
rect 43904 370942 43956 370948
rect 43916 364426 43944 370942
rect 44008 364614 44036 379442
rect 44088 374944 44140 374950
rect 44088 374886 44140 374892
rect 43996 364608 44048 364614
rect 43996 364550 44048 364556
rect 43916 364398 44036 364426
rect 43904 364336 43956 364342
rect 43904 364278 43956 364284
rect 43916 358358 43944 364278
rect 44008 360194 44036 364398
rect 43996 360188 44048 360194
rect 43996 360130 44048 360136
rect 43904 358352 43956 358358
rect 43904 358294 43956 358300
rect 44100 345030 44128 374886
rect 44088 345024 44140 345030
rect 44088 344966 44140 344972
rect 43812 344140 43864 344146
rect 43812 344082 43864 344088
rect 43904 342644 43956 342650
rect 43904 342586 43956 342592
rect 43720 341488 43772 341494
rect 43720 341430 43772 341436
rect 41788 341420 41840 341426
rect 41788 341362 41840 341368
rect 43536 341420 43588 341426
rect 43536 341362 43588 341368
rect 41786 341320 41842 341329
rect 41786 341255 41842 341264
rect 41510 341048 41566 341057
rect 41510 340983 41566 340992
rect 29918 339824 29974 339833
rect 29918 339759 29974 339768
rect 33046 339824 33102 339833
rect 33046 339759 33102 339768
rect 29932 330041 29960 339759
rect 30102 339008 30158 339017
rect 30102 338943 30158 338952
rect 30010 338600 30066 338609
rect 30010 338535 30066 338544
rect 29918 330032 29974 330041
rect 29918 329967 29974 329976
rect 30024 329905 30052 338535
rect 30116 330177 30144 338943
rect 30194 338192 30250 338201
rect 30194 338127 30250 338136
rect 30102 330168 30158 330177
rect 30102 330103 30158 330112
rect 30208 330070 30236 338127
rect 30286 337784 30342 337793
rect 30286 337719 30342 337728
rect 30300 330342 30328 337719
rect 30288 330336 30340 330342
rect 30288 330278 30340 330284
rect 33060 330274 33088 339759
rect 41800 339522 41828 341255
rect 41788 339516 41840 339522
rect 41788 339458 41840 339464
rect 43352 339516 43404 339522
rect 43352 339458 43404 339464
rect 41510 336152 41566 336161
rect 41510 336087 41566 336096
rect 41418 334928 41474 334937
rect 41418 334863 41474 334872
rect 41432 331158 41460 334863
rect 41524 331226 41552 336087
rect 41786 336016 41842 336025
rect 41786 335951 41842 335960
rect 41602 335336 41658 335345
rect 41602 335271 41658 335280
rect 41512 331220 41564 331226
rect 41512 331162 41564 331168
rect 41420 331152 41472 331158
rect 41420 331094 41472 331100
rect 33048 330268 33100 330274
rect 33048 330210 33100 330216
rect 30196 330064 30248 330070
rect 30196 330006 30248 330012
rect 30010 329896 30066 329905
rect 30010 329831 30066 329840
rect 41616 329390 41644 335271
rect 41694 334520 41750 334529
rect 41694 334455 41750 334464
rect 41708 330954 41736 334455
rect 41696 330948 41748 330954
rect 41696 330890 41748 330896
rect 41800 329458 41828 335951
rect 41878 334384 41934 334393
rect 41878 334319 41934 334328
rect 41892 333169 41920 334319
rect 41878 333160 41934 333169
rect 41878 333095 41880 333104
rect 41932 333095 41934 333104
rect 41880 333066 41932 333072
rect 42708 331220 42760 331226
rect 42708 331162 42760 331168
rect 42248 330336 42300 330342
rect 42248 330278 42300 330284
rect 41788 329452 41840 329458
rect 41788 329394 41840 329400
rect 41604 329384 41656 329390
rect 41604 329326 41656 329332
rect 42168 326210 42196 326264
rect 42260 326210 42288 330278
rect 42340 330268 42392 330274
rect 42340 330210 42392 330216
rect 42168 326182 42288 326210
rect 42352 324442 42380 330210
rect 42168 324306 42196 324428
rect 42260 324414 42380 324442
rect 42260 324306 42288 324414
rect 42168 324278 42288 324306
rect 42182 323734 42288 323762
rect 42064 323128 42116 323134
rect 42064 323070 42116 323076
rect 42076 322592 42104 323070
rect 42260 322046 42288 323734
rect 42720 323134 42748 331162
rect 43168 331152 43220 331158
rect 43168 331094 43220 331100
rect 43076 329384 43128 329390
rect 43076 329326 43128 329332
rect 43088 323202 43116 329326
rect 43076 323196 43128 323202
rect 43076 323138 43128 323144
rect 42708 323128 42760 323134
rect 43180 323082 43208 331094
rect 43260 329452 43312 329458
rect 43260 329394 43312 329400
rect 42708 323070 42760 323076
rect 43088 323054 43208 323082
rect 42708 322992 42760 322998
rect 42708 322934 42760 322940
rect 42248 322040 42300 322046
rect 42248 321982 42300 321988
rect 42182 321898 42380 321926
rect 42248 321836 42300 321842
rect 42248 321778 42300 321784
rect 42156 321632 42208 321638
rect 42156 321574 42208 321580
rect 42168 321368 42196 321574
rect 42260 320739 42288 321778
rect 42182 320711 42288 320739
rect 42248 320612 42300 320618
rect 42248 320554 42300 320560
rect 42260 320090 42288 320554
rect 42182 320062 42288 320090
rect 42248 320000 42300 320006
rect 42248 319942 42300 319948
rect 42260 319546 42288 319942
rect 42182 319518 42288 319546
rect 42352 317422 42380 321898
rect 42720 318782 42748 322934
rect 43088 320618 43116 323054
rect 43272 322946 43300 329394
rect 43180 322918 43300 322946
rect 43180 321842 43208 322918
rect 43260 322040 43312 322046
rect 43260 321982 43312 321988
rect 43168 321836 43220 321842
rect 43168 321778 43220 321784
rect 43076 320612 43128 320618
rect 43076 320554 43128 320560
rect 43272 318782 43300 321982
rect 42432 318776 42484 318782
rect 42432 318718 42484 318724
rect 42708 318776 42760 318782
rect 42708 318718 42760 318724
rect 43260 318776 43312 318782
rect 43260 318718 43312 318724
rect 42340 317416 42392 317422
rect 42340 317358 42392 317364
rect 42444 317059 42472 318718
rect 42182 317031 42472 317059
rect 42430 316432 42486 316441
rect 42182 316390 42430 316418
rect 42430 316367 42486 316376
rect 41786 316296 41842 316305
rect 41786 316231 41842 316240
rect 41800 315757 41828 316231
rect 42154 315480 42210 315489
rect 42154 315415 42210 315424
rect 42168 315180 42196 315415
rect 41970 313848 42026 313857
rect 41970 313783 42026 313792
rect 41984 313344 42012 313783
rect 41786 313032 41842 313041
rect 41786 312967 41842 312976
rect 41800 312732 41828 312967
rect 42154 312352 42210 312361
rect 42154 312287 42210 312296
rect 42168 312052 42196 312287
rect 42076 306338 42104 311508
rect 42064 306332 42116 306338
rect 42064 306274 42116 306280
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41970 301336 42026 301345
rect 41970 301271 42026 301280
rect 27526 300928 27582 300937
rect 27526 300863 27582 300872
rect 27540 289814 27568 300863
rect 41878 300520 41934 300529
rect 41878 300455 41934 300464
rect 41788 300144 41840 300150
rect 41786 300112 41788 300121
rect 41840 300112 41842 300121
rect 41786 300047 41842 300056
rect 41788 300008 41840 300014
rect 41788 299950 41840 299956
rect 41800 299305 41828 299950
rect 41786 299296 41842 299305
rect 41786 299231 41842 299240
rect 41788 299124 41840 299130
rect 41788 299066 41840 299072
rect 41800 298489 41828 299066
rect 41786 298480 41842 298489
rect 41786 298415 41842 298424
rect 41786 298072 41842 298081
rect 41786 298007 41842 298016
rect 41800 297362 41828 298007
rect 41788 297356 41840 297362
rect 41788 297298 41840 297304
rect 41786 297256 41842 297265
rect 41786 297191 41842 297200
rect 35806 296440 35862 296449
rect 35806 296375 35862 296384
rect 27528 289808 27580 289814
rect 27528 289750 27580 289756
rect 35820 287026 35848 296375
rect 41800 296274 41828 297191
rect 41788 296268 41840 296274
rect 41788 296210 41840 296216
rect 41694 295080 41750 295089
rect 41694 295015 41750 295024
rect 35808 287020 35860 287026
rect 35808 286962 35860 286968
rect 41708 285802 41736 295015
rect 41786 294808 41842 294817
rect 41786 294743 41842 294752
rect 41800 292074 41828 294743
rect 41892 292466 41920 300455
rect 41984 292534 42012 301271
rect 42062 299704 42118 299713
rect 42062 299639 42118 299648
rect 42076 299402 42104 299639
rect 42064 299396 42116 299402
rect 42064 299338 42116 299344
rect 43260 299396 43312 299402
rect 43260 299338 43312 299344
rect 42430 298888 42486 298897
rect 42430 298823 42486 298832
rect 42340 295384 42392 295390
rect 42340 295326 42392 295332
rect 42062 293992 42118 294001
rect 42062 293927 42118 293936
rect 42076 293690 42104 293927
rect 42064 293684 42116 293690
rect 42064 293626 42116 293632
rect 42062 293584 42118 293593
rect 42062 293519 42118 293528
rect 42076 293486 42104 293519
rect 42064 293480 42116 293486
rect 42064 293422 42116 293428
rect 42062 293176 42118 293185
rect 42062 293111 42118 293120
rect 41972 292528 42024 292534
rect 41972 292470 42024 292476
rect 41880 292460 41932 292466
rect 41880 292402 41932 292408
rect 41878 292360 41934 292369
rect 41878 292295 41880 292304
rect 41932 292295 41934 292304
rect 41880 292266 41932 292272
rect 41800 292046 41920 292074
rect 41786 291136 41842 291145
rect 41786 291071 41788 291080
rect 41840 291071 41842 291080
rect 41788 291042 41840 291048
rect 41786 290728 41842 290737
rect 41786 290663 41788 290672
rect 41840 290663 41842 290672
rect 41788 290634 41840 290640
rect 41786 289912 41842 289921
rect 41786 289847 41788 289856
rect 41840 289847 41842 289856
rect 41788 289818 41840 289824
rect 41696 285796 41748 285802
rect 41696 285738 41748 285744
rect 41892 283830 41920 292046
rect 41970 291952 42026 291961
rect 41970 291887 42026 291896
rect 41984 286890 42012 291887
rect 41972 286884 42024 286890
rect 41972 286826 42024 286832
rect 42076 286210 42104 293111
rect 42154 292768 42210 292777
rect 42154 292703 42210 292712
rect 42168 286958 42196 292703
rect 42248 287020 42300 287026
rect 42248 286962 42300 286968
rect 42156 286952 42208 286958
rect 42156 286894 42208 286900
rect 42064 286204 42116 286210
rect 42064 286146 42116 286152
rect 41880 283824 41932 283830
rect 41880 283766 41932 283772
rect 41880 283620 41932 283626
rect 41880 283562 41932 283568
rect 41892 283045 41920 283562
rect 42260 281738 42288 286962
rect 42168 281710 42288 281738
rect 42168 281180 42196 281710
rect 42352 280582 42380 295326
rect 42444 285666 42472 298823
rect 43076 292324 43128 292330
rect 43076 292266 43128 292272
rect 42706 291544 42762 291553
rect 42706 291479 42762 291488
rect 42432 285660 42484 285666
rect 42432 285602 42484 285608
rect 42182 280554 42380 280582
rect 42340 280492 42392 280498
rect 42340 280434 42392 280440
rect 42248 280424 42300 280430
rect 42248 280366 42300 280372
rect 42156 279880 42208 279886
rect 42156 279822 42208 279828
rect 42168 279344 42196 279822
rect 42260 278746 42288 280366
rect 42182 278718 42288 278746
rect 42064 278452 42116 278458
rect 42064 278394 42116 278400
rect 42076 278188 42104 278394
rect 42156 277908 42208 277914
rect 42156 277850 42208 277856
rect 42168 277508 42196 277850
rect 42352 276910 42380 280434
rect 42720 278458 42748 291479
rect 43088 284170 43116 292266
rect 43168 286204 43220 286210
rect 43168 286146 43220 286152
rect 43076 284164 43128 284170
rect 43076 284106 43128 284112
rect 43076 281648 43128 281654
rect 43076 281590 43128 281596
rect 42708 278452 42760 278458
rect 42708 278394 42760 278400
rect 42182 276882 42380 276910
rect 42340 276820 42392 276826
rect 42340 276762 42392 276768
rect 42352 276366 42380 276762
rect 42168 276298 42196 276352
rect 42260 276338 42380 276366
rect 42260 276298 42288 276338
rect 42168 276270 42288 276298
rect 42432 275596 42484 275602
rect 42432 275538 42484 275544
rect 42444 273850 42472 275538
rect 42182 273822 42472 273850
rect 42432 273760 42484 273766
rect 42432 273702 42484 273708
rect 42444 273238 42472 273702
rect 42168 273170 42196 273224
rect 42260 273210 42472 273238
rect 42260 273170 42288 273210
rect 42168 273142 42288 273170
rect 43088 273154 43116 281590
rect 43180 279886 43208 286146
rect 43168 279880 43220 279886
rect 43168 279822 43220 279828
rect 42432 273148 42484 273154
rect 42432 273090 42484 273096
rect 43076 273148 43128 273154
rect 43076 273090 43128 273096
rect 42444 272558 42472 273090
rect 42182 272530 42472 272558
rect 41786 272368 41842 272377
rect 41786 272303 41842 272312
rect 41800 272000 41828 272303
rect 42432 271856 42484 271862
rect 42432 271798 42484 271804
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 41970 269784 42026 269793
rect 41970 269719 42026 269728
rect 41984 269521 42012 269719
rect 41786 269376 41842 269385
rect 41786 269311 41842 269320
rect 41800 268872 41828 269311
rect 42444 268342 42472 271798
rect 42182 268314 42472 268342
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 43272 258874 43300 299338
rect 43364 299130 43392 339458
rect 43444 330948 43496 330954
rect 43444 330890 43496 330896
rect 43456 321638 43484 330890
rect 43444 321632 43496 321638
rect 43444 321574 43496 321580
rect 43548 300014 43576 341362
rect 43628 330064 43680 330070
rect 43628 330006 43680 330012
rect 43640 320006 43668 330006
rect 43628 320000 43680 320006
rect 43628 319942 43680 319948
rect 43916 300150 43944 342586
rect 43904 300144 43956 300150
rect 43904 300086 43956 300092
rect 43536 300008 43588 300014
rect 43536 299950 43588 299956
rect 43352 299124 43404 299130
rect 43352 299066 43404 299072
rect 43628 297356 43680 297362
rect 43628 297298 43680 297304
rect 43536 292664 43588 292670
rect 43536 292606 43588 292612
rect 43444 286952 43496 286958
rect 43444 286894 43496 286900
rect 43352 286884 43404 286890
rect 43352 286826 43404 286832
rect 43364 280498 43392 286826
rect 43352 280492 43404 280498
rect 43352 280434 43404 280440
rect 43456 277914 43484 286894
rect 43548 280430 43576 292606
rect 43536 280424 43588 280430
rect 43536 280366 43588 280372
rect 43444 277908 43496 277914
rect 43444 277850 43496 277856
rect 41788 258868 41840 258874
rect 41788 258810 41840 258816
rect 43260 258868 43312 258874
rect 43260 258810 43312 258816
rect 41510 257952 41566 257961
rect 41510 257887 41566 257896
rect 41524 256766 41552 257887
rect 41604 257576 41656 257582
rect 41602 257544 41604 257553
rect 41656 257544 41658 257553
rect 41602 257479 41658 257488
rect 41800 256873 41828 258810
rect 41880 257712 41932 257718
rect 41878 257680 41880 257689
rect 41932 257680 41934 257689
rect 41878 257615 41934 257624
rect 41786 256864 41842 256873
rect 41786 256799 41842 256808
rect 41512 256760 41564 256766
rect 41512 256702 41564 256708
rect 41878 256456 41934 256465
rect 41878 256391 41934 256400
rect 41512 256352 41564 256358
rect 41510 256320 41512 256329
rect 41564 256320 41566 256329
rect 41510 256255 41566 256264
rect 41512 255740 41564 255746
rect 41512 255682 41564 255688
rect 41524 255513 41552 255682
rect 41510 255504 41566 255513
rect 41510 255439 41566 255448
rect 41512 254924 41564 254930
rect 41512 254866 41564 254872
rect 41524 254697 41552 254866
rect 41786 254824 41842 254833
rect 41786 254759 41842 254768
rect 41510 254688 41566 254697
rect 41510 254623 41566 254632
rect 41800 253978 41828 254759
rect 41892 254182 41920 256391
rect 43640 255746 43668 297298
rect 43812 296268 43864 296274
rect 43812 296210 43864 296216
rect 43824 295334 43852 296210
rect 43824 295306 43944 295334
rect 43812 285796 43864 285802
rect 43812 285738 43864 285744
rect 43720 285660 43772 285666
rect 43720 285602 43772 285608
rect 43732 256358 43760 285602
rect 43824 276826 43852 285738
rect 43812 276820 43864 276826
rect 43812 276762 43864 276768
rect 43720 256352 43772 256358
rect 43720 256294 43772 256300
rect 43628 255740 43680 255746
rect 43628 255682 43680 255688
rect 43916 254930 43944 295306
rect 43996 293684 44048 293690
rect 43996 293626 44048 293632
rect 44008 284306 44036 293626
rect 44088 293480 44140 293486
rect 44088 293422 44140 293428
rect 44100 284458 44128 293422
rect 44100 284430 44220 284458
rect 43996 284300 44048 284306
rect 43996 284242 44048 284248
rect 44192 284186 44220 284430
rect 44272 284300 44324 284306
rect 44272 284242 44324 284248
rect 43996 284164 44048 284170
rect 43996 284106 44048 284112
rect 44100 284158 44220 284186
rect 44008 275602 44036 284106
rect 43996 275596 44048 275602
rect 43996 275538 44048 275544
rect 44100 273766 44128 284158
rect 44284 281654 44312 284242
rect 44272 281648 44324 281654
rect 44272 281590 44324 281596
rect 44088 273760 44140 273766
rect 44088 273702 44140 273708
rect 43904 254924 43956 254930
rect 43904 254866 43956 254872
rect 41880 254176 41932 254182
rect 41880 254118 41932 254124
rect 43904 254176 43956 254182
rect 43904 254118 43956 254124
rect 41880 254040 41932 254046
rect 41878 254008 41880 254017
rect 43628 254040 43680 254046
rect 41932 254008 41934 254017
rect 41788 253972 41840 253978
rect 43628 253982 43680 253988
rect 41878 253943 41934 253952
rect 43168 253972 43220 253978
rect 41788 253914 41840 253920
rect 43168 253914 43220 253920
rect 42062 253600 42118 253609
rect 42062 253535 42118 253544
rect 41694 253056 41750 253065
rect 41694 252991 41750 253000
rect 41142 251424 41198 251433
rect 41142 251359 41198 251368
rect 35806 251016 35862 251025
rect 35806 250951 35862 250960
rect 35820 242486 35848 250951
rect 38474 250608 38530 250617
rect 38474 250543 38530 250552
rect 38488 242554 38516 250543
rect 38566 250200 38622 250209
rect 38566 250135 38622 250144
rect 38580 242622 38608 250135
rect 38568 242616 38620 242622
rect 38568 242558 38620 242564
rect 38476 242548 38528 242554
rect 38476 242490 38528 242496
rect 35808 242480 35860 242486
rect 35808 242422 35860 242428
rect 41156 240990 41184 251359
rect 41234 249792 41290 249801
rect 41234 249727 41290 249736
rect 41248 242758 41276 249727
rect 41602 248976 41658 248985
rect 41602 248911 41658 248920
rect 41418 248568 41474 248577
rect 41418 248503 41474 248512
rect 41326 248160 41382 248169
rect 41326 248095 41382 248104
rect 41340 242894 41368 248095
rect 41328 242888 41380 242894
rect 41328 242830 41380 242836
rect 41432 242826 41460 248503
rect 41510 247752 41566 247761
rect 41510 247687 41512 247696
rect 41564 247687 41566 247696
rect 41512 247658 41564 247664
rect 41510 247344 41566 247353
rect 41510 247279 41512 247288
rect 41564 247279 41566 247288
rect 41512 247250 41564 247256
rect 41510 246528 41566 246537
rect 41510 246463 41512 246472
rect 41564 246463 41566 246472
rect 41512 246434 41564 246440
rect 41420 242820 41472 242826
rect 41420 242762 41472 242768
rect 41236 242752 41288 242758
rect 41236 242694 41288 242700
rect 41616 242690 41644 248911
rect 41708 245614 41736 252991
rect 41878 252784 41934 252793
rect 41878 252719 41934 252728
rect 41786 251968 41842 251977
rect 41786 251903 41842 251912
rect 41696 245608 41748 245614
rect 41696 245550 41748 245556
rect 41800 244662 41828 251903
rect 41892 245138 41920 252719
rect 41970 252376 42026 252385
rect 41970 252311 42026 252320
rect 41880 245132 41932 245138
rect 41880 245074 41932 245080
rect 41788 244656 41840 244662
rect 41788 244598 41840 244604
rect 41604 242684 41656 242690
rect 41604 242626 41656 242632
rect 41984 242321 42012 252311
rect 41970 242312 42026 242321
rect 41970 242247 42026 242256
rect 42076 242185 42104 253535
rect 42338 249520 42394 249529
rect 42338 249455 42394 249464
rect 42248 242752 42300 242758
rect 42248 242694 42300 242700
rect 42062 242176 42118 242185
rect 42062 242111 42118 242120
rect 41144 240984 41196 240990
rect 41144 240926 41196 240932
rect 41788 240372 41840 240378
rect 41788 240314 41840 240320
rect 41800 239836 41828 240314
rect 42156 238536 42208 238542
rect 42156 238478 42208 238484
rect 42168 238000 42196 238478
rect 42260 236178 42288 242694
rect 42182 236150 42288 236178
rect 42248 236088 42300 236094
rect 42248 236030 42300 236036
rect 42260 234983 42288 236030
rect 42182 234955 42288 234983
rect 42352 234342 42380 249455
rect 42708 245608 42760 245614
rect 42708 245550 42760 245556
rect 42720 238542 42748 245550
rect 43076 242820 43128 242826
rect 43076 242762 43128 242768
rect 42708 238536 42760 238542
rect 42708 238478 42760 238484
rect 42182 234314 42380 234342
rect 43088 234258 43116 242762
rect 42340 234252 42392 234258
rect 42340 234194 42392 234200
rect 43076 234252 43128 234258
rect 43076 234194 43128 234200
rect 42352 233695 42380 234194
rect 42182 233667 42380 233695
rect 42156 233368 42208 233374
rect 42156 233310 42208 233316
rect 42168 233104 42196 233310
rect 42432 232348 42484 232354
rect 42432 232290 42484 232296
rect 42444 230670 42472 232290
rect 42182 230642 42472 230670
rect 42432 230580 42484 230586
rect 42432 230522 42484 230528
rect 42156 230376 42208 230382
rect 42156 230318 42208 230324
rect 42168 229976 42196 230318
rect 42444 229378 42472 230522
rect 42182 229350 42472 229378
rect 42430 228848 42486 228857
rect 42182 228806 42430 228834
rect 42430 228783 42486 228792
rect 42430 228712 42486 228721
rect 42430 228647 42486 228656
rect 42444 226998 42472 228647
rect 42168 226930 42196 226984
rect 42260 226970 42472 226998
rect 42260 226930 42288 226970
rect 42168 226902 42288 226930
rect 42156 226704 42208 226710
rect 42156 226646 42208 226652
rect 42168 226304 42196 226646
rect 42430 225720 42486 225729
rect 42182 225678 42430 225706
rect 42430 225655 42486 225664
rect 42432 225616 42484 225622
rect 42432 225558 42484 225564
rect 42444 225162 42472 225558
rect 42168 225026 42196 225148
rect 42260 225134 42472 225162
rect 42260 225026 42288 225134
rect 42168 224998 42288 225026
rect 24952 217524 25004 217530
rect 24952 217466 25004 217472
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 24860 215416 24912 215422
rect 24860 215358 24912 215364
rect 24872 203697 24900 215358
rect 24964 204513 24992 217466
rect 25136 215484 25188 215490
rect 25136 215426 25188 215432
rect 25148 204921 25176 215426
rect 41512 215144 41564 215150
rect 41510 215112 41512 215121
rect 41564 215112 41566 215121
rect 41510 215047 41566 215056
rect 41512 214736 41564 214742
rect 41510 214704 41512 214713
rect 41564 214704 41566 214713
rect 41510 214639 41566 214648
rect 41512 214328 41564 214334
rect 41510 214296 41512 214305
rect 41564 214296 41566 214305
rect 41510 214231 41566 214240
rect 41512 214124 41564 214130
rect 41512 214066 41564 214072
rect 41524 213897 41552 214066
rect 41510 213888 41566 213897
rect 41510 213823 41566 213832
rect 33048 213648 33100 213654
rect 33048 213590 33100 213596
rect 32956 213580 33008 213586
rect 32956 213522 33008 213528
rect 32864 213512 32916 213518
rect 32864 213454 32916 213460
rect 32876 211041 32904 213454
rect 32968 211857 32996 213522
rect 33060 212673 33088 213590
rect 41510 213480 41566 213489
rect 41510 213415 41512 213424
rect 41564 213415 41566 213424
rect 41512 213386 41564 213392
rect 33046 212664 33102 212673
rect 33046 212599 33102 212608
rect 43180 212294 43208 253914
rect 43536 245132 43588 245138
rect 43536 245074 43588 245080
rect 43352 244656 43404 244662
rect 43352 244598 43404 244604
rect 43260 242888 43312 242894
rect 43260 242830 43312 242836
rect 43272 236094 43300 242830
rect 43260 236088 43312 236094
rect 43260 236030 43312 236036
rect 43364 233374 43392 244598
rect 43444 242684 43496 242690
rect 43444 242626 43496 242632
rect 43352 233368 43404 233374
rect 43352 233310 43404 233316
rect 43456 232354 43484 242626
rect 43548 238105 43576 245074
rect 43534 238096 43590 238105
rect 43534 238031 43590 238040
rect 43536 237992 43588 237998
rect 43536 237934 43588 237940
rect 43444 232348 43496 232354
rect 43444 232290 43496 232296
rect 43548 214130 43576 237934
rect 43536 214124 43588 214130
rect 43536 214066 43588 214072
rect 41512 212288 41564 212294
rect 41510 212256 41512 212265
rect 43168 212288 43220 212294
rect 41564 212256 41566 212265
rect 43168 212230 43220 212236
rect 41510 212191 41566 212200
rect 43640 212158 43668 253982
rect 43720 242616 43772 242622
rect 43720 242558 43772 242564
rect 43732 230382 43760 242558
rect 43812 242548 43864 242554
rect 43812 242490 43864 242496
rect 43824 230586 43852 242490
rect 43916 237998 43944 254118
rect 43996 242480 44048 242486
rect 43996 242422 44048 242428
rect 43904 237992 43956 237998
rect 43904 237934 43956 237940
rect 43812 230580 43864 230586
rect 43812 230522 43864 230528
rect 43720 230376 43772 230382
rect 43720 230318 43772 230324
rect 44008 226710 44036 242422
rect 43996 226704 44048 226710
rect 43996 226646 44048 226652
rect 45480 219706 45508 805938
rect 45572 789274 45600 816818
rect 45560 789268 45612 789274
rect 45560 789210 45612 789216
rect 48240 786622 48268 817226
rect 48228 786616 48280 786622
rect 48228 786558 48280 786564
rect 51000 786554 51028 817634
rect 58256 800488 58308 800494
rect 58256 800430 58308 800436
rect 58268 790945 58296 800430
rect 655520 792192 655572 792198
rect 655520 792134 655572 792140
rect 58254 790936 58310 790945
rect 58254 790871 58310 790880
rect 58164 789404 58216 789410
rect 58164 789346 58216 789352
rect 58176 788497 58204 789346
rect 58532 789336 58584 789342
rect 58530 789304 58532 789313
rect 58584 789304 58586 789313
rect 58440 789268 58492 789274
rect 58530 789239 58586 789248
rect 58440 789210 58492 789216
rect 58162 788488 58218 788497
rect 58162 788423 58218 788432
rect 58452 787409 58480 789210
rect 58438 787400 58494 787409
rect 58438 787335 58494 787344
rect 58440 786616 58492 786622
rect 58440 786558 58492 786564
rect 50988 786548 51040 786554
rect 50988 786490 51040 786496
rect 58452 784961 58480 786558
rect 58532 786548 58584 786554
rect 58532 786490 58584 786496
rect 58544 786185 58572 786490
rect 58530 786176 58586 786185
rect 58530 786111 58586 786120
rect 58438 784952 58494 784961
rect 58438 784887 58494 784896
rect 655426 778424 655482 778433
rect 655426 778359 655482 778368
rect 654968 775532 655020 775538
rect 654968 775474 655020 775480
rect 50988 774444 51040 774450
rect 50988 774386 51040 774392
rect 48228 773900 48280 773906
rect 48228 773842 48280 773848
rect 45744 773628 45796 773634
rect 45744 773570 45796 773576
rect 45652 767372 45704 767378
rect 45652 767314 45704 767320
rect 45560 762884 45612 762890
rect 45560 762826 45612 762832
rect 45468 219700 45520 219706
rect 45468 219642 45520 219648
rect 45572 219638 45600 762826
rect 45664 277370 45692 767314
rect 45756 745210 45784 773570
rect 45744 745204 45796 745210
rect 45744 745146 45796 745152
rect 48240 742422 48268 773842
rect 48228 742416 48280 742422
rect 48228 742358 48280 742364
rect 51000 742354 51028 774386
rect 654980 773537 655008 775474
rect 654966 773528 655022 773537
rect 654966 773463 655022 773472
rect 59268 756288 59320 756294
rect 59268 756230 59320 756236
rect 58440 747924 58492 747930
rect 58440 747866 58492 747872
rect 58452 747697 58480 747866
rect 58438 747688 58494 747697
rect 58438 747623 58494 747632
rect 59280 746473 59308 756230
rect 59266 746464 59322 746473
rect 59266 746399 59322 746408
rect 58440 745272 58492 745278
rect 58440 745214 58492 745220
rect 58452 744977 58480 745214
rect 58532 745204 58584 745210
rect 58532 745146 58584 745152
rect 58438 744968 58494 744977
rect 58438 744903 58494 744912
rect 58544 744161 58572 745146
rect 58530 744152 58586 744161
rect 58530 744087 58586 744096
rect 58440 742416 58492 742422
rect 57978 742384 58034 742393
rect 50988 742348 51040 742354
rect 58440 742358 58492 742364
rect 57978 742319 57980 742328
rect 50988 742290 51040 742296
rect 58032 742319 58034 742328
rect 57980 742290 58032 742296
rect 58452 741849 58480 742358
rect 58438 741840 58494 741849
rect 58438 741775 58494 741784
rect 654324 737044 654376 737050
rect 654324 736986 654376 736992
rect 50988 731060 51040 731066
rect 50988 731002 51040 731008
rect 48228 730652 48280 730658
rect 48228 730594 48280 730600
rect 45836 730244 45888 730250
rect 45836 730186 45888 730192
rect 45744 719636 45796 719642
rect 45744 719578 45796 719584
rect 45652 277364 45704 277370
rect 45652 277306 45704 277312
rect 45652 247308 45704 247314
rect 45652 247250 45704 247256
rect 45560 219632 45612 219638
rect 45560 219574 45612 219580
rect 45664 216646 45692 247250
rect 45756 219570 45784 719578
rect 45848 701010 45876 730186
rect 45836 701004 45888 701010
rect 45836 700946 45888 700952
rect 48240 698290 48268 730594
rect 51000 700942 51028 731002
rect 654336 730289 654364 736986
rect 654322 730280 654378 730289
rect 654322 730215 654378 730224
rect 655440 715018 655468 778359
rect 655532 775577 655560 792134
rect 656532 783896 656584 783902
rect 656532 783838 656584 783844
rect 655794 777064 655850 777073
rect 655794 776999 655850 777008
rect 655610 775976 655666 775985
rect 655610 775911 655666 775920
rect 655518 775568 655574 775577
rect 655518 775503 655574 775512
rect 655518 734360 655574 734369
rect 655518 734295 655574 734304
rect 655428 715012 655480 715018
rect 655428 714954 655480 714960
rect 59360 714876 59412 714882
rect 59360 714818 59412 714824
rect 59268 712156 59320 712162
rect 59268 712098 59320 712104
rect 58532 703860 58584 703866
rect 58532 703802 58584 703808
rect 58544 702137 58572 703802
rect 59280 703361 59308 712098
rect 59372 704449 59400 714818
rect 59358 704440 59414 704449
rect 59358 704375 59414 704384
rect 59266 703352 59322 703361
rect 59266 703287 59322 703296
rect 58530 702128 58586 702137
rect 58530 702063 58586 702072
rect 58256 701004 58308 701010
rect 58256 700946 58308 700952
rect 50988 700936 51040 700942
rect 50988 700878 51040 700884
rect 58268 700777 58296 700946
rect 58532 700936 58584 700942
rect 58532 700878 58584 700884
rect 58254 700768 58310 700777
rect 58254 700703 58310 700712
rect 58544 699689 58572 700878
rect 58530 699680 58586 699689
rect 58530 699615 58586 699624
rect 48228 698284 48280 698290
rect 48228 698226 48280 698232
rect 58532 698284 58584 698290
rect 58532 698226 58584 698232
rect 58544 698193 58572 698226
rect 58530 698184 58586 698193
rect 58530 698119 58586 698128
rect 654232 692912 654284 692918
rect 654232 692854 654284 692860
rect 654140 690056 654192 690062
rect 654140 689998 654192 690004
rect 50988 688084 51040 688090
rect 50988 688026 51040 688032
rect 48228 687676 48280 687682
rect 48228 687618 48280 687624
rect 45928 687336 45980 687342
rect 45928 687278 45980 687284
rect 45836 676524 45888 676530
rect 45836 676466 45888 676472
rect 45744 219564 45796 219570
rect 45744 219506 45796 219512
rect 45848 219502 45876 676466
rect 45940 659598 45968 687278
rect 45928 659592 45980 659598
rect 45928 659534 45980 659540
rect 48240 656878 48268 687618
rect 48228 656872 48280 656878
rect 48228 656814 48280 656820
rect 51000 656810 51028 688026
rect 654152 684457 654180 689998
rect 654244 685817 654272 692854
rect 655426 687304 655482 687313
rect 655426 687239 655482 687248
rect 654230 685808 654286 685817
rect 654230 685743 654286 685752
rect 654138 684448 654194 684457
rect 654138 684383 654194 684392
rect 60648 670880 60700 670886
rect 60648 670822 60700 670828
rect 60660 661201 60688 670822
rect 60646 661192 60702 661201
rect 60646 661127 60702 661136
rect 58440 659728 58492 659734
rect 58440 659670 58492 659676
rect 58452 658889 58480 659670
rect 58532 659660 58584 659666
rect 58532 659602 58584 659608
rect 58544 659569 58572 659602
rect 58624 659592 58676 659598
rect 58530 659560 58586 659569
rect 58624 659534 58676 659540
rect 58530 659495 58586 659504
rect 58438 658880 58494 658889
rect 58438 658815 58494 658824
rect 58636 657665 58664 659534
rect 58622 657656 58678 657665
rect 58622 657591 58678 657600
rect 58072 656872 58124 656878
rect 58072 656814 58124 656820
rect 50988 656804 51040 656810
rect 50988 656746 51040 656752
rect 58084 655353 58112 656814
rect 58440 656804 58492 656810
rect 58440 656746 58492 656752
rect 58452 656577 58480 656746
rect 58438 656568 58494 656577
rect 58438 656503 58494 656512
rect 58070 655344 58126 655353
rect 58070 655279 58126 655288
rect 654416 648644 654468 648650
rect 654416 648586 654468 648592
rect 50988 644700 51040 644706
rect 50988 644642 51040 644648
rect 48228 644292 48280 644298
rect 48228 644234 48280 644240
rect 46020 644088 46072 644094
rect 46020 644030 46072 644036
rect 45928 633276 45980 633282
rect 45928 633218 45980 633224
rect 45836 219496 45888 219502
rect 45836 219438 45888 219444
rect 45940 219434 45968 633218
rect 46032 615466 46060 644030
rect 46020 615460 46072 615466
rect 46020 615402 46072 615408
rect 48240 612746 48268 644234
rect 48228 612740 48280 612746
rect 48228 612682 48280 612688
rect 51000 612678 51028 644642
rect 654428 639441 654456 648586
rect 654414 639432 654470 639441
rect 654414 639367 654470 639376
rect 58532 626612 58584 626618
rect 58532 626554 58584 626560
rect 58164 618248 58216 618254
rect 58164 618190 58216 618196
rect 58176 617817 58204 618190
rect 58162 617808 58218 617817
rect 58162 617743 58218 617752
rect 58544 616865 58572 626554
rect 655440 623898 655468 687239
rect 655532 670818 655560 734295
rect 655624 715154 655652 775911
rect 655702 731504 655758 731513
rect 655702 731439 655758 731448
rect 655612 715148 655664 715154
rect 655612 715090 655664 715096
rect 655610 688256 655666 688265
rect 655610 688191 655666 688200
rect 655520 670812 655572 670818
rect 655520 670754 655572 670760
rect 655518 643240 655574 643249
rect 655518 643175 655574 643184
rect 655428 623892 655480 623898
rect 655428 623834 655480 623840
rect 58530 616856 58586 616865
rect 58530 616791 58586 616800
rect 58532 615528 58584 615534
rect 58530 615496 58532 615505
rect 58584 615496 58586 615505
rect 58164 615460 58216 615466
rect 58530 615431 58586 615440
rect 58164 615402 58216 615408
rect 58176 614553 58204 615402
rect 58162 614544 58218 614553
rect 58162 614479 58218 614488
rect 655428 612876 655480 612882
rect 655428 612818 655480 612824
rect 58348 612740 58400 612746
rect 58348 612682 58400 612688
rect 50988 612672 51040 612678
rect 50988 612614 51040 612620
rect 58360 612105 58388 612682
rect 58532 612672 58584 612678
rect 58530 612640 58532 612649
rect 58584 612640 58586 612649
rect 58530 612575 58586 612584
rect 58346 612096 58402 612105
rect 58346 612031 58402 612040
rect 655244 601792 655296 601798
rect 655244 601734 655296 601740
rect 50988 601724 51040 601730
rect 50988 601666 51040 601672
rect 48228 601316 48280 601322
rect 48228 601258 48280 601264
rect 46112 600908 46164 600914
rect 46112 600850 46164 600856
rect 46020 590028 46072 590034
rect 46020 589970 46072 589976
rect 46032 230994 46060 589970
rect 46124 571334 46152 600850
rect 46112 571328 46164 571334
rect 46112 571270 46164 571276
rect 48240 568546 48268 601258
rect 51000 571266 51028 601666
rect 655256 594289 655284 601734
rect 655440 595377 655468 612818
rect 655426 595368 655482 595377
rect 655426 595303 655482 595312
rect 655242 594280 655298 594289
rect 655242 594215 655298 594224
rect 58532 585200 58584 585206
rect 58532 585142 58584 585148
rect 58544 574841 58572 585142
rect 59268 582616 59320 582622
rect 59268 582558 59320 582564
rect 58530 574832 58586 574841
rect 58530 574767 58586 574776
rect 59280 573617 59308 582558
rect 655532 579834 655560 643175
rect 655624 624034 655652 688191
rect 655716 668098 655744 731439
rect 655808 715290 655836 776999
rect 656544 774761 656572 783838
rect 656530 774752 656586 774761
rect 656530 774687 656586 774696
rect 655980 747992 656032 747998
rect 655980 747934 656032 747940
rect 655886 732728 655942 732737
rect 655886 732663 655942 732672
rect 655796 715284 655848 715290
rect 655796 715226 655848 715232
rect 655794 689480 655850 689489
rect 655794 689415 655850 689424
rect 655704 668092 655756 668098
rect 655704 668034 655756 668040
rect 655704 656940 655756 656946
rect 655704 656882 655756 656888
rect 655716 640257 655744 656882
rect 655702 640248 655758 640257
rect 655702 640183 655758 640192
rect 655808 624170 655836 689415
rect 655900 670954 655928 732663
rect 655992 731377 656020 747934
rect 656072 736976 656124 736982
rect 656072 736918 656124 736924
rect 655978 731368 656034 731377
rect 655978 731303 656034 731312
rect 656084 728657 656112 736918
rect 656070 728648 656126 728657
rect 656070 728583 656126 728592
rect 655980 703928 656032 703934
rect 655980 703870 656032 703876
rect 655992 687041 656020 703870
rect 655978 687032 656034 687041
rect 655978 686967 656034 686976
rect 655888 670948 655940 670954
rect 655888 670890 655940 670896
rect 656440 645924 656492 645930
rect 656440 645866 656492 645872
rect 655886 641880 655942 641889
rect 655886 641815 655942 641824
rect 655796 624164 655848 624170
rect 655796 624106 655848 624112
rect 655612 624028 655664 624034
rect 655612 623970 655664 623976
rect 655612 601724 655664 601730
rect 655612 601666 655664 601672
rect 655624 593065 655652 601666
rect 655702 596592 655758 596601
rect 655702 596527 655758 596536
rect 655610 593056 655666 593065
rect 655610 592991 655666 593000
rect 655520 579828 655572 579834
rect 655520 579770 655572 579776
rect 60648 574116 60700 574122
rect 60648 574058 60700 574064
rect 59266 573608 59322 573617
rect 59266 573543 59322 573552
rect 60660 572393 60688 574058
rect 60646 572384 60702 572393
rect 60646 572319 60702 572328
rect 58072 571328 58124 571334
rect 58072 571270 58124 571276
rect 50988 571260 51040 571266
rect 50988 571202 51040 571208
rect 58084 571033 58112 571270
rect 58348 571260 58400 571266
rect 58348 571202 58400 571208
rect 58070 571024 58126 571033
rect 58070 570959 58126 570968
rect 58360 570081 58388 571202
rect 58346 570072 58402 570081
rect 58346 570007 58402 570016
rect 48228 568540 48280 568546
rect 48228 568482 48280 568488
rect 58256 568540 58308 568546
rect 58256 568482 58308 568488
rect 58268 568313 58296 568482
rect 58254 568304 58310 568313
rect 58254 568239 58310 568248
rect 50988 558340 51040 558346
rect 50988 558282 51040 558288
rect 48320 557932 48372 557938
rect 48320 557874 48372 557880
rect 46112 557592 46164 557598
rect 46112 557534 46164 557540
rect 46124 529922 46152 557534
rect 48228 546916 48280 546922
rect 48228 546858 48280 546864
rect 46112 529916 46164 529922
rect 46112 529858 46164 529864
rect 46112 430092 46164 430098
rect 46112 430034 46164 430040
rect 46124 400178 46152 430034
rect 46112 400172 46164 400178
rect 46112 400114 46164 400120
rect 46112 386844 46164 386850
rect 46112 386786 46164 386792
rect 46124 358766 46152 386786
rect 46112 358760 46164 358766
rect 46112 358702 46164 358708
rect 46112 343460 46164 343466
rect 46112 343402 46164 343408
rect 46124 314634 46152 343402
rect 46112 314628 46164 314634
rect 46112 314570 46164 314576
rect 46296 287088 46348 287094
rect 46296 287030 46348 287036
rect 46204 278860 46256 278866
rect 46204 278802 46256 278808
rect 46112 278792 46164 278798
rect 46112 278734 46164 278740
rect 46020 230988 46072 230994
rect 46020 230930 46072 230936
rect 45928 219428 45980 219434
rect 45928 219370 45980 219376
rect 45652 216640 45704 216646
rect 45652 216582 45704 216588
rect 46124 214742 46152 278734
rect 46216 215150 46244 278802
rect 46308 257582 46336 287030
rect 46296 257576 46348 257582
rect 46296 257518 46348 257524
rect 46296 247716 46348 247722
rect 46296 247658 46348 247664
rect 46308 216714 46336 247658
rect 48240 230858 48268 546858
rect 48332 527134 48360 557874
rect 48320 527128 48372 527134
rect 48320 527070 48372 527076
rect 51000 527066 51028 558282
rect 654232 557592 654284 557598
rect 654232 557534 654284 557540
rect 654140 554804 654192 554810
rect 654140 554746 654192 554752
rect 654152 548593 654180 554746
rect 654244 549273 654272 557534
rect 655426 553344 655482 553353
rect 655426 553279 655482 553288
rect 654230 549264 654286 549273
rect 654230 549199 654286 549208
rect 654138 548584 654194 548593
rect 654138 548519 654194 548528
rect 59268 541068 59320 541074
rect 59268 541010 59320 541016
rect 59280 530641 59308 541010
rect 59452 541000 59504 541006
rect 59452 540942 59504 540948
rect 59464 531729 59492 540942
rect 59450 531720 59506 531729
rect 59450 531655 59506 531664
rect 59266 530632 59322 530641
rect 59266 530567 59322 530576
rect 58532 529984 58584 529990
rect 58532 529926 58584 529932
rect 58348 529916 58400 529922
rect 58348 529858 58400 529864
rect 58360 528193 58388 529858
rect 58544 529417 58572 529926
rect 58530 529408 58586 529417
rect 58530 529343 58586 529352
rect 58346 528184 58402 528193
rect 58346 528119 58402 528128
rect 58072 527128 58124 527134
rect 58072 527070 58124 527076
rect 50988 527060 51040 527066
rect 50988 527002 51040 527008
rect 57980 527060 58032 527066
rect 57980 527002 58032 527008
rect 57992 526969 58020 527002
rect 57978 526960 58034 526969
rect 57978 526895 58034 526904
rect 58084 525881 58112 527070
rect 58070 525872 58126 525881
rect 58070 525807 58126 525816
rect 655440 491434 655468 553279
rect 655610 552120 655666 552129
rect 655610 552055 655666 552064
rect 655518 551032 655574 551041
rect 655518 550967 655574 550976
rect 655532 491570 655560 550967
rect 655624 491706 655652 552055
rect 655716 535634 655744 596527
rect 655794 595504 655850 595513
rect 655794 595439 655850 595448
rect 655704 535628 655756 535634
rect 655704 535570 655756 535576
rect 655808 532914 655836 595439
rect 655900 579970 655928 641815
rect 656070 640656 656126 640665
rect 656070 640591 656126 640600
rect 655978 597816 656034 597825
rect 655978 597751 656034 597760
rect 655888 579964 655940 579970
rect 655888 579906 655940 579912
rect 655888 568676 655940 568682
rect 655888 568618 655940 568624
rect 655900 550905 655928 568618
rect 655886 550896 655942 550905
rect 655886 550831 655942 550840
rect 655992 535770 656020 597751
rect 656084 580106 656112 640591
rect 656452 638217 656480 645866
rect 656438 638208 656494 638217
rect 656438 638143 656494 638152
rect 656072 580100 656124 580106
rect 656072 580042 656124 580048
rect 655980 535764 656032 535770
rect 655980 535706 656032 535712
rect 655796 532908 655848 532914
rect 655796 532850 655848 532856
rect 655612 491700 655664 491706
rect 655612 491642 655664 491648
rect 655520 491564 655572 491570
rect 655520 491506 655572 491512
rect 655428 491428 655480 491434
rect 655428 491370 655480 491376
rect 50988 430908 51040 430914
rect 50988 430850 51040 430856
rect 48412 430500 48464 430506
rect 48412 430442 48464 430448
rect 48320 419484 48372 419490
rect 48320 419426 48372 419432
rect 48332 230926 48360 419426
rect 48424 400110 48452 430442
rect 48412 400104 48464 400110
rect 48412 400046 48464 400052
rect 51000 400042 51028 430850
rect 58440 405680 58492 405686
rect 58440 405622 58492 405628
rect 58452 404161 58480 405622
rect 58438 404152 58494 404161
rect 58438 404087 58494 404096
rect 655704 403164 655756 403170
rect 655704 403106 655756 403112
rect 655520 403096 655572 403102
rect 655520 403038 655572 403044
rect 655428 403028 655480 403034
rect 655428 402970 655480 402976
rect 58532 402960 58584 402966
rect 58530 402928 58532 402937
rect 58584 402928 58586 402937
rect 58530 402863 58586 402872
rect 60370 400752 60426 400761
rect 60370 400687 60426 400696
rect 58440 400172 58492 400178
rect 58440 400114 58492 400120
rect 58348 400104 58400 400110
rect 58452 400081 58480 400114
rect 58348 400046 58400 400052
rect 58438 400072 58494 400081
rect 50988 400036 51040 400042
rect 50988 399978 51040 399984
rect 58360 398313 58388 400046
rect 58438 400007 58494 400016
rect 58532 400036 58584 400042
rect 58532 399978 58584 399984
rect 58544 399401 58572 399978
rect 58530 399392 58586 399401
rect 58530 399327 58586 399336
rect 58346 398304 58402 398313
rect 58346 398239 58402 398248
rect 60384 394670 60412 400687
rect 60372 394664 60424 394670
rect 60372 394606 60424 394612
rect 50988 387524 51040 387530
rect 50988 387466 51040 387472
rect 48504 387116 48556 387122
rect 48504 387058 48556 387064
rect 48412 376100 48464 376106
rect 48412 376042 48464 376048
rect 48320 230920 48372 230926
rect 48320 230862 48372 230868
rect 48228 230852 48280 230858
rect 48228 230794 48280 230800
rect 48424 230586 48452 376042
rect 48516 356046 48544 387058
rect 48504 356040 48556 356046
rect 48504 355982 48556 355988
rect 51000 355978 51028 387466
rect 654508 372564 654560 372570
rect 654508 372506 654560 372512
rect 654520 370977 654548 372506
rect 655440 372201 655468 402970
rect 655532 374513 655560 403038
rect 655518 374504 655574 374513
rect 655518 374439 655574 374448
rect 655716 373289 655744 403106
rect 655702 373280 655758 373289
rect 655702 373215 655758 373224
rect 655426 372192 655482 372201
rect 655426 372127 655482 372136
rect 654506 370968 654562 370977
rect 654506 370903 654562 370912
rect 58164 361548 58216 361554
rect 58164 361490 58216 361496
rect 58176 360913 58204 361490
rect 58532 361344 58584 361350
rect 58532 361286 58584 361292
rect 58162 360904 58218 360913
rect 58162 360839 58218 360848
rect 58544 359825 58572 361286
rect 58530 359816 58586 359825
rect 58530 359751 58586 359760
rect 58532 358760 58584 358766
rect 58532 358702 58584 358708
rect 57978 357504 58034 357513
rect 57978 357439 58034 357448
rect 50988 355972 51040 355978
rect 50988 355914 51040 355920
rect 57992 350538 58020 357439
rect 58544 357377 58572 358702
rect 58530 357368 58586 357377
rect 58530 357303 58586 357312
rect 655520 356448 655572 356454
rect 655520 356390 655572 356396
rect 655428 356312 655480 356318
rect 655428 356254 655480 356260
rect 58440 356040 58492 356046
rect 58440 355982 58492 355988
rect 58452 355065 58480 355982
rect 58532 355972 58584 355978
rect 58532 355914 58584 355920
rect 58544 355881 58572 355914
rect 58530 355872 58586 355881
rect 58530 355807 58586 355816
rect 58438 355056 58494 355065
rect 58438 354991 58494 355000
rect 57980 350532 58032 350538
rect 57980 350474 58032 350480
rect 50988 344276 51040 344282
rect 50988 344218 51040 344224
rect 48504 343868 48556 343874
rect 48504 343810 48556 343816
rect 48516 311846 48544 343810
rect 48596 333124 48648 333130
rect 48596 333066 48648 333072
rect 48504 311840 48556 311846
rect 48504 311782 48556 311788
rect 48504 281580 48556 281586
rect 48504 281522 48556 281528
rect 48412 230580 48464 230586
rect 48412 230522 48464 230528
rect 46296 216708 46348 216714
rect 46296 216650 46348 216656
rect 46204 215144 46256 215150
rect 46204 215086 46256 215092
rect 46112 214736 46164 214742
rect 46112 214678 46164 214684
rect 41512 212152 41564 212158
rect 41512 212094 41564 212100
rect 43628 212152 43680 212158
rect 43628 212094 43680 212100
rect 32954 211848 33010 211857
rect 32954 211783 33010 211792
rect 41524 211449 41552 212094
rect 41510 211440 41566 211449
rect 41510 211375 41566 211384
rect 32862 211032 32918 211041
rect 32862 210967 32918 210976
rect 30010 210216 30066 210225
rect 30010 210151 30066 210160
rect 25134 204912 25190 204921
rect 25134 204847 25190 204856
rect 24950 204504 25006 204513
rect 24950 204439 25006 204448
rect 24858 203688 24914 203697
rect 24858 203623 24914 203632
rect 30024 200161 30052 210151
rect 30194 209808 30250 209817
rect 30194 209743 30250 209752
rect 30102 209400 30158 209409
rect 30102 209335 30158 209344
rect 30116 200297 30144 209335
rect 30208 200666 30236 209743
rect 41510 208992 41566 209001
rect 41510 208927 41566 208936
rect 38014 208584 38070 208593
rect 38014 208519 38070 208528
rect 30286 208176 30342 208185
rect 30286 208111 30342 208120
rect 30196 200660 30248 200666
rect 30196 200602 30248 200608
rect 30300 200530 30328 208111
rect 38028 201482 38056 208519
rect 41524 208282 41552 208927
rect 41512 208276 41564 208282
rect 41512 208218 41564 208224
rect 43352 208276 43404 208282
rect 43352 208218 43404 208224
rect 38106 207768 38162 207777
rect 38106 207703 38162 207712
rect 38016 201476 38068 201482
rect 38016 201418 38068 201424
rect 38120 201385 38148 207703
rect 41510 207360 41566 207369
rect 41510 207295 41512 207304
rect 41564 207295 41566 207304
rect 41512 207266 41564 207272
rect 41786 207224 41842 207233
rect 41786 207159 41788 207168
rect 41840 207159 41842 207168
rect 41788 207130 41840 207136
rect 41418 206544 41474 206553
rect 41418 206479 41474 206488
rect 41432 201414 41460 206479
rect 41694 206136 41750 206145
rect 41694 206071 41750 206080
rect 41602 205320 41658 205329
rect 41602 205255 41658 205264
rect 41510 204912 41566 204921
rect 41510 204847 41566 204856
rect 41420 201408 41472 201414
rect 38106 201376 38162 201385
rect 41420 201350 41472 201356
rect 38106 201311 38162 201320
rect 30288 200524 30340 200530
rect 30288 200466 30340 200472
rect 30102 200288 30158 200297
rect 30102 200223 30158 200232
rect 30010 200152 30066 200161
rect 30010 200087 30066 200096
rect 41524 198830 41552 204847
rect 41616 199170 41644 205255
rect 41604 199164 41656 199170
rect 41604 199106 41656 199112
rect 41708 199034 41736 206071
rect 41786 206000 41842 206009
rect 41786 205935 41842 205944
rect 41696 199028 41748 199034
rect 41696 198970 41748 198976
rect 41800 198966 41828 205935
rect 43076 201408 43128 201414
rect 43076 201350 43128 201356
rect 42708 200660 42760 200666
rect 42708 200602 42760 200608
rect 42248 200524 42300 200530
rect 42248 200466 42300 200472
rect 41788 198960 41840 198966
rect 41788 198902 41840 198908
rect 41512 198824 41564 198830
rect 41512 198766 41564 198772
rect 42260 196670 42288 200466
rect 42340 198824 42392 198830
rect 42340 198766 42392 198772
rect 42182 196642 42288 196670
rect 42248 196580 42300 196586
rect 42248 196522 42300 196528
rect 42260 194834 42288 196522
rect 42182 194806 42288 194834
rect 42064 193520 42116 193526
rect 42064 193462 42116 193468
rect 42076 192984 42104 193462
rect 42352 191774 42380 198766
rect 42720 196586 42748 200602
rect 42708 196580 42760 196586
rect 42708 196522 42760 196528
rect 43088 193526 43116 201350
rect 43168 199164 43220 199170
rect 43168 199106 43220 199112
rect 43076 193520 43128 193526
rect 43076 193462 43128 193468
rect 42182 191746 42380 191774
rect 43180 191690 43208 199106
rect 43260 199028 43312 199034
rect 43260 198970 43312 198976
rect 42340 191684 42392 191690
rect 42340 191626 42392 191632
rect 43168 191684 43220 191690
rect 43168 191626 43220 191632
rect 42064 191480 42116 191486
rect 42064 191422 42116 191428
rect 42076 191148 42104 191422
rect 42352 190482 42380 191626
rect 43272 191486 43300 198970
rect 43260 191480 43312 191486
rect 43260 191422 43312 191428
rect 42182 190454 42380 190482
rect 42248 190188 42300 190194
rect 42248 190130 42300 190136
rect 42156 190120 42208 190126
rect 42156 190062 42208 190068
rect 42168 189924 42196 190062
rect 42156 187876 42208 187882
rect 42156 187818 42208 187824
rect 42168 187445 42196 187818
rect 42156 187196 42208 187202
rect 42156 187138 42208 187144
rect 42168 186796 42196 187138
rect 42168 186130 42196 186184
rect 42260 186130 42288 190130
rect 43364 189174 43392 208218
rect 43444 207324 43496 207330
rect 43444 207266 43496 207272
rect 43456 190194 43484 207266
rect 43720 207188 43772 207194
rect 43720 207130 43772 207136
rect 43536 201476 43588 201482
rect 43536 201418 43588 201424
rect 43444 190188 43496 190194
rect 43444 190130 43496 190136
rect 43548 190126 43576 201418
rect 43628 198960 43680 198966
rect 43628 198902 43680 198908
rect 43536 190120 43588 190126
rect 43536 190062 43588 190068
rect 42432 189168 42484 189174
rect 42432 189110 42484 189116
rect 43352 189168 43404 189174
rect 43352 189110 43404 189116
rect 42168 186102 42288 186130
rect 42444 185619 42472 189110
rect 43640 187882 43668 198902
rect 43628 187876 43680 187882
rect 43628 187818 43680 187824
rect 43732 187202 43760 207130
rect 43720 187196 43772 187202
rect 43720 187138 43772 187144
rect 42182 185591 42472 185619
rect 41878 184240 41934 184249
rect 41878 184175 41934 184184
rect 41892 183765 41920 184175
rect 41786 183424 41842 183433
rect 41786 183359 41842 183368
rect 41800 183124 41828 183359
rect 41786 183016 41842 183025
rect 41786 182951 41842 182960
rect 41800 182477 41828 182951
rect 48516 182170 48544 281522
rect 48608 230790 48636 333066
rect 51000 314566 51028 344218
rect 655440 328273 655468 356254
rect 655532 329905 655560 356390
rect 655612 356244 655664 356250
rect 655612 356186 655664 356192
rect 655518 329896 655574 329905
rect 655518 329831 655574 329840
rect 655426 328264 655482 328273
rect 655426 328199 655482 328208
rect 655624 327457 655652 356186
rect 655980 335368 656032 335374
rect 655980 335310 656032 335316
rect 655610 327448 655666 327457
rect 655610 327383 655666 327392
rect 655992 325689 656020 335310
rect 655978 325680 656034 325689
rect 655978 325615 656034 325624
rect 58532 318776 58584 318782
rect 58532 318718 58584 318724
rect 58072 317416 58124 317422
rect 58544 317393 58572 318718
rect 58072 317358 58124 317364
rect 58530 317384 58586 317393
rect 58084 316577 58112 317358
rect 58530 317319 58586 317328
rect 58070 316568 58126 316577
rect 58070 316503 58126 316512
rect 58346 314800 58402 314809
rect 58346 314735 58402 314744
rect 50988 314560 51040 314566
rect 50988 314502 51040 314508
rect 58164 314560 58216 314566
rect 58164 314502 58216 314508
rect 58176 313041 58204 314502
rect 58162 313032 58218 313041
rect 58162 312967 58218 312976
rect 58360 306338 58388 314735
rect 58532 314628 58584 314634
rect 58532 314570 58584 314576
rect 58544 314129 58572 314570
rect 58530 314120 58586 314129
rect 58530 314055 58586 314064
rect 655428 312112 655480 312118
rect 655428 312054 655480 312060
rect 58532 311840 58584 311846
rect 58530 311808 58532 311817
rect 58584 311808 58586 311817
rect 58530 311743 58586 311752
rect 58348 306332 58400 306338
rect 58348 306274 58400 306280
rect 655440 300801 655468 312054
rect 655704 312044 655756 312050
rect 655704 311986 655756 311992
rect 655520 311976 655572 311982
rect 655520 311918 655572 311924
rect 655532 303385 655560 311918
rect 655518 303376 655574 303385
rect 655518 303311 655574 303320
rect 655716 302161 655744 311986
rect 655702 302152 655758 302161
rect 655702 302087 655758 302096
rect 655426 300792 655482 300801
rect 655426 300727 655482 300736
rect 655058 298752 655114 298761
rect 655058 298687 655114 298696
rect 655072 298178 655100 298687
rect 655060 298172 655112 298178
rect 655060 298114 655112 298120
rect 656070 297528 656126 297537
rect 656070 297463 656126 297472
rect 655886 296304 655942 296313
rect 655886 296239 655942 296248
rect 58530 295488 58586 295497
rect 58530 295423 58586 295432
rect 58544 295390 58572 295423
rect 58532 295384 58584 295390
rect 58532 295326 58584 295332
rect 58438 293992 58494 294001
rect 58438 293927 58494 293936
rect 655702 293992 655758 294001
rect 655702 293927 655758 293936
rect 58452 292670 58480 293927
rect 59266 292768 59322 292777
rect 59266 292703 59322 292712
rect 655518 292768 655574 292777
rect 655518 292703 655574 292712
rect 58440 292664 58492 292670
rect 58440 292606 58492 292612
rect 57980 292528 58032 292534
rect 57980 292470 58032 292476
rect 57992 291553 58020 292470
rect 58532 292460 58584 292466
rect 58532 292402 58584 292408
rect 58544 292369 58572 292402
rect 58530 292360 58586 292369
rect 58530 292295 58586 292304
rect 57978 291544 58034 291553
rect 57978 291479 58034 291488
rect 51080 291100 51132 291106
rect 51080 291042 51132 291048
rect 48780 289876 48832 289882
rect 48780 289818 48832 289824
rect 48688 287156 48740 287162
rect 48688 287098 48740 287104
rect 48596 230784 48648 230790
rect 48596 230726 48648 230732
rect 48700 225622 48728 287098
rect 48792 230518 48820 289818
rect 50988 281648 51040 281654
rect 50988 281590 51040 281596
rect 48872 246492 48924 246498
rect 48872 246434 48924 246440
rect 48780 230512 48832 230518
rect 48780 230454 48832 230460
rect 48884 230450 48912 246434
rect 48872 230444 48924 230450
rect 48872 230386 48924 230392
rect 48688 225616 48740 225622
rect 48688 225558 48740 225564
rect 51000 214334 51028 281590
rect 51092 230654 51120 291042
rect 51172 290692 51224 290698
rect 51172 290634 51224 290640
rect 51184 230722 51212 290634
rect 57980 289808 58032 289814
rect 57978 289776 57980 289785
rect 58032 289776 58034 289785
rect 57978 289711 58034 289720
rect 58162 288008 58218 288017
rect 58162 287943 58218 287952
rect 58176 287162 58204 287943
rect 58530 287192 58586 287201
rect 58164 287156 58216 287162
rect 58530 287127 58586 287136
rect 58164 287098 58216 287104
rect 58544 287094 58572 287127
rect 58532 287088 58584 287094
rect 58532 287030 58584 287036
rect 57978 285696 58034 285705
rect 57978 285631 58034 285640
rect 57992 284850 58020 285631
rect 56508 284844 56560 284850
rect 56508 284786 56560 284792
rect 57980 284844 58032 284850
rect 57980 284786 58032 284792
rect 51264 284368 51316 284374
rect 51264 284310 51316 284316
rect 51276 257718 51304 284310
rect 51264 257712 51316 257718
rect 51264 257654 51316 257660
rect 56520 256766 56548 284786
rect 58530 284472 58586 284481
rect 58530 284407 58586 284416
rect 58544 284374 58572 284407
rect 58532 284368 58584 284374
rect 58532 284310 58584 284316
rect 58530 283248 58586 283257
rect 58530 283183 58586 283192
rect 58254 282160 58310 282169
rect 58254 282095 58310 282104
rect 58268 281654 58296 282095
rect 58256 281648 58308 281654
rect 58256 281590 58308 281596
rect 58544 281586 58572 283183
rect 58532 281580 58584 281586
rect 58532 281522 58584 281528
rect 58162 280936 58218 280945
rect 58162 280871 58218 280880
rect 58176 278866 58204 280871
rect 58254 279712 58310 279721
rect 58254 279647 58310 279656
rect 58164 278860 58216 278866
rect 58164 278802 58216 278808
rect 58268 278798 58296 279647
rect 58256 278792 58308 278798
rect 58256 278734 58308 278740
rect 59280 271862 59308 292703
rect 654506 289232 654562 289241
rect 654506 289167 654562 289176
rect 654520 288590 654548 289167
rect 654508 288584 654560 288590
rect 654508 288526 654560 288532
rect 654874 288008 654930 288017
rect 654874 287943 654930 287952
rect 654888 287094 654916 287943
rect 654876 287088 654928 287094
rect 654876 287030 654928 287036
rect 655426 285696 655482 285705
rect 655426 285631 655482 285640
rect 655440 284986 655468 285631
rect 655428 284980 655480 284986
rect 655428 284922 655480 284928
rect 654874 284744 654930 284753
rect 654874 284679 654876 284688
rect 654928 284679 654930 284688
rect 654876 284650 654928 284656
rect 655426 283248 655482 283257
rect 655426 283183 655482 283192
rect 654690 280936 654746 280945
rect 654690 280871 654746 280880
rect 654704 280226 654732 280871
rect 654692 280220 654744 280226
rect 654692 280162 654744 280168
rect 654874 279984 654930 279993
rect 654874 279919 654930 279928
rect 654888 279002 654916 279919
rect 654876 278996 654928 279002
rect 654876 278938 654928 278944
rect 59268 271856 59320 271862
rect 59268 271798 59320 271804
rect 65904 269142 65932 278052
rect 67100 271862 67128 278052
rect 67088 271856 67140 271862
rect 67088 271798 67140 271804
rect 65892 269136 65944 269142
rect 65892 269078 65944 269084
rect 68204 266354 68232 278052
rect 69400 271833 69428 278052
rect 69386 271824 69442 271833
rect 69386 271759 69442 271768
rect 70596 269113 70624 278052
rect 71792 270706 71820 278052
rect 71780 270700 71832 270706
rect 71780 270642 71832 270648
rect 70582 269104 70638 269113
rect 70582 269039 70638 269048
rect 72988 266490 73016 278052
rect 74184 267986 74212 278052
rect 75380 269278 75408 278052
rect 75368 269272 75420 269278
rect 76484 269249 76512 278052
rect 77680 271998 77708 278052
rect 77668 271992 77720 271998
rect 77668 271934 77720 271940
rect 78876 269385 78904 278052
rect 80072 272105 80100 278052
rect 81268 272241 81296 278052
rect 81254 272232 81310 272241
rect 81254 272167 81310 272176
rect 80058 272096 80114 272105
rect 80058 272031 80114 272040
rect 78862 269376 78918 269385
rect 82464 269346 82492 278052
rect 83660 271969 83688 278052
rect 84764 272377 84792 278052
rect 84750 272368 84806 272377
rect 84750 272303 84806 272312
rect 83646 271960 83702 271969
rect 83646 271895 83702 271904
rect 85960 269657 85988 278052
rect 85946 269648 86002 269657
rect 85946 269583 86002 269592
rect 87156 269521 87184 278052
rect 88352 272270 88380 278052
rect 89548 272474 89576 278052
rect 90744 272513 90772 278052
rect 90730 272504 90786 272513
rect 89536 272468 89588 272474
rect 90730 272439 90786 272448
rect 89536 272410 89588 272416
rect 88340 272264 88392 272270
rect 88340 272206 88392 272212
rect 87142 269512 87198 269521
rect 87142 269447 87198 269456
rect 91848 269414 91876 278052
rect 93044 269793 93072 278052
rect 93030 269784 93086 269793
rect 93030 269719 93086 269728
rect 94240 269482 94268 278052
rect 95436 272649 95464 278052
rect 95422 272640 95478 272649
rect 95422 272575 95478 272584
rect 96632 272066 96660 278052
rect 97828 272134 97856 278052
rect 97816 272128 97868 272134
rect 97816 272070 97868 272076
rect 96620 272060 96672 272066
rect 96620 272002 96672 272008
rect 99024 269929 99052 278052
rect 99010 269920 99066 269929
rect 99010 269855 99066 269864
rect 100128 269550 100156 278052
rect 101324 269686 101352 278052
rect 102520 272202 102548 278052
rect 103716 272785 103744 278052
rect 104912 272921 104940 278052
rect 104898 272912 104954 272921
rect 104898 272847 104954 272856
rect 103702 272776 103758 272785
rect 103702 272711 103758 272720
rect 102508 272196 102560 272202
rect 102508 272138 102560 272144
rect 106108 270065 106136 278052
rect 107212 270201 107240 278052
rect 108408 270337 108436 278052
rect 109604 273057 109632 278052
rect 110800 273193 110828 278052
rect 110786 273184 110842 273193
rect 110786 273119 110842 273128
rect 109590 273048 109646 273057
rect 109590 272983 109646 272992
rect 111996 272406 112024 278052
rect 111984 272400 112036 272406
rect 111984 272342 112036 272348
rect 108394 270328 108450 270337
rect 108394 270263 108450 270272
rect 107198 270192 107254 270201
rect 107198 270127 107254 270136
rect 106094 270056 106150 270065
rect 106094 269991 106150 270000
rect 101312 269680 101364 269686
rect 101312 269622 101364 269628
rect 100116 269544 100168 269550
rect 100116 269486 100168 269492
rect 94228 269476 94280 269482
rect 94228 269418 94280 269424
rect 91836 269408 91888 269414
rect 91836 269350 91888 269356
rect 78862 269311 78918 269320
rect 82452 269340 82504 269346
rect 82452 269282 82504 269288
rect 75368 269214 75420 269220
rect 76470 269240 76526 269249
rect 76470 269175 76526 269184
rect 74172 267980 74224 267986
rect 74172 267922 74224 267928
rect 72976 266484 73028 266490
rect 72976 266426 73028 266432
rect 113192 266422 113220 278052
rect 114388 270473 114416 278052
rect 114374 270464 114430 270473
rect 114374 270399 114430 270408
rect 115492 269618 115520 278052
rect 115480 269612 115532 269618
rect 115480 269554 115532 269560
rect 116688 266558 116716 278052
rect 117884 272338 117912 278052
rect 119080 272678 119108 278052
rect 119068 272672 119120 272678
rect 119068 272614 119120 272620
rect 117872 272332 117924 272338
rect 117872 272274 117924 272280
rect 120276 271697 120304 278052
rect 120262 271688 120318 271697
rect 120262 271623 120318 271632
rect 121472 268977 121500 278052
rect 122576 269754 122604 278052
rect 122564 269748 122616 269754
rect 122564 269690 122616 269696
rect 121458 268968 121514 268977
rect 121458 268903 121514 268912
rect 123772 266626 123800 278052
rect 124968 271561 124996 278052
rect 126164 272610 126192 278052
rect 126152 272604 126204 272610
rect 126152 272546 126204 272552
rect 127360 271794 127388 278052
rect 127348 271788 127400 271794
rect 127348 271730 127400 271736
rect 124954 271552 125010 271561
rect 124954 271487 125010 271496
rect 128556 269822 128584 278052
rect 129660 269890 129688 278052
rect 130856 269958 130884 278052
rect 132052 271289 132080 278052
rect 132038 271280 132094 271289
rect 132038 271215 132094 271224
rect 133248 271153 133276 278052
rect 134444 271425 134472 278052
rect 134430 271416 134486 271425
rect 134430 271351 134486 271360
rect 133234 271144 133290 271153
rect 133234 271079 133290 271088
rect 135640 270230 135668 278052
rect 135628 270224 135680 270230
rect 135628 270166 135680 270172
rect 136836 270094 136864 278052
rect 136824 270088 136876 270094
rect 136824 270030 136876 270036
rect 137940 270026 137968 278052
rect 139136 272814 139164 278052
rect 139124 272808 139176 272814
rect 139124 272750 139176 272756
rect 140332 272678 140360 278052
rect 141528 272746 141556 278052
rect 141516 272740 141568 272746
rect 141516 272682 141568 272688
rect 140320 272672 140372 272678
rect 140320 272614 140372 272620
rect 142724 270162 142752 278052
rect 143920 270298 143948 278052
rect 145116 270366 145144 278052
rect 146220 272882 146248 278052
rect 147416 273018 147444 278052
rect 147404 273012 147456 273018
rect 147404 272954 147456 272960
rect 146208 272876 146260 272882
rect 146208 272818 146260 272824
rect 148612 270434 148640 278052
rect 149808 272950 149836 278052
rect 149796 272944 149848 272950
rect 149796 272886 149848 272892
rect 151004 270570 151032 278052
rect 152200 273086 152228 278052
rect 152188 273080 152240 273086
rect 152188 273022 152240 273028
rect 150992 270564 151044 270570
rect 150992 270506 151044 270512
rect 148600 270428 148652 270434
rect 148600 270370 148652 270376
rect 145104 270360 145156 270366
rect 145104 270302 145156 270308
rect 143908 270292 143960 270298
rect 143908 270234 143960 270240
rect 142712 270156 142764 270162
rect 142712 270098 142764 270104
rect 137928 270020 137980 270026
rect 137928 269962 137980 269968
rect 130844 269952 130896 269958
rect 130844 269894 130896 269900
rect 129648 269884 129700 269890
rect 129648 269826 129700 269832
rect 128544 269816 128596 269822
rect 128544 269758 128596 269764
rect 153396 269074 153424 278052
rect 154500 273222 154528 278052
rect 154488 273216 154540 273222
rect 154488 273158 154540 273164
rect 153384 269068 153436 269074
rect 153384 269010 153436 269016
rect 155696 268938 155724 278052
rect 156892 271930 156920 278052
rect 156880 271924 156932 271930
rect 156880 271866 156932 271872
rect 158088 269006 158116 278052
rect 159284 271726 159312 278052
rect 159272 271720 159324 271726
rect 159272 271662 159324 271668
rect 158076 269000 158128 269006
rect 158076 268942 158128 268948
rect 155684 268932 155736 268938
rect 155684 268874 155736 268880
rect 160480 268870 160508 278052
rect 161584 271590 161612 278052
rect 161572 271584 161624 271590
rect 161572 271526 161624 271532
rect 160468 268864 160520 268870
rect 160468 268806 160520 268812
rect 162780 268734 162808 278052
rect 163976 271658 164004 278052
rect 163964 271652 164016 271658
rect 163964 271594 164016 271600
rect 165172 268802 165200 278052
rect 166368 271386 166396 278052
rect 166356 271380 166408 271386
rect 166356 271322 166408 271328
rect 165160 268796 165212 268802
rect 165160 268738 165212 268744
rect 162768 268728 162820 268734
rect 162768 268670 162820 268676
rect 167564 268666 167592 278052
rect 168760 271454 168788 278052
rect 168748 271448 168800 271454
rect 168748 271390 168800 271396
rect 167552 268660 167604 268666
rect 167552 268602 167604 268608
rect 169864 268598 169892 278052
rect 171060 271522 171088 278052
rect 171048 271516 171100 271522
rect 171048 271458 171100 271464
rect 169852 268592 169904 268598
rect 169852 268534 169904 268540
rect 172256 268530 172284 278052
rect 173452 271318 173480 278052
rect 173440 271312 173492 271318
rect 173440 271254 173492 271260
rect 172244 268524 172296 268530
rect 172244 268466 172296 268472
rect 174648 268462 174676 278052
rect 175844 271182 175872 278052
rect 176844 273148 176896 273154
rect 176844 273090 176896 273096
rect 176856 271930 176884 273090
rect 176948 271930 176976 278052
rect 177120 272468 177172 272474
rect 177120 272410 177172 272416
rect 176844 271924 176896 271930
rect 176844 271866 176896 271872
rect 176936 271924 176988 271930
rect 176936 271866 176988 271872
rect 175832 271176 175884 271182
rect 175832 271118 175884 271124
rect 174636 268456 174688 268462
rect 174636 268398 174688 268404
rect 177132 268054 177160 272410
rect 178144 271250 178172 278052
rect 178132 271244 178184 271250
rect 178132 271186 178184 271192
rect 179340 270774 179368 278052
rect 180536 271046 180564 278052
rect 180524 271040 180576 271046
rect 180524 270982 180576 270988
rect 179328 270768 179380 270774
rect 179328 270710 179380 270716
rect 181732 268394 181760 278052
rect 181720 268388 181772 268394
rect 181720 268330 181772 268336
rect 182928 268190 182956 278052
rect 184124 270910 184152 278052
rect 185228 272270 185256 278052
rect 184940 272264 184992 272270
rect 184940 272206 184992 272212
rect 185216 272264 185268 272270
rect 185216 272206 185268 272212
rect 184112 270904 184164 270910
rect 184112 270846 184164 270852
rect 184112 270768 184164 270774
rect 184112 270710 184164 270716
rect 184124 268326 184152 270710
rect 184952 268841 184980 272206
rect 186424 271114 186452 278052
rect 186412 271108 186464 271114
rect 186412 271050 186464 271056
rect 187620 270978 187648 278052
rect 187700 272536 187752 272542
rect 187700 272478 187752 272484
rect 187608 270972 187660 270978
rect 187608 270914 187660 270920
rect 187712 270774 187740 272478
rect 187700 270768 187752 270774
rect 187700 270710 187752 270716
rect 184938 268832 184994 268841
rect 184938 268767 184994 268776
rect 184112 268320 184164 268326
rect 184112 268262 184164 268268
rect 182916 268184 182968 268190
rect 182916 268126 182968 268132
rect 188816 268122 188844 278052
rect 189908 271788 189960 271794
rect 189908 271730 189960 271736
rect 189920 270638 189948 271730
rect 190012 270842 190040 278052
rect 191208 271862 191236 278052
rect 191196 271856 191248 271862
rect 191196 271798 191248 271804
rect 190000 270836 190052 270842
rect 190000 270778 190052 270784
rect 189908 270632 189960 270638
rect 189908 270574 189960 270580
rect 192404 270570 192432 278052
rect 193508 272610 193536 278052
rect 193496 272604 193548 272610
rect 193496 272546 193548 272552
rect 193220 271992 193272 271998
rect 193220 271934 193272 271940
rect 193128 271924 193180 271930
rect 193128 271866 193180 271872
rect 192484 271788 192536 271794
rect 192484 271730 192536 271736
rect 192392 270564 192444 270570
rect 192392 270506 192444 270512
rect 192392 269136 192444 269142
rect 192392 269078 192444 269084
rect 188804 268116 188856 268122
rect 188804 268058 188856 268064
rect 177120 268048 177172 268054
rect 177120 267990 177172 267996
rect 123760 266620 123812 266626
rect 123760 266562 123812 266568
rect 116676 266552 116728 266558
rect 116676 266494 116728 266500
rect 113180 266416 113232 266422
rect 113180 266358 113232 266364
rect 68192 266348 68244 266354
rect 68192 266290 68244 266296
rect 192404 264316 192432 269078
rect 192496 264330 192524 271730
rect 193140 267918 193168 271866
rect 193232 268258 193260 271934
rect 194704 271930 194732 278052
rect 194692 271924 194744 271930
rect 194692 271866 194744 271872
rect 193678 271824 193734 271833
rect 193678 271759 193734 271768
rect 193220 268252 193272 268258
rect 193220 268194 193272 268200
rect 193128 267912 193180 267918
rect 193128 267854 193180 267860
rect 193220 266348 193272 266354
rect 193220 266290 193272 266296
rect 192496 264302 192786 264330
rect 193232 264316 193260 266290
rect 193692 264316 193720 271759
rect 194600 270700 194652 270706
rect 194600 270642 194652 270648
rect 194138 269104 194194 269113
rect 194138 269039 194194 269048
rect 194152 264316 194180 269039
rect 194612 264316 194640 270642
rect 195428 269272 195480 269278
rect 195428 269214 195480 269220
rect 195060 266484 195112 266490
rect 195060 266426 195112 266432
rect 195072 264316 195100 266426
rect 195440 264316 195468 269214
rect 195900 269142 195928 278052
rect 196898 272096 196954 272105
rect 196898 272031 196954 272040
rect 195978 269240 196034 269249
rect 195978 269175 196034 269184
rect 195888 269136 195940 269142
rect 195888 269078 195940 269084
rect 195888 267980 195940 267986
rect 195888 267922 195940 267928
rect 195900 264316 195928 267922
rect 195992 264330 196020 269175
rect 196348 268252 196400 268258
rect 196348 268194 196400 268200
rect 196360 264974 196388 268194
rect 196360 264946 196480 264974
rect 196452 264330 196480 264946
rect 196912 264330 196940 272031
rect 197096 269210 197124 278052
rect 197268 272536 197320 272542
rect 197268 272478 197320 272484
rect 197280 272270 197308 272478
rect 197268 272264 197320 272270
rect 197268 272206 197320 272212
rect 198094 272232 198150 272241
rect 198094 272167 198150 272176
rect 197176 270632 197228 270638
rect 197176 270574 197228 270580
rect 197084 269204 197136 269210
rect 197084 269146 197136 269152
rect 197188 267782 197216 270574
rect 197726 269376 197782 269385
rect 197726 269311 197782 269320
rect 197268 268184 197320 268190
rect 197268 268126 197320 268132
rect 197280 267986 197308 268126
rect 197268 267980 197320 267986
rect 197268 267922 197320 267928
rect 197176 267776 197228 267782
rect 197176 267718 197228 267724
rect 195992 264302 196374 264330
rect 196452 264302 196834 264330
rect 196912 264302 197294 264330
rect 197740 264316 197768 269311
rect 198108 264316 198136 272167
rect 198292 271998 198320 278052
rect 199106 272368 199162 272377
rect 199106 272303 199162 272312
rect 198832 272128 198884 272134
rect 198832 272070 198884 272076
rect 198740 272060 198792 272066
rect 198740 272002 198792 272008
rect 198280 271992 198332 271998
rect 198280 271934 198332 271940
rect 198752 269385 198780 272002
rect 198738 269376 198794 269385
rect 198556 269340 198608 269346
rect 198738 269311 198794 269320
rect 198556 269282 198608 269288
rect 198568 264316 198596 269282
rect 198844 268122 198872 272070
rect 198832 268116 198884 268122
rect 198832 268058 198884 268064
rect 199120 264330 199148 272303
rect 199382 271960 199438 271969
rect 199382 271895 199438 271904
rect 199042 264302 199148 264330
rect 199396 264330 199424 271895
rect 199488 270774 199516 278052
rect 200592 271794 200620 278052
rect 201592 272400 201644 272406
rect 201592 272342 201644 272348
rect 201500 272196 201552 272202
rect 201500 272138 201552 272144
rect 200580 271788 200632 271794
rect 200580 271730 200632 271736
rect 199476 270768 199528 270774
rect 199476 270710 199528 270716
rect 199934 269648 199990 269657
rect 199934 269583 199990 269592
rect 199396 264302 199502 264330
rect 199948 264316 199976 269583
rect 200394 269512 200450 269521
rect 200394 269447 200450 269456
rect 200408 264316 200436 269447
rect 201222 268832 201278 268841
rect 201222 268767 201278 268776
rect 200764 268048 200816 268054
rect 200764 267990 200816 267996
rect 200776 264316 200804 267990
rect 201236 264316 201264 268767
rect 201512 268054 201540 272138
rect 201500 268048 201552 268054
rect 201500 267990 201552 267996
rect 201604 267850 201632 272342
rect 201788 270706 201816 278052
rect 201958 272504 202014 272513
rect 201958 272439 202014 272448
rect 201776 270700 201828 270706
rect 201776 270642 201828 270648
rect 201592 267844 201644 267850
rect 201592 267786 201644 267792
rect 201972 264330 202000 272439
rect 202984 272066 203012 278052
rect 203522 272640 203578 272649
rect 203522 272575 203578 272584
rect 203616 272604 203668 272610
rect 202972 272060 203024 272066
rect 202972 272002 203024 272008
rect 203062 269784 203118 269793
rect 203062 269719 203118 269728
rect 202604 269476 202656 269482
rect 202604 269418 202656 269424
rect 202144 269408 202196 269414
rect 202144 269350 202196 269356
rect 201710 264302 202000 264330
rect 202156 264316 202184 269350
rect 202616 264316 202644 269418
rect 203076 264316 203104 269719
rect 203536 264316 203564 272575
rect 203616 272546 203668 272552
rect 203628 269278 203656 272546
rect 204180 272134 204208 278052
rect 205376 272202 205404 278052
rect 206466 272912 206522 272921
rect 206466 272847 206522 272856
rect 205364 272196 205416 272202
rect 205364 272138 205416 272144
rect 204168 272128 204220 272134
rect 204168 272070 204220 272076
rect 204810 269920 204866 269929
rect 204810 269855 204866 269864
rect 204350 269376 204406 269385
rect 204350 269311 204406 269320
rect 203616 269272 203668 269278
rect 203616 269214 203668 269220
rect 203892 268116 203944 268122
rect 203892 268058 203944 268064
rect 203904 264316 203932 268058
rect 204364 264316 204392 269311
rect 204824 264316 204852 269855
rect 205272 269680 205324 269686
rect 205272 269622 205324 269628
rect 205284 264316 205312 269622
rect 205732 269544 205784 269550
rect 205732 269486 205784 269492
rect 205744 264316 205772 269486
rect 206192 268048 206244 268054
rect 206192 267990 206244 267996
rect 206204 264316 206232 267990
rect 206480 264330 206508 272847
rect 206572 269346 206600 278052
rect 206742 273048 206798 273057
rect 206742 272983 206798 272992
rect 206560 269340 206612 269346
rect 206560 269282 206612 269288
rect 206560 268048 206612 268054
rect 206560 267990 206612 267996
rect 206572 267782 206600 267990
rect 206756 267850 206784 272983
rect 207386 272776 207442 272785
rect 207386 272711 207442 272720
rect 206836 272468 206888 272474
rect 206836 272410 206888 272416
rect 206848 267918 206876 272410
rect 206836 267912 206888 267918
rect 206836 267854 206888 267860
rect 206744 267844 206796 267850
rect 206744 267786 206796 267792
rect 206560 267776 206612 267782
rect 206560 267718 206612 267724
rect 207400 264330 207428 272711
rect 207768 270638 207796 278052
rect 207664 270632 207716 270638
rect 207664 270574 207716 270580
rect 207756 270632 207808 270638
rect 207756 270574 207808 270580
rect 207676 270502 207704 270574
rect 207572 270496 207624 270502
rect 207572 270438 207624 270444
rect 207664 270496 207716 270502
rect 207664 270438 207716 270444
rect 207478 270056 207534 270065
rect 207478 269991 207534 270000
rect 206480 264302 206586 264330
rect 207046 264302 207428 264330
rect 207492 264316 207520 269991
rect 207584 267782 207612 270438
rect 207938 270328 207994 270337
rect 207938 270263 207994 270272
rect 207572 267776 207624 267782
rect 207572 267718 207624 267724
rect 207952 264316 207980 270263
rect 208398 270192 208454 270201
rect 208398 270127 208454 270136
rect 208412 264316 208440 270127
rect 208872 269414 208900 278052
rect 209410 273184 209466 273193
rect 209410 273119 209466 273128
rect 208860 269408 208912 269414
rect 208860 269350 208912 269356
rect 209228 267980 209280 267986
rect 209228 267922 209280 267928
rect 208860 267844 208912 267850
rect 208860 267786 208912 267792
rect 208872 264316 208900 267786
rect 209240 264316 209268 267922
rect 209424 264330 209452 273119
rect 209688 272264 209740 272270
rect 209688 272206 209740 272212
rect 209700 267986 209728 272206
rect 210068 269482 210096 278052
rect 211068 273216 211120 273222
rect 211068 273158 211120 273164
rect 210976 273148 211028 273154
rect 210976 273090 211028 273096
rect 210988 272338 211016 273090
rect 211080 272542 211108 273158
rect 211264 273086 211292 278052
rect 211252 273080 211304 273086
rect 211252 273022 211304 273028
rect 211068 272536 211120 272542
rect 211068 272478 211120 272484
rect 210976 272332 211028 272338
rect 210976 272274 211028 272280
rect 212354 271688 212410 271697
rect 212354 271623 212410 271632
rect 210698 270464 210754 270473
rect 210698 270399 210754 270408
rect 210608 269612 210660 269618
rect 210608 269554 210660 269560
rect 210056 269476 210108 269482
rect 210056 269418 210108 269424
rect 209688 267980 209740 267986
rect 209688 267922 209740 267928
rect 210148 266416 210200 266422
rect 210148 266358 210200 266364
rect 209424 264302 209714 264330
rect 210160 264316 210188 266358
rect 210620 264316 210648 269554
rect 210712 264330 210740 270399
rect 212368 269328 212396 271623
rect 212460 269550 212488 278052
rect 213276 269748 213328 269754
rect 213276 269690 213328 269696
rect 212448 269544 212500 269550
rect 212448 269486 212500 269492
rect 212368 269300 212580 269328
rect 212356 267980 212408 267986
rect 212356 267922 212408 267928
rect 211896 267912 211948 267918
rect 211896 267854 211948 267860
rect 211528 266552 211580 266558
rect 211528 266494 211580 266500
rect 210712 264302 211094 264330
rect 211540 264316 211568 266494
rect 211908 264316 211936 267854
rect 212368 264316 212396 267922
rect 212552 264330 212580 269300
rect 212552 264302 212842 264330
rect 213288 264316 213316 269690
rect 213656 267986 213684 278052
rect 214852 272950 214880 278052
rect 214748 272944 214800 272950
rect 214748 272886 214800 272892
rect 214840 272944 214892 272950
rect 214840 272886 214892 272892
rect 214760 272610 214788 272886
rect 214748 272604 214800 272610
rect 214748 272546 214800 272552
rect 215022 271552 215078 271561
rect 215022 271487 215078 271496
rect 214656 270496 214708 270502
rect 214656 270438 214708 270444
rect 213734 268968 213790 268977
rect 213734 268903 213790 268912
rect 213644 267980 213696 267986
rect 213644 267922 213696 267928
rect 213748 264316 213776 268903
rect 214196 266620 214248 266626
rect 214196 266562 214248 266568
rect 214208 264316 214236 266562
rect 214668 264316 214696 270438
rect 215036 264316 215064 271487
rect 215208 270632 215260 270638
rect 215208 270574 215260 270580
rect 215220 269686 215248 270574
rect 215852 269884 215904 269890
rect 215852 269826 215904 269832
rect 215208 269680 215260 269686
rect 215208 269622 215260 269628
rect 215484 268048 215536 268054
rect 215484 267990 215536 267996
rect 215496 264316 215524 267990
rect 215864 264330 215892 269826
rect 215956 269754 215984 278052
rect 216864 269952 216916 269958
rect 216864 269894 216916 269900
rect 216404 269816 216456 269822
rect 216404 269758 216456 269764
rect 215944 269748 215996 269754
rect 215944 269690 215996 269696
rect 215864 264302 215970 264330
rect 216416 264316 216444 269758
rect 216876 264316 216904 269894
rect 217152 269618 217180 278052
rect 217968 273080 218020 273086
rect 217968 273022 218020 273028
rect 217690 271280 217746 271289
rect 217690 271215 217746 271224
rect 217322 271144 217378 271153
rect 217322 271079 217378 271088
rect 217140 269612 217192 269618
rect 217140 269554 217192 269560
rect 217336 264316 217364 271079
rect 217704 264316 217732 271215
rect 217980 269822 218008 273022
rect 218150 271416 218206 271425
rect 218150 271351 218206 271360
rect 217968 269816 218020 269822
rect 217968 269758 218020 269764
rect 218164 264316 218192 271351
rect 218348 270638 218376 278052
rect 218336 270632 218388 270638
rect 218336 270574 218388 270580
rect 219544 270230 219572 278052
rect 220452 272944 220504 272950
rect 220452 272886 220504 272892
rect 220360 272808 220412 272814
rect 220360 272750 220412 272756
rect 219992 272672 220044 272678
rect 219992 272614 220044 272620
rect 219072 270224 219124 270230
rect 219072 270166 219124 270172
rect 219532 270224 219584 270230
rect 219532 270166 219584 270172
rect 218612 270088 218664 270094
rect 218612 270030 218664 270036
rect 218624 264316 218652 270030
rect 219084 264316 219112 270166
rect 219532 270020 219584 270026
rect 219532 269962 219584 269968
rect 219544 264316 219572 269962
rect 220004 264316 220032 272614
rect 220372 264316 220400 272750
rect 220464 269890 220492 272886
rect 220740 270026 220768 278052
rect 221188 272740 221240 272746
rect 221188 272682 221240 272688
rect 220728 270020 220780 270026
rect 220728 269962 220780 269968
rect 220452 269884 220504 269890
rect 220452 269826 220504 269832
rect 221200 264330 221228 272682
rect 221280 270292 221332 270298
rect 221280 270234 221332 270240
rect 220846 264302 221228 264330
rect 221292 264316 221320 270234
rect 221936 270162 221964 278052
rect 222660 273012 222712 273018
rect 222660 272954 222712 272960
rect 222200 270360 222252 270366
rect 222200 270302 222252 270308
rect 221740 270156 221792 270162
rect 221740 270098 221792 270104
rect 221924 270156 221976 270162
rect 221924 270098 221976 270104
rect 221752 264316 221780 270098
rect 222212 264316 222240 270302
rect 222672 264316 222700 272954
rect 223028 272876 223080 272882
rect 223028 272818 223080 272824
rect 223040 264316 223068 272818
rect 223132 269958 223160 278052
rect 224040 271380 224092 271386
rect 224040 271322 224092 271328
rect 223396 270632 223448 270638
rect 223396 270574 223448 270580
rect 223212 270428 223264 270434
rect 223212 270370 223264 270376
rect 223120 269952 223172 269958
rect 223120 269894 223172 269900
rect 223224 264330 223252 270370
rect 223408 270094 223436 270574
rect 223396 270088 223448 270094
rect 223396 270030 223448 270036
rect 224052 267782 224080 271322
rect 224236 270366 224264 278052
rect 224500 273216 224552 273222
rect 224500 273158 224552 273164
rect 224408 272604 224460 272610
rect 224408 272546 224460 272552
rect 224224 270360 224276 270366
rect 224224 270302 224276 270308
rect 223948 267776 224000 267782
rect 223948 267718 224000 267724
rect 224040 267776 224092 267782
rect 224040 267718 224092 267724
rect 223224 264302 223514 264330
rect 223960 264316 223988 267718
rect 224420 264316 224448 272546
rect 224512 264330 224540 273158
rect 225328 272536 225380 272542
rect 225328 272478 225380 272484
rect 224512 264302 224894 264330
rect 225340 264316 225368 272478
rect 225432 270298 225460 278052
rect 226628 270638 226656 278052
rect 227076 272332 227128 272338
rect 227076 272274 227128 272280
rect 226616 270632 226668 270638
rect 226616 270574 226668 270580
rect 225420 270292 225472 270298
rect 225420 270234 225472 270240
rect 225788 269068 225840 269074
rect 225788 269010 225840 269016
rect 225800 264316 225828 269010
rect 226616 269000 226668 269006
rect 226616 268942 226668 268948
rect 226156 268932 226208 268938
rect 226156 268874 226208 268880
rect 226168 264316 226196 268874
rect 226628 264316 226656 268942
rect 227088 264316 227116 272274
rect 227536 271720 227588 271726
rect 227536 271662 227588 271668
rect 227444 270904 227496 270910
rect 227444 270846 227496 270852
rect 227456 267918 227484 270846
rect 227444 267912 227496 267918
rect 227444 267854 227496 267860
rect 227548 264316 227576 271662
rect 227824 271386 227852 278052
rect 229020 272542 229048 278052
rect 229008 272536 229060 272542
rect 229008 272478 229060 272484
rect 230216 272338 230244 278052
rect 230204 272332 230256 272338
rect 230204 272274 230256 272280
rect 229744 271652 229796 271658
rect 229744 271594 229796 271600
rect 227996 271584 228048 271590
rect 227996 271526 228048 271532
rect 227812 271380 227864 271386
rect 227812 271322 227864 271328
rect 227628 271312 227680 271318
rect 227628 271254 227680 271260
rect 227640 270502 227668 271254
rect 227812 271040 227864 271046
rect 227812 270982 227864 270988
rect 227628 270496 227680 270502
rect 227628 270438 227680 270444
rect 227824 267986 227852 270982
rect 227812 267980 227864 267986
rect 227812 267922 227864 267928
rect 228008 264316 228036 271526
rect 229284 271516 229336 271522
rect 229284 271458 229336 271464
rect 229100 271176 229152 271182
rect 229100 271118 229152 271124
rect 229112 269346 229140 271118
rect 229296 270434 229324 271458
rect 229284 270428 229336 270434
rect 229284 270370 229336 270376
rect 229008 269340 229060 269346
rect 229008 269282 229060 269288
rect 229100 269340 229152 269346
rect 229100 269282 229152 269288
rect 229020 269074 229048 269282
rect 229008 269068 229060 269074
rect 229008 269010 229060 269016
rect 228456 268864 228508 268870
rect 228456 268806 228508 268812
rect 228468 264316 228496 268806
rect 229284 268796 229336 268802
rect 229284 268738 229336 268744
rect 228824 268728 228876 268734
rect 228824 268670 228876 268676
rect 228836 264316 228864 268670
rect 229296 264316 229324 268738
rect 229756 264316 229784 271594
rect 230388 271448 230440 271454
rect 230388 271390 230440 271396
rect 229836 270836 229888 270842
rect 229836 270778 229888 270784
rect 229848 268734 229876 270778
rect 229836 268728 229888 268734
rect 229836 268670 229888 268676
rect 230204 267776 230256 267782
rect 230204 267718 230256 267724
rect 230216 264316 230244 267718
rect 230400 264330 230428 271390
rect 231320 271318 231348 278052
rect 232516 272746 232544 278052
rect 233712 272882 233740 278052
rect 234908 272950 234936 278052
rect 234896 272944 234948 272950
rect 234896 272886 234948 272892
rect 233700 272876 233752 272882
rect 233700 272818 233752 272824
rect 236104 272814 236132 278052
rect 236092 272808 236144 272814
rect 236092 272750 236144 272756
rect 232504 272740 232556 272746
rect 232504 272682 232556 272688
rect 237300 272474 237328 278052
rect 232044 272468 232096 272474
rect 232044 272410 232096 272416
rect 237288 272468 237340 272474
rect 237288 272410 237340 272416
rect 231308 271312 231360 271318
rect 231308 271254 231360 271260
rect 231860 271244 231912 271250
rect 231860 271186 231912 271192
rect 230756 270972 230808 270978
rect 230756 270914 230808 270920
rect 230768 267782 230796 270914
rect 231124 268660 231176 268666
rect 231124 268602 231176 268608
rect 230756 267776 230808 267782
rect 230756 267718 230808 267724
rect 230400 264302 230690 264330
rect 231136 264316 231164 268602
rect 231492 268592 231544 268598
rect 231492 268534 231544 268540
rect 231504 264316 231532 268534
rect 231872 267850 231900 271186
rect 231952 271108 232004 271114
rect 231952 271050 232004 271056
rect 231964 268666 231992 271050
rect 232056 269006 232084 272410
rect 238496 272270 238524 278052
rect 238484 272264 238536 272270
rect 238484 272206 238536 272212
rect 239496 271856 239548 271862
rect 239496 271798 239548 271804
rect 232872 270496 232924 270502
rect 232872 270438 232924 270444
rect 232412 270428 232464 270434
rect 232412 270370 232464 270376
rect 232044 269000 232096 269006
rect 232044 268942 232096 268948
rect 231952 268660 232004 268666
rect 231952 268602 232004 268608
rect 231952 268524 232004 268530
rect 231952 268466 232004 268472
rect 231860 267844 231912 267850
rect 231860 267786 231912 267792
rect 231964 264316 231992 268466
rect 232424 264316 232452 270370
rect 232884 264316 232912 270438
rect 233332 269340 233384 269346
rect 233332 269282 233384 269288
rect 233344 264316 233372 269282
rect 237748 269000 237800 269006
rect 237748 268942 237800 268948
rect 237288 268660 237340 268666
rect 237288 268602 237340 268608
rect 233792 268456 233844 268462
rect 233792 268398 233844 268404
rect 233804 264316 233832 268398
rect 236460 268388 236512 268394
rect 236460 268330 236512 268336
rect 234620 268320 234672 268326
rect 234620 268262 234672 268268
rect 234160 268116 234212 268122
rect 234160 268058 234212 268064
rect 234172 264316 234200 268058
rect 234632 264316 234660 268262
rect 236000 268184 236052 268190
rect 236000 268126 236052 268132
rect 235540 267980 235592 267986
rect 235540 267922 235592 267928
rect 235080 267844 235132 267850
rect 235080 267786 235132 267792
rect 235092 264316 235120 267786
rect 235552 264316 235580 267922
rect 236012 264316 236040 268126
rect 236472 264316 236500 268330
rect 236920 267912 236972 267918
rect 236920 267854 236972 267860
rect 236932 264316 236960 267854
rect 237300 264316 237328 268602
rect 237760 264316 237788 268942
rect 238668 268728 238720 268734
rect 238668 268670 238720 268676
rect 238208 267776 238260 267782
rect 238208 267718 238260 267724
rect 238220 264316 238248 267718
rect 238680 264316 238708 268670
rect 239128 268252 239180 268258
rect 239128 268194 239180 268200
rect 239140 264316 239168 268194
rect 239508 264330 239536 271798
rect 239600 271726 239628 278052
rect 240796 273018 240824 278052
rect 240784 273012 240836 273018
rect 240784 272954 240836 272960
rect 240140 272128 240192 272134
rect 240140 272070 240192 272076
rect 239588 271720 239640 271726
rect 239588 271662 239640 271668
rect 239956 270564 240008 270570
rect 239956 270506 240008 270512
rect 239508 264302 239614 264330
rect 239968 264316 239996 270506
rect 240152 268598 240180 272070
rect 240876 271924 240928 271930
rect 240876 271866 240928 271872
rect 240416 269272 240468 269278
rect 240416 269214 240468 269220
rect 240140 268592 240192 268598
rect 240140 268534 240192 268540
rect 240428 264316 240456 269214
rect 240888 264316 240916 271866
rect 241992 271522 242020 278052
rect 243188 273086 243216 278052
rect 243176 273080 243228 273086
rect 243176 273022 243228 273028
rect 244004 272060 244056 272066
rect 244004 272002 244056 272008
rect 242256 271992 242308 271998
rect 242256 271934 242308 271940
rect 241980 271516 242032 271522
rect 241980 271458 242032 271464
rect 241796 269204 241848 269210
rect 241796 269146 241848 269152
rect 241336 269136 241388 269142
rect 241336 269078 241388 269084
rect 241348 264316 241376 269078
rect 241808 264316 241836 269146
rect 242268 264316 242296 271934
rect 243268 271788 243320 271794
rect 243268 271730 243320 271736
rect 242624 270768 242676 270774
rect 242624 270710 242676 270716
rect 242636 264316 242664 270710
rect 243280 264330 243308 271730
rect 243544 270700 243596 270706
rect 243544 270642 243596 270648
rect 243110 264302 243308 264330
rect 243556 264316 243584 270642
rect 244016 264316 244044 272002
rect 244384 271998 244412 278052
rect 244924 272196 244976 272202
rect 244924 272138 244976 272144
rect 244372 271992 244424 271998
rect 244372 271934 244424 271940
rect 244464 268592 244516 268598
rect 244464 268534 244516 268540
rect 244476 264316 244504 268534
rect 244936 264316 244964 272138
rect 245580 271658 245608 278052
rect 245568 271652 245620 271658
rect 245568 271594 245620 271600
rect 246776 271182 246804 278052
rect 247880 271862 247908 278052
rect 247868 271856 247920 271862
rect 247868 271798 247920 271804
rect 249076 271794 249104 278052
rect 249064 271788 249116 271794
rect 249064 271730 249116 271736
rect 250272 271318 250300 278052
rect 251468 271726 251496 278052
rect 251456 271720 251508 271726
rect 251456 271662 251508 271668
rect 251180 271652 251232 271658
rect 251180 271594 251232 271600
rect 250260 271312 250312 271318
rect 250260 271254 250312 271260
rect 246764 271176 246816 271182
rect 246764 271118 246816 271124
rect 251192 271046 251220 271594
rect 251272 271516 251324 271522
rect 251272 271458 251324 271464
rect 251284 271114 251312 271458
rect 252664 271386 252692 278052
rect 253756 272536 253808 272542
rect 253756 272478 253808 272484
rect 253388 271448 253440 271454
rect 253388 271390 253440 271396
rect 252652 271380 252704 271386
rect 252652 271322 252704 271328
rect 251272 271108 251324 271114
rect 251272 271050 251324 271056
rect 251180 271040 251232 271046
rect 251180 270982 251232 270988
rect 252928 270632 252980 270638
rect 252928 270574 252980 270580
rect 252008 270360 252060 270366
rect 252008 270302 252060 270308
rect 250260 270224 250312 270230
rect 250260 270166 250312 270172
rect 249800 270088 249852 270094
rect 249800 270030 249852 270036
rect 248420 269884 248472 269890
rect 248420 269826 248472 269832
rect 247132 269816 247184 269822
rect 247132 269758 247184 269764
rect 245752 269680 245804 269686
rect 245752 269622 245804 269628
rect 245292 269068 245344 269074
rect 245292 269010 245344 269016
rect 245304 264316 245332 269010
rect 245764 264316 245792 269622
rect 246672 269476 246724 269482
rect 246672 269418 246724 269424
rect 246212 269408 246264 269414
rect 246212 269350 246264 269356
rect 246224 264316 246252 269350
rect 246684 264316 246712 269418
rect 247144 264316 247172 269758
rect 247592 269544 247644 269550
rect 247592 269486 247644 269492
rect 247604 264316 247632 269486
rect 248052 268048 248104 268054
rect 248052 267990 248104 267996
rect 248064 264316 248092 267990
rect 248432 264316 248460 269826
rect 248880 269748 248932 269754
rect 248880 269690 248932 269696
rect 248892 264316 248920 269690
rect 249340 269612 249392 269618
rect 249340 269554 249392 269560
rect 249352 264316 249380 269554
rect 249812 264316 249840 270030
rect 250272 264316 250300 270166
rect 251088 270156 251140 270162
rect 251088 270098 251140 270104
rect 250720 270020 250772 270026
rect 250720 269962 250772 269968
rect 250732 264316 250760 269962
rect 251100 264316 251128 270098
rect 251548 269952 251600 269958
rect 251548 269894 251600 269900
rect 251560 264316 251588 269894
rect 252020 264316 252048 270302
rect 252468 270292 252520 270298
rect 252468 270234 252520 270240
rect 252480 264316 252508 270234
rect 252940 264316 252968 270574
rect 253400 264316 253428 271390
rect 253768 264316 253796 272478
rect 253860 271658 253888 278052
rect 254216 272332 254268 272338
rect 254216 272274 254268 272280
rect 253848 271652 253900 271658
rect 253848 271594 253900 271600
rect 254228 264316 254256 272274
rect 254964 271454 254992 278052
rect 256056 272944 256108 272950
rect 256056 272886 256108 272892
rect 255596 272876 255648 272882
rect 255596 272818 255648 272824
rect 255136 272740 255188 272746
rect 255136 272682 255188 272688
rect 254952 271448 255004 271454
rect 254952 271390 255004 271396
rect 254676 271244 254728 271250
rect 254676 271186 254728 271192
rect 254688 264316 254716 271186
rect 255148 264316 255176 272682
rect 255608 264316 255636 272818
rect 256068 264316 256096 272886
rect 256160 270706 256188 278052
rect 256424 272808 256476 272814
rect 256424 272750 256476 272756
rect 256148 270700 256200 270706
rect 256148 270642 256200 270648
rect 256436 264316 256464 272750
rect 256884 272468 256936 272474
rect 256884 272410 256936 272416
rect 256896 264316 256924 272410
rect 257252 272264 257304 272270
rect 257252 272206 257304 272212
rect 257264 264330 257292 272206
rect 257356 271590 257384 278052
rect 258264 273012 258316 273018
rect 258264 272954 258316 272960
rect 257344 271584 257396 271590
rect 257344 271526 257396 271532
rect 257804 271516 257856 271522
rect 257804 271458 257856 271464
rect 257264 264302 257370 264330
rect 257816 264316 257844 271458
rect 258276 264316 258304 272954
rect 258552 271522 258580 278052
rect 259748 273086 259776 278052
rect 260944 273154 260972 278052
rect 260932 273148 260984 273154
rect 260932 273090 260984 273096
rect 259184 273080 259236 273086
rect 259184 273022 259236 273028
rect 259736 273080 259788 273086
rect 259736 273022 259788 273028
rect 258540 271516 258592 271522
rect 258540 271458 258592 271464
rect 258724 271108 258776 271114
rect 258724 271050 258776 271056
rect 258736 264316 258764 271050
rect 259196 264316 259224 273022
rect 262140 271998 262168 278052
rect 263244 273222 263272 278052
rect 263232 273216 263284 273222
rect 263232 273158 263284 273164
rect 259552 271992 259604 271998
rect 259552 271934 259604 271940
rect 262128 271992 262180 271998
rect 262128 271934 262180 271940
rect 259564 264316 259592 271934
rect 264440 271862 264468 278052
rect 265440 273080 265492 273086
rect 265440 273022 265492 273028
rect 260932 271856 260984 271862
rect 260932 271798 260984 271804
rect 264428 271856 264480 271862
rect 264428 271798 264480 271804
rect 260472 271176 260524 271182
rect 260472 271118 260524 271124
rect 260012 271040 260064 271046
rect 260012 270982 260064 270988
rect 260024 264316 260052 270982
rect 260484 264316 260512 271118
rect 260944 264316 260972 271798
rect 261392 271788 261444 271794
rect 261392 271730 261444 271736
rect 261404 264316 261432 271730
rect 262220 271720 262272 271726
rect 262220 271662 262272 271668
rect 261852 271312 261904 271318
rect 261852 271254 261904 271260
rect 261864 264316 261892 271254
rect 262232 264316 262260 271662
rect 263140 271652 263192 271658
rect 263140 271594 263192 271600
rect 262864 271380 262916 271386
rect 262864 271322 262916 271328
rect 262876 264330 262904 271322
rect 262706 264302 262904 264330
rect 263152 264316 263180 271594
rect 264520 271584 264572 271590
rect 264520 271526 264572 271532
rect 263600 271448 263652 271454
rect 263600 271390 263652 271396
rect 263612 264316 263640 271390
rect 264060 270700 264112 270706
rect 264060 270642 264112 270648
rect 264072 264316 264100 270642
rect 264532 264316 264560 271526
rect 264888 271516 264940 271522
rect 264888 271458 264940 271464
rect 264900 264316 264928 271458
rect 265452 264330 265480 273022
rect 265636 270502 265664 278052
rect 266728 273216 266780 273222
rect 266728 273158 266780 273164
rect 265808 273148 265860 273154
rect 265808 273090 265860 273096
rect 265624 270496 265676 270502
rect 265624 270438 265676 270444
rect 265374 264302 265480 264330
rect 265820 264316 265848 273090
rect 266268 271992 266320 271998
rect 266268 271934 266320 271940
rect 266280 264316 266308 271934
rect 266740 264316 266768 273158
rect 266832 271522 266860 278052
rect 268042 278038 268516 278066
rect 267188 271856 267240 271862
rect 267188 271798 267240 271804
rect 266820 271516 266872 271522
rect 266820 271458 266872 271464
rect 267200 264316 267228 271798
rect 268016 271516 268068 271522
rect 268016 271458 268068 271464
rect 267556 270496 267608 270502
rect 267556 270438 267608 270444
rect 267568 264316 267596 270438
rect 268028 264316 268056 271458
rect 268488 264316 268516 278038
rect 268948 278038 269146 278066
rect 268948 264316 268976 278038
rect 270328 270502 270356 278052
rect 269396 270496 269448 270502
rect 269396 270438 269448 270444
rect 270316 270496 270368 270502
rect 270316 270438 270368 270444
rect 270684 270496 270736 270502
rect 270684 270438 270736 270444
rect 269408 264316 269436 270438
rect 269856 268524 269908 268530
rect 269856 268466 269908 268472
rect 269868 264316 269896 268466
rect 270316 268184 270368 268190
rect 270316 268126 270368 268132
rect 270328 264316 270356 268126
rect 270696 264316 270724 270438
rect 271144 270428 271196 270434
rect 271144 270370 271196 270376
rect 271156 264316 271184 270370
rect 271524 268530 271552 278052
rect 271604 270360 271656 270366
rect 271604 270302 271656 270308
rect 271512 268524 271564 268530
rect 271512 268466 271564 268472
rect 271616 264316 271644 270302
rect 272064 270292 272116 270298
rect 272064 270234 272116 270240
rect 272076 264316 272104 270234
rect 272524 270224 272576 270230
rect 272524 270166 272576 270172
rect 272536 264316 272564 270166
rect 272720 268190 272748 278052
rect 273916 270502 273944 278052
rect 273904 270496 273956 270502
rect 273904 270438 273956 270444
rect 274272 270496 274324 270502
rect 274272 270438 274324 270444
rect 272984 270156 273036 270162
rect 272984 270098 273036 270104
rect 272708 268184 272760 268190
rect 272708 268126 272760 268132
rect 272996 264316 273024 270098
rect 273720 270088 273772 270094
rect 273720 270030 273772 270036
rect 273732 264330 273760 270030
rect 273812 270020 273864 270026
rect 273812 269962 273864 269968
rect 273378 264302 273760 264330
rect 273824 264316 273852 269962
rect 274284 264316 274312 270438
rect 275112 270434 275140 278052
rect 275100 270428 275152 270434
rect 275100 270370 275152 270376
rect 276216 270366 276244 278052
rect 276204 270360 276256 270366
rect 276204 270302 276256 270308
rect 277412 270298 277440 278052
rect 277492 270428 277544 270434
rect 277492 270370 277544 270376
rect 277400 270292 277452 270298
rect 277400 270234 277452 270240
rect 275652 269476 275704 269482
rect 275652 269418 275704 269424
rect 274732 268320 274784 268326
rect 274732 268262 274784 268268
rect 274744 264316 274772 268262
rect 275192 268252 275244 268258
rect 275192 268194 275244 268200
rect 275204 264316 275232 268194
rect 275664 264316 275692 269418
rect 276940 269340 276992 269346
rect 276940 269282 276992 269288
rect 276480 268388 276532 268394
rect 276480 268330 276532 268336
rect 276296 267912 276348 267918
rect 276296 267854 276348 267860
rect 276308 264330 276336 267854
rect 276046 264302 276336 264330
rect 276492 264316 276520 268330
rect 276952 264316 276980 269282
rect 277504 264330 277532 270370
rect 277860 270360 277912 270366
rect 277860 270302 277912 270308
rect 277426 264302 277532 264330
rect 277872 264316 277900 270302
rect 278608 270230 278636 278052
rect 278688 270292 278740 270298
rect 278688 270234 278740 270240
rect 278596 270224 278648 270230
rect 278596 270166 278648 270172
rect 278320 269884 278372 269890
rect 278320 269826 278372 269832
rect 278332 264316 278360 269826
rect 278700 264316 278728 270234
rect 279148 270224 279200 270230
rect 279148 270166 279200 270172
rect 279160 264316 279188 270166
rect 279804 270162 279832 278052
rect 279792 270156 279844 270162
rect 279792 270098 279844 270104
rect 281000 270094 281028 278052
rect 280988 270088 281040 270094
rect 280988 270030 281040 270036
rect 282196 270026 282224 278052
rect 283392 270502 283420 278052
rect 284208 272264 284260 272270
rect 284208 272206 284260 272212
rect 283380 270496 283432 270502
rect 283380 270438 283432 270444
rect 282552 270292 282604 270298
rect 282552 270234 282604 270240
rect 282368 270088 282420 270094
rect 282368 270030 282420 270036
rect 282184 270020 282236 270026
rect 282184 269962 282236 269968
rect 279608 269952 279660 269958
rect 279608 269894 279660 269900
rect 279620 264316 279648 269894
rect 282380 269890 282408 270030
rect 282368 269884 282420 269890
rect 282368 269826 282420 269832
rect 282460 269884 282512 269890
rect 282460 269826 282512 269832
rect 280528 269816 280580 269822
rect 280528 269758 280580 269764
rect 280068 269748 280120 269754
rect 280068 269690 280120 269696
rect 280080 264316 280108 269690
rect 280540 264316 280568 269758
rect 281816 269680 281868 269686
rect 281816 269622 281868 269628
rect 281448 269612 281500 269618
rect 281448 269554 281500 269560
rect 280988 269544 281040 269550
rect 280988 269486 281040 269492
rect 281000 264316 281028 269486
rect 281460 264316 281488 269554
rect 281828 264316 281856 269622
rect 282472 269482 282500 269826
rect 282460 269476 282512 269482
rect 282460 269418 282512 269424
rect 282276 269408 282328 269414
rect 282276 269350 282328 269356
rect 282288 264316 282316 269350
rect 282564 269346 282592 270234
rect 282736 269476 282788 269482
rect 282736 269418 282788 269424
rect 282552 269340 282604 269346
rect 282552 269282 282604 269288
rect 282748 264316 282776 269418
rect 283656 269340 283708 269346
rect 283656 269282 283708 269288
rect 283196 269272 283248 269278
rect 283196 269214 283248 269220
rect 283208 264316 283236 269214
rect 283668 264316 283696 269282
rect 284220 264330 284248 272206
rect 284496 268326 284524 278052
rect 285404 271380 285456 271386
rect 285404 271322 285456 271328
rect 284944 269204 284996 269210
rect 284944 269146 284996 269152
rect 284576 269136 284628 269142
rect 284576 269078 284628 269084
rect 284484 268320 284536 268326
rect 284484 268262 284536 268268
rect 284588 264330 284616 269078
rect 284142 264302 284248 264330
rect 284510 264302 284616 264330
rect 284956 264316 284984 269146
rect 285416 264316 285444 271322
rect 285692 268258 285720 278052
rect 285864 272196 285916 272202
rect 285864 272138 285916 272144
rect 285680 268252 285732 268258
rect 285680 268194 285732 268200
rect 285876 264316 285904 272138
rect 286692 272060 286744 272066
rect 286692 272002 286744 272008
rect 286600 271992 286652 271998
rect 286600 271934 286652 271940
rect 286612 264330 286640 271934
rect 286350 264302 286640 264330
rect 286704 264330 286732 272002
rect 286888 269890 286916 278052
rect 287612 271448 287664 271454
rect 287612 271390 287664 271396
rect 287152 271312 287204 271318
rect 287152 271254 287204 271260
rect 286876 269884 286928 269890
rect 286876 269826 286928 269832
rect 286704 264302 286810 264330
rect 287164 264316 287192 271254
rect 287624 264316 287652 271390
rect 288084 267918 288112 278052
rect 288164 272400 288216 272406
rect 288164 272342 288216 272348
rect 288072 267912 288124 267918
rect 288072 267854 288124 267860
rect 288176 264330 288204 272342
rect 288532 272128 288584 272134
rect 288532 272070 288584 272076
rect 288098 264302 288204 264330
rect 288544 264316 288572 272070
rect 289176 271924 289228 271930
rect 289176 271866 289228 271872
rect 289188 264330 289216 271866
rect 289280 268394 289308 278052
rect 289636 271856 289688 271862
rect 289636 271798 289688 271804
rect 289268 268388 289320 268394
rect 289268 268330 289320 268336
rect 289648 264330 289676 271798
rect 290280 271652 290332 271658
rect 290280 271594 290332 271600
rect 289820 271516 289872 271522
rect 289820 271458 289872 271464
rect 289018 264302 289216 264330
rect 289478 264302 289676 264330
rect 289832 264316 289860 271458
rect 290292 264316 290320 271594
rect 290476 270298 290504 278052
rect 291200 271720 291252 271726
rect 291200 271662 291252 271668
rect 290740 271584 290792 271590
rect 290740 271526 290792 271532
rect 290464 270292 290516 270298
rect 290464 270234 290516 270240
rect 290752 264316 290780 271526
rect 291212 264316 291240 271662
rect 291580 270434 291608 278052
rect 292120 273216 292172 273222
rect 292120 273158 292172 273164
rect 292028 271788 292080 271794
rect 292028 271730 292080 271736
rect 291568 270428 291620 270434
rect 291568 270370 291620 270376
rect 292040 264330 292068 271730
rect 291686 264302 292068 264330
rect 292132 264316 292160 273158
rect 292580 272264 292632 272270
rect 292580 272206 292632 272212
rect 292592 264316 292620 272206
rect 292776 270230 292804 278052
rect 293868 273148 293920 273154
rect 293868 273090 293920 273096
rect 293408 272604 293460 272610
rect 293408 272546 293460 272552
rect 292764 270224 292816 270230
rect 292764 270166 292816 270172
rect 292948 269068 293000 269074
rect 292948 269010 293000 269016
rect 292960 264316 292988 269010
rect 293420 264316 293448 272546
rect 293880 264316 293908 273090
rect 293972 270094 294000 278052
rect 294880 272876 294932 272882
rect 294880 272818 294932 272824
rect 294328 270496 294380 270502
rect 294328 270438 294380 270444
rect 293960 270088 294012 270094
rect 293960 270030 294012 270036
rect 294340 264316 294368 270438
rect 294892 264330 294920 272818
rect 295064 272808 295116 272814
rect 295064 272750 295116 272756
rect 294814 264302 294920 264330
rect 295076 264330 295104 272750
rect 295168 270162 295196 278052
rect 296076 273080 296128 273086
rect 296076 273022 296128 273028
rect 295616 270428 295668 270434
rect 295616 270370 295668 270376
rect 295156 270156 295208 270162
rect 295156 270098 295208 270104
rect 295076 264302 295274 264330
rect 295628 264316 295656 270370
rect 296088 264316 296116 273022
rect 296364 270026 296392 278052
rect 297456 270360 297508 270366
rect 297456 270302 297508 270308
rect 296996 270292 297048 270298
rect 296996 270234 297048 270240
rect 296352 270020 296404 270026
rect 296352 269962 296404 269968
rect 296536 268728 296588 268734
rect 296536 268670 296588 268676
rect 296548 264316 296576 268670
rect 297008 264316 297036 270234
rect 297468 264316 297496 270302
rect 297560 269958 297588 278052
rect 298284 270224 298336 270230
rect 298284 270166 298336 270172
rect 297548 269952 297600 269958
rect 297548 269894 297600 269900
rect 297916 268864 297968 268870
rect 297916 268806 297968 268812
rect 297928 264316 297956 268806
rect 298296 264316 298324 270166
rect 298756 269754 298784 278052
rect 298836 270156 298888 270162
rect 298836 270098 298888 270104
rect 298744 269748 298796 269754
rect 298744 269690 298796 269696
rect 298848 264330 298876 270098
rect 299860 269822 299888 278052
rect 300584 270088 300636 270094
rect 300584 270030 300636 270036
rect 300124 270020 300176 270026
rect 300124 269962 300176 269968
rect 299848 269816 299900 269822
rect 299848 269758 299900 269764
rect 299204 268932 299256 268938
rect 299204 268874 299256 268880
rect 298770 264302 298876 264330
rect 299216 264316 299244 268874
rect 299664 267232 299716 267238
rect 299664 267174 299716 267180
rect 299676 264316 299704 267174
rect 300136 264316 300164 269962
rect 300596 264316 300624 270030
rect 301056 269550 301084 278052
rect 301872 273012 301924 273018
rect 301872 272954 301924 272960
rect 301412 269952 301464 269958
rect 301412 269894 301464 269900
rect 301044 269544 301096 269550
rect 301044 269486 301096 269492
rect 300952 267164 301004 267170
rect 300952 267106 301004 267112
rect 300964 264316 300992 267106
rect 301424 264316 301452 269894
rect 301884 264316 301912 272954
rect 302252 269618 302280 278052
rect 302792 269816 302844 269822
rect 302792 269758 302844 269764
rect 302240 269612 302292 269618
rect 302240 269554 302292 269560
rect 302332 267096 302384 267102
rect 302332 267038 302384 267044
rect 302344 264316 302372 267038
rect 302804 264316 302832 269758
rect 303448 269686 303476 278052
rect 303528 272944 303580 272950
rect 303528 272886 303580 272892
rect 303436 269680 303488 269686
rect 303436 269622 303488 269628
rect 303540 264330 303568 272886
rect 304080 271244 304132 271250
rect 304080 271186 304132 271192
rect 303712 267028 303764 267034
rect 303712 266970 303764 266976
rect 303278 264302 303568 264330
rect 303724 264316 303752 266970
rect 304092 264316 304120 271186
rect 304540 269612 304592 269618
rect 304540 269554 304592 269560
rect 304552 264316 304580 269554
rect 304644 269414 304672 278052
rect 305840 269482 305868 278052
rect 306748 272672 306800 272678
rect 306748 272614 306800 272620
rect 306288 272468 306340 272474
rect 306288 272410 306340 272416
rect 305828 269476 305880 269482
rect 305828 269418 305880 269424
rect 304632 269408 304684 269414
rect 304632 269350 304684 269356
rect 305460 269000 305512 269006
rect 305460 268942 305512 268948
rect 305000 266960 305052 266966
rect 305000 266902 305052 266908
rect 305012 264316 305040 266902
rect 305472 264316 305500 268942
rect 306300 264330 306328 272410
rect 306380 266892 306432 266898
rect 306380 266834 306432 266840
rect 305946 264302 306328 264330
rect 306392 264316 306420 266834
rect 306760 264316 306788 272614
rect 307036 269278 307064 278052
rect 307208 272536 307260 272542
rect 307208 272478 307260 272484
rect 307024 269272 307076 269278
rect 307024 269214 307076 269220
rect 307220 264316 307248 272478
rect 308140 269346 308168 278052
rect 309336 272338 309364 278052
rect 309324 272332 309376 272338
rect 309324 272274 309376 272280
rect 309876 272332 309928 272338
rect 309876 272274 309928 272280
rect 308220 269884 308272 269890
rect 308220 269826 308272 269832
rect 308128 269340 308180 269346
rect 308128 269282 308180 269288
rect 307668 266824 307720 266830
rect 307668 266766 307720 266772
rect 307680 264316 307708 266766
rect 308232 264330 308260 269826
rect 308588 269476 308640 269482
rect 308588 269418 308640 269424
rect 308154 264302 308260 264330
rect 308600 264316 308628 269418
rect 309416 268252 309468 268258
rect 309416 268194 309468 268200
rect 309048 266756 309100 266762
rect 309048 266698 309100 266704
rect 309060 264316 309088 266698
rect 309428 264316 309456 268194
rect 309888 264316 309916 272274
rect 310532 269142 310560 278052
rect 310796 269748 310848 269754
rect 310796 269690 310848 269696
rect 310520 269136 310572 269142
rect 310520 269078 310572 269084
rect 310336 266688 310388 266694
rect 310336 266630 310388 266636
rect 310348 264316 310376 266630
rect 310808 264316 310836 269690
rect 311256 269408 311308 269414
rect 311256 269350 311308 269356
rect 311268 264316 311296 269350
rect 311728 269210 311756 278052
rect 312924 271386 312952 278052
rect 314120 272202 314148 278052
rect 314108 272196 314160 272202
rect 314108 272138 314160 272144
rect 315224 271998 315252 278052
rect 316420 272066 316448 278052
rect 317512 274848 317564 274854
rect 317512 274790 317564 274796
rect 316408 272060 316460 272066
rect 316408 272002 316460 272008
rect 317328 272060 317380 272066
rect 317328 272002 317380 272008
rect 315212 271992 315264 271998
rect 315212 271934 315264 271940
rect 312912 271380 312964 271386
rect 312912 271322 312964 271328
rect 315212 271380 315264 271386
rect 315212 271322 315264 271328
rect 313188 270632 313240 270638
rect 313188 270574 313240 270580
rect 311716 269204 311768 269210
rect 311716 269146 311768 269152
rect 313200 268734 313228 270574
rect 313464 269680 313516 269686
rect 313464 269622 313516 269628
rect 313188 268728 313240 268734
rect 313188 268670 313240 268676
rect 312084 268660 312136 268666
rect 312084 268602 312136 268608
rect 311716 266620 311768 266626
rect 311716 266562 311768 266568
rect 311728 264316 311756 266562
rect 312096 264316 312124 268602
rect 312544 268524 312596 268530
rect 312544 268466 312596 268472
rect 312556 264316 312584 268466
rect 313004 266552 313056 266558
rect 313004 266494 313056 266500
rect 313016 264316 313044 266494
rect 313476 264316 313504 269622
rect 313924 269340 313976 269346
rect 313924 269282 313976 269288
rect 313936 264316 313964 269282
rect 314844 267776 314896 267782
rect 314844 267718 314896 267724
rect 314384 265260 314436 265266
rect 314384 265202 314436 265208
rect 314396 264316 314424 265202
rect 314856 264316 314884 267718
rect 315224 264316 315252 271322
rect 317236 270768 317288 270774
rect 317236 270710 317288 270716
rect 316132 269544 316184 269550
rect 316132 269486 316184 269492
rect 315672 266416 315724 266422
rect 315672 266358 315724 266364
rect 315684 264316 315712 266358
rect 316144 264316 316172 269486
rect 317248 268870 317276 270710
rect 317236 268864 317288 268870
rect 317236 268806 317288 268812
rect 316592 268796 316644 268802
rect 316592 268738 316644 268744
rect 316604 264316 316632 268738
rect 317340 268530 317368 272002
rect 317328 268524 317380 268530
rect 317328 268466 317380 268472
rect 317052 266348 317104 266354
rect 317052 266290 317104 266296
rect 317064 264316 317092 266290
rect 317524 264316 317552 274790
rect 317616 271318 317644 278052
rect 318812 271454 318840 278052
rect 320008 272406 320036 278052
rect 320180 274780 320232 274786
rect 320180 274722 320232 274728
rect 319996 272400 320048 272406
rect 319996 272342 320048 272348
rect 318800 271448 318852 271454
rect 318800 271390 318852 271396
rect 317604 271312 317656 271318
rect 317604 271254 317656 271260
rect 317880 271312 317932 271318
rect 317880 271254 317932 271260
rect 317892 264316 317920 271254
rect 319904 270700 319956 270706
rect 319904 270642 319956 270648
rect 319260 269272 319312 269278
rect 319260 269214 319312 269220
rect 318800 267844 318852 267850
rect 318800 267786 318852 267792
rect 318340 265328 318392 265334
rect 318340 265270 318392 265276
rect 318352 264316 318380 265270
rect 318812 264316 318840 267786
rect 319272 264316 319300 269214
rect 319916 268938 319944 270642
rect 319904 268932 319956 268938
rect 319904 268874 319956 268880
rect 319720 265396 319772 265402
rect 319720 265338 319772 265344
rect 319732 264316 319760 265338
rect 320192 264316 320220 274722
rect 321008 274712 321060 274718
rect 321008 274654 321060 274660
rect 320548 271992 320600 271998
rect 320548 271934 320600 271940
rect 320560 264316 320588 271934
rect 321020 264316 321048 274654
rect 321204 272134 321232 278052
rect 322296 272536 322348 272542
rect 322296 272478 322348 272484
rect 322308 272406 322336 272478
rect 322296 272400 322348 272406
rect 322296 272342 322348 272348
rect 321192 272128 321244 272134
rect 321192 272070 321244 272076
rect 322400 271930 322428 278052
rect 322572 274644 322624 274650
rect 322572 274586 322624 274592
rect 322388 271924 322440 271930
rect 322388 271866 322440 271872
rect 321928 269136 321980 269142
rect 321928 269078 321980 269084
rect 321468 268116 321520 268122
rect 321468 268058 321520 268064
rect 321480 264316 321508 268058
rect 321940 264316 321968 269078
rect 322584 264330 322612 274586
rect 322848 272400 322900 272406
rect 322848 272342 322900 272348
rect 322664 271448 322716 271454
rect 322664 271390 322716 271396
rect 322676 267782 322704 271390
rect 322860 268666 322888 272342
rect 323504 271862 323532 278052
rect 323676 273624 323728 273630
rect 323676 273566 323728 273572
rect 323492 271856 323544 271862
rect 323492 271798 323544 271804
rect 323584 271856 323636 271862
rect 323584 271798 323636 271804
rect 322848 268660 322900 268666
rect 322848 268602 322900 268608
rect 322664 267776 322716 267782
rect 322664 267718 322716 267724
rect 322848 265464 322900 265470
rect 322848 265406 322900 265412
rect 322414 264302 322612 264330
rect 322860 264316 322888 265406
rect 323596 264330 323624 271798
rect 323242 264302 323624 264330
rect 323688 264316 323716 273566
rect 324228 272740 324280 272746
rect 324228 272682 324280 272688
rect 324240 271250 324268 272682
rect 324700 271522 324728 278052
rect 325056 273828 325108 273834
rect 325056 273770 325108 273776
rect 324688 271516 324740 271522
rect 324688 271458 324740 271464
rect 324228 271244 324280 271250
rect 324228 271186 324280 271192
rect 324596 268184 324648 268190
rect 324596 268126 324648 268132
rect 324136 265532 324188 265538
rect 324136 265474 324188 265480
rect 324148 264316 324176 265474
rect 324608 264316 324636 268126
rect 325068 264316 325096 273770
rect 325516 273760 325568 273766
rect 325516 273702 325568 273708
rect 325528 264316 325556 273702
rect 325896 271658 325924 278052
rect 326344 273692 326396 273698
rect 326344 273634 326396 273640
rect 325884 271652 325936 271658
rect 325884 271594 325936 271600
rect 325976 270972 326028 270978
rect 325976 270914 326028 270920
rect 325792 270904 325844 270910
rect 325792 270846 325844 270852
rect 325700 270836 325752 270842
rect 325700 270778 325752 270784
rect 325712 269006 325740 270778
rect 325700 269000 325752 269006
rect 325700 268942 325752 268948
rect 325804 268258 325832 270846
rect 325792 268252 325844 268258
rect 325792 268194 325844 268200
rect 325988 264316 326016 270914
rect 326356 264316 326384 273634
rect 327092 271590 327120 278052
rect 327724 273964 327776 273970
rect 327724 273906 327776 273912
rect 327080 271584 327132 271590
rect 327080 271526 327132 271532
rect 327264 268252 327316 268258
rect 327264 268194 327316 268200
rect 326804 267980 326856 267986
rect 326804 267922 326856 267928
rect 326816 264316 326844 267922
rect 327276 264316 327304 268194
rect 327736 264316 327764 273906
rect 328288 271726 328316 278052
rect 329012 273896 329064 273902
rect 329012 273838 329064 273844
rect 328276 271720 328328 271726
rect 328276 271662 328328 271668
rect 328644 271040 328696 271046
rect 328644 270982 328696 270988
rect 328184 265600 328236 265606
rect 328184 265542 328236 265548
rect 328196 264316 328224 265542
rect 328656 264316 328684 270982
rect 329024 264316 329052 273838
rect 329484 271794 329512 278052
rect 330392 274100 330444 274106
rect 330392 274042 330444 274048
rect 329472 271788 329524 271794
rect 329472 271730 329524 271736
rect 329472 271108 329524 271114
rect 329472 271050 329524 271056
rect 329484 264316 329512 271050
rect 329932 268932 329984 268938
rect 329932 268874 329984 268880
rect 329944 264316 329972 268874
rect 330404 264316 330432 274042
rect 330588 273222 330616 278052
rect 331680 274032 331732 274038
rect 331680 273974 331732 273980
rect 330852 273556 330904 273562
rect 330852 273498 330904 273504
rect 330576 273216 330628 273222
rect 330576 273158 330628 273164
rect 330864 264316 330892 273498
rect 331312 272196 331364 272202
rect 331312 272138 331364 272144
rect 331324 264316 331352 272138
rect 331692 264316 331720 273974
rect 331784 272270 331812 278052
rect 331772 272264 331824 272270
rect 331772 272206 331824 272212
rect 332324 272128 332376 272134
rect 332324 272070 332376 272076
rect 332232 272060 332284 272066
rect 332232 272002 332284 272008
rect 332140 271992 332192 271998
rect 332140 271934 332192 271940
rect 332152 271318 332180 271934
rect 332244 271386 332272 272002
rect 332336 271454 332364 272070
rect 332324 271448 332376 271454
rect 332324 271390 332376 271396
rect 332232 271380 332284 271386
rect 332232 271322 332284 271328
rect 332140 271312 332192 271318
rect 332140 271254 332192 271260
rect 332980 269210 333008 278052
rect 333060 274168 333112 274174
rect 333060 274110 333112 274116
rect 332968 269204 333020 269210
rect 332968 269146 333020 269152
rect 332600 269068 332652 269074
rect 332600 269010 332652 269016
rect 332140 268388 332192 268394
rect 332140 268330 332192 268336
rect 332152 264316 332180 268330
rect 332612 264316 332640 269010
rect 333072 264316 333100 274110
rect 334176 272610 334204 278052
rect 334348 274304 334400 274310
rect 334348 274246 334400 274252
rect 334164 272604 334216 272610
rect 334164 272546 334216 272552
rect 333980 271244 334032 271250
rect 333980 271186 334032 271192
rect 333152 269272 333204 269278
rect 333152 269214 333204 269220
rect 333164 268802 333192 269214
rect 333152 268796 333204 268802
rect 333152 268738 333204 268744
rect 333520 265668 333572 265674
rect 333520 265610 333572 265616
rect 333532 264316 333560 265610
rect 333992 264316 334020 271186
rect 334360 264316 334388 274246
rect 335372 273154 335400 278052
rect 336096 274372 336148 274378
rect 336096 274314 336148 274320
rect 335360 273148 335412 273154
rect 335360 273090 335412 273096
rect 334808 271176 334860 271182
rect 334808 271118 334860 271124
rect 334820 264316 334848 271118
rect 335268 268524 335320 268530
rect 335268 268466 335320 268472
rect 335280 264316 335308 268466
rect 336108 264330 336136 274314
rect 336568 270502 336596 278052
rect 337108 274440 337160 274446
rect 337108 274382 337160 274388
rect 336648 272604 336700 272610
rect 336648 272546 336700 272552
rect 336556 270496 336608 270502
rect 336556 270438 336608 270444
rect 336464 268320 336516 268326
rect 336464 268262 336516 268268
rect 336476 264330 336504 268262
rect 335754 264302 336136 264330
rect 336214 264302 336504 264330
rect 336660 264316 336688 272546
rect 337120 264316 337148 274382
rect 337764 272882 337792 278052
rect 338396 274508 338448 274514
rect 338396 274450 338448 274456
rect 337752 272876 337804 272882
rect 337752 272818 337804 272824
rect 337476 271312 337528 271318
rect 337476 271254 337528 271260
rect 337488 264316 337516 271254
rect 337936 268592 337988 268598
rect 337936 268534 337988 268540
rect 337948 264316 337976 268534
rect 338408 264316 338436 274450
rect 338868 272814 338896 278052
rect 338856 272808 338908 272814
rect 338856 272750 338908 272756
rect 339224 271380 339276 271386
rect 339224 271322 339276 271328
rect 338856 268456 338908 268462
rect 338856 268398 338908 268404
rect 338868 264316 338896 268398
rect 339236 264330 339264 271322
rect 340064 270434 340092 278052
rect 341064 274576 341116 274582
rect 341064 274518 341116 274524
rect 340052 270428 340104 270434
rect 340052 270370 340104 270376
rect 340604 268728 340656 268734
rect 340604 268670 340656 268676
rect 340144 268660 340196 268666
rect 340144 268602 340196 268608
rect 339776 265736 339828 265742
rect 339776 265678 339828 265684
rect 339236 264302 339342 264330
rect 339788 264316 339816 265678
rect 340156 264316 340184 268602
rect 340616 264316 340644 268670
rect 341076 264316 341104 274518
rect 341260 273086 341288 278052
rect 341248 273080 341300 273086
rect 341248 273022 341300 273028
rect 342168 272808 342220 272814
rect 342168 272750 342220 272756
rect 342076 271448 342128 271454
rect 342076 271390 342128 271396
rect 342088 264974 342116 271390
rect 341904 264946 342116 264974
rect 341904 264330 341932 264946
rect 342180 264330 342208 272750
rect 342456 270638 342484 278052
rect 342536 276004 342588 276010
rect 342536 275946 342588 275952
rect 342444 270632 342496 270638
rect 342444 270574 342496 270580
rect 342548 264330 342576 275946
rect 343652 270298 343680 278052
rect 344192 271516 344244 271522
rect 344192 271458 344244 271464
rect 343640 270292 343692 270298
rect 343640 270234 343692 270240
rect 343272 268116 343324 268122
rect 343272 268058 343324 268064
rect 342812 267776 342864 267782
rect 342812 267718 342864 267724
rect 341550 264302 341932 264330
rect 342010 264302 342208 264330
rect 342470 264302 342576 264330
rect 342824 264316 342852 267718
rect 343284 264316 343312 268058
rect 343732 265804 343784 265810
rect 343732 265746 343784 265752
rect 343744 264316 343772 265746
rect 344204 264316 344232 271458
rect 344848 270366 344876 278052
rect 345112 275936 345164 275942
rect 345112 275878 345164 275884
rect 344928 273148 344980 273154
rect 344928 273090 344980 273096
rect 344836 270360 344888 270366
rect 344836 270302 344888 270308
rect 344940 264330 344968 273090
rect 344678 264302 344968 264330
rect 345124 264316 345152 275878
rect 345952 270774 345980 278052
rect 346400 275800 346452 275806
rect 346400 275742 346452 275748
rect 345940 270768 345992 270774
rect 345940 270710 345992 270716
rect 345480 269000 345532 269006
rect 345480 268942 345532 268948
rect 345492 264316 345520 268942
rect 345940 268864 345992 268870
rect 345940 268806 345992 268812
rect 345952 264316 345980 268806
rect 346412 264316 346440 275742
rect 346860 271584 346912 271590
rect 346860 271526 346912 271532
rect 346872 264316 346900 271526
rect 347148 270230 347176 278052
rect 347780 275868 347832 275874
rect 347780 275810 347832 275816
rect 347504 272876 347556 272882
rect 347504 272818 347556 272824
rect 347136 270224 347188 270230
rect 347136 270166 347188 270172
rect 347516 264330 347544 272818
rect 347346 264302 347544 264330
rect 347792 264316 347820 275810
rect 348344 270162 348372 278052
rect 349540 270706 349568 278052
rect 350172 271720 350224 271726
rect 350172 271662 350224 271668
rect 349620 271652 349672 271658
rect 349620 271594 349672 271600
rect 349528 270700 349580 270706
rect 349528 270642 349580 270648
rect 349068 270428 349120 270434
rect 349068 270370 349120 270376
rect 348608 270224 348660 270230
rect 348608 270166 348660 270172
rect 348332 270156 348384 270162
rect 348332 270098 348384 270104
rect 348240 268796 348292 268802
rect 348240 268738 348292 268744
rect 348148 268388 348200 268394
rect 348148 268330 348200 268336
rect 348160 267918 348188 268330
rect 348148 267912 348200 267918
rect 348148 267854 348200 267860
rect 348252 264316 348280 268738
rect 348620 264316 348648 270166
rect 348792 270156 348844 270162
rect 348792 270098 348844 270104
rect 348804 269958 348832 270098
rect 348792 269952 348844 269958
rect 348792 269894 348844 269900
rect 349080 269822 349108 270370
rect 349068 269816 349120 269822
rect 349068 269758 349120 269764
rect 349068 265872 349120 265878
rect 349068 265814 349120 265820
rect 349080 264316 349108 265814
rect 349632 264330 349660 271594
rect 350184 264330 350212 271662
rect 350736 267238 350764 278052
rect 351564 278038 351946 278066
rect 351276 270496 351328 270502
rect 351276 270438 351328 270444
rect 350908 270360 350960 270366
rect 350908 270302 350960 270308
rect 350724 267232 350776 267238
rect 350724 267174 350776 267180
rect 350264 265940 350316 265946
rect 350264 265882 350316 265888
rect 349554 264302 349660 264330
rect 350014 264302 350212 264330
rect 350276 264330 350304 265882
rect 350276 264302 350474 264330
rect 350920 264316 350948 270302
rect 351288 264316 351316 270438
rect 351564 270026 351592 278038
rect 351644 275732 351696 275738
rect 351644 275674 351696 275680
rect 351552 270020 351604 270026
rect 351552 269962 351604 269968
rect 351656 264330 351684 275674
rect 351920 274304 351972 274310
rect 351748 274252 351920 274258
rect 351748 274246 351972 274252
rect 351748 274230 351960 274246
rect 351748 274174 351776 274230
rect 351736 274168 351788 274174
rect 351736 274110 351788 274116
rect 351828 274168 351880 274174
rect 351828 274110 351880 274116
rect 351840 273562 351868 274110
rect 351828 273556 351880 273562
rect 351828 273498 351880 273504
rect 352656 273216 352708 273222
rect 352656 273158 352708 273164
rect 352196 271788 352248 271794
rect 352196 271730 352248 271736
rect 351920 270224 351972 270230
rect 351920 270166 351972 270172
rect 351932 269890 351960 270166
rect 351920 269884 351972 269890
rect 351920 269826 351972 269832
rect 351828 269680 351880 269686
rect 352012 269680 352064 269686
rect 351880 269628 352012 269634
rect 351828 269622 352064 269628
rect 351840 269606 352052 269622
rect 351736 269068 351788 269074
rect 351736 269010 351788 269016
rect 351748 268394 351776 269010
rect 351920 268932 351972 268938
rect 351920 268874 351972 268880
rect 351736 268388 351788 268394
rect 351736 268330 351788 268336
rect 351932 268326 351960 268874
rect 352104 268864 352156 268870
rect 352104 268806 352156 268812
rect 351828 268320 351880 268326
rect 351828 268262 351880 268268
rect 351920 268320 351972 268326
rect 351920 268262 351972 268268
rect 351840 268122 351868 268262
rect 352116 268138 352144 268806
rect 351736 268116 351788 268122
rect 351736 268058 351788 268064
rect 351828 268116 351880 268122
rect 351828 268058 351880 268064
rect 351932 268110 352144 268138
rect 351748 268002 351776 268058
rect 351932 268002 351960 268110
rect 351748 267974 351960 268002
rect 351656 264302 351762 264330
rect 352208 264316 352236 271730
rect 352472 269612 352524 269618
rect 352472 269554 352524 269560
rect 352484 268802 352512 269554
rect 352472 268796 352524 268802
rect 352472 268738 352524 268744
rect 352564 268796 352616 268802
rect 352564 268738 352616 268744
rect 352576 267782 352604 268738
rect 352564 267776 352616 267782
rect 352564 267718 352616 267724
rect 352668 264316 352696 273158
rect 353128 270094 353156 278052
rect 353208 275664 353260 275670
rect 353208 275606 353260 275612
rect 353116 270088 353168 270094
rect 353116 270030 353168 270036
rect 353220 264330 353248 275606
rect 353576 270224 353628 270230
rect 353576 270166 353628 270172
rect 353142 264302 353248 264330
rect 353588 264316 353616 270166
rect 353944 270088 353996 270094
rect 353944 270030 353996 270036
rect 353956 264316 353984 270030
rect 354232 267170 354260 278052
rect 355322 271144 355378 271153
rect 355322 271079 355378 271088
rect 354864 270836 354916 270842
rect 354864 270778 354916 270784
rect 354220 267164 354272 267170
rect 354220 267106 354272 267112
rect 354404 266008 354456 266014
rect 354404 265950 354456 265956
rect 354416 264316 354444 265950
rect 354876 264316 354904 270778
rect 355336 264316 355364 271079
rect 355428 270162 355456 278052
rect 356060 273080 356112 273086
rect 356060 273022 356112 273028
rect 356072 270434 356100 273022
rect 356624 273018 356652 278052
rect 357072 275596 357124 275602
rect 357072 275538 357124 275544
rect 356612 273012 356664 273018
rect 356612 272954 356664 272960
rect 356060 270428 356112 270434
rect 356060 270370 356112 270376
rect 355416 270156 355468 270162
rect 355416 270098 355468 270104
rect 356244 270088 356296 270094
rect 356244 270030 356296 270036
rect 355784 266076 355836 266082
rect 355784 266018 355836 266024
rect 355796 264316 355824 266018
rect 356256 264316 356284 270030
rect 356610 268696 356666 268705
rect 356610 268631 356666 268640
rect 356624 264316 356652 268631
rect 357084 264316 357112 275538
rect 357530 271280 357586 271289
rect 357530 271215 357586 271224
rect 357544 264316 357572 271215
rect 357820 267102 357848 278052
rect 358832 278038 359030 278066
rect 358452 275528 358504 275534
rect 358452 275470 358504 275476
rect 357990 271416 358046 271425
rect 357990 271351 358046 271360
rect 357808 267096 357860 267102
rect 357808 267038 357860 267044
rect 358004 264316 358032 271351
rect 358464 264316 358492 275470
rect 358832 273086 358860 278038
rect 358820 273080 358872 273086
rect 358820 273022 358872 273028
rect 358912 273080 358964 273086
rect 358912 273022 358964 273028
rect 358924 270842 358952 273022
rect 360212 272950 360240 278052
rect 361120 275460 361172 275466
rect 361120 275402 361172 275408
rect 360568 273012 360620 273018
rect 360568 272954 360620 272960
rect 360200 272944 360252 272950
rect 360200 272886 360252 272892
rect 358912 270836 358964 270842
rect 358912 270778 358964 270784
rect 358912 270428 358964 270434
rect 358912 270370 358964 270376
rect 358924 264316 358952 270370
rect 359370 268832 359426 268841
rect 359370 268767 359426 268776
rect 359384 264316 359412 268767
rect 359740 266144 359792 266150
rect 359740 266086 359792 266092
rect 359752 264316 359780 266086
rect 360580 264330 360608 272954
rect 360658 271552 360714 271561
rect 360658 271487 360714 271496
rect 360226 264302 360608 264330
rect 360672 264316 360700 271487
rect 360844 270768 360896 270774
rect 360844 270710 360896 270716
rect 360856 270026 360884 270710
rect 360844 270020 360896 270026
rect 360844 269962 360896 269968
rect 361132 264316 361160 275402
rect 361408 267034 361436 278052
rect 362512 272746 362540 278052
rect 363144 272944 363196 272950
rect 363144 272886 363196 272892
rect 362500 272740 362552 272746
rect 362500 272682 362552 272688
rect 362592 272740 362644 272746
rect 362592 272682 362644 272688
rect 362604 272474 362632 272682
rect 362592 272468 362644 272474
rect 362592 272410 362644 272416
rect 362868 272468 362920 272474
rect 362868 272410 362920 272416
rect 362880 272202 362908 272410
rect 362868 272196 362920 272202
rect 362868 272138 362920 272144
rect 362868 270496 362920 270502
rect 362868 270438 362920 270444
rect 361580 270020 361632 270026
rect 361580 269962 361632 269968
rect 361396 267028 361448 267034
rect 361396 266970 361448 266976
rect 361592 264316 361620 269962
rect 362880 269890 362908 270438
rect 362868 269884 362920 269890
rect 362868 269826 362920 269832
rect 361672 269612 361724 269618
rect 361672 269554 361724 269560
rect 362868 269612 362920 269618
rect 362868 269554 362920 269560
rect 361684 269074 361712 269554
rect 361672 269068 361724 269074
rect 361672 269010 361724 269016
rect 362038 268968 362094 268977
rect 362038 268903 362094 268912
rect 362052 264316 362080 268903
rect 362880 267918 362908 269554
rect 362868 267912 362920 267918
rect 362868 267854 362920 267860
rect 362408 266212 362460 266218
rect 362408 266154 362460 266160
rect 362420 264316 362448 266154
rect 363156 264330 363184 272886
rect 363326 271688 363382 271697
rect 363326 271623 363382 271632
rect 362894 264302 363184 264330
rect 363340 264316 363368 271623
rect 363708 269754 363736 278052
rect 363788 275392 363840 275398
rect 363788 275334 363840 275340
rect 363696 269748 363748 269754
rect 363696 269690 363748 269696
rect 363800 264316 363828 275334
rect 364340 270564 364392 270570
rect 364340 270506 364392 270512
rect 364246 270464 364302 270473
rect 364246 270399 364302 270408
rect 364260 264316 364288 270399
rect 364352 269958 364380 270506
rect 364340 269952 364392 269958
rect 364340 269894 364392 269900
rect 364708 269952 364760 269958
rect 364708 269894 364760 269900
rect 364720 264316 364748 269894
rect 364904 266966 364932 278052
rect 365994 273184 366050 273193
rect 365994 273119 366050 273128
rect 365534 273048 365590 273057
rect 365534 272983 365590 272992
rect 364892 266960 364944 266966
rect 364892 266902 364944 266908
rect 365076 266280 365128 266286
rect 365076 266222 365128 266228
rect 365088 264316 365116 266222
rect 365548 264316 365576 272983
rect 366008 264316 366036 273119
rect 366100 270706 366128 278052
rect 366456 275324 366508 275330
rect 366456 275266 366508 275272
rect 366088 270700 366140 270706
rect 366088 270642 366140 270648
rect 366468 264316 366496 275266
rect 367296 272542 367324 278052
rect 367284 272536 367336 272542
rect 367284 272478 367336 272484
rect 367100 272196 367152 272202
rect 367100 272138 367152 272144
rect 366914 270328 366970 270337
rect 366914 270263 366970 270272
rect 366928 264316 366956 270263
rect 367112 269686 367140 272138
rect 367376 269884 367428 269890
rect 367376 269826 367428 269832
rect 367100 269680 367152 269686
rect 367100 269622 367152 269628
rect 367388 264316 367416 269826
rect 368204 267912 368256 267918
rect 368204 267854 368256 267860
rect 367744 267708 367796 267714
rect 367744 267650 367796 267656
rect 367756 264316 367784 267650
rect 368216 264316 368244 267854
rect 368492 266898 368520 278052
rect 369124 273488 369176 273494
rect 369124 273430 369176 273436
rect 368662 272912 368718 272921
rect 368662 272847 368718 272856
rect 368480 266892 368532 266898
rect 368480 266834 368532 266840
rect 368676 264316 368704 272847
rect 369136 264316 369164 273430
rect 369596 272678 369624 278052
rect 370792 272746 370820 278052
rect 371792 275256 371844 275262
rect 371792 275198 371844 275204
rect 370870 272776 370926 272785
rect 370780 272740 370832 272746
rect 370870 272711 370926 272720
rect 370780 272682 370832 272688
rect 369584 272672 369636 272678
rect 369584 272614 369636 272620
rect 369676 272672 369728 272678
rect 369676 272614 369728 272620
rect 369582 270192 369638 270201
rect 369582 270127 369638 270136
rect 369596 264316 369624 270127
rect 369688 267918 369716 272614
rect 369860 270700 369912 270706
rect 369860 270642 369912 270648
rect 369676 267912 369728 267918
rect 369676 267854 369728 267860
rect 369872 267850 369900 270642
rect 370044 269816 370096 269822
rect 370044 269758 370096 269764
rect 369860 267844 369912 267850
rect 369860 267786 369912 267792
rect 370056 264316 370084 269758
rect 370504 267640 370556 267646
rect 370504 267582 370556 267588
rect 370516 264316 370544 267582
rect 370884 264316 370912 272711
rect 371330 272640 371386 272649
rect 371330 272575 371386 272584
rect 371344 264316 371372 272575
rect 371804 264316 371832 275198
rect 371988 266830 372016 278052
rect 373184 270774 373212 278052
rect 373998 272504 374054 272513
rect 373998 272439 374054 272448
rect 373172 270768 373224 270774
rect 373172 270710 373224 270716
rect 372250 270056 372306 270065
rect 372250 269991 372306 270000
rect 371976 266824 372028 266830
rect 371976 266766 372028 266772
rect 372264 264316 372292 269991
rect 372712 269748 372764 269754
rect 372712 269690 372764 269696
rect 372724 264316 372752 269690
rect 373172 267572 373224 267578
rect 373172 267514 373224 267520
rect 373184 264316 373212 267514
rect 373540 267504 373592 267510
rect 373540 267446 373592 267452
rect 373552 264316 373580 267446
rect 374012 264316 374040 272439
rect 374380 269482 374408 278052
rect 375590 278038 375788 278066
rect 375288 275188 375340 275194
rect 375288 275130 375340 275136
rect 374368 269476 374420 269482
rect 374368 269418 374420 269424
rect 374460 267436 374512 267442
rect 374460 267378 374512 267384
rect 374472 264316 374500 267378
rect 375300 264330 375328 275130
rect 375656 272740 375708 272746
rect 375656 272682 375708 272688
rect 375564 270768 375616 270774
rect 375564 270710 375616 270716
rect 375380 270632 375432 270638
rect 375380 270574 375432 270580
rect 375392 269550 375420 270574
rect 375472 269680 375524 269686
rect 375472 269622 375524 269628
rect 375380 269544 375432 269550
rect 375380 269486 375432 269492
rect 375484 264330 375512 269622
rect 375576 268054 375604 270710
rect 375668 269414 375696 272682
rect 375656 269408 375708 269414
rect 375656 269350 375708 269356
rect 375564 268048 375616 268054
rect 375564 267990 375616 267996
rect 375760 266762 375788 278038
rect 376772 270910 376800 278052
rect 377772 275120 377824 275126
rect 377772 275062 377824 275068
rect 376760 270904 376812 270910
rect 376760 270846 376812 270852
rect 376668 267844 376720 267850
rect 376668 267786 376720 267792
rect 376208 267368 376260 267374
rect 376208 267310 376260 267316
rect 375840 267300 375892 267306
rect 375840 267242 375892 267248
rect 375748 266756 375800 266762
rect 375748 266698 375800 266704
rect 374946 264302 375328 264330
rect 375406 264302 375512 264330
rect 375852 264316 375880 267242
rect 376220 264316 376248 267310
rect 376680 264316 376708 267786
rect 377128 267232 377180 267238
rect 377128 267174 377180 267180
rect 377140 264316 377168 267174
rect 377784 264330 377812 275062
rect 377876 272338 377904 278052
rect 377864 272332 377916 272338
rect 377864 272274 377916 272280
rect 377864 269544 377916 269550
rect 377864 269486 377916 269492
rect 377614 264302 377812 264330
rect 377876 264330 377904 269486
rect 378508 267164 378560 267170
rect 378508 267106 378560 267112
rect 377876 264302 378074 264330
rect 378520 264316 378548 267106
rect 378876 267096 378928 267102
rect 378876 267038 378928 267044
rect 378888 264316 378916 267038
rect 379072 266694 379100 278052
rect 379336 272536 379388 272542
rect 379336 272478 379388 272484
rect 379060 266688 379112 266694
rect 379060 266630 379112 266636
rect 379348 264316 379376 272478
rect 380268 270570 380296 278052
rect 380348 274984 380400 274990
rect 380348 274926 380400 274932
rect 380256 270564 380308 270570
rect 380256 270506 380308 270512
rect 379796 267028 379848 267034
rect 379796 266970 379848 266976
rect 379808 264316 379836 266970
rect 380360 264330 380388 274926
rect 381464 272746 381492 278052
rect 381452 272740 381504 272746
rect 381452 272682 381504 272688
rect 381360 270836 381412 270842
rect 381360 270778 381412 270784
rect 380714 269920 380770 269929
rect 380714 269855 380770 269864
rect 380282 264302 380388 264330
rect 380728 264316 380756 269855
rect 381372 267986 381400 270778
rect 382004 268048 382056 268054
rect 382004 267990 382056 267996
rect 381360 267980 381412 267986
rect 381360 267922 381412 267928
rect 381636 266960 381688 266966
rect 381636 266902 381688 266908
rect 381176 266892 381228 266898
rect 381176 266834 381228 266840
rect 381188 264316 381216 266834
rect 381648 264316 381676 266902
rect 382016 264316 382044 267990
rect 382464 266824 382516 266830
rect 382464 266766 382516 266772
rect 382476 264316 382504 266766
rect 382660 266626 382688 278052
rect 383292 274916 383344 274922
rect 383292 274858 383344 274864
rect 382648 266620 382700 266626
rect 382648 266562 382700 266568
rect 383304 264330 383332 274858
rect 383856 272406 383884 278052
rect 384960 272474 384988 278052
rect 385590 274136 385646 274145
rect 385590 274071 385646 274080
rect 384948 272468 385000 272474
rect 384948 272410 385000 272416
rect 383844 272400 383896 272406
rect 383844 272342 383896 272348
rect 384672 272400 384724 272406
rect 384672 272342 384724 272348
rect 383382 269784 383438 269793
rect 383382 269719 383438 269728
rect 382950 264302 383332 264330
rect 383396 264316 383424 269719
rect 384304 266756 384356 266762
rect 384304 266698 384356 266704
rect 383844 266688 383896 266694
rect 383844 266630 383896 266636
rect 383856 264316 383884 266630
rect 384316 264316 384344 266698
rect 384684 264316 384712 272342
rect 385132 266620 385184 266626
rect 385132 266562 385184 266568
rect 385144 264316 385172 266562
rect 385604 264316 385632 274071
rect 385684 270904 385736 270910
rect 385684 270846 385736 270852
rect 385696 269618 385724 270846
rect 385684 269612 385736 269618
rect 385684 269554 385736 269560
rect 386052 269408 386104 269414
rect 386052 269350 386104 269356
rect 386064 264316 386092 269350
rect 386156 266558 386184 278052
rect 386420 272468 386472 272474
rect 386420 272410 386472 272416
rect 386432 268054 386460 272410
rect 387352 272202 387380 278052
rect 388258 274272 388314 274281
rect 388258 274207 388314 274216
rect 387430 272368 387486 272377
rect 387430 272303 387486 272312
rect 387340 272196 387392 272202
rect 387340 272138 387392 272144
rect 386420 268048 386472 268054
rect 386420 267990 386472 267996
rect 386970 267064 387026 267073
rect 386970 266999 387026 267008
rect 386144 266552 386196 266558
rect 386144 266494 386196 266500
rect 386512 266552 386564 266558
rect 386512 266494 386564 266500
rect 386524 264316 386552 266494
rect 386880 266348 386932 266354
rect 386880 266290 386932 266296
rect 386892 265266 386920 266290
rect 386880 265260 386932 265266
rect 386880 265202 386932 265208
rect 386984 264316 387012 266999
rect 387444 264330 387472 272303
rect 387798 267200 387854 267209
rect 387798 267135 387854 267144
rect 387366 264302 387472 264330
rect 387812 264316 387840 267135
rect 388272 264316 388300 274207
rect 388548 269346 388576 278052
rect 388536 269340 388588 269346
rect 388536 269282 388588 269288
rect 388720 269340 388772 269346
rect 388720 269282 388772 269288
rect 388732 264316 388760 269282
rect 389638 266928 389694 266937
rect 389638 266863 389694 266872
rect 389180 266484 389232 266490
rect 389180 266426 389232 266432
rect 389192 264316 389220 266426
rect 389652 264316 389680 266863
rect 389744 265198 389772 278052
rect 390652 275256 390704 275262
rect 390652 275198 390704 275204
rect 390468 274780 390520 274786
rect 390468 274722 390520 274728
rect 390480 273562 390508 274722
rect 390468 273556 390520 273562
rect 390468 273498 390520 273504
rect 390664 273494 390692 275198
rect 390652 273488 390704 273494
rect 390652 273430 390704 273436
rect 390008 272332 390060 272338
rect 390008 272274 390060 272280
rect 389732 265192 389784 265198
rect 389732 265134 389784 265140
rect 390020 264316 390048 272274
rect 390940 272134 390968 278052
rect 391018 274408 391074 274417
rect 391018 274343 391074 274352
rect 390928 272128 390980 272134
rect 390928 272070 390980 272076
rect 390466 266792 390522 266801
rect 390466 266727 390522 266736
rect 390480 264316 390508 266727
rect 391032 264330 391060 274343
rect 391940 272740 391992 272746
rect 391940 272682 391992 272688
rect 391388 269408 391440 269414
rect 391388 269350 391440 269356
rect 390954 264302 391060 264330
rect 391400 264316 391428 269350
rect 391952 267850 391980 272682
rect 392136 272066 392164 278052
rect 392768 272196 392820 272202
rect 392768 272138 392820 272144
rect 392124 272060 392176 272066
rect 392124 272002 392176 272008
rect 391940 267844 391992 267850
rect 391940 267786 391992 267792
rect 391846 266656 391902 266665
rect 391846 266591 391902 266600
rect 391860 264316 391888 266591
rect 392308 266416 392360 266422
rect 392308 266358 392360 266364
rect 392320 264316 392348 266358
rect 392780 264316 392808 272138
rect 393134 266520 393190 266529
rect 393134 266455 393190 266464
rect 393148 264316 393176 266455
rect 393240 266354 393268 278052
rect 394436 270638 394464 278052
rect 394974 275904 395030 275913
rect 394974 275839 395030 275848
rect 394424 270632 394476 270638
rect 394424 270574 394476 270580
rect 394056 269340 394108 269346
rect 394056 269282 394108 269288
rect 393594 267336 393650 267345
rect 393594 267271 393650 267280
rect 393228 266348 393280 266354
rect 393228 266290 393280 266296
rect 393608 264316 393636 267271
rect 394068 264316 394096 269282
rect 394514 266384 394570 266393
rect 394514 266319 394570 266328
rect 394528 264316 394556 266319
rect 394988 264316 395016 275839
rect 395434 272232 395490 272241
rect 395434 272167 395490 272176
rect 395448 264316 395476 272167
rect 395632 269278 395660 278052
rect 395620 269272 395672 269278
rect 395620 269214 395672 269220
rect 396724 269272 396776 269278
rect 396724 269214 396776 269220
rect 396262 267472 396318 267481
rect 396262 267407 396318 267416
rect 395804 266348 395856 266354
rect 395804 266290 395856 266296
rect 395816 264316 395844 266290
rect 396276 264316 396304 267407
rect 396736 264316 396764 269214
rect 396828 265266 396856 278052
rect 397366 275768 397422 275777
rect 397366 275703 397422 275712
rect 396816 265260 396868 265266
rect 396816 265202 396868 265208
rect 397380 264330 397408 275703
rect 398024 274854 398052 278052
rect 398470 275632 398526 275641
rect 398470 275567 398526 275576
rect 398012 274848 398064 274854
rect 398012 274790 398064 274796
rect 397644 274780 397696 274786
rect 397644 274722 397696 274728
rect 397210 264302 397408 264330
rect 397656 264316 397684 274722
rect 398104 272128 398156 272134
rect 398104 272070 398156 272076
rect 398116 264316 398144 272070
rect 398484 264316 398512 275567
rect 399220 271998 399248 278052
rect 399850 275224 399906 275233
rect 399850 275159 399906 275168
rect 399208 271992 399260 271998
rect 399208 271934 399260 271940
rect 399390 269648 399446 269657
rect 399390 269583 399446 269592
rect 398930 267608 398986 267617
rect 398930 267543 398986 267552
rect 398944 264316 398972 267543
rect 399404 264316 399432 269583
rect 399864 264316 399892 275159
rect 400324 265334 400352 278052
rect 400402 275496 400458 275505
rect 400402 275431 400458 275440
rect 400312 265328 400364 265334
rect 400312 265270 400364 265276
rect 400416 264330 400444 275431
rect 401138 275360 401194 275369
rect 401138 275295 401194 275304
rect 400772 270632 400824 270638
rect 400772 270574 400824 270580
rect 400338 264302 400444 264330
rect 400784 264316 400812 270574
rect 401152 264316 401180 275295
rect 401520 270706 401548 278052
rect 402610 275088 402666 275097
rect 402610 275023 402666 275032
rect 401508 270700 401560 270706
rect 401508 270642 401560 270648
rect 402060 269204 402112 269210
rect 402060 269146 402112 269152
rect 401324 269136 401376 269142
rect 401324 269078 401376 269084
rect 401336 268190 401364 269078
rect 401324 268184 401376 268190
rect 401324 268126 401376 268132
rect 401600 265328 401652 265334
rect 401600 265270 401652 265276
rect 401612 264316 401640 265270
rect 402072 264316 402100 269146
rect 402624 264330 402652 275023
rect 402716 269142 402744 278052
rect 402980 274780 403032 274786
rect 402980 274722 403032 274728
rect 402704 269136 402756 269142
rect 402704 269078 402756 269084
rect 402546 264302 402652 264330
rect 402992 264316 403020 274722
rect 403438 272096 403494 272105
rect 403438 272031 403494 272040
rect 403452 264316 403480 272031
rect 403912 265402 403940 278052
rect 403990 274952 404046 274961
rect 403990 274887 404046 274896
rect 403900 265396 403952 265402
rect 403900 265338 403952 265344
rect 404004 264330 404032 274887
rect 405108 273562 405136 278052
rect 405186 274816 405242 274825
rect 405186 274751 405242 274760
rect 405096 273556 405148 273562
rect 405096 273498 405148 273504
rect 404726 269512 404782 269521
rect 404726 269447 404782 269456
rect 404268 265396 404320 265402
rect 404268 265338 404320 265344
rect 403926 264302 404032 264330
rect 404280 264316 404308 265338
rect 404740 264316 404768 269447
rect 405200 264316 405228 274751
rect 406108 272060 406160 272066
rect 406108 272002 406160 272008
rect 405462 267744 405518 267753
rect 405462 267679 405518 267688
rect 405476 264330 405504 267679
rect 405476 264302 405674 264330
rect 406120 264316 406148 272002
rect 406304 271930 406332 278052
rect 407500 274718 407528 278052
rect 407488 274712 407540 274718
rect 406934 274680 406990 274689
rect 407488 274654 407540 274660
rect 406934 274615 406990 274624
rect 406568 273556 406620 273562
rect 406568 273498 406620 273504
rect 406292 271924 406344 271930
rect 406292 271866 406344 271872
rect 406580 264316 406608 273498
rect 406948 264316 406976 274615
rect 408130 274544 408186 274553
rect 408130 274479 408186 274488
rect 407394 269376 407450 269385
rect 407394 269311 407450 269320
rect 407408 264316 407436 269311
rect 408144 264330 408172 274479
rect 408604 270774 408632 278052
rect 409236 274712 409288 274718
rect 409236 274654 409288 274660
rect 408774 271960 408830 271969
rect 408774 271895 408830 271904
rect 408592 270768 408644 270774
rect 408592 270710 408644 270716
rect 408314 266248 408370 266257
rect 408314 266183 408370 266192
rect 407882 264302 408172 264330
rect 408328 264316 408356 266183
rect 408788 264316 408816 271895
rect 409248 264316 409276 274654
rect 409604 271992 409656 271998
rect 409604 271934 409656 271940
rect 409616 264316 409644 271934
rect 409800 268190 409828 278052
rect 410996 274650 411024 278052
rect 410984 274644 411036 274650
rect 410984 274586 411036 274592
rect 411444 271924 411496 271930
rect 411444 271866 411496 271872
rect 410522 271824 410578 271833
rect 410522 271759 410578 271768
rect 410064 269136 410116 269142
rect 410064 269078 410116 269084
rect 409788 268184 409840 268190
rect 409788 268126 409840 268132
rect 410076 264316 410104 269078
rect 410536 264316 410564 271759
rect 410798 269240 410854 269249
rect 410798 269175 410854 269184
rect 410812 264330 410840 269175
rect 410812 264302 411010 264330
rect 411456 264316 411484 271866
rect 411902 269104 411958 269113
rect 411902 269039 411958 269048
rect 411916 264316 411944 269039
rect 412192 265470 412220 278052
rect 413388 271862 413416 278052
rect 414584 273630 414612 278052
rect 414572 273624 414624 273630
rect 414572 273566 414624 273572
rect 413836 272060 413888 272066
rect 413836 272002 413888 272008
rect 413376 271856 413428 271862
rect 413376 271798 413428 271804
rect 413848 270638 413876 272002
rect 413836 270632 413888 270638
rect 413836 270574 413888 270580
rect 415780 265538 415808 278052
rect 416884 268054 416912 278052
rect 418080 273834 418108 278052
rect 418068 273828 418120 273834
rect 418068 273770 418120 273776
rect 419276 273766 419304 278052
rect 419264 273760 419316 273766
rect 419264 273702 419316 273708
rect 420472 270978 420500 278052
rect 421668 273698 421696 278052
rect 421656 273692 421708 273698
rect 421656 273634 421708 273640
rect 420460 270972 420512 270978
rect 420460 270914 420512 270920
rect 420828 270972 420880 270978
rect 420828 270914 420880 270920
rect 420840 268122 420868 270914
rect 422864 270842 422892 278052
rect 422852 270836 422904 270842
rect 422852 270778 422904 270784
rect 423968 268258 423996 278052
rect 425164 273970 425192 278052
rect 425152 273964 425204 273970
rect 425152 273906 425204 273912
rect 423956 268252 424008 268258
rect 423956 268194 424008 268200
rect 420828 268116 420880 268122
rect 420828 268058 420880 268064
rect 416872 268048 416924 268054
rect 416872 267990 416924 267996
rect 426360 265606 426388 278052
rect 427556 271046 427584 278052
rect 428752 273902 428780 278052
rect 429108 274712 429160 274718
rect 429108 274654 429160 274660
rect 428740 273896 428792 273902
rect 428740 273838 428792 273844
rect 429120 273562 429148 274654
rect 429108 273556 429160 273562
rect 429108 273498 429160 273504
rect 429948 271114 429976 278052
rect 429936 271108 429988 271114
rect 429936 271050 429988 271056
rect 427544 271040 427596 271046
rect 427544 270982 427596 270988
rect 431144 268326 431172 278052
rect 432248 274038 432276 278052
rect 433444 274106 433472 278052
rect 433432 274100 433484 274106
rect 433432 274042 433484 274048
rect 432236 274032 432288 274038
rect 432236 273974 432288 273980
rect 434640 272270 434668 278052
rect 435836 273970 435864 278052
rect 435824 273964 435876 273970
rect 435824 273906 435876 273912
rect 434628 272264 434680 272270
rect 434628 272206 434680 272212
rect 436100 272264 436152 272270
rect 436100 272206 436152 272212
rect 431132 268320 431184 268326
rect 431132 268262 431184 268268
rect 436112 266257 436140 272206
rect 437032 270910 437060 278052
rect 437020 270904 437072 270910
rect 437020 270846 437072 270852
rect 438228 268394 438256 278052
rect 439332 274310 439360 278052
rect 439320 274304 439372 274310
rect 439320 274246 439372 274252
rect 438216 268388 438268 268394
rect 438216 268330 438268 268336
rect 436098 266248 436154 266257
rect 436098 266183 436154 266192
rect 440528 265674 440556 278052
rect 441724 271250 441752 278052
rect 442920 274174 442948 278052
rect 442908 274168 442960 274174
rect 442908 274110 442960 274116
rect 441712 271244 441764 271250
rect 441712 271186 441764 271192
rect 444116 271182 444144 278052
rect 444104 271176 444156 271182
rect 444104 271118 444156 271124
rect 442540 271108 442592 271114
rect 442540 271050 442592 271056
rect 442552 268462 442580 271050
rect 445312 268530 445340 278052
rect 446508 274378 446536 278052
rect 446496 274372 446548 274378
rect 446496 274314 446548 274320
rect 447612 270978 447640 278052
rect 448808 272610 448836 278052
rect 450004 274446 450032 278052
rect 449992 274440 450044 274446
rect 449992 274382 450044 274388
rect 448796 272604 448848 272610
rect 448796 272546 448848 272552
rect 448888 272604 448940 272610
rect 448888 272546 448940 272552
rect 447600 270972 447652 270978
rect 447600 270914 447652 270920
rect 445300 268524 445352 268530
rect 445300 268466 445352 268472
rect 442540 268456 442592 268462
rect 442540 268398 442592 268404
rect 440516 265668 440568 265674
rect 440516 265610 440568 265616
rect 426348 265600 426400 265606
rect 426348 265542 426400 265548
rect 415768 265532 415820 265538
rect 415768 265474 415820 265480
rect 412180 265464 412232 265470
rect 412180 265406 412232 265412
rect 448900 265402 448928 272546
rect 451200 271182 451228 278052
rect 451188 271176 451240 271182
rect 451188 271118 451240 271124
rect 452396 268598 452424 278052
rect 453592 274514 453620 278052
rect 453580 274508 453632 274514
rect 453580 274450 453632 274456
rect 452660 271448 452712 271454
rect 452660 271390 452712 271396
rect 452672 268666 452700 271390
rect 454696 271114 454724 278052
rect 455892 271250 455920 278052
rect 455880 271244 455932 271250
rect 455880 271186 455932 271192
rect 454684 271108 454736 271114
rect 454684 271050 454736 271056
rect 452660 268660 452712 268666
rect 452660 268602 452712 268608
rect 452384 268592 452436 268598
rect 452384 268534 452436 268540
rect 457088 265742 457116 278052
rect 458284 271454 458312 278052
rect 458272 271448 458324 271454
rect 458272 271390 458324 271396
rect 459480 268734 459508 278052
rect 460676 274582 460704 278052
rect 460664 274576 460716 274582
rect 460664 274518 460716 274524
rect 461872 271318 461900 278052
rect 462976 272814 463004 278052
rect 464172 276010 464200 278052
rect 464160 276004 464212 276010
rect 464160 275946 464212 275952
rect 462964 272808 463016 272814
rect 462964 272750 463016 272756
rect 463332 272808 463384 272814
rect 463332 272750 463384 272756
rect 461860 271312 461912 271318
rect 461860 271254 461912 271260
rect 459468 268728 459520 268734
rect 459468 268670 459520 268676
rect 457076 265736 457128 265742
rect 457076 265678 457128 265684
rect 448888 265396 448940 265402
rect 448888 265338 448940 265344
rect 463344 265334 463372 272750
rect 465368 268802 465396 278052
rect 466564 268870 466592 278052
rect 466552 268864 466604 268870
rect 466552 268806 466604 268812
rect 465356 268796 465408 268802
rect 465356 268738 465408 268744
rect 467760 265810 467788 278052
rect 468956 271522 468984 278052
rect 470152 273154 470180 278052
rect 471256 275942 471284 278052
rect 471244 275936 471296 275942
rect 471244 275878 471296 275884
rect 470140 273148 470192 273154
rect 470140 273090 470192 273096
rect 471980 273148 472032 273154
rect 471980 273090 472032 273096
rect 468944 271516 468996 271522
rect 468944 271458 468996 271464
rect 471992 267617 472020 273090
rect 472452 269006 472480 278052
rect 472440 269000 472492 269006
rect 472440 268942 472492 268948
rect 473648 268938 473676 278052
rect 474844 275806 474872 278052
rect 474832 275800 474884 275806
rect 474832 275742 474884 275748
rect 476040 271590 476068 278052
rect 477236 272882 477264 278052
rect 478340 275874 478368 278052
rect 478328 275868 478380 275874
rect 478328 275810 478380 275816
rect 477224 272876 477276 272882
rect 477224 272818 477276 272824
rect 477316 272876 477368 272882
rect 477316 272818 477368 272824
rect 476028 271584 476080 271590
rect 476028 271526 476080 271532
rect 473636 268932 473688 268938
rect 473636 268874 473688 268880
rect 477328 267753 477356 272818
rect 479536 269074 479564 278052
rect 480732 270502 480760 278052
rect 480720 270496 480772 270502
rect 480720 270438 480772 270444
rect 479524 269068 479576 269074
rect 479524 269010 479576 269016
rect 477314 267744 477370 267753
rect 477314 267679 477370 267688
rect 471978 267608 472034 267617
rect 471978 267543 472034 267552
rect 481928 265878 481956 278052
rect 483124 271658 483152 278052
rect 484320 271726 484348 278052
rect 484308 271720 484360 271726
rect 484308 271662 484360 271668
rect 483112 271652 483164 271658
rect 483112 271594 483164 271600
rect 485516 265946 485544 278052
rect 485688 271720 485740 271726
rect 485688 271662 485740 271668
rect 485700 267481 485728 271662
rect 486620 270298 486648 278052
rect 487816 270366 487844 278052
rect 489012 275738 489040 278052
rect 489000 275732 489052 275738
rect 489000 275674 489052 275680
rect 490208 271794 490236 278052
rect 491404 273222 491432 278052
rect 492600 275670 492628 278052
rect 492588 275664 492640 275670
rect 492588 275606 492640 275612
rect 491392 273216 491444 273222
rect 491392 273158 491444 273164
rect 491484 273216 491536 273222
rect 491484 273158 491536 273164
rect 490196 271788 490248 271794
rect 490196 271730 490248 271736
rect 491496 270434 491524 273158
rect 491484 270428 491536 270434
rect 491484 270370 491536 270376
rect 487804 270360 487856 270366
rect 487804 270302 487856 270308
rect 486608 270292 486660 270298
rect 486608 270234 486660 270240
rect 493704 270230 493732 278052
rect 493692 270224 493744 270230
rect 493692 270166 493744 270172
rect 494900 270162 494928 278052
rect 494888 270156 494940 270162
rect 494888 270098 494940 270104
rect 485686 267472 485742 267481
rect 485686 267407 485742 267416
rect 496096 266014 496124 278052
rect 497292 273086 497320 278052
rect 497280 273080 497332 273086
rect 497280 273022 497332 273028
rect 497924 273080 497976 273086
rect 497924 273022 497976 273028
rect 497936 267345 497964 273022
rect 498488 271153 498516 278052
rect 498474 271144 498530 271153
rect 498474 271079 498530 271088
rect 497922 267336 497978 267345
rect 497922 267271 497978 267280
rect 499684 266082 499712 278052
rect 500880 270094 500908 278052
rect 500868 270088 500920 270094
rect 500868 270030 500920 270036
rect 501984 268705 502012 278052
rect 503180 275602 503208 278052
rect 503168 275596 503220 275602
rect 503168 275538 503220 275544
rect 504376 271289 504404 278052
rect 505572 271425 505600 278052
rect 506768 275534 506796 278052
rect 506756 275528 506808 275534
rect 506756 275470 506808 275476
rect 507964 273222 507992 278052
rect 507952 273216 508004 273222
rect 507952 273158 508004 273164
rect 505558 271416 505614 271425
rect 505558 271351 505614 271360
rect 504362 271280 504418 271289
rect 504362 271215 504418 271224
rect 509068 268841 509096 278052
rect 509054 268832 509110 268841
rect 509054 268767 509110 268776
rect 501970 268696 502026 268705
rect 501970 268631 502026 268640
rect 510264 266150 510292 278052
rect 511460 273018 511488 278052
rect 511448 273012 511500 273018
rect 511448 272954 511500 272960
rect 512656 271561 512684 278052
rect 513852 275466 513880 278052
rect 513840 275460 513892 275466
rect 513840 275402 513892 275408
rect 512642 271552 512698 271561
rect 512642 271487 512698 271496
rect 515048 270026 515076 278052
rect 515036 270020 515088 270026
rect 515036 269962 515088 269968
rect 516244 268977 516272 278052
rect 516230 268968 516286 268977
rect 516230 268903 516286 268912
rect 517348 266218 517376 278052
rect 518544 272950 518572 278052
rect 518532 272944 518584 272950
rect 518532 272886 518584 272892
rect 519740 271697 519768 278052
rect 520936 275398 520964 278052
rect 520924 275392 520976 275398
rect 520924 275334 520976 275340
rect 519726 271688 519782 271697
rect 519726 271623 519782 271632
rect 522132 270473 522160 278052
rect 522118 270464 522174 270473
rect 522118 270399 522174 270408
rect 523328 269958 523356 278052
rect 523316 269952 523368 269958
rect 523316 269894 523368 269900
rect 524524 266286 524552 278052
rect 525628 273057 525656 278052
rect 526824 273193 526852 278052
rect 528020 275330 528048 278052
rect 528008 275324 528060 275330
rect 528008 275266 528060 275272
rect 526810 273184 526866 273193
rect 526810 273119 526866 273128
rect 525614 273048 525670 273057
rect 525614 272983 525670 272992
rect 529216 270337 529244 278052
rect 529202 270328 529258 270337
rect 529202 270263 529258 270272
rect 530412 269890 530440 278052
rect 530400 269884 530452 269890
rect 530400 269826 530452 269832
rect 531608 267714 531636 278052
rect 532712 272678 532740 278052
rect 533908 272921 533936 278052
rect 535104 275262 535132 278052
rect 535092 275256 535144 275262
rect 535092 275198 535144 275204
rect 533894 272912 533950 272921
rect 533894 272847 533950 272856
rect 532700 272672 532752 272678
rect 532700 272614 532752 272620
rect 536300 270201 536328 278052
rect 536286 270192 536342 270201
rect 536286 270127 536342 270136
rect 537496 269822 537524 278052
rect 537484 269816 537536 269822
rect 537484 269758 537536 269764
rect 531596 267708 531648 267714
rect 531596 267650 531648 267656
rect 538692 267646 538720 278052
rect 539888 272785 539916 278052
rect 539874 272776 539930 272785
rect 539874 272711 539930 272720
rect 540992 272649 541020 278052
rect 542188 275194 542216 278052
rect 542176 275188 542228 275194
rect 542176 275130 542228 275136
rect 540978 272640 541034 272649
rect 540978 272575 541034 272584
rect 543384 270065 543412 278052
rect 543370 270056 543426 270065
rect 543370 269991 543426 270000
rect 544580 269754 544608 278052
rect 544568 269748 544620 269754
rect 544568 269690 544620 269696
rect 538680 267640 538732 267646
rect 538680 267582 538732 267588
rect 545776 267578 545804 278052
rect 545764 267572 545816 267578
rect 545764 267514 545816 267520
rect 546972 267510 547000 278052
rect 548076 272513 548104 278052
rect 548062 272504 548118 272513
rect 548062 272439 548118 272448
rect 546960 267504 547012 267510
rect 546960 267446 547012 267452
rect 549272 267442 549300 278052
rect 550468 275126 550496 278052
rect 550456 275120 550508 275126
rect 550456 275062 550508 275068
rect 551664 269686 551692 278052
rect 551652 269680 551704 269686
rect 551652 269622 551704 269628
rect 549260 267436 549312 267442
rect 549260 267378 549312 267384
rect 552860 267306 552888 278052
rect 554056 267374 554084 278052
rect 555252 272746 555280 278052
rect 555240 272740 555292 272746
rect 555240 272682 555292 272688
rect 554044 267368 554096 267374
rect 554044 267310 554096 267316
rect 552848 267300 552900 267306
rect 552848 267242 552900 267248
rect 556356 267238 556384 278052
rect 557552 275058 557580 278052
rect 557540 275052 557592 275058
rect 557540 274994 557592 275000
rect 558748 269618 558776 278052
rect 558736 269612 558788 269618
rect 558736 269554 558788 269560
rect 556344 267232 556396 267238
rect 556344 267174 556396 267180
rect 559944 267170 559972 278052
rect 559932 267164 559984 267170
rect 559932 267106 559984 267112
rect 561140 267102 561168 278052
rect 562336 272542 562364 278052
rect 562324 272536 562376 272542
rect 562324 272478 562376 272484
rect 561128 267096 561180 267102
rect 561128 267038 561180 267044
rect 563440 267034 563468 278052
rect 564636 274990 564664 278052
rect 564624 274984 564676 274990
rect 564624 274926 564676 274932
rect 565832 269929 565860 278052
rect 565818 269920 565874 269929
rect 565818 269855 565874 269864
rect 563428 267028 563480 267034
rect 563428 266970 563480 266976
rect 567028 266898 567056 278052
rect 568224 266966 568252 278052
rect 569420 272474 569448 278052
rect 569408 272468 569460 272474
rect 569408 272410 569460 272416
rect 568212 266960 568264 266966
rect 568212 266902 568264 266908
rect 567016 266892 567068 266898
rect 567016 266834 567068 266840
rect 570616 266830 570644 278052
rect 571720 274922 571748 278052
rect 571708 274916 571760 274922
rect 571708 274858 571760 274864
rect 572916 269793 572944 278052
rect 572902 269784 572958 269793
rect 572902 269719 572958 269728
rect 570604 266824 570656 266830
rect 570604 266766 570656 266772
rect 574112 266694 574140 278052
rect 575308 266762 575336 278052
rect 576504 272406 576532 278052
rect 576492 272400 576544 272406
rect 576492 272342 576544 272348
rect 575296 266756 575348 266762
rect 575296 266698 575348 266704
rect 574100 266688 574152 266694
rect 574100 266630 574152 266636
rect 577700 266626 577728 278052
rect 578896 274145 578924 278052
rect 578882 274136 578938 274145
rect 578882 274071 578938 274080
rect 580000 269550 580028 278052
rect 579988 269544 580040 269550
rect 579988 269486 580040 269492
rect 577688 266620 577740 266626
rect 577688 266562 577740 266568
rect 581196 266558 581224 278052
rect 582392 267073 582420 278052
rect 583588 272377 583616 278052
rect 583574 272368 583630 272377
rect 583574 272303 583630 272312
rect 584784 267209 584812 278052
rect 585980 274281 586008 278052
rect 585966 274272 586022 274281
rect 585966 274207 586022 274216
rect 587084 269482 587112 278052
rect 587072 269476 587124 269482
rect 587072 269418 587124 269424
rect 584770 267200 584826 267209
rect 584770 267135 584826 267144
rect 582378 267064 582434 267073
rect 582378 266999 582434 267008
rect 581184 266552 581236 266558
rect 581184 266494 581236 266500
rect 588280 266490 588308 278052
rect 589476 266937 589504 278052
rect 590672 272338 590700 278052
rect 590660 272332 590712 272338
rect 590660 272274 590712 272280
rect 589462 266928 589518 266937
rect 589462 266863 589518 266872
rect 591868 266801 591896 278052
rect 593064 274417 593092 278052
rect 593050 274408 593106 274417
rect 593050 274343 593106 274352
rect 594260 269414 594288 278052
rect 594248 269408 594300 269414
rect 594248 269350 594300 269356
rect 591854 266792 591910 266801
rect 591854 266727 591910 266736
rect 595364 266665 595392 278052
rect 595350 266656 595406 266665
rect 595350 266591 595406 266600
rect 588268 266484 588320 266490
rect 588268 266426 588320 266432
rect 596560 266422 596588 278052
rect 597756 272202 597784 278052
rect 597744 272196 597796 272202
rect 597744 272138 597796 272144
rect 598952 266529 598980 278052
rect 600148 273086 600176 278052
rect 600136 273080 600188 273086
rect 600136 273022 600188 273028
rect 601344 269346 601372 278052
rect 601332 269340 601384 269346
rect 601332 269282 601384 269288
rect 598938 266520 598994 266529
rect 598938 266455 598994 266464
rect 596548 266416 596600 266422
rect 602448 266393 602476 278052
rect 603644 275913 603672 278052
rect 603630 275904 603686 275913
rect 603630 275839 603686 275848
rect 604840 272241 604868 278052
rect 604826 272232 604882 272241
rect 604826 272167 604882 272176
rect 596548 266358 596600 266364
rect 602434 266384 602490 266393
rect 606036 266354 606064 278052
rect 607232 271726 607260 278052
rect 607220 271720 607272 271726
rect 607220 271662 607272 271668
rect 608428 269278 608456 278052
rect 609624 275777 609652 278052
rect 609610 275768 609666 275777
rect 609610 275703 609666 275712
rect 610728 274854 610756 278052
rect 610716 274848 610768 274854
rect 610716 274790 610768 274796
rect 611924 272134 611952 278052
rect 613120 275641 613148 278052
rect 613106 275632 613162 275641
rect 613106 275567 613162 275576
rect 614316 273154 614344 278052
rect 614304 273148 614356 273154
rect 614304 273090 614356 273096
rect 611912 272128 611964 272134
rect 611912 272070 611964 272076
rect 615512 269657 615540 278052
rect 616708 275233 616736 278052
rect 617812 275505 617840 278052
rect 617798 275496 617854 275505
rect 617798 275431 617854 275440
rect 616694 275224 616750 275233
rect 616694 275159 616750 275168
rect 619008 272066 619036 278052
rect 620204 275369 620232 278052
rect 620190 275360 620246 275369
rect 620190 275295 620246 275304
rect 621400 272814 621428 278052
rect 621388 272808 621440 272814
rect 621388 272750 621440 272756
rect 618996 272060 619048 272066
rect 618996 272002 619048 272008
rect 615498 269648 615554 269657
rect 615498 269583 615554 269592
rect 608416 269272 608468 269278
rect 608416 269214 608468 269220
rect 622596 269210 622624 278052
rect 623792 275097 623820 278052
rect 623778 275088 623834 275097
rect 623778 275023 623834 275032
rect 624988 274786 625016 278052
rect 624976 274780 625028 274786
rect 624976 274722 625028 274728
rect 626092 272105 626120 278052
rect 627288 274961 627316 278052
rect 627274 274952 627330 274961
rect 627274 274887 627330 274896
rect 628484 272610 628512 278052
rect 628472 272604 628524 272610
rect 628472 272546 628524 272552
rect 626078 272096 626134 272105
rect 626078 272031 626134 272040
rect 629680 269521 629708 278052
rect 630876 274825 630904 278052
rect 630862 274816 630918 274825
rect 630862 274751 630918 274760
rect 632072 272882 632100 278052
rect 632060 272876 632112 272882
rect 632060 272818 632112 272824
rect 633268 271998 633296 278052
rect 634372 274718 634400 278052
rect 634360 274712 634412 274718
rect 635568 274689 635596 278052
rect 634360 274654 634412 274660
rect 635554 274680 635610 274689
rect 635554 274615 635610 274624
rect 633256 271992 633308 271998
rect 633256 271934 633308 271940
rect 629666 269512 629722 269521
rect 629666 269447 629722 269456
rect 636764 269385 636792 278052
rect 637960 274553 637988 278052
rect 637946 274544 638002 274553
rect 637946 274479 638002 274488
rect 639156 272270 639184 278052
rect 639144 272264 639196 272270
rect 639144 272206 639196 272212
rect 640352 271969 640380 278052
rect 641456 274650 641484 278052
rect 641444 274644 641496 274650
rect 641444 274586 641496 274592
rect 640338 271960 640394 271969
rect 642652 271930 642680 278052
rect 640338 271895 640394 271904
rect 642640 271924 642692 271930
rect 642640 271866 642692 271872
rect 636750 269376 636806 269385
rect 636750 269311 636806 269320
rect 622584 269204 622636 269210
rect 622584 269146 622636 269152
rect 643848 269142 643876 278052
rect 645044 271833 645072 278052
rect 645030 271824 645086 271833
rect 645030 271759 645086 271768
rect 646240 269249 646268 278052
rect 647436 271862 647464 278052
rect 647424 271856 647476 271862
rect 647424 271798 647476 271804
rect 646226 269240 646282 269249
rect 646226 269175 646282 269184
rect 643836 269136 643888 269142
rect 648632 269113 648660 278052
rect 643836 269078 643888 269084
rect 648618 269104 648674 269113
rect 648618 269039 648674 269048
rect 602434 266319 602490 266328
rect 606024 266348 606076 266354
rect 606024 266290 606076 266296
rect 524512 266280 524564 266286
rect 524512 266222 524564 266228
rect 517336 266212 517388 266218
rect 517336 266154 517388 266160
rect 510252 266144 510304 266150
rect 510252 266086 510304 266092
rect 499672 266076 499724 266082
rect 499672 266018 499724 266024
rect 496084 266008 496136 266014
rect 496084 265950 496136 265956
rect 485504 265940 485556 265946
rect 485504 265882 485556 265888
rect 481916 265872 481968 265878
rect 481916 265814 481968 265820
rect 467748 265804 467800 265810
rect 467748 265746 467800 265752
rect 463332 265328 463384 265334
rect 463332 265270 463384 265276
rect 573060 262329 573088 262338
rect 573044 262320 573104 262329
rect 573044 262251 573104 262260
rect 572234 259193 572262 259198
rect 572218 259184 572278 259193
rect 572218 259115 572278 259124
rect 184938 258632 184994 258641
rect 184938 258567 184994 258576
rect 56508 256760 56560 256766
rect 56508 256702 56560 256708
rect 184952 253994 184980 258567
rect 571410 255912 571438 255930
rect 571385 255852 571394 255912
rect 571454 255852 571463 255912
rect 184860 253966 184980 253994
rect 184860 246498 184888 253966
rect 416778 252784 416834 252793
rect 416778 252719 416834 252728
rect 416792 251258 416820 252719
rect 416780 251252 416832 251258
rect 416780 251194 416832 251200
rect 567108 251252 567160 251258
rect 567108 251194 567160 251200
rect 416778 249520 416834 249529
rect 416778 249455 416834 249464
rect 416792 248470 416820 249455
rect 416780 248464 416832 248470
rect 416780 248406 416832 248412
rect 187606 248024 187662 248033
rect 187606 247959 187662 247968
rect 180708 246492 180760 246498
rect 180708 246434 180760 246440
rect 184848 246492 184900 246498
rect 184848 246434 184900 246440
rect 177948 237380 178000 237386
rect 177948 237322 178000 237328
rect 177960 232558 177988 237322
rect 74448 232552 74500 232558
rect 74448 232494 74500 232500
rect 177948 232552 178000 232558
rect 177948 232494 178000 232500
rect 51172 230716 51224 230722
rect 51172 230658 51224 230664
rect 51080 230648 51132 230654
rect 51080 230590 51132 230596
rect 74460 229158 74488 232494
rect 74448 229152 74500 229158
rect 74448 229094 74500 229100
rect 63500 229084 63552 229090
rect 63500 229026 63552 229032
rect 156972 229084 157024 229090
rect 156972 229026 157024 229032
rect 62762 227896 62818 227905
rect 62762 227831 62818 227840
rect 57610 227760 57666 227769
rect 52736 227724 52788 227730
rect 57610 227695 57666 227704
rect 52736 227666 52788 227672
rect 52748 217410 52776 227666
rect 56046 227624 56102 227633
rect 56046 227559 56102 227568
rect 55126 224904 55182 224913
rect 55126 224839 55182 224848
rect 53564 222352 53616 222358
rect 53564 222294 53616 222300
rect 53576 217410 53604 222294
rect 54390 222184 54446 222193
rect 54390 222119 54446 222128
rect 54404 217410 54432 222119
rect 55140 217410 55168 224839
rect 56060 217410 56088 227559
rect 56874 225040 56930 225049
rect 56874 224975 56930 224984
rect 56888 217410 56916 224975
rect 57624 217410 57652 227695
rect 60280 224936 60332 224942
rect 60280 224878 60332 224884
rect 57980 223644 58032 223650
rect 57980 223586 58032 223592
rect 52440 217382 52776 217410
rect 53268 217382 53604 217410
rect 54096 217382 54432 217410
rect 54924 217382 55168 217410
rect 55752 217382 56088 217410
rect 56580 217382 56916 217410
rect 57408 217382 57652 217410
rect 57992 216850 58020 223586
rect 59452 222216 59504 222222
rect 59452 222158 59504 222164
rect 58624 219768 58676 219774
rect 58624 219710 58676 219716
rect 58636 217410 58664 219710
rect 59464 217410 59492 222158
rect 60292 217410 60320 224878
rect 61106 222320 61162 222329
rect 61106 222255 61162 222264
rect 61936 222284 61988 222290
rect 61120 217410 61148 222255
rect 61936 222226 61988 222232
rect 61948 217410 61976 222226
rect 62776 217410 62804 227831
rect 63406 225176 63462 225185
rect 63406 225111 63462 225120
rect 63420 217410 63448 225111
rect 63512 223650 63540 229026
rect 152832 229016 152884 229022
rect 93030 228984 93086 228993
rect 152832 228958 152884 228964
rect 93030 228919 93086 228928
rect 84658 228848 84714 228857
rect 84658 228783 84714 228792
rect 82726 228440 82782 228449
rect 82726 228375 82782 228384
rect 76286 228304 76342 228313
rect 76286 228239 76342 228248
rect 69478 228168 69534 228177
rect 69478 228103 69534 228112
rect 64512 227860 64564 227866
rect 64512 227802 64564 227808
rect 63500 223644 63552 223650
rect 63500 223586 63552 223592
rect 64524 217410 64552 227802
rect 65340 227792 65392 227798
rect 65340 227734 65392 227740
rect 65352 217410 65380 227734
rect 66994 225312 67050 225321
rect 66994 225247 67050 225256
rect 66166 222456 66222 222465
rect 66166 222391 66222 222400
rect 66180 217410 66208 222391
rect 67008 217410 67036 225247
rect 67822 222592 67878 222601
rect 67822 222527 67878 222536
rect 67836 217410 67864 222527
rect 68652 222420 68704 222426
rect 68652 222362 68704 222368
rect 68664 217410 68692 222362
rect 69492 217410 69520 228103
rect 71226 228032 71282 228041
rect 71226 227967 71282 227976
rect 70398 225448 70454 225457
rect 70398 225383 70454 225392
rect 70412 217410 70440 225383
rect 71240 217410 71268 227967
rect 72056 227928 72108 227934
rect 72056 227870 72108 227876
rect 72068 217410 72096 227870
rect 73712 225004 73764 225010
rect 73712 224946 73764 224952
rect 72884 222488 72936 222494
rect 72884 222430 72936 222436
rect 72896 217410 72924 222430
rect 73724 217410 73752 224946
rect 74446 222728 74502 222737
rect 74446 222663 74502 222672
rect 74460 217410 74488 222663
rect 75368 222556 75420 222562
rect 75368 222498 75420 222504
rect 75380 217410 75408 222498
rect 76300 217410 76328 228239
rect 78772 227996 78824 228002
rect 78772 227938 78824 227944
rect 77114 225584 77170 225593
rect 77114 225519 77170 225528
rect 77128 217410 77156 225519
rect 77944 222964 77996 222970
rect 77944 222906 77996 222912
rect 77956 217410 77984 222906
rect 78784 217410 78812 227938
rect 80426 225720 80482 225729
rect 80426 225655 80482 225664
rect 79598 222864 79654 222873
rect 79598 222799 79654 222808
rect 79612 217410 79640 222799
rect 80440 217410 80468 225655
rect 81254 223000 81310 223009
rect 81254 222935 81310 222944
rect 81268 217410 81296 222935
rect 82176 222624 82228 222630
rect 82176 222566 82228 222572
rect 82188 217410 82216 222566
rect 82740 217410 82768 228375
rect 83830 225856 83886 225865
rect 83830 225791 83886 225800
rect 83844 217410 83872 225791
rect 84672 217410 84700 228783
rect 88062 228712 88118 228721
rect 88062 228647 88118 228656
rect 86314 228576 86370 228585
rect 86314 228511 86370 228520
rect 85488 222692 85540 222698
rect 85488 222634 85540 222640
rect 85500 217410 85528 222634
rect 86328 217410 86356 228511
rect 87144 223508 87196 223514
rect 87144 223450 87196 223456
rect 87156 217410 87184 223450
rect 88076 217410 88104 228647
rect 92202 225992 92258 226001
rect 92202 225927 92258 225936
rect 90548 225344 90600 225350
rect 90548 225286 90600 225292
rect 88892 225072 88944 225078
rect 88892 225014 88944 225020
rect 88904 217410 88932 225014
rect 89718 223136 89774 223145
rect 89718 223071 89774 223080
rect 89732 217410 89760 223071
rect 90560 217410 90588 225286
rect 91376 222760 91428 222766
rect 91376 222702 91428 222708
rect 91388 217410 91416 222702
rect 92216 217410 92244 225927
rect 93044 217410 93072 228919
rect 150256 228880 150308 228886
rect 150256 228822 150308 228828
rect 121184 228812 121236 228818
rect 121184 228754 121236 228760
rect 108212 228064 108264 228070
rect 108212 228006 108264 228012
rect 94778 227488 94834 227497
rect 94778 227423 94834 227432
rect 93768 222080 93820 222086
rect 93768 222022 93820 222028
rect 93780 217410 93808 222022
rect 94792 217410 94820 227423
rect 99838 227352 99894 227361
rect 99838 227287 99894 227296
rect 98918 226264 98974 226273
rect 98918 226199 98974 226208
rect 97262 226128 97318 226137
rect 97262 226063 97318 226072
rect 95608 225140 95660 225146
rect 95608 225082 95660 225088
rect 95620 217410 95648 225082
rect 96434 223272 96490 223281
rect 96434 223207 96490 223216
rect 96448 217410 96476 223207
rect 97276 217410 97304 226063
rect 98090 223408 98146 223417
rect 98090 223343 98146 223352
rect 98104 217410 98132 223343
rect 98932 217410 98960 226199
rect 99852 217410 99880 227287
rect 101494 227216 101550 227225
rect 101494 227151 101550 227160
rect 100668 225208 100720 225214
rect 100668 225150 100720 225156
rect 100680 217410 100708 225150
rect 101508 217410 101536 227151
rect 106554 227080 106610 227089
rect 106554 227015 106610 227024
rect 105728 225480 105780 225486
rect 105728 225422 105780 225428
rect 103980 225276 104032 225282
rect 103980 225218 104032 225224
rect 102046 224768 102102 224777
rect 102046 224703 102102 224712
rect 102060 217410 102088 224703
rect 103150 222048 103206 222057
rect 103150 221983 103206 221992
rect 103164 217410 103192 221983
rect 103992 217410 104020 225218
rect 104806 223544 104862 223553
rect 104806 223479 104862 223488
rect 104820 217410 104848 223479
rect 105740 217410 105768 225422
rect 106568 217410 106596 227015
rect 107384 225412 107436 225418
rect 107384 225354 107436 225360
rect 107396 217410 107424 225354
rect 108224 217410 108252 228006
rect 113086 226944 113142 226953
rect 113086 226879 113142 226888
rect 109038 224632 109094 224641
rect 109038 224567 109094 224576
rect 109052 217410 109080 224567
rect 110694 224496 110750 224505
rect 110694 224431 110750 224440
rect 109866 221912 109922 221921
rect 109866 221847 109922 221856
rect 109880 217410 109908 221847
rect 110708 217410 110736 224431
rect 112442 224224 112498 224233
rect 112442 224159 112498 224168
rect 111614 221776 111670 221785
rect 111614 221711 111670 221720
rect 111628 217410 111656 221711
rect 112456 217410 112484 224159
rect 113100 217410 113128 226879
rect 114926 226808 114982 226817
rect 114926 226743 114982 226752
rect 114100 225616 114152 225622
rect 114100 225558 114152 225564
rect 114112 217410 114140 225558
rect 114940 217410 114968 226743
rect 119160 225752 119212 225758
rect 119160 225694 119212 225700
rect 117504 225548 117556 225554
rect 117504 225490 117556 225496
rect 115754 224360 115810 224369
rect 115754 224295 115810 224304
rect 115768 217410 115796 224295
rect 116584 222896 116636 222902
rect 116584 222838 116636 222844
rect 116596 217410 116624 222838
rect 117516 217410 117544 225490
rect 118330 221640 118386 221649
rect 118330 221575 118386 221584
rect 118344 217410 118372 221575
rect 119172 217410 119200 225694
rect 120814 224088 120870 224097
rect 120814 224023 120870 224032
rect 119988 222828 120040 222834
rect 119988 222770 120040 222776
rect 120000 217410 120028 222770
rect 120828 217410 120856 224023
rect 121196 222970 121224 228754
rect 146024 228676 146076 228682
rect 146024 228618 146076 228624
rect 145196 228608 145248 228614
rect 145196 228550 145248 228556
rect 138480 228540 138532 228546
rect 138480 228482 138532 228488
rect 136824 228404 136876 228410
rect 136824 228346 136876 228352
rect 130108 228336 130160 228342
rect 130108 228278 130160 228284
rect 125048 228268 125100 228274
rect 125048 228210 125100 228216
rect 123392 228132 123444 228138
rect 123392 228074 123444 228080
rect 121184 222964 121236 222970
rect 121184 222906 121236 222912
rect 121366 221504 121422 221513
rect 121366 221439 121422 221448
rect 121380 217410 121408 221439
rect 122472 219836 122524 219842
rect 122472 219778 122524 219784
rect 122484 217410 122512 219778
rect 123404 217410 123432 228074
rect 124128 225684 124180 225690
rect 124128 225626 124180 225632
rect 124140 217410 124168 225626
rect 125060 217410 125088 228210
rect 127532 225820 127584 225826
rect 127532 225762 127584 225768
rect 126704 222964 126756 222970
rect 126704 222906 126756 222912
rect 125876 219904 125928 219910
rect 125876 219846 125928 219852
rect 125888 217410 125916 219846
rect 126716 217410 126744 222906
rect 127544 217410 127572 225762
rect 128360 223032 128412 223038
rect 128360 222974 128412 222980
rect 128372 217410 128400 222974
rect 129280 219972 129332 219978
rect 129280 219914 129332 219920
rect 129292 217410 129320 219914
rect 130120 217410 130148 228278
rect 131764 228200 131816 228206
rect 131764 228142 131816 228148
rect 130936 225956 130988 225962
rect 130936 225898 130988 225904
rect 130948 217410 130976 225898
rect 131776 217410 131804 228142
rect 134248 225888 134300 225894
rect 134248 225830 134300 225836
rect 133420 223100 133472 223106
rect 133420 223042 133472 223048
rect 132408 220040 132460 220046
rect 132408 219982 132460 219988
rect 132420 217410 132448 219982
rect 133432 217410 133460 223042
rect 134260 217410 134288 225830
rect 135168 223168 135220 223174
rect 135168 223110 135220 223116
rect 135180 217410 135208 223110
rect 135996 220108 136048 220114
rect 135996 220050 136048 220056
rect 136008 217410 136036 220050
rect 136836 217410 136864 228346
rect 137652 226024 137704 226030
rect 137652 225966 137704 225972
rect 137664 217410 137692 225966
rect 138492 217410 138520 228482
rect 143448 228472 143500 228478
rect 143448 228414 143500 228420
rect 141056 226092 141108 226098
rect 141056 226034 141108 226040
rect 140136 223236 140188 223242
rect 140136 223178 140188 223184
rect 139308 220176 139360 220182
rect 139308 220118 139360 220124
rect 139320 217410 139348 220118
rect 140148 217410 140176 223178
rect 141068 217410 141096 226034
rect 141884 223304 141936 223310
rect 141884 223246 141936 223252
rect 141896 217410 141924 223246
rect 142712 220244 142764 220250
rect 142712 220186 142764 220192
rect 142724 217410 142752 220186
rect 143460 217410 143488 228414
rect 144368 226228 144420 226234
rect 144368 226170 144420 226176
rect 144380 217410 144408 226170
rect 145208 217410 145236 228550
rect 146036 217410 146064 228618
rect 147772 226160 147824 226166
rect 147772 226102 147824 226108
rect 146944 223372 146996 223378
rect 146944 223314 146996 223320
rect 146956 217410 146984 223314
rect 147784 217410 147812 226102
rect 148600 223440 148652 223446
rect 148600 223382 148652 223388
rect 148612 217410 148640 223382
rect 149428 221332 149480 221338
rect 149428 221274 149480 221280
rect 149440 217410 149468 221274
rect 150268 217410 150296 228822
rect 151728 228744 151780 228750
rect 151728 228686 151780 228692
rect 151084 224868 151136 224874
rect 151084 224810 151136 224816
rect 151096 217410 151124 224810
rect 151740 217410 151768 228686
rect 152844 217410 152872 228958
rect 156144 228948 156196 228954
rect 156144 228890 156196 228896
rect 154488 226296 154540 226302
rect 154488 226238 154540 226244
rect 153660 223576 153712 223582
rect 153660 223518 153712 223524
rect 153672 217410 153700 223518
rect 154500 217410 154528 226238
rect 155408 224052 155460 224058
rect 155408 223994 155460 224000
rect 155316 222148 155368 222154
rect 155316 222090 155368 222096
rect 155328 217410 155356 222090
rect 155420 222086 155448 223994
rect 155408 222080 155460 222086
rect 155408 222022 155460 222028
rect 156156 217410 156184 228890
rect 156984 217410 157012 229026
rect 158720 227656 158772 227662
rect 158720 227598 158772 227604
rect 157800 224800 157852 224806
rect 157800 224742 157852 224748
rect 157812 217410 157840 224742
rect 158732 217410 158760 227598
rect 165436 227588 165488 227594
rect 165436 227530 165488 227536
rect 162768 227520 162820 227526
rect 162768 227462 162820 227468
rect 161204 224732 161256 224738
rect 161204 224674 161256 224680
rect 160376 222080 160428 222086
rect 160376 222022 160428 222028
rect 159548 221468 159600 221474
rect 159548 221410 159600 221416
rect 159560 217410 159588 221410
rect 160388 217410 160416 222022
rect 161216 217410 161244 224674
rect 162032 222012 162084 222018
rect 162032 221954 162084 221960
rect 162044 217410 162072 221954
rect 162780 217410 162808 227462
rect 163688 227452 163740 227458
rect 163688 227394 163740 227400
rect 163700 217410 163728 227394
rect 164608 224596 164660 224602
rect 164608 224538 164660 224544
rect 164620 217410 164648 224538
rect 165448 217410 165476 227530
rect 167092 227384 167144 227390
rect 167092 227326 167144 227332
rect 166264 221808 166316 221814
rect 166264 221750 166316 221756
rect 166276 217410 166304 221750
rect 167104 217410 167132 227326
rect 173624 227316 173676 227322
rect 173624 227258 173676 227264
rect 169576 227248 169628 227254
rect 169576 227190 169628 227196
rect 167920 224664 167972 224670
rect 167920 224606 167972 224612
rect 167932 217410 167960 224606
rect 168748 221876 168800 221882
rect 168748 221818 168800 221824
rect 168760 217410 168788 221818
rect 169588 217410 169616 227190
rect 172152 227180 172204 227186
rect 172152 227122 172204 227128
rect 170956 224528 171008 224534
rect 170956 224470 171008 224476
rect 169668 223644 169720 223650
rect 169668 223586 169720 223592
rect 58328 217382 58664 217410
rect 59156 217382 59492 217410
rect 59984 217382 60320 217410
rect 60812 217382 61148 217410
rect 61640 217382 61976 217410
rect 62468 217382 62804 217410
rect 63296 217382 63448 217410
rect 64216 217382 64552 217410
rect 65044 217382 65380 217410
rect 65872 217382 66208 217410
rect 66700 217382 67036 217410
rect 67528 217382 67864 217410
rect 68356 217382 68692 217410
rect 69184 217382 69520 217410
rect 70104 217382 70440 217410
rect 70932 217382 71268 217410
rect 71760 217382 72096 217410
rect 72588 217382 72924 217410
rect 73416 217382 73752 217410
rect 74244 217382 74488 217410
rect 75072 217382 75408 217410
rect 75992 217382 76328 217410
rect 76820 217382 77156 217410
rect 77648 217382 77984 217410
rect 78476 217382 78812 217410
rect 79304 217382 79640 217410
rect 80132 217382 80468 217410
rect 80960 217382 81296 217410
rect 81880 217382 82216 217410
rect 82708 217382 82768 217410
rect 83536 217382 83872 217410
rect 84364 217382 84700 217410
rect 85192 217382 85528 217410
rect 86020 217382 86356 217410
rect 86848 217382 87184 217410
rect 87768 217382 88104 217410
rect 88596 217382 88932 217410
rect 89424 217382 89760 217410
rect 90252 217382 90588 217410
rect 91080 217382 91416 217410
rect 91908 217382 92244 217410
rect 92736 217382 93072 217410
rect 93656 217382 93808 217410
rect 94484 217382 94820 217410
rect 95312 217382 95648 217410
rect 96140 217382 96476 217410
rect 96968 217382 97304 217410
rect 97796 217382 98132 217410
rect 98624 217382 98960 217410
rect 99544 217382 99880 217410
rect 100372 217382 100708 217410
rect 101200 217382 101536 217410
rect 102028 217382 102088 217410
rect 102856 217382 103192 217410
rect 103684 217382 104020 217410
rect 104512 217382 104848 217410
rect 105432 217382 105768 217410
rect 106260 217382 106596 217410
rect 107088 217382 107424 217410
rect 107916 217382 108252 217410
rect 108744 217382 109080 217410
rect 109572 217382 109908 217410
rect 110400 217382 110736 217410
rect 111320 217382 111656 217410
rect 112148 217382 112484 217410
rect 112976 217382 113128 217410
rect 113804 217382 114140 217410
rect 114632 217382 114968 217410
rect 115460 217382 115796 217410
rect 116288 217382 116624 217410
rect 117208 217382 117544 217410
rect 118036 217382 118372 217410
rect 118864 217382 119200 217410
rect 119692 217382 120028 217410
rect 120520 217382 120856 217410
rect 121348 217382 121408 217410
rect 122176 217382 122512 217410
rect 123096 217382 123432 217410
rect 123924 217382 124168 217410
rect 124752 217382 125088 217410
rect 125580 217382 125916 217410
rect 126408 217382 126744 217410
rect 127236 217382 127572 217410
rect 128064 217382 128400 217410
rect 128984 217382 129320 217410
rect 129812 217382 130148 217410
rect 130640 217382 130976 217410
rect 131468 217382 131804 217410
rect 132296 217382 132448 217410
rect 133124 217382 133460 217410
rect 133952 217382 134288 217410
rect 134872 217382 135208 217410
rect 135700 217382 136036 217410
rect 136528 217382 136864 217410
rect 137356 217382 137692 217410
rect 138184 217382 138520 217410
rect 139012 217382 139348 217410
rect 139840 217382 140176 217410
rect 140760 217382 141096 217410
rect 141588 217382 141924 217410
rect 142416 217382 142752 217410
rect 143244 217382 143488 217410
rect 144072 217382 144408 217410
rect 144900 217382 145236 217410
rect 145728 217382 146064 217410
rect 146648 217382 146984 217410
rect 147476 217382 147812 217410
rect 148304 217382 148640 217410
rect 149132 217382 149468 217410
rect 149960 217382 150296 217410
rect 150788 217382 151124 217410
rect 151616 217382 151768 217410
rect 152536 217382 152872 217410
rect 153364 217382 153700 217410
rect 154192 217382 154528 217410
rect 155020 217382 155356 217410
rect 155848 217382 156184 217410
rect 156676 217382 157012 217410
rect 157504 217382 157840 217410
rect 158424 217382 158760 217410
rect 159252 217382 159588 217410
rect 160080 217382 160416 217410
rect 160908 217382 161244 217410
rect 161736 217382 162072 217410
rect 162564 217382 162808 217410
rect 163392 217382 163728 217410
rect 164312 217382 164648 217410
rect 165140 217382 165476 217410
rect 165968 217382 166304 217410
rect 166796 217382 167132 217410
rect 167624 217382 167960 217410
rect 168452 217382 168788 217410
rect 169280 217382 169616 217410
rect 52184 216844 52236 216850
rect 52184 216786 52236 216792
rect 57980 216844 58032 216850
rect 57980 216786 58032 216792
rect 50988 214328 51040 214334
rect 50988 214270 51040 214276
rect 42156 182164 42208 182170
rect 42156 182106 42208 182112
rect 48504 182164 48556 182170
rect 48504 182106 48556 182112
rect 42168 181900 42196 182106
rect 52196 53922 52224 216786
rect 169680 216782 169708 223586
rect 170496 221944 170548 221950
rect 170496 221886 170548 221892
rect 170508 217410 170536 221886
rect 170200 217382 170536 217410
rect 170968 217410 170996 224470
rect 171048 223780 171100 223786
rect 171048 223722 171100 223728
rect 171060 223514 171088 223722
rect 171048 223508 171100 223514
rect 171048 223450 171100 223456
rect 172164 217410 172192 227122
rect 172980 221196 173032 221202
rect 172980 221138 173032 221144
rect 172992 217410 173020 221138
rect 173636 217410 173664 227258
rect 176384 227112 176436 227118
rect 176384 227054 176436 227060
rect 174636 224460 174688 224466
rect 174636 224402 174688 224408
rect 174648 217410 174676 224402
rect 175464 223508 175516 223514
rect 175464 223450 175516 223456
rect 175476 217410 175504 223450
rect 176396 217410 176424 227054
rect 180524 226976 180576 226982
rect 180524 226918 180576 226924
rect 178040 224324 178092 224330
rect 178040 224266 178092 224272
rect 177212 221740 177264 221746
rect 177212 221682 177264 221688
rect 177224 217410 177252 221682
rect 178052 217410 178080 224266
rect 178868 221400 178920 221406
rect 178868 221342 178920 221348
rect 178880 217410 178908 221342
rect 179696 221264 179748 221270
rect 179696 221206 179748 221212
rect 179708 217410 179736 221206
rect 180536 217410 180564 226918
rect 180720 223650 180748 246434
rect 184940 237448 184992 237454
rect 184938 237416 184940 237425
rect 184992 237416 184994 237425
rect 184938 237351 184994 237360
rect 181904 227044 181956 227050
rect 181904 226986 181956 226992
rect 181352 224392 181404 224398
rect 181352 224334 181404 224340
rect 180708 223644 180760 223650
rect 180708 223586 180760 223592
rect 181364 217410 181392 224334
rect 181916 221406 181944 226986
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 184756 224256 184808 224262
rect 184756 224198 184808 224204
rect 182180 223644 182232 223650
rect 182180 223586 182232 223592
rect 182192 222358 182220 223586
rect 182180 222352 182232 222358
rect 182180 222294 182232 222300
rect 183928 221672 183980 221678
rect 183928 221614 183980 221620
rect 182088 221604 182140 221610
rect 182088 221546 182140 221552
rect 181904 221400 181956 221406
rect 181904 221342 181956 221348
rect 181996 221400 182048 221406
rect 181996 221342 182048 221348
rect 182008 221202 182036 221342
rect 181996 221196 182048 221202
rect 181996 221138 182048 221144
rect 182100 217410 182128 221546
rect 183100 221196 183152 221202
rect 183100 221138 183152 221144
rect 183112 217410 183140 221138
rect 183940 217410 183968 221614
rect 184768 217410 184796 224198
rect 185596 217410 185624 226850
rect 186412 226772 186464 226778
rect 186412 226714 186464 226720
rect 186424 217410 186452 226714
rect 187240 222352 187292 222358
rect 187240 222294 187292 222300
rect 187252 217410 187280 222294
rect 170968 217382 171028 217410
rect 171856 217382 172192 217410
rect 172684 217382 173020 217410
rect 173512 217382 173664 217410
rect 174340 217382 174676 217410
rect 175168 217382 175504 217410
rect 176088 217382 176424 217410
rect 176916 217382 177252 217410
rect 177744 217382 178080 217410
rect 178572 217382 178908 217410
rect 179400 217382 179736 217410
rect 180228 217382 180564 217410
rect 181056 217382 181392 217410
rect 181976 217382 182128 217410
rect 182804 217382 183140 217410
rect 183632 217382 183968 217410
rect 184460 217382 184796 217410
rect 185288 217382 185624 217410
rect 186116 217382 186452 217410
rect 186944 217382 187280 217410
rect 187620 216782 187648 247959
rect 416778 246392 416834 246401
rect 416778 246327 416834 246336
rect 416792 245682 416820 246327
rect 416780 245676 416832 245682
rect 416780 245618 416832 245624
rect 564348 245676 564400 245682
rect 564348 245618 564400 245624
rect 418066 243128 418122 243137
rect 418066 243063 418122 243072
rect 190368 226840 190420 226846
rect 190368 226782 190420 226788
rect 188160 224188 188212 224194
rect 188160 224130 188212 224136
rect 188172 217410 188200 224130
rect 190276 223916 190328 223922
rect 190276 223858 190328 223864
rect 188988 221536 189040 221542
rect 188988 221478 189040 221484
rect 189000 217410 189028 221478
rect 190288 221338 190316 223858
rect 190276 221332 190328 221338
rect 190276 221274 190328 221280
rect 189816 221128 189868 221134
rect 189816 221070 189868 221076
rect 189828 217410 189856 221070
rect 190380 217410 190408 226782
rect 191472 224120 191524 224126
rect 191472 224062 191524 224068
rect 191484 217410 191512 224062
rect 192312 223650 192340 231676
rect 192588 224913 192616 231676
rect 192956 227730 192984 231676
rect 192944 227724 192996 227730
rect 192944 227666 192996 227672
rect 193036 227724 193088 227730
rect 193036 227666 193088 227672
rect 192944 226704 192996 226710
rect 192944 226646 192996 226652
rect 192574 224904 192630 224913
rect 192574 224839 192630 224848
rect 192300 223644 192352 223650
rect 192300 223586 192352 223592
rect 192852 222692 192904 222698
rect 192852 222634 192904 222640
rect 192300 221060 192352 221066
rect 192300 221002 192352 221008
rect 192312 217410 192340 221002
rect 192864 220998 192892 222634
rect 192852 220992 192904 220998
rect 192852 220934 192904 220940
rect 192956 217410 192984 226646
rect 193048 221066 193076 227666
rect 193128 222624 193180 222630
rect 193128 222566 193180 222572
rect 193140 222494 193168 222566
rect 193128 222488 193180 222494
rect 193128 222430 193180 222436
rect 193220 222488 193272 222494
rect 193220 222430 193272 222436
rect 193232 222222 193260 222430
rect 193220 222216 193272 222222
rect 193324 222193 193352 231676
rect 193416 228002 193628 228018
rect 193404 227996 193628 228002
rect 193456 227990 193628 227996
rect 193404 227938 193456 227944
rect 193600 227934 193628 227990
rect 193588 227928 193640 227934
rect 193588 227870 193640 227876
rect 193692 225049 193720 231676
rect 193784 231662 194074 231690
rect 193678 225040 193734 225049
rect 193678 224975 193734 224984
rect 193220 222158 193272 222164
rect 193310 222184 193366 222193
rect 193310 222119 193366 222128
rect 193036 221060 193088 221066
rect 193036 221002 193088 221008
rect 193784 219774 193812 231662
rect 194428 227633 194456 231676
rect 194796 227769 194824 231676
rect 194782 227760 194838 227769
rect 194782 227695 194838 227704
rect 194414 227624 194470 227633
rect 194414 227559 194470 227568
rect 195164 224942 195192 231676
rect 195152 224936 195204 224942
rect 195152 224878 195204 224884
rect 194876 223712 194928 223718
rect 194876 223654 194928 223660
rect 194048 222216 194100 222222
rect 194048 222158 194100 222164
rect 193772 219768 193824 219774
rect 193772 219710 193824 219716
rect 194060 217410 194088 222158
rect 194888 217410 194916 223654
rect 195440 222290 195468 231676
rect 195808 222494 195836 231676
rect 195796 222488 195848 222494
rect 195796 222430 195848 222436
rect 196176 222329 196204 231676
rect 196544 225185 196572 231676
rect 196912 227798 196940 231676
rect 197280 227905 197308 231676
rect 197266 227896 197322 227905
rect 197648 227866 197676 231676
rect 197266 227831 197322 227840
rect 197636 227860 197688 227866
rect 197636 227802 197688 227808
rect 196900 227792 196952 227798
rect 196900 227734 196952 227740
rect 197360 227792 197412 227798
rect 197360 227734 197412 227740
rect 196530 225176 196586 225185
rect 196530 225111 196586 225120
rect 197268 222760 197320 222766
rect 197268 222702 197320 222708
rect 196162 222320 196218 222329
rect 195428 222284 195480 222290
rect 195428 222226 195480 222232
rect 195704 222284 195756 222290
rect 196162 222255 196218 222264
rect 195704 222226 195756 222232
rect 195716 217410 195744 222226
rect 197280 220998 197308 222702
rect 197268 220992 197320 220998
rect 197268 220934 197320 220940
rect 196532 220856 196584 220862
rect 196532 220798 196584 220804
rect 196544 217410 196572 220798
rect 197372 217410 197400 227734
rect 197820 226500 197872 226506
rect 197820 226442 197872 226448
rect 197832 225350 197860 226442
rect 197820 225344 197872 225350
rect 198016 225321 198044 231676
rect 198188 225344 198240 225350
rect 197820 225286 197872 225292
rect 198002 225312 198058 225321
rect 198188 225286 198240 225292
rect 198002 225247 198058 225256
rect 197452 225208 197504 225214
rect 197452 225150 197504 225156
rect 197464 224058 197492 225150
rect 197452 224052 197504 224058
rect 197452 223994 197504 224000
rect 198200 217410 198228 225286
rect 198292 222426 198320 231676
rect 198660 222465 198688 231676
rect 198752 231662 199042 231690
rect 198752 222601 198780 231662
rect 199016 227928 199068 227934
rect 199016 227870 199068 227876
rect 198738 222592 198794 222601
rect 198738 222527 198794 222536
rect 198646 222456 198702 222465
rect 198280 222420 198332 222426
rect 198646 222391 198702 222400
rect 198280 222362 198332 222368
rect 199028 217410 199056 227870
rect 199396 225457 199424 231676
rect 199764 228002 199792 231676
rect 200132 228177 200160 231676
rect 200118 228168 200174 228177
rect 200118 228103 200174 228112
rect 200500 228041 200528 231676
rect 200486 228032 200542 228041
rect 199752 227996 199804 228002
rect 200486 227967 200542 227976
rect 199752 227938 199804 227944
rect 199382 225448 199438 225457
rect 199382 225383 199438 225392
rect 200868 225010 200896 231676
rect 200856 225004 200908 225010
rect 200856 224946 200908 224952
rect 201144 222562 201172 231676
rect 201512 226334 201540 231676
rect 201328 226306 201540 226334
rect 201328 222630 201356 226306
rect 201408 224936 201460 224942
rect 201408 224878 201460 224884
rect 201316 222624 201368 222630
rect 201316 222566 201368 222572
rect 201132 222556 201184 222562
rect 201132 222498 201184 222504
rect 200764 222420 200816 222426
rect 200764 222362 200816 222368
rect 199936 221332 199988 221338
rect 199936 221274 199988 221280
rect 199948 217410 199976 221274
rect 200776 217410 200804 222362
rect 201420 217410 201448 224878
rect 201880 222737 201908 231676
rect 202248 225593 202276 231676
rect 202616 227866 202644 231676
rect 202984 228313 203012 231676
rect 203352 228818 203380 231676
rect 203340 228812 203392 228818
rect 203340 228754 203392 228760
rect 202970 228304 203026 228313
rect 202970 228239 203026 228248
rect 203248 227996 203300 228002
rect 203248 227938 203300 227944
rect 202604 227860 202656 227866
rect 202604 227802 202656 227808
rect 202234 225584 202290 225593
rect 202234 225519 202290 225528
rect 201866 222728 201922 222737
rect 201866 222663 201922 222672
rect 202420 222488 202472 222494
rect 202420 222430 202472 222436
rect 202432 217410 202460 222430
rect 203260 217410 203288 227938
rect 203720 225729 203748 231676
rect 203706 225720 203762 225729
rect 203706 225655 203762 225664
rect 203996 222698 204024 231676
rect 204378 231662 204484 231690
rect 204076 227860 204128 227866
rect 204076 227802 204128 227808
rect 203984 222692 204036 222698
rect 203984 222634 204036 222640
rect 204088 217410 204116 227802
rect 204260 223984 204312 223990
rect 204260 223926 204312 223932
rect 204272 220862 204300 223926
rect 204456 222873 204484 231662
rect 204732 223009 204760 231676
rect 205100 225865 205128 231676
rect 205086 225856 205142 225865
rect 205086 225791 205142 225800
rect 204718 223000 204774 223009
rect 204718 222935 204774 222944
rect 204442 222864 204498 222873
rect 204442 222799 204498 222808
rect 205468 221066 205496 231676
rect 205836 228449 205864 231676
rect 206204 228857 206232 231676
rect 206190 228848 206246 228857
rect 206190 228783 206246 228792
rect 205822 228440 205878 228449
rect 205822 228375 205878 228384
rect 206572 223786 206600 231676
rect 206848 226334 206876 231676
rect 207216 228585 207244 231676
rect 207584 228721 207612 231676
rect 207570 228712 207626 228721
rect 207570 228647 207626 228656
rect 207202 228576 207258 228585
rect 207202 228511 207258 228520
rect 207952 226506 207980 231676
rect 207940 226500 207992 226506
rect 207940 226442 207992 226448
rect 206756 226306 206876 226334
rect 206756 225078 206784 226306
rect 208320 226001 208348 231676
rect 208306 225992 208362 226001
rect 208306 225927 208362 225936
rect 208308 225208 208360 225214
rect 208308 225150 208360 225156
rect 206744 225072 206796 225078
rect 206928 225072 206980 225078
rect 206744 225014 206796 225020
rect 206848 225020 206928 225026
rect 206848 225014 206980 225020
rect 206848 224998 206968 225014
rect 206560 223780 206612 223786
rect 206560 223722 206612 223728
rect 205824 222556 205876 222562
rect 205824 222498 205876 222504
rect 205456 221060 205508 221066
rect 205456 221002 205508 221008
rect 204260 220856 204312 220862
rect 204260 220798 204312 220804
rect 204904 220856 204956 220862
rect 204904 220798 204956 220804
rect 204916 217410 204944 220798
rect 205836 217410 205864 222498
rect 206652 221060 206704 221066
rect 206652 221002 206704 221008
rect 206664 217410 206692 221002
rect 206848 220862 206876 224998
rect 207020 224936 207072 224942
rect 206940 224884 207020 224890
rect 206940 224878 207072 224884
rect 206940 224862 207060 224878
rect 206940 223718 206968 224862
rect 206928 223712 206980 223718
rect 206928 223654 206980 223660
rect 207480 222760 207532 222766
rect 207480 222702 207532 222708
rect 206836 220856 206888 220862
rect 206836 220798 206888 220804
rect 207492 217410 207520 222702
rect 208320 217410 208348 225150
rect 208688 223145 208716 231676
rect 208674 223136 208730 223145
rect 208674 223071 208730 223080
rect 209056 220998 209084 231676
rect 209424 223854 209452 231676
rect 209596 228812 209648 228818
rect 209596 228754 209648 228760
rect 209412 223848 209464 223854
rect 209412 223790 209464 223796
rect 209136 222624 209188 222630
rect 209136 222566 209188 222572
rect 209044 220992 209096 220998
rect 209044 220934 209096 220940
rect 209148 217410 209176 222566
rect 187864 217382 188200 217410
rect 188692 217382 189028 217410
rect 189520 217382 189856 217410
rect 190348 217382 190408 217410
rect 191176 217382 191512 217410
rect 192004 217382 192340 217410
rect 192832 217382 192984 217410
rect 193752 217382 194088 217410
rect 194580 217382 194916 217410
rect 195408 217382 195744 217410
rect 196236 217382 196572 217410
rect 197064 217382 197400 217410
rect 197892 217382 198228 217410
rect 198720 217382 199056 217410
rect 199640 217382 199976 217410
rect 200468 217382 200804 217410
rect 201296 217382 201448 217410
rect 202124 217382 202460 217410
rect 202952 217382 203288 217410
rect 203780 217382 204116 217410
rect 204608 217382 204944 217410
rect 205528 217382 205864 217410
rect 206356 217382 206692 217410
rect 207184 217382 207520 217410
rect 208012 217382 208348 217410
rect 208840 217382 209176 217410
rect 209608 217410 209636 228754
rect 209700 225146 209728 231676
rect 210068 228993 210096 231676
rect 210054 228984 210110 228993
rect 210054 228919 210110 228928
rect 210436 227497 210464 231676
rect 210698 227624 210754 227633
rect 210698 227559 210754 227568
rect 210422 227488 210478 227497
rect 210422 227423 210478 227432
rect 209688 225140 209740 225146
rect 209688 225082 209740 225088
rect 209688 223780 209740 223786
rect 209688 223722 209740 223728
rect 209700 221474 209728 223722
rect 209688 221468 209740 221474
rect 209688 221410 209740 221416
rect 210712 217410 210740 227559
rect 210804 226137 210832 231676
rect 211172 226273 211200 231676
rect 211158 226264 211214 226273
rect 211158 226199 211214 226208
rect 210790 226128 210846 226137
rect 210790 226063 210846 226072
rect 211540 223281 211568 231676
rect 211712 225208 211764 225214
rect 211712 225150 211764 225156
rect 211526 223272 211582 223281
rect 211526 223207 211582 223216
rect 211724 217410 211752 225150
rect 211908 223417 211936 231676
rect 212276 224058 212304 231676
rect 212354 227760 212410 227769
rect 212354 227695 212410 227704
rect 212264 224052 212316 224058
rect 212264 223994 212316 224000
rect 211894 223408 211950 223417
rect 211894 223343 211950 223352
rect 212368 217410 212396 227695
rect 212552 224777 212580 231676
rect 212920 227361 212948 231676
rect 212906 227352 212962 227361
rect 212906 227287 212962 227296
rect 213288 227225 213316 231676
rect 213274 227216 213330 227225
rect 213274 227151 213330 227160
rect 213656 225282 213684 231676
rect 214024 225486 214052 231676
rect 214012 225480 214064 225486
rect 214012 225422 214064 225428
rect 213644 225276 213696 225282
rect 213644 225218 213696 225224
rect 212538 224768 212594 224777
rect 212538 224703 212594 224712
rect 214288 224052 214340 224058
rect 214288 223994 214340 224000
rect 214300 221270 214328 223994
rect 214392 222057 214420 231676
rect 214760 223553 214788 231676
rect 215128 225418 215156 231676
rect 215116 225412 215168 225418
rect 215116 225354 215168 225360
rect 215024 225276 215076 225282
rect 215024 225218 215076 225224
rect 214746 223544 214802 223553
rect 214746 223479 214802 223488
rect 214378 222048 214434 222057
rect 214378 221983 214434 221992
rect 214288 221264 214340 221270
rect 214288 221206 214340 221212
rect 213368 220992 213420 220998
rect 213368 220934 213420 220940
rect 213380 217410 213408 220934
rect 213874 217660 213926 217666
rect 213874 217602 213926 217608
rect 209608 217382 209668 217410
rect 210496 217382 210740 217410
rect 211416 217382 211752 217410
rect 212244 217382 212396 217410
rect 213072 217382 213408 217410
rect 213886 217396 213914 217602
rect 215036 217410 215064 225218
rect 215404 224641 215432 231676
rect 215772 227089 215800 231676
rect 216140 228070 216168 231676
rect 216128 228064 216180 228070
rect 216128 228006 216180 228012
rect 215758 227080 215814 227089
rect 215758 227015 215814 227024
rect 215390 224632 215446 224641
rect 215390 224567 215446 224576
rect 216508 224505 216536 231676
rect 216680 228064 216732 228070
rect 216680 228006 216732 228012
rect 216494 224496 216550 224505
rect 216494 224431 216550 224440
rect 216220 223848 216272 223854
rect 216220 223790 216272 223796
rect 215208 223712 215260 223718
rect 215208 223654 215260 223660
rect 215220 221406 215248 223654
rect 215852 222692 215904 222698
rect 215852 222634 215904 222640
rect 215208 221400 215260 221406
rect 215208 221342 215260 221348
rect 215864 217410 215892 222634
rect 216232 221202 216260 223790
rect 216220 221196 216272 221202
rect 216220 221138 216272 221144
rect 216692 217410 216720 228006
rect 216876 224233 216904 231676
rect 216862 224224 216918 224233
rect 216862 224159 216918 224168
rect 217244 221921 217272 231676
rect 217336 231662 217626 231690
rect 217230 221912 217286 221921
rect 217230 221847 217286 221856
rect 217336 221785 217364 231662
rect 217598 227896 217654 227905
rect 217598 227831 217654 227840
rect 217322 221776 217378 221785
rect 217322 221711 217378 221720
rect 217612 217410 217640 227831
rect 217980 225622 218008 231676
rect 217968 225616 218020 225622
rect 217968 225558 218020 225564
rect 218256 224369 218284 231676
rect 218624 226953 218652 231676
rect 218610 226944 218666 226953
rect 218610 226879 218666 226888
rect 218992 226817 219020 231676
rect 219254 228168 219310 228177
rect 219254 228103 219310 228112
rect 218978 226808 219034 226817
rect 218978 226743 219034 226752
rect 218428 225480 218480 225486
rect 218428 225422 218480 225428
rect 218242 224360 218298 224369
rect 218242 224295 218298 224304
rect 218440 217410 218468 225422
rect 219268 217410 219296 228103
rect 219360 225554 219388 231676
rect 219728 225758 219756 231676
rect 219716 225752 219768 225758
rect 219716 225694 219768 225700
rect 219348 225548 219400 225554
rect 219348 225490 219400 225496
rect 220096 222902 220124 231676
rect 220084 222896 220136 222902
rect 220084 222838 220136 222844
rect 219992 222148 220044 222154
rect 219992 222090 220044 222096
rect 220084 222148 220136 222154
rect 220084 222090 220136 222096
rect 220004 221542 220032 222090
rect 219992 221536 220044 221542
rect 219992 221478 220044 221484
rect 219900 221468 219952 221474
rect 219900 221410 219952 221416
rect 219912 217666 219940 221410
rect 219900 217660 219952 217666
rect 219900 217602 219952 217608
rect 220096 217410 220124 222090
rect 220464 221649 220492 231676
rect 220726 228032 220782 228041
rect 220726 227967 220782 227976
rect 220636 225752 220688 225758
rect 220636 225694 220688 225700
rect 220450 221640 220506 221649
rect 220450 221575 220506 221584
rect 220648 221134 220676 225694
rect 220636 221128 220688 221134
rect 220636 221070 220688 221076
rect 220740 217410 220768 227967
rect 220832 224097 220860 231676
rect 220818 224088 220874 224097
rect 220818 224023 220874 224032
rect 221108 219842 221136 231676
rect 221476 222834 221504 231676
rect 221740 225480 221792 225486
rect 221740 225422 221792 225428
rect 221464 222828 221516 222834
rect 221464 222770 221516 222776
rect 221096 219836 221148 219842
rect 221096 219778 221148 219784
rect 221752 217410 221780 225422
rect 221844 221513 221872 231676
rect 222212 225690 222240 231676
rect 222304 231662 222594 231690
rect 222200 225684 222252 225690
rect 222200 225626 222252 225632
rect 222108 223576 222160 223582
rect 222106 223544 222108 223553
rect 222160 223544 222162 223553
rect 222106 223479 222162 223488
rect 221830 221504 221886 221513
rect 221830 221439 221886 221448
rect 222304 219910 222332 231662
rect 222948 228138 222976 231676
rect 223316 228274 223344 231676
rect 223304 228268 223356 228274
rect 223304 228210 223356 228216
rect 222936 228132 222988 228138
rect 222936 228074 222988 228080
rect 223488 228132 223540 228138
rect 223488 228074 223540 228080
rect 222568 222828 222620 222834
rect 222568 222770 222620 222776
rect 222292 219904 222344 219910
rect 222292 219846 222344 219852
rect 222580 217410 222608 222770
rect 223500 217410 223528 228074
rect 223684 225826 223712 231676
rect 223776 231662 223974 231690
rect 224052 231662 224342 231690
rect 223672 225820 223724 225826
rect 223672 225762 223724 225768
rect 223776 219978 223804 231662
rect 223856 223440 223908 223446
rect 223856 223382 223908 223388
rect 223868 222902 223896 223382
rect 224052 222970 224080 231662
rect 224408 223576 224460 223582
rect 224408 223518 224460 223524
rect 224132 223372 224184 223378
rect 224420 223360 224448 223518
rect 224184 223332 224448 223360
rect 224132 223314 224184 223320
rect 224696 223038 224724 231676
rect 225064 225962 225092 231676
rect 225052 225956 225104 225962
rect 225052 225898 225104 225904
rect 225144 225412 225196 225418
rect 225144 225354 225196 225360
rect 224684 223032 224736 223038
rect 224684 222974 224736 222980
rect 224040 222964 224092 222970
rect 224040 222906 224092 222912
rect 223856 222896 223908 222902
rect 223856 222838 223908 222844
rect 224316 222896 224368 222902
rect 224316 222838 224368 222844
rect 223764 219972 223816 219978
rect 223764 219914 223816 219920
rect 224328 217410 224356 222838
rect 225156 217410 225184 225354
rect 225432 220046 225460 231676
rect 225800 228342 225828 231676
rect 225788 228336 225840 228342
rect 225788 228278 225840 228284
rect 225970 228304 226026 228313
rect 225970 228239 226026 228248
rect 225420 220040 225472 220046
rect 225420 219982 225472 219988
rect 225984 217410 226012 228239
rect 226168 228206 226196 231676
rect 226156 228200 226208 228206
rect 226156 228142 226208 228148
rect 226536 225894 226564 231676
rect 226628 231662 226826 231690
rect 226524 225888 226576 225894
rect 226524 225830 226576 225836
rect 226628 220114 226656 231662
rect 227180 223106 227208 231676
rect 227444 223440 227496 223446
rect 227444 223382 227496 223388
rect 227168 223100 227220 223106
rect 227168 223042 227220 223048
rect 227456 221950 227484 223382
rect 227548 223174 227576 231676
rect 227720 228268 227772 228274
rect 227720 228210 227772 228216
rect 227628 223304 227680 223310
rect 227628 223246 227680 223252
rect 227536 223168 227588 223174
rect 227536 223110 227588 223116
rect 227640 222358 227668 223246
rect 227628 222352 227680 222358
rect 227628 222294 227680 222300
rect 227444 221944 227496 221950
rect 227444 221886 227496 221892
rect 226800 221264 226852 221270
rect 226800 221206 226852 221212
rect 226616 220108 226668 220114
rect 226616 220050 226668 220056
rect 226812 217410 226840 221206
rect 227732 218054 227760 228210
rect 227916 226030 227944 231676
rect 227904 226024 227956 226030
rect 227904 225966 227956 225972
rect 227810 223544 227866 223553
rect 227810 223479 227866 223488
rect 227824 223174 227852 223479
rect 227812 223168 227864 223174
rect 227812 223110 227864 223116
rect 228284 220182 228312 231676
rect 228652 228410 228680 231676
rect 229020 228546 229048 231676
rect 229008 228540 229060 228546
rect 229008 228482 229060 228488
rect 228640 228404 228692 228410
rect 228640 228346 228692 228352
rect 229284 228404 229336 228410
rect 229284 228346 229336 228352
rect 228456 225616 228508 225622
rect 228456 225558 228508 225564
rect 228272 220176 228324 220182
rect 228272 220118 228324 220124
rect 227640 218026 227760 218054
rect 227640 217410 227668 218026
rect 228468 217410 228496 225558
rect 229296 217410 229324 228346
rect 229388 226098 229416 231676
rect 229376 226092 229428 226098
rect 229376 226034 229428 226040
rect 229664 220250 229692 231676
rect 230032 223242 230060 231676
rect 230400 223378 230428 231676
rect 230768 226234 230796 231676
rect 231136 228682 231164 231676
rect 231124 228676 231176 228682
rect 231124 228618 231176 228624
rect 231504 228478 231532 231676
rect 231872 228614 231900 231676
rect 231860 228608 231912 228614
rect 231860 228550 231912 228556
rect 231492 228472 231544 228478
rect 231492 228414 231544 228420
rect 231676 228200 231728 228206
rect 231676 228142 231728 228148
rect 230756 226228 230808 226234
rect 230756 226170 230808 226176
rect 230388 223372 230440 223378
rect 230388 223314 230440 223320
rect 230020 223236 230072 223242
rect 230020 223178 230072 223184
rect 231032 223100 231084 223106
rect 231032 223042 231084 223048
rect 230204 221060 230256 221066
rect 230204 221002 230256 221008
rect 229652 220244 229704 220250
rect 229652 220186 229704 220192
rect 230216 217410 230244 221002
rect 231044 217410 231072 223042
rect 231688 217410 231716 228142
rect 232240 226166 232268 231676
rect 232228 226160 232280 226166
rect 232228 226102 232280 226108
rect 231860 225684 231912 225690
rect 231860 225626 231912 225632
rect 231872 221338 231900 225626
rect 232516 223922 232544 231676
rect 232504 223916 232556 223922
rect 232504 223858 232556 223864
rect 232884 223582 232912 231676
rect 232872 223576 232924 223582
rect 232872 223518 232924 223524
rect 233252 223038 233280 231676
rect 233620 224874 233648 231676
rect 233988 229022 234016 231676
rect 233976 229016 234028 229022
rect 233976 228958 234028 228964
rect 234356 228886 234384 231676
rect 234344 228880 234396 228886
rect 234344 228822 234396 228828
rect 234724 228750 234752 231676
rect 234712 228744 234764 228750
rect 234712 228686 234764 228692
rect 234802 228576 234858 228585
rect 234802 228511 234858 228520
rect 234618 228440 234674 228449
rect 234618 228375 234674 228384
rect 233608 224868 233660 224874
rect 233608 224810 233660 224816
rect 233240 223032 233292 223038
rect 233240 222974 233292 222980
rect 232688 222964 232740 222970
rect 232688 222906 232740 222912
rect 231860 221332 231912 221338
rect 231860 221274 231912 221280
rect 232700 217410 232728 222906
rect 234632 222154 234660 228375
rect 234712 226636 234764 226642
rect 234712 226578 234764 226584
rect 234620 222148 234672 222154
rect 234620 222090 234672 222096
rect 234344 221808 234396 221814
rect 234344 221750 234396 221756
rect 233516 220856 233568 220862
rect 233516 220798 233568 220804
rect 233528 217410 233556 220798
rect 234356 217410 234384 221750
rect 234724 221134 234752 226578
rect 234712 221128 234764 221134
rect 234712 221070 234764 221076
rect 234816 220998 234844 228511
rect 235092 226302 235120 231676
rect 235368 228954 235396 231676
rect 235356 228948 235408 228954
rect 235356 228890 235408 228896
rect 235264 228472 235316 228478
rect 235264 228414 235316 228420
rect 235080 226296 235132 226302
rect 235080 226238 235132 226244
rect 234804 220992 234856 220998
rect 234804 220934 234856 220940
rect 235276 217410 235304 228414
rect 235736 223174 235764 231676
rect 235828 231662 236118 231690
rect 235724 223168 235776 223174
rect 235724 223110 235776 223116
rect 235828 221542 235856 231662
rect 236472 224806 236500 231676
rect 236460 224800 236512 224806
rect 236460 224742 236512 224748
rect 236840 223786 236868 231676
rect 237208 229090 237236 231676
rect 237196 229084 237248 229090
rect 237196 229026 237248 229032
rect 237576 227662 237604 231676
rect 237564 227656 237616 227662
rect 237564 227598 237616 227604
rect 237944 224738 237972 231676
rect 238220 227526 238248 231676
rect 238312 231662 238602 231690
rect 238208 227520 238260 227526
rect 238208 227462 238260 227468
rect 237932 224732 237984 224738
rect 237932 224674 237984 224680
rect 236828 223780 236880 223786
rect 236828 223722 236880 223728
rect 237748 223372 237800 223378
rect 237748 223314 237800 223320
rect 236092 223032 236144 223038
rect 236092 222974 236144 222980
rect 235816 221536 235868 221542
rect 235816 221478 235868 221484
rect 236104 217410 236132 222974
rect 236920 221332 236972 221338
rect 236920 221274 236972 221280
rect 236932 217410 236960 221274
rect 237760 217410 237788 223314
rect 238312 222086 238340 231662
rect 238484 228608 238536 228614
rect 238484 228550 238536 228556
rect 238300 222080 238352 222086
rect 238300 222022 238352 222028
rect 238496 220862 238524 228550
rect 238576 228336 238628 228342
rect 238576 228278 238628 228284
rect 238484 220856 238536 220862
rect 238484 220798 238536 220804
rect 238588 217410 238616 228278
rect 238956 222018 238984 231676
rect 239324 224602 239352 231676
rect 239312 224596 239364 224602
rect 239312 224538 239364 224544
rect 239404 223236 239456 223242
rect 239404 223178 239456 223184
rect 238944 222012 238996 222018
rect 238944 221954 238996 221960
rect 239416 217410 239444 223178
rect 239692 221882 239720 231676
rect 239864 229016 239916 229022
rect 239864 228958 239916 228964
rect 239680 221876 239732 221882
rect 239680 221818 239732 221824
rect 239876 221270 239904 228958
rect 239956 228880 240008 228886
rect 239956 228822 240008 228828
rect 239864 221264 239916 221270
rect 239864 221206 239916 221212
rect 239968 221066 239996 228822
rect 240060 227458 240088 231676
rect 240324 228948 240376 228954
rect 240324 228890 240376 228896
rect 240140 228540 240192 228546
rect 240140 228482 240192 228488
rect 240048 227452 240100 227458
rect 240048 227394 240100 227400
rect 239956 221060 240008 221066
rect 239956 221002 240008 221008
rect 240152 220946 240180 228482
rect 240336 221338 240364 228890
rect 240428 227594 240456 231676
rect 240416 227588 240468 227594
rect 240416 227530 240468 227536
rect 240796 224670 240824 231676
rect 241072 227254 241100 231676
rect 241440 227390 241468 231676
rect 241428 227384 241480 227390
rect 241428 227326 241480 227332
rect 241060 227248 241112 227254
rect 241060 227190 241112 227196
rect 240784 224664 240836 224670
rect 240784 224606 240836 224612
rect 241152 223576 241204 223582
rect 241152 223518 241204 223524
rect 240324 221332 240376 221338
rect 240324 221274 240376 221280
rect 240060 220918 240180 220946
rect 240060 217410 240088 220918
rect 241164 217410 241192 223518
rect 241808 221950 241836 231676
rect 241980 228744 242032 228750
rect 241980 228686 242032 228692
rect 241796 221944 241848 221950
rect 241796 221886 241848 221892
rect 241992 217410 242020 228686
rect 242176 224534 242204 231676
rect 242164 224528 242216 224534
rect 242164 224470 242216 224476
rect 242544 223718 242572 231676
rect 242532 223712 242584 223718
rect 242532 223654 242584 223660
rect 242912 223446 242940 231676
rect 243280 227186 243308 231676
rect 243372 231662 243662 231690
rect 243268 227180 243320 227186
rect 243268 227122 243320 227128
rect 243372 224466 243400 231662
rect 243636 227656 243688 227662
rect 243636 227598 243688 227604
rect 243360 224460 243412 224466
rect 243360 224402 243412 224408
rect 242900 223440 242952 223446
rect 242900 223382 242952 223388
rect 242808 223168 242860 223174
rect 242808 223110 242860 223116
rect 242820 217410 242848 223110
rect 243648 217410 243676 227598
rect 243924 227118 243952 231676
rect 244292 227322 244320 231676
rect 244280 227316 244332 227322
rect 244280 227258 244332 227264
rect 243912 227112 243964 227118
rect 243912 227054 243964 227060
rect 244660 223514 244688 231676
rect 245028 224330 245056 231676
rect 245292 228676 245344 228682
rect 245292 228618 245344 228624
rect 245016 224324 245068 224330
rect 245016 224266 245068 224272
rect 244648 223508 244700 223514
rect 244648 223450 244700 223456
rect 244464 222080 244516 222086
rect 244464 222022 244516 222028
rect 244476 217410 244504 222022
rect 245304 217410 245332 228618
rect 245396 224058 245424 231676
rect 245660 226500 245712 226506
rect 245660 226442 245712 226448
rect 245384 224052 245436 224058
rect 245384 223994 245436 224000
rect 245672 222766 245700 226442
rect 245660 222760 245712 222766
rect 245660 222702 245712 222708
rect 245764 221746 245792 231676
rect 245842 228848 245898 228857
rect 245842 228783 245898 228792
rect 245752 221740 245804 221746
rect 245752 221682 245804 221688
rect 245856 221474 245884 228783
rect 246132 227050 246160 231676
rect 246120 227044 246172 227050
rect 246120 226986 246172 226992
rect 246500 224398 246528 231676
rect 246488 224392 246540 224398
rect 246488 224334 246540 224340
rect 246776 223854 246804 231676
rect 247144 226982 247172 231676
rect 247132 226976 247184 226982
rect 247132 226918 247184 226924
rect 247040 226568 247092 226574
rect 247040 226510 247092 226516
rect 246764 223848 246816 223854
rect 246764 223790 246816 223796
rect 245844 221468 245896 221474
rect 245844 221410 245896 221416
rect 246120 221196 246172 221202
rect 246120 221138 246172 221144
rect 246132 217410 246160 221138
rect 247052 217410 247080 226510
rect 247512 221542 247540 231676
rect 247880 224262 247908 231676
rect 248248 226778 248276 231676
rect 248340 231662 248630 231690
rect 248236 226772 248288 226778
rect 248236 226714 248288 226720
rect 247868 224256 247920 224262
rect 247868 224198 247920 224204
rect 248340 221678 248368 231662
rect 248696 227520 248748 227526
rect 248696 227462 248748 227468
rect 248604 227384 248656 227390
rect 248604 227326 248656 227332
rect 248420 227248 248472 227254
rect 248420 227190 248472 227196
rect 248432 221814 248460 227190
rect 248512 227044 248564 227050
rect 248512 226986 248564 226992
rect 248524 222902 248552 226986
rect 248616 223106 248644 227326
rect 248604 223100 248656 223106
rect 248604 223042 248656 223048
rect 248512 222896 248564 222902
rect 248512 222838 248564 222844
rect 248420 221808 248472 221814
rect 248420 221750 248472 221756
rect 248328 221672 248380 221678
rect 248328 221614 248380 221620
rect 247500 221536 247552 221542
rect 247500 221478 247552 221484
rect 247868 221332 247920 221338
rect 247868 221274 247920 221280
rect 247880 217410 247908 221274
rect 248708 217410 248736 227462
rect 248984 226914 249012 231676
rect 248972 226908 249024 226914
rect 248972 226850 249024 226856
rect 249352 224194 249380 231676
rect 249628 225758 249656 231676
rect 249616 225752 249668 225758
rect 249616 225694 249668 225700
rect 249340 224188 249392 224194
rect 249340 224130 249392 224136
rect 249996 223310 250024 231676
rect 250088 231662 250378 231690
rect 249984 223304 250036 223310
rect 249984 223246 250036 223252
rect 249524 221468 249576 221474
rect 249524 221410 249576 221416
rect 249536 217410 249564 221410
rect 250088 221406 250116 231662
rect 250352 227588 250404 227594
rect 250352 227530 250404 227536
rect 250076 221400 250128 221406
rect 250076 221342 250128 221348
rect 250364 217410 250392 227530
rect 250732 224126 250760 231676
rect 251100 226710 251128 231676
rect 251468 226846 251496 231676
rect 251836 227730 251864 231676
rect 251824 227724 251876 227730
rect 251824 227666 251876 227672
rect 252008 227452 252060 227458
rect 252008 227394 252060 227400
rect 251456 226840 251508 226846
rect 251456 226782 251508 226788
rect 251088 226704 251140 226710
rect 251088 226646 251140 226652
rect 250720 224120 250772 224126
rect 250720 224062 250772 224068
rect 251088 221400 251140 221406
rect 251088 221342 251140 221348
rect 251100 217410 251128 221342
rect 252020 217410 252048 227394
rect 252204 224942 252232 231676
rect 252192 224936 252244 224942
rect 252192 224878 252244 224884
rect 252480 223990 252508 231676
rect 252468 223984 252520 223990
rect 252468 223926 252520 223932
rect 252848 222222 252876 231676
rect 252928 227180 252980 227186
rect 252928 227122 252980 227128
rect 252940 223378 252968 227122
rect 252928 223372 252980 223378
rect 252928 223314 252980 223320
rect 253216 222290 253244 231676
rect 253584 225350 253612 231676
rect 253664 227724 253716 227730
rect 253664 227666 253716 227672
rect 253572 225344 253624 225350
rect 253572 225286 253624 225292
rect 253204 222284 253256 222290
rect 253204 222226 253256 222232
rect 252836 222216 252888 222222
rect 252836 222158 252888 222164
rect 252928 221264 252980 221270
rect 252928 221206 252980 221212
rect 252940 217410 252968 221206
rect 253676 217410 253704 227666
rect 253756 227316 253808 227322
rect 253756 227258 253808 227264
rect 253768 223582 253796 227258
rect 253952 225690 253980 231676
rect 254320 227798 254348 231676
rect 254688 227934 254716 231676
rect 254676 227928 254728 227934
rect 254676 227870 254728 227876
rect 254308 227792 254360 227798
rect 254308 227734 254360 227740
rect 254676 226364 254728 226370
rect 254676 226306 254728 226312
rect 253940 225684 253992 225690
rect 253940 225626 253992 225632
rect 253756 223576 253808 223582
rect 253756 223518 253808 223524
rect 254688 222970 254716 226306
rect 255056 225010 255084 231676
rect 255332 228002 255360 231676
rect 255320 227996 255372 228002
rect 255320 227938 255372 227944
rect 255228 227112 255280 227118
rect 255228 227054 255280 227060
rect 255044 225004 255096 225010
rect 255044 224946 255096 224952
rect 254676 222964 254728 222970
rect 254676 222906 254728 222912
rect 254584 222284 254636 222290
rect 254584 222226 254636 222232
rect 254596 217410 254624 222226
rect 255240 221338 255268 227054
rect 255596 226976 255648 226982
rect 255596 226918 255648 226924
rect 255412 226840 255464 226846
rect 255412 226782 255464 226788
rect 255424 223038 255452 226782
rect 255608 223242 255636 226918
rect 255596 223236 255648 223242
rect 255596 223178 255648 223184
rect 255412 223032 255464 223038
rect 255412 222974 255464 222980
rect 255700 222426 255728 231676
rect 256068 222494 256096 231676
rect 256148 227792 256200 227798
rect 256148 227734 256200 227740
rect 256056 222488 256108 222494
rect 256056 222430 256108 222436
rect 255688 222420 255740 222426
rect 255688 222362 255740 222368
rect 255412 222216 255464 222222
rect 255412 222158 255464 222164
rect 255228 221332 255280 221338
rect 255228 221274 255280 221280
rect 255424 217410 255452 222158
rect 256160 222086 256188 227734
rect 256436 225078 256464 231676
rect 256698 228984 256754 228993
rect 256698 228919 256754 228928
rect 256608 227928 256660 227934
rect 256608 227870 256660 227876
rect 256424 225072 256476 225078
rect 256424 225014 256476 225020
rect 256148 222080 256200 222086
rect 256148 222022 256200 222028
rect 256620 221406 256648 227870
rect 256712 222698 256740 228919
rect 256804 226642 256832 231676
rect 256976 229084 257028 229090
rect 256976 229026 257028 229032
rect 256792 226636 256844 226642
rect 256792 226578 256844 226584
rect 256988 222834 257016 229026
rect 257172 227866 257200 231676
rect 257160 227860 257212 227866
rect 257160 227802 257212 227808
rect 257068 222896 257120 222902
rect 257068 222838 257120 222844
rect 256976 222828 257028 222834
rect 256976 222770 257028 222776
rect 256700 222692 256752 222698
rect 256700 222634 256752 222640
rect 256608 221400 256660 221406
rect 256608 221342 256660 221348
rect 256240 221332 256292 221338
rect 256240 221274 256292 221280
rect 256252 217410 256280 221274
rect 257080 217410 257108 222838
rect 257540 222562 257568 231676
rect 257712 227996 257764 228002
rect 257712 227938 257764 227944
rect 257528 222556 257580 222562
rect 257528 222498 257580 222504
rect 257724 221474 257752 227938
rect 257908 225146 257936 231676
rect 258184 228818 258212 231676
rect 258172 228812 258224 228818
rect 258172 228754 258224 228760
rect 258264 228812 258316 228818
rect 258264 228754 258316 228760
rect 257896 225140 257948 225146
rect 257896 225082 257948 225088
rect 257896 222488 257948 222494
rect 257896 222430 257948 222436
rect 257712 221468 257764 221474
rect 257712 221410 257764 221416
rect 257908 217410 257936 222430
rect 258276 221270 258304 228754
rect 258448 226908 258500 226914
rect 258448 226850 258500 226856
rect 258264 221264 258316 221270
rect 258264 221206 258316 221212
rect 258460 221202 258488 226850
rect 258552 226506 258580 231676
rect 258540 226500 258592 226506
rect 258540 226442 258592 226448
rect 258920 222630 258948 231676
rect 259288 225214 259316 231676
rect 259656 228585 259684 231676
rect 259642 228576 259698 228585
rect 259642 228511 259698 228520
rect 259644 227860 259696 227866
rect 259644 227802 259696 227808
rect 259368 226704 259420 226710
rect 259368 226646 259420 226652
rect 259276 225208 259328 225214
rect 259276 225150 259328 225156
rect 259380 223174 259408 226646
rect 259368 223168 259420 223174
rect 259368 223110 259420 223116
rect 258908 222624 258960 222630
rect 258908 222566 258960 222572
rect 259368 222352 259420 222358
rect 259368 222294 259420 222300
rect 258816 221604 258868 221610
rect 258816 221546 258868 221552
rect 258448 221196 258500 221202
rect 258448 221138 258500 221144
rect 258828 217410 258856 221546
rect 259380 217410 259408 222294
rect 259656 221338 259684 227802
rect 260024 227633 260052 231676
rect 260392 227769 260420 231676
rect 260378 227760 260434 227769
rect 260378 227695 260434 227704
rect 260010 227624 260066 227633
rect 260010 227559 260066 227568
rect 260760 225282 260788 231676
rect 261036 228070 261064 231676
rect 261404 228857 261432 231676
rect 261772 228993 261800 231676
rect 261758 228984 261814 228993
rect 261758 228919 261814 228928
rect 261390 228848 261446 228857
rect 261390 228783 261446 228792
rect 261024 228064 261076 228070
rect 261024 228006 261076 228012
rect 262140 225554 262168 231676
rect 262508 228449 262536 231676
rect 262494 228440 262550 228449
rect 262494 228375 262550 228384
rect 262876 227905 262904 231676
rect 263244 228177 263272 231676
rect 263230 228168 263286 228177
rect 263230 228103 263286 228112
rect 262862 227896 262918 227905
rect 262862 227831 262918 227840
rect 262128 225548 262180 225554
rect 262128 225490 262180 225496
rect 263612 225486 263640 231676
rect 263888 228138 263916 231676
rect 263876 228132 263928 228138
rect 263876 228074 263928 228080
rect 264256 228041 264284 231676
rect 264624 229090 264652 231676
rect 264612 229084 264664 229090
rect 264612 229026 264664 229032
rect 264704 229084 264756 229090
rect 264704 229026 264756 229032
rect 264242 228032 264298 228041
rect 264242 227967 264298 227976
rect 264716 226574 264744 229026
rect 264704 226568 264756 226574
rect 264704 226510 264756 226516
rect 263600 225480 263652 225486
rect 263600 225422 263652 225428
rect 264992 225418 265020 231676
rect 265360 229022 265388 231676
rect 265348 229016 265400 229022
rect 265348 228958 265400 228964
rect 265728 227050 265756 231676
rect 266096 228313 266124 231676
rect 266082 228304 266138 228313
rect 266082 228239 266138 228248
rect 265716 227044 265768 227050
rect 265716 226986 265768 226992
rect 266464 225622 266492 231676
rect 266740 228886 266768 231676
rect 266728 228880 266780 228886
rect 266728 228822 266780 228828
rect 267108 228274 267136 231676
rect 267476 228410 267504 231676
rect 267464 228404 267516 228410
rect 267464 228346 267516 228352
rect 267096 228268 267148 228274
rect 267096 228210 267148 228216
rect 267844 228206 267872 231676
rect 268212 228614 268240 231676
rect 268200 228608 268252 228614
rect 268200 228550 268252 228556
rect 267832 228200 267884 228206
rect 267832 228142 267884 228148
rect 268580 227390 268608 231676
rect 268568 227384 268620 227390
rect 268568 227326 268620 227332
rect 268948 226370 268976 231676
rect 269316 228478 269344 231676
rect 269592 228954 269620 231676
rect 269580 228948 269632 228954
rect 269580 228890 269632 228896
rect 269304 228472 269356 228478
rect 269304 228414 269356 228420
rect 269960 227254 269988 231676
rect 269948 227248 270000 227254
rect 269948 227190 270000 227196
rect 270328 226846 270356 231676
rect 270696 228342 270724 231676
rect 271064 228546 271092 231676
rect 271052 228540 271104 228546
rect 271052 228482 271104 228488
rect 270684 228336 270736 228342
rect 270684 228278 270736 228284
rect 271432 227186 271460 231676
rect 271420 227180 271472 227186
rect 271420 227122 271472 227128
rect 271800 226982 271828 231676
rect 272168 228750 272196 231676
rect 272156 228744 272208 228750
rect 272156 228686 272208 228692
rect 272444 227662 272472 231676
rect 272432 227656 272484 227662
rect 272432 227598 272484 227604
rect 272812 227322 272840 231676
rect 272800 227316 272852 227322
rect 272800 227258 272852 227264
rect 271788 226976 271840 226982
rect 271788 226918 271840 226924
rect 270316 226840 270368 226846
rect 270316 226782 270368 226788
rect 273180 226710 273208 231676
rect 273548 228682 273576 231676
rect 273916 229090 273944 231676
rect 273904 229084 273956 229090
rect 273904 229026 273956 229032
rect 273536 228676 273588 228682
rect 273536 228618 273588 228624
rect 274284 227798 274312 231676
rect 274272 227792 274324 227798
rect 274272 227734 274324 227740
rect 274652 226914 274680 231676
rect 275020 227526 275048 231676
rect 275296 227594 275324 231676
rect 275284 227588 275336 227594
rect 275284 227530 275336 227536
rect 275008 227520 275060 227526
rect 275008 227462 275060 227468
rect 275664 227118 275692 231676
rect 276032 228002 276060 231676
rect 276020 227996 276072 228002
rect 276020 227938 276072 227944
rect 276400 227458 276428 231676
rect 276768 227730 276796 231676
rect 277136 227934 277164 231676
rect 277504 228818 277532 231676
rect 277492 228812 277544 228818
rect 277492 228754 277544 228760
rect 277124 227928 277176 227934
rect 277124 227870 277176 227876
rect 276756 227724 276808 227730
rect 276756 227666 276808 227672
rect 276388 227452 276440 227458
rect 276388 227394 276440 227400
rect 275652 227112 275704 227118
rect 275652 227054 275704 227060
rect 274640 226908 274692 226914
rect 274640 226850 274692 226856
rect 273168 226704 273220 226710
rect 273168 226646 273220 226652
rect 268936 226364 268988 226370
rect 268936 226306 268988 226312
rect 266452 225616 266504 225622
rect 266452 225558 266504 225564
rect 264980 225412 265032 225418
rect 264980 225354 265032 225360
rect 260748 225276 260800 225282
rect 260748 225218 260800 225224
rect 273076 223372 273128 223378
rect 273076 223314 273128 223320
rect 271420 223100 271472 223106
rect 271420 223042 271472 223048
rect 263784 222964 263836 222970
rect 263784 222906 263836 222912
rect 261300 222828 261352 222834
rect 261300 222770 261352 222776
rect 260472 222692 260524 222698
rect 260472 222634 260524 222640
rect 259644 221332 259696 221338
rect 259644 221274 259696 221280
rect 260484 217410 260512 222634
rect 261312 217410 261340 222770
rect 262956 222624 263008 222630
rect 262956 222566 263008 222572
rect 262128 222556 262180 222562
rect 262128 222498 262180 222504
rect 262140 217410 262168 222498
rect 262968 217410 262996 222566
rect 263796 217410 263824 222906
rect 266360 222760 266412 222766
rect 266360 222702 266412 222708
rect 264612 221672 264664 221678
rect 264612 221614 264664 221620
rect 264624 217410 264652 221614
rect 265532 221060 265584 221066
rect 265532 221002 265584 221008
rect 265544 217410 265572 221002
rect 266372 217410 266400 222702
rect 269672 222148 269724 222154
rect 269672 222090 269724 222096
rect 268844 221468 268896 221474
rect 268844 221410 268896 221416
rect 267188 221400 267240 221406
rect 267188 221342 267240 221348
rect 267200 217410 267228 221342
rect 268016 220992 268068 220998
rect 268016 220934 268068 220940
rect 268028 217410 268056 220934
rect 268856 217410 268884 221410
rect 269684 217410 269712 222090
rect 270408 221264 270460 221270
rect 270408 221206 270460 221212
rect 270420 217410 270448 221206
rect 271432 217410 271460 223042
rect 272248 222420 272300 222426
rect 272248 222362 272300 222368
rect 272260 217410 272288 222362
rect 273088 217410 273116 223314
rect 274732 223168 274784 223174
rect 274732 223110 274784 223116
rect 273904 221536 273956 221542
rect 273904 221478 273956 221484
rect 273916 217410 273944 221478
rect 274744 217410 274772 223110
rect 277872 222222 277900 231676
rect 278148 222902 278176 231676
rect 278136 222896 278188 222902
rect 278136 222838 278188 222844
rect 278516 222290 278544 231676
rect 278884 227866 278912 231676
rect 278872 227860 278924 227866
rect 278872 227802 278924 227808
rect 278688 223576 278740 223582
rect 278688 223518 278740 223524
rect 278504 222284 278556 222290
rect 278504 222226 278556 222232
rect 277860 222216 277912 222222
rect 277860 222158 277912 222164
rect 275560 221944 275612 221950
rect 275560 221886 275612 221892
rect 275572 217410 275600 221886
rect 278136 221808 278188 221814
rect 278136 221750 278188 221756
rect 276480 221196 276532 221202
rect 276480 221138 276532 221144
rect 276492 217410 276520 221138
rect 277308 221128 277360 221134
rect 277308 221070 277360 221076
rect 277320 217410 277348 221070
rect 278148 217410 278176 221750
rect 278700 217410 278728 223518
rect 279252 221610 279280 231676
rect 279620 222698 279648 231676
rect 279608 222692 279660 222698
rect 279608 222634 279660 222640
rect 279988 222494 280016 231676
rect 279976 222488 280028 222494
rect 279976 222430 280028 222436
rect 280356 222358 280384 231676
rect 280724 222562 280752 231676
rect 281000 222970 281028 231676
rect 280988 222964 281040 222970
rect 280988 222906 281040 222912
rect 281368 222834 281396 231676
rect 281356 222828 281408 222834
rect 281356 222770 281408 222776
rect 281736 222630 281764 231676
rect 281724 222624 281776 222630
rect 281724 222566 281776 222572
rect 280712 222556 280764 222562
rect 280712 222498 280764 222504
rect 280344 222352 280396 222358
rect 280344 222294 280396 222300
rect 281448 221740 281500 221746
rect 281448 221682 281500 221688
rect 279240 221604 279292 221610
rect 279240 221546 279292 221552
rect 280620 221332 280672 221338
rect 280620 221274 280672 221280
rect 279792 220924 279844 220930
rect 279792 220866 279844 220872
rect 279804 217410 279832 220866
rect 280632 217410 280660 221274
rect 281460 217410 281488 221682
rect 282104 221066 282132 231676
rect 282472 221406 282500 231676
rect 282840 221678 282868 231676
rect 283208 222766 283236 231676
rect 283196 222760 283248 222766
rect 283196 222702 283248 222708
rect 283196 222556 283248 222562
rect 283196 222498 283248 222504
rect 282828 221672 282880 221678
rect 282828 221614 282880 221620
rect 282460 221400 282512 221406
rect 282460 221342 282512 221348
rect 282092 221060 282144 221066
rect 282092 221002 282144 221008
rect 282368 221060 282420 221066
rect 282368 221002 282420 221008
rect 282380 217410 282408 221002
rect 283208 217410 283236 222498
rect 283576 221474 283604 231676
rect 283564 221468 283616 221474
rect 283564 221410 283616 221416
rect 283852 221270 283880 231676
rect 283932 221604 283984 221610
rect 283932 221546 283984 221552
rect 283840 221264 283892 221270
rect 283840 221206 283892 221212
rect 283944 217410 283972 221546
rect 284220 220998 284248 231676
rect 284588 222154 284616 231676
rect 284956 222630 284984 231676
rect 284944 222624 284996 222630
rect 284944 222566 284996 222572
rect 284576 222148 284628 222154
rect 284576 222090 284628 222096
rect 285324 221542 285352 231676
rect 285692 222902 285720 231676
rect 286060 223378 286088 231676
rect 286048 223372 286100 223378
rect 286048 223314 286100 223320
rect 285680 222896 285732 222902
rect 285680 222838 285732 222844
rect 286428 221950 286456 231676
rect 286416 221944 286468 221950
rect 286416 221886 286468 221892
rect 285312 221536 285364 221542
rect 285312 221478 285364 221484
rect 286508 221536 286560 221542
rect 286508 221478 286560 221484
rect 284852 221264 284904 221270
rect 284852 221206 284904 221212
rect 284208 220992 284260 220998
rect 284208 220934 284260 220940
rect 284864 217410 284892 221206
rect 285680 220992 285732 220998
rect 285680 220934 285732 220940
rect 285692 217410 285720 220934
rect 286520 217410 286548 221478
rect 286704 221134 286732 231676
rect 287072 223174 287100 231676
rect 287060 223168 287112 223174
rect 287060 223110 287112 223116
rect 287440 221202 287468 231676
rect 287808 223582 287836 231676
rect 287796 223576 287848 223582
rect 287796 223518 287848 223524
rect 288176 221338 288204 231676
rect 288544 221814 288572 231676
rect 288532 221808 288584 221814
rect 288532 221750 288584 221756
rect 288256 221468 288308 221474
rect 288256 221410 288308 221416
rect 288164 221332 288216 221338
rect 288164 221274 288216 221280
rect 287428 221196 287480 221202
rect 287428 221138 287480 221144
rect 286692 221128 286744 221134
rect 286692 221070 286744 221076
rect 287336 221060 287388 221066
rect 287336 221002 287388 221008
rect 287348 217410 287376 221002
rect 288268 217410 288296 221410
rect 288912 220930 288940 231676
rect 289084 221400 289136 221406
rect 289084 221342 289136 221348
rect 288900 220924 288952 220930
rect 288900 220866 288952 220872
rect 289096 217410 289124 221342
rect 289280 221134 289308 231676
rect 289556 221610 289584 231676
rect 289924 221746 289952 231676
rect 290292 222562 290320 231676
rect 290280 222556 290332 222562
rect 290280 222498 290332 222504
rect 289912 221740 289964 221746
rect 289912 221682 289964 221688
rect 289544 221604 289596 221610
rect 289544 221546 289596 221552
rect 289728 221332 289780 221338
rect 289728 221274 289780 221280
rect 289268 221128 289320 221134
rect 289268 221070 289320 221076
rect 289740 217410 289768 221274
rect 290660 220998 290688 231676
rect 290740 229016 290792 229022
rect 290740 228958 290792 228964
rect 290648 220992 290700 220998
rect 290648 220934 290700 220940
rect 290752 217410 290780 228958
rect 291028 221066 291056 231676
rect 291396 221270 291424 231676
rect 291764 221542 291792 231676
rect 291752 221536 291804 221542
rect 291752 221478 291804 221484
rect 292132 221406 292160 231676
rect 292408 229022 292436 231676
rect 292396 229016 292448 229022
rect 292396 228958 292448 228964
rect 292776 221474 292804 231676
rect 292764 221468 292816 221474
rect 292764 221410 292816 221416
rect 292120 221400 292172 221406
rect 292120 221342 292172 221348
rect 292396 221400 292448 221406
rect 292396 221342 292448 221348
rect 291384 221264 291436 221270
rect 291384 221206 291436 221212
rect 291568 221264 291620 221270
rect 291568 221206 291620 221212
rect 291016 221060 291068 221066
rect 291016 221002 291068 221008
rect 291580 217410 291608 221206
rect 292408 217410 292436 221342
rect 293144 221338 293172 231676
rect 293224 229016 293276 229022
rect 293224 228958 293276 228964
rect 293132 221332 293184 221338
rect 293132 221274 293184 221280
rect 293236 217410 293264 228958
rect 293512 221406 293540 231676
rect 293500 221400 293552 221406
rect 293500 221342 293552 221348
rect 293880 217410 293908 231676
rect 294248 221270 294276 231676
rect 294616 229022 294644 231676
rect 294998 231662 295196 231690
rect 294604 229016 294656 229022
rect 294604 228958 294656 228964
rect 295168 226334 295196 231662
rect 295260 227322 295288 231676
rect 295248 227316 295300 227322
rect 295248 227258 295300 227264
rect 295168 226306 295380 226334
rect 294972 221332 295024 221338
rect 294972 221274 295024 221280
rect 294236 221264 294288 221270
rect 294236 221206 294288 221212
rect 294984 217410 295012 221274
rect 214728 217382 215064 217410
rect 215556 217382 215892 217410
rect 216384 217382 216720 217410
rect 217304 217382 217640 217410
rect 218132 217382 218468 217410
rect 218960 217382 219296 217410
rect 219788 217382 220124 217410
rect 220616 217382 220768 217410
rect 221444 217382 221780 217410
rect 222272 217382 222608 217410
rect 223192 217382 223528 217410
rect 224020 217382 224356 217410
rect 224848 217382 225184 217410
rect 225676 217382 226012 217410
rect 226504 217382 226840 217410
rect 227332 217382 227668 217410
rect 228160 217382 228496 217410
rect 229080 217382 229324 217410
rect 229908 217382 230244 217410
rect 230736 217382 231072 217410
rect 231564 217382 231716 217410
rect 232392 217382 232728 217410
rect 233220 217382 233556 217410
rect 234048 217382 234384 217410
rect 234968 217382 235304 217410
rect 235796 217382 236132 217410
rect 236624 217382 236960 217410
rect 237452 217382 237788 217410
rect 238280 217382 238616 217410
rect 239108 217382 239444 217410
rect 239936 217382 240088 217410
rect 240856 217382 241192 217410
rect 241684 217382 242020 217410
rect 242512 217382 242848 217410
rect 243340 217382 243676 217410
rect 244168 217382 244504 217410
rect 244996 217382 245332 217410
rect 245824 217382 246160 217410
rect 246744 217382 247080 217410
rect 247572 217382 247908 217410
rect 248400 217382 248736 217410
rect 249228 217382 249564 217410
rect 250056 217382 250392 217410
rect 250884 217382 251128 217410
rect 251712 217382 252048 217410
rect 252632 217382 252968 217410
rect 253460 217382 253704 217410
rect 254288 217382 254624 217410
rect 255116 217382 255452 217410
rect 255944 217382 256280 217410
rect 256772 217382 257108 217410
rect 257600 217382 257936 217410
rect 258520 217382 258856 217410
rect 259348 217382 259408 217410
rect 260176 217382 260512 217410
rect 261004 217382 261340 217410
rect 261832 217382 262168 217410
rect 262660 217382 262996 217410
rect 263488 217382 263824 217410
rect 264408 217382 264652 217410
rect 265236 217382 265572 217410
rect 266064 217382 266400 217410
rect 266892 217382 267228 217410
rect 267720 217382 268056 217410
rect 268548 217382 268884 217410
rect 269376 217382 269712 217410
rect 270296 217382 270448 217410
rect 271124 217382 271460 217410
rect 271952 217382 272288 217410
rect 272780 217382 273116 217410
rect 273608 217382 273944 217410
rect 274436 217382 274772 217410
rect 275264 217382 275600 217410
rect 276184 217382 276520 217410
rect 277012 217382 277348 217410
rect 277840 217382 278176 217410
rect 278668 217382 278728 217410
rect 279496 217382 279832 217410
rect 280324 217382 280660 217410
rect 281152 217382 281488 217410
rect 282072 217382 282408 217410
rect 282900 217382 283236 217410
rect 283728 217382 283972 217410
rect 284556 217382 284892 217410
rect 285384 217382 285720 217410
rect 286212 217382 286548 217410
rect 287040 217382 287376 217410
rect 287960 217382 288296 217410
rect 288788 217382 289124 217410
rect 289616 217382 289768 217410
rect 290444 217382 290780 217410
rect 291272 217382 291608 217410
rect 292100 217382 292436 217410
rect 292928 217382 293264 217410
rect 293848 217382 293908 217410
rect 294676 217382 295012 217410
rect 295352 217410 295380 226306
rect 295628 221338 295656 231676
rect 295616 221332 295668 221338
rect 295616 221274 295668 221280
rect 295996 217410 296024 231676
rect 296364 229090 296392 231676
rect 296352 229084 296404 229090
rect 296352 229026 296404 229032
rect 296732 228274 296760 231676
rect 297114 231662 297404 231690
rect 296720 228268 296772 228274
rect 296720 228210 296772 228216
rect 296812 227316 296864 227322
rect 296812 227258 296864 227264
rect 296824 217410 296852 227258
rect 297376 226334 297404 231662
rect 297468 229022 297496 231676
rect 297456 229016 297508 229022
rect 297456 228958 297508 228964
rect 297836 227322 297864 231676
rect 297824 227316 297876 227322
rect 297824 227258 297876 227264
rect 298112 226710 298140 231676
rect 298494 231662 298784 231690
rect 298468 229084 298520 229090
rect 298468 229026 298520 229032
rect 298100 226704 298152 226710
rect 298100 226646 298152 226652
rect 297376 226306 297588 226334
rect 297560 217410 297588 226306
rect 298480 217410 298508 229026
rect 298756 228410 298784 231662
rect 298848 228750 298876 231676
rect 298836 228744 298888 228750
rect 298836 228686 298888 228692
rect 298744 228404 298796 228410
rect 298744 228346 298796 228352
rect 299216 226778 299244 231676
rect 299388 229016 299440 229022
rect 299388 228958 299440 228964
rect 299204 226772 299256 226778
rect 299204 226714 299256 226720
rect 299400 217410 299428 228958
rect 299584 226846 299612 231676
rect 299572 226840 299624 226846
rect 299572 226782 299624 226788
rect 299952 226370 299980 231676
rect 300216 228268 300268 228274
rect 300216 228210 300268 228216
rect 299940 226364 299992 226370
rect 299940 226306 299992 226312
rect 300228 217410 300256 228210
rect 300320 226642 300348 231676
rect 300688 226914 300716 231676
rect 300964 227390 300992 231676
rect 301044 228404 301096 228410
rect 301044 228346 301096 228352
rect 300952 227384 301004 227390
rect 300952 227326 301004 227332
rect 300676 226908 300728 226914
rect 300676 226850 300728 226856
rect 300308 226636 300360 226642
rect 300308 226578 300360 226584
rect 301056 217410 301084 228346
rect 301332 226574 301360 231676
rect 301700 227934 301728 231676
rect 301688 227928 301740 227934
rect 301688 227870 301740 227876
rect 302068 227798 302096 231676
rect 302056 227792 302108 227798
rect 302056 227734 302108 227740
rect 302436 227390 302464 231676
rect 302700 228744 302752 228750
rect 302700 228686 302752 228692
rect 302424 227384 302476 227390
rect 302424 227326 302476 227332
rect 301872 227316 301924 227322
rect 301872 227258 301924 227264
rect 301320 226568 301372 226574
rect 301320 226510 301372 226516
rect 301884 217410 301912 227258
rect 302712 217410 302740 228686
rect 302804 228274 302832 231676
rect 302792 228268 302844 228274
rect 302792 228210 302844 228216
rect 303172 228002 303200 231676
rect 303160 227996 303212 228002
rect 303160 227938 303212 227944
rect 303540 227254 303568 231676
rect 303528 227248 303580 227254
rect 303528 227190 303580 227196
rect 303620 226704 303672 226710
rect 303620 226646 303672 226652
rect 303632 217410 303660 226646
rect 303816 226506 303844 231676
rect 304184 229022 304212 231676
rect 304172 229016 304224 229022
rect 304172 228958 304224 228964
rect 304552 228954 304580 231676
rect 304540 228948 304592 228954
rect 304540 228890 304592 228896
rect 303804 226500 303856 226506
rect 303804 226442 303856 226448
rect 304920 226438 304948 231676
rect 305288 228750 305316 231676
rect 305656 228886 305684 231676
rect 305644 228880 305696 228886
rect 305644 228822 305696 228828
rect 306024 228818 306052 231676
rect 306012 228812 306064 228818
rect 306012 228754 306064 228760
rect 305276 228744 305328 228750
rect 305276 228686 305328 228692
rect 306392 227458 306420 231676
rect 306668 229090 306696 231676
rect 306656 229084 306708 229090
rect 306656 229026 306708 229032
rect 307036 227594 307064 231676
rect 307404 228614 307432 231676
rect 307392 228608 307444 228614
rect 307392 228550 307444 228556
rect 307772 228546 307800 231676
rect 307760 228540 307812 228546
rect 307760 228482 307812 228488
rect 308140 228410 308168 231676
rect 308128 228404 308180 228410
rect 308128 228346 308180 228352
rect 308508 227662 308536 231676
rect 308876 228682 308904 231676
rect 308864 228676 308916 228682
rect 308864 228618 308916 228624
rect 309244 228206 309272 231676
rect 309520 228342 309548 231676
rect 309508 228336 309560 228342
rect 309508 228278 309560 228284
rect 309232 228200 309284 228206
rect 309232 228142 309284 228148
rect 309416 227928 309468 227934
rect 309416 227870 309468 227876
rect 308496 227656 308548 227662
rect 308496 227598 308548 227604
rect 307024 227588 307076 227594
rect 307024 227530 307076 227536
rect 306380 227452 306432 227458
rect 306380 227394 306432 227400
rect 308588 226908 308640 226914
rect 308588 226850 308640 226856
rect 306932 226840 306984 226846
rect 306932 226782 306984 226788
rect 305276 226772 305328 226778
rect 305276 226714 305328 226720
rect 304908 226432 304960 226438
rect 304908 226374 304960 226380
rect 304356 226364 304408 226370
rect 304356 226306 304408 226312
rect 304368 217410 304396 226306
rect 305288 217410 305316 226714
rect 306380 226636 306432 226642
rect 306380 226578 306432 226584
rect 306392 217410 306420 226578
rect 306944 217410 306972 226782
rect 307760 226568 307812 226574
rect 307760 226510 307812 226516
rect 307772 217410 307800 226510
rect 308600 217410 308628 226850
rect 309428 217410 309456 227870
rect 309888 226370 309916 231676
rect 310256 228478 310284 231676
rect 310244 228472 310296 228478
rect 310244 228414 310296 228420
rect 310624 227934 310652 231676
rect 310612 227928 310664 227934
rect 310612 227870 310664 227876
rect 310244 227316 310296 227322
rect 310244 227258 310296 227264
rect 309876 226364 309928 226370
rect 309876 226306 309928 226312
rect 310256 217410 310284 227258
rect 310992 222358 311020 231676
rect 311164 228268 311216 228274
rect 311164 228210 311216 228216
rect 310980 222352 311032 222358
rect 310980 222294 311032 222300
rect 311176 217410 311204 228210
rect 311360 228070 311388 231676
rect 311728 228138 311756 231676
rect 311716 228132 311768 228138
rect 311716 228074 311768 228080
rect 311348 228064 311400 228070
rect 311348 228006 311400 228012
rect 311992 227792 312044 227798
rect 311992 227734 312044 227740
rect 312004 217410 312032 227734
rect 312096 227050 312124 231676
rect 312084 227044 312136 227050
rect 312084 226986 312136 226992
rect 312372 221270 312400 231676
rect 312740 227798 312768 231676
rect 312820 227996 312872 228002
rect 312820 227938 312872 227944
rect 312728 227792 312780 227798
rect 312728 227734 312780 227740
rect 312360 221264 312412 221270
rect 312360 221206 312412 221212
rect 312832 217410 312860 227938
rect 313108 221134 313136 231676
rect 313476 225282 313504 231676
rect 313648 227384 313700 227390
rect 313648 227326 313700 227332
rect 313464 225276 313516 225282
rect 313464 225218 313516 225224
rect 313096 221128 313148 221134
rect 313096 221070 313148 221076
rect 313660 217410 313688 227326
rect 313844 221406 313872 231676
rect 314212 222222 314240 231676
rect 314200 222216 314252 222222
rect 314200 222158 314252 222164
rect 314580 221542 314608 231676
rect 314660 229016 314712 229022
rect 314660 228958 314712 228964
rect 314568 221536 314620 221542
rect 314568 221478 314620 221484
rect 313832 221400 313884 221406
rect 313832 221342 313884 221348
rect 314672 217410 314700 228958
rect 314948 225214 314976 231676
rect 314936 225208 314988 225214
rect 314936 225150 314988 225156
rect 315224 221474 315252 231676
rect 315304 227248 315356 227254
rect 315304 227190 315356 227196
rect 315212 221468 315264 221474
rect 315212 221410 315264 221416
rect 315316 217410 315344 227190
rect 315592 221338 315620 231676
rect 315960 227866 315988 231676
rect 316132 228948 316184 228954
rect 316132 228890 316184 228896
rect 315948 227860 316000 227866
rect 315948 227802 316000 227808
rect 315580 221332 315632 221338
rect 315580 221274 315632 221280
rect 316144 217410 316172 228890
rect 316224 228676 316276 228682
rect 316224 228618 316276 228624
rect 316236 228206 316264 228618
rect 316224 228200 316276 228206
rect 316224 228142 316276 228148
rect 316328 225078 316356 231676
rect 316316 225072 316368 225078
rect 316316 225014 316368 225020
rect 316696 221950 316724 231676
rect 316684 221944 316736 221950
rect 316684 221886 316736 221892
rect 317064 221678 317092 231676
rect 317432 227118 317460 231676
rect 317420 227112 317472 227118
rect 317420 227054 317472 227060
rect 317420 226500 317472 226506
rect 317420 226442 317472 226448
rect 317052 221672 317104 221678
rect 317052 221614 317104 221620
rect 317432 217410 317460 226442
rect 317800 225146 317828 231676
rect 317880 228880 317932 228886
rect 317880 228822 317932 228828
rect 317788 225140 317840 225146
rect 317788 225082 317840 225088
rect 295352 217382 295504 217410
rect 295996 217382 296332 217410
rect 296824 217382 297160 217410
rect 297560 217382 297988 217410
rect 298480 217382 298816 217410
rect 299400 217382 299736 217410
rect 300228 217382 300564 217410
rect 301056 217382 301392 217410
rect 301884 217382 302220 217410
rect 302712 217382 303048 217410
rect 303632 217382 303876 217410
rect 304368 217382 304704 217410
rect 305288 217382 305624 217410
rect 306392 217382 306452 217410
rect 306944 217382 307280 217410
rect 307772 217382 308108 217410
rect 308600 217382 308936 217410
rect 309428 217382 309764 217410
rect 310256 217382 310592 217410
rect 311176 217382 311512 217410
rect 312004 217382 312340 217410
rect 312832 217382 313168 217410
rect 313660 217382 313996 217410
rect 314672 217382 314824 217410
rect 315316 217382 315652 217410
rect 316144 217382 316480 217410
rect 317400 217382 317460 217410
rect 317892 217410 317920 228822
rect 318076 221746 318104 231676
rect 318064 221740 318116 221746
rect 318064 221682 318116 221688
rect 318444 221610 318472 231676
rect 318812 227798 318840 231676
rect 318800 227792 318852 227798
rect 318800 227734 318852 227740
rect 318708 226432 318760 226438
rect 318708 226374 318760 226380
rect 318432 221604 318484 221610
rect 318432 221546 318484 221552
rect 318720 217410 318748 226374
rect 319180 225010 319208 231676
rect 319562 231662 319852 231690
rect 319536 228812 319588 228818
rect 319536 228754 319588 228760
rect 319168 225004 319220 225010
rect 319168 224946 319220 224952
rect 319548 217410 319576 228754
rect 319824 222086 319852 231662
rect 319812 222080 319864 222086
rect 319812 222022 319864 222028
rect 319916 221814 319944 231676
rect 320284 227730 320312 231676
rect 320364 228744 320416 228750
rect 320364 228686 320416 228692
rect 320272 227724 320324 227730
rect 320272 227666 320324 227672
rect 319904 221808 319956 221814
rect 319904 221750 319956 221756
rect 320376 217410 320404 228686
rect 320652 227526 320680 231676
rect 320640 227520 320692 227526
rect 320640 227462 320692 227468
rect 320928 222154 320956 231676
rect 321192 227588 321244 227594
rect 321192 227530 321244 227536
rect 320916 222148 320968 222154
rect 320916 222090 320968 222096
rect 321204 217410 321232 227530
rect 321296 221882 321324 231676
rect 321664 229022 321692 231676
rect 321652 229016 321704 229022
rect 321652 228958 321704 228964
rect 322032 228750 322060 231676
rect 322020 228744 322072 228750
rect 322020 228686 322072 228692
rect 322020 227452 322072 227458
rect 322020 227394 322072 227400
rect 321284 221876 321336 221882
rect 321284 221818 321336 221824
rect 322032 217410 322060 227394
rect 322400 223514 322428 231676
rect 322388 223508 322440 223514
rect 322388 223450 322440 223456
rect 322768 222018 322796 231676
rect 322940 228608 322992 228614
rect 322940 228550 322992 228556
rect 322756 222012 322808 222018
rect 322756 221954 322808 221960
rect 322952 217410 322980 228550
rect 323136 227458 323164 231676
rect 323124 227452 323176 227458
rect 323124 227394 323176 227400
rect 323504 226846 323532 231676
rect 323492 226840 323544 226846
rect 323492 226782 323544 226788
rect 323780 223446 323808 231676
rect 323860 229084 323912 229090
rect 323860 229026 323912 229032
rect 323768 223440 323820 223446
rect 323768 223382 323820 223388
rect 323872 217410 323900 229026
rect 324148 223582 324176 231676
rect 324136 223576 324188 223582
rect 324136 223518 324188 223524
rect 324516 223378 324544 231676
rect 324596 227656 324648 227662
rect 324596 227598 324648 227604
rect 324504 223372 324556 223378
rect 324504 223314 324556 223320
rect 324608 217410 324636 227598
rect 324884 223038 324912 231676
rect 324872 223032 324924 223038
rect 324872 222974 324924 222980
rect 325252 222834 325280 231676
rect 325620 223310 325648 231676
rect 325700 228540 325752 228546
rect 325700 228482 325752 228488
rect 325608 223304 325660 223310
rect 325608 223246 325660 223252
rect 325240 222828 325292 222834
rect 325240 222770 325292 222776
rect 325712 217410 325740 228482
rect 325988 227322 326016 231676
rect 326252 228200 326304 228206
rect 326252 228142 326304 228148
rect 325976 227316 326028 227322
rect 325976 227258 326028 227264
rect 326264 217410 326292 228142
rect 326356 223106 326384 231676
rect 326344 223100 326396 223106
rect 326344 223042 326396 223048
rect 326632 222970 326660 231676
rect 327000 223242 327028 231676
rect 327080 228404 327132 228410
rect 327080 228346 327132 228352
rect 326988 223236 327040 223242
rect 326988 223178 327040 223184
rect 326620 222964 326672 222970
rect 326620 222906 326672 222912
rect 327092 217410 327120 228346
rect 327368 222902 327396 231676
rect 327356 222896 327408 222902
rect 327356 222838 327408 222844
rect 327736 222494 327764 231676
rect 327908 226364 327960 226370
rect 327908 226306 327960 226312
rect 327724 222488 327776 222494
rect 327724 222430 327776 222436
rect 327920 217410 327948 226306
rect 328104 222766 328132 231676
rect 328472 223174 328500 231676
rect 328840 228682 328868 231676
rect 328828 228676 328880 228682
rect 328828 228618 328880 228624
rect 329208 228546 329236 231676
rect 329196 228540 329248 228546
rect 329196 228482 329248 228488
rect 328828 228268 328880 228274
rect 328828 228210 328880 228216
rect 328460 223168 328512 223174
rect 328460 223110 328512 223116
rect 328092 222760 328144 222766
rect 328092 222702 328144 222708
rect 328840 217410 328868 228210
rect 329484 222698 329512 231676
rect 329656 228472 329708 228478
rect 329656 228414 329708 228420
rect 329472 222692 329524 222698
rect 329472 222634 329524 222640
rect 329668 217410 329696 228414
rect 329852 222630 329880 231676
rect 329840 222624 329892 222630
rect 329840 222566 329892 222572
rect 330220 221202 330248 231676
rect 330484 228336 330536 228342
rect 330484 228278 330536 228284
rect 330208 221196 330260 221202
rect 330208 221138 330260 221144
rect 330496 217410 330524 228278
rect 330588 226506 330616 231676
rect 330576 226500 330628 226506
rect 330576 226442 330628 226448
rect 330956 223009 330984 231676
rect 331338 231662 331628 231690
rect 331312 228064 331364 228070
rect 331312 228006 331364 228012
rect 330942 223000 330998 223009
rect 330942 222935 330998 222944
rect 331324 217410 331352 228006
rect 331600 222562 331628 231662
rect 331692 226370 331720 231676
rect 332060 227390 332088 231676
rect 332140 227996 332192 228002
rect 332140 227938 332192 227944
rect 332048 227384 332100 227390
rect 332048 227326 332100 227332
rect 331680 226364 331732 226370
rect 331680 226306 331732 226312
rect 331588 222556 331640 222562
rect 331588 222498 331640 222504
rect 332152 217410 332180 227938
rect 332336 222601 332364 231676
rect 332322 222592 332378 222601
rect 332322 222527 332378 222536
rect 332704 222426 332732 231676
rect 332968 228132 333020 228138
rect 332968 228074 333020 228080
rect 332692 222420 332744 222426
rect 332692 222362 332744 222368
rect 332980 217410 333008 228074
rect 333072 222873 333100 231676
rect 333440 228410 333468 231676
rect 333428 228404 333480 228410
rect 333428 228346 333480 228352
rect 333058 222864 333114 222873
rect 333058 222799 333114 222808
rect 333808 222465 333836 231676
rect 333794 222456 333850 222465
rect 333794 222391 333850 222400
rect 334176 222358 334204 231676
rect 334544 222737 334572 231676
rect 334912 228342 334940 231676
rect 334900 228336 334952 228342
rect 334900 228278 334952 228284
rect 334716 227928 334768 227934
rect 334716 227870 334768 227876
rect 334530 222728 334586 222737
rect 334530 222663 334586 222672
rect 333980 222352 334032 222358
rect 333980 222294 334032 222300
rect 334164 222352 334216 222358
rect 334164 222294 334216 222300
rect 333992 217410 334020 222294
rect 334728 217410 334756 227870
rect 335188 224942 335216 231676
rect 335570 231662 335860 231690
rect 335544 227044 335596 227050
rect 335544 226986 335596 226992
rect 335176 224936 335228 224942
rect 335176 224878 335228 224884
rect 335556 217410 335584 226986
rect 335832 221921 335860 231662
rect 335924 222329 335952 231676
rect 336292 228138 336320 231676
rect 336660 228614 336688 231676
rect 336648 228608 336700 228614
rect 336648 228550 336700 228556
rect 337028 228274 337056 231676
rect 337016 228268 337068 228274
rect 337016 228210 337068 228216
rect 336280 228132 336332 228138
rect 336280 228074 336332 228080
rect 335910 222320 335966 222329
rect 337396 222290 337424 231676
rect 337764 228818 337792 231676
rect 338040 229090 338068 231676
rect 338028 229084 338080 229090
rect 338028 229026 338080 229032
rect 337752 228812 337804 228818
rect 337752 228754 337804 228760
rect 338408 228002 338436 231676
rect 338396 227996 338448 228002
rect 338396 227938 338448 227944
rect 338120 227860 338172 227866
rect 338120 227802 338172 227808
rect 337660 227112 337712 227118
rect 337660 227054 337712 227060
rect 335910 222255 335966 222264
rect 337384 222284 337436 222290
rect 337384 222226 337436 222232
rect 335818 221912 335874 221921
rect 335818 221847 335874 221856
rect 337672 221270 337700 227054
rect 338132 222222 338160 227802
rect 338028 222216 338080 222222
rect 338028 222158 338080 222164
rect 338120 222216 338172 222222
rect 338776 222193 338804 231676
rect 339144 228206 339172 231676
rect 339132 228200 339184 228206
rect 339132 228142 339184 228148
rect 339512 227662 339540 231676
rect 339592 227792 339644 227798
rect 339592 227734 339644 227740
rect 339500 227656 339552 227662
rect 339500 227598 339552 227604
rect 338856 225276 338908 225282
rect 338856 225218 338908 225224
rect 338120 222158 338172 222164
rect 338762 222184 338818 222193
rect 337200 221264 337252 221270
rect 337200 221206 337252 221212
rect 337660 221264 337712 221270
rect 337660 221206 337712 221212
rect 336740 221128 336792 221134
rect 336740 221070 336792 221076
rect 336752 217410 336780 221070
rect 317892 217382 318228 217410
rect 318720 217382 319056 217410
rect 319548 217382 319884 217410
rect 320376 217382 320712 217410
rect 321204 217382 321540 217410
rect 322032 217382 322368 217410
rect 322952 217382 323288 217410
rect 323872 217382 324116 217410
rect 324608 217382 324944 217410
rect 325712 217382 325772 217410
rect 326264 217382 326600 217410
rect 327092 217382 327428 217410
rect 327920 217382 328256 217410
rect 328840 217382 329176 217410
rect 329668 217382 330004 217410
rect 330496 217382 330832 217410
rect 331324 217382 331660 217410
rect 332152 217382 332488 217410
rect 332980 217382 333316 217410
rect 333992 217382 334144 217410
rect 334728 217382 335064 217410
rect 335556 217382 335892 217410
rect 336720 217382 336780 217410
rect 337212 217410 337240 221206
rect 338040 217410 338068 222158
rect 338762 222119 338818 222128
rect 338868 217410 338896 225218
rect 339604 221202 339632 227734
rect 339880 225418 339908 231676
rect 340248 226030 340276 231676
rect 340616 227866 340644 231676
rect 340696 229016 340748 229022
rect 340696 228958 340748 228964
rect 340604 227860 340656 227866
rect 340604 227802 340656 227808
rect 340236 226024 340288 226030
rect 340236 225966 340288 225972
rect 339868 225412 339920 225418
rect 339868 225354 339920 225360
rect 339684 221536 339736 221542
rect 339684 221478 339736 221484
rect 339592 221196 339644 221202
rect 339592 221138 339644 221144
rect 339696 217410 339724 221478
rect 340708 221406 340736 228958
rect 340892 228886 340920 231676
rect 340880 228880 340932 228886
rect 340880 228822 340932 228828
rect 341260 228070 341288 231676
rect 341248 228064 341300 228070
rect 341248 228006 341300 228012
rect 341628 227934 341656 231676
rect 341616 227928 341668 227934
rect 341616 227870 341668 227876
rect 341996 227798 342024 231676
rect 342364 229022 342392 231676
rect 342352 229016 342404 229022
rect 342352 228958 342404 228964
rect 342732 228954 342760 231676
rect 342720 228948 342772 228954
rect 342720 228890 342772 228896
rect 341984 227792 342036 227798
rect 341984 227734 342036 227740
rect 341524 227724 341576 227730
rect 341524 227666 341576 227672
rect 340604 221400 340656 221406
rect 340604 221342 340656 221348
rect 340696 221400 340748 221406
rect 340696 221342 340748 221348
rect 340616 217410 340644 221342
rect 341536 221338 341564 227666
rect 343100 225554 343128 231676
rect 343088 225548 343140 225554
rect 343088 225490 343140 225496
rect 342444 225208 342496 225214
rect 342444 225150 342496 225156
rect 341432 221332 341484 221338
rect 341432 221274 341484 221280
rect 341524 221332 341576 221338
rect 341524 221274 341576 221280
rect 341444 217410 341472 221274
rect 342456 217410 342484 225150
rect 343088 222216 343140 222222
rect 343088 222158 343140 222164
rect 343100 217410 343128 222158
rect 343468 219094 343496 231676
rect 343744 227594 343772 231676
rect 343732 227588 343784 227594
rect 343732 227530 343784 227536
rect 344008 227452 344060 227458
rect 344008 227394 344060 227400
rect 344020 221474 344048 227394
rect 344112 224262 344140 231676
rect 344480 227730 344508 231676
rect 344468 227724 344520 227730
rect 344468 227666 344520 227672
rect 344100 224256 344152 224262
rect 344100 224198 344152 224204
rect 343916 221468 343968 221474
rect 343916 221410 343968 221416
rect 344008 221468 344060 221474
rect 344008 221410 344060 221416
rect 343456 219088 343508 219094
rect 343456 219030 343508 219036
rect 343928 217410 343956 221410
rect 344848 219162 344876 231676
rect 345112 227316 345164 227322
rect 345112 227258 345164 227264
rect 345020 221672 345072 221678
rect 345020 221614 345072 221620
rect 344836 219156 344888 219162
rect 344836 219098 344888 219104
rect 345032 217410 345060 221614
rect 345124 221542 345152 227258
rect 345216 226778 345244 231676
rect 345204 226772 345256 226778
rect 345204 226714 345256 226720
rect 345584 226334 345612 231676
rect 345952 230110 345980 231676
rect 345940 230104 345992 230110
rect 345940 230046 345992 230052
rect 345940 228676 345992 228682
rect 345940 228618 345992 228624
rect 345584 226306 345704 226334
rect 345572 225072 345624 225078
rect 345572 225014 345624 225020
rect 345112 221536 345164 221542
rect 345112 221478 345164 221484
rect 345584 217410 345612 225014
rect 345676 224194 345704 226306
rect 345664 224188 345716 224194
rect 345664 224130 345716 224136
rect 345952 221678 345980 228618
rect 345940 221672 345992 221678
rect 345940 221614 345992 221620
rect 346320 219230 346348 231676
rect 346596 224466 346624 231676
rect 346584 224460 346636 224466
rect 346584 224402 346636 224408
rect 346964 224330 346992 231676
rect 347332 227458 347360 231676
rect 347320 227452 347372 227458
rect 347320 227394 347372 227400
rect 347412 226364 347464 226370
rect 347412 226306 347464 226312
rect 346952 224324 347004 224330
rect 346952 224266 347004 224272
rect 347424 221950 347452 226306
rect 347320 221944 347372 221950
rect 347320 221886 347372 221892
rect 347412 221944 347464 221950
rect 347412 221886 347464 221892
rect 346492 221264 346544 221270
rect 346492 221206 346544 221212
rect 346308 219224 346360 219230
rect 346308 219166 346360 219172
rect 346504 217410 346532 221206
rect 347332 217410 347360 221886
rect 347700 219366 347728 231676
rect 348068 224534 348096 231676
rect 348056 224528 348108 224534
rect 348056 224470 348108 224476
rect 348436 224398 348464 231676
rect 348804 230178 348832 231676
rect 348792 230172 348844 230178
rect 348792 230114 348844 230120
rect 348976 225140 349028 225146
rect 348976 225082 349028 225088
rect 348424 224392 348476 224398
rect 348424 224334 348476 224340
rect 348148 221604 348200 221610
rect 348148 221546 348200 221552
rect 347688 219360 347740 219366
rect 347688 219302 347740 219308
rect 348160 217410 348188 221546
rect 348988 217410 349016 225082
rect 349172 219298 349200 231676
rect 349448 224806 349476 231676
rect 349816 225214 349844 231676
rect 350184 230246 350212 231676
rect 350172 230240 350224 230246
rect 350172 230182 350224 230188
rect 349804 225208 349856 225214
rect 349804 225150 349856 225156
rect 349436 224800 349488 224806
rect 349436 224742 349488 224748
rect 349804 221196 349856 221202
rect 349804 221138 349856 221144
rect 349160 219292 349212 219298
rect 349160 219234 349212 219240
rect 349816 217410 349844 221138
rect 350552 220794 350580 231676
rect 350920 224874 350948 231676
rect 350908 224868 350960 224874
rect 350908 224810 350960 224816
rect 351288 224602 351316 231676
rect 351656 230042 351684 231676
rect 351644 230036 351696 230042
rect 351644 229978 351696 229984
rect 352024 226334 352052 231676
rect 352024 226306 352144 226334
rect 351276 224596 351328 224602
rect 351276 224538 351328 224544
rect 351920 222420 351972 222426
rect 351920 222362 351972 222368
rect 352012 222420 352064 222426
rect 352012 222362 352064 222368
rect 351932 222290 351960 222362
rect 351920 222284 351972 222290
rect 351920 222226 351972 222232
rect 351460 221808 351512 221814
rect 351460 221750 351512 221756
rect 350632 221740 350684 221746
rect 350632 221682 350684 221688
rect 350540 220788 350592 220794
rect 350540 220730 350592 220736
rect 350644 217410 350672 221682
rect 351472 217410 351500 221750
rect 352024 221134 352052 222362
rect 352012 221128 352064 221134
rect 352012 221070 352064 221076
rect 352116 220726 352144 226306
rect 352300 226166 352328 231676
rect 352288 226160 352340 226166
rect 352288 226102 352340 226108
rect 352380 225004 352432 225010
rect 352380 224946 352432 224952
rect 352104 220720 352156 220726
rect 352104 220662 352156 220668
rect 352392 217410 352420 224946
rect 352668 224738 352696 231676
rect 353036 229906 353064 231676
rect 353024 229900 353076 229906
rect 353024 229842 353076 229848
rect 352656 224732 352708 224738
rect 352656 224674 352708 224680
rect 353300 221332 353352 221338
rect 353300 221274 353352 221280
rect 353312 217410 353340 221274
rect 353404 220658 353432 231676
rect 353772 226234 353800 231676
rect 354140 226302 354168 231676
rect 354508 229974 354536 231676
rect 354890 231662 355088 231690
rect 354496 229968 354548 229974
rect 354496 229910 354548 229916
rect 354128 226296 354180 226302
rect 354128 226238 354180 226244
rect 353760 226228 353812 226234
rect 353760 226170 353812 226176
rect 354036 222080 354088 222086
rect 354036 222022 354088 222028
rect 353392 220652 353444 220658
rect 353392 220594 353444 220600
rect 354048 217410 354076 222022
rect 354864 221876 354916 221882
rect 354864 221818 354916 221824
rect 354876 217410 354904 221818
rect 355060 220590 355088 231662
rect 355152 225350 355180 231676
rect 355520 226098 355548 231676
rect 355888 226914 355916 231676
rect 356060 227520 356112 227526
rect 356060 227462 356112 227468
rect 355876 226908 355928 226914
rect 355876 226850 355928 226856
rect 355508 226092 355560 226098
rect 355508 226034 355560 226040
rect 355140 225344 355192 225350
rect 355140 225286 355192 225292
rect 355048 220584 355100 220590
rect 355048 220526 355100 220532
rect 356072 217410 356100 227462
rect 356256 220522 356284 231676
rect 356624 225962 356652 231676
rect 356612 225956 356664 225962
rect 356612 225898 356664 225904
rect 356992 225146 357020 231676
rect 357360 229838 357388 231676
rect 357348 229832 357400 229838
rect 357348 229774 357400 229780
rect 356980 225140 357032 225146
rect 356980 225082 357032 225088
rect 357348 222148 357400 222154
rect 357348 222090 357400 222096
rect 356520 221400 356572 221406
rect 356520 221342 356572 221348
rect 356244 220516 356296 220522
rect 356244 220458 356296 220464
rect 337212 217382 337548 217410
rect 338040 217382 338376 217410
rect 338868 217382 339204 217410
rect 339696 217382 340032 217410
rect 340616 217382 340952 217410
rect 341444 217382 341780 217410
rect 342456 217382 342608 217410
rect 343100 217382 343436 217410
rect 343928 217382 344264 217410
rect 345032 217382 345092 217410
rect 345584 217382 345920 217410
rect 346504 217382 346840 217410
rect 347332 217382 347668 217410
rect 348160 217382 348496 217410
rect 348988 217382 349324 217410
rect 349816 217382 350152 217410
rect 350644 217382 350980 217410
rect 351472 217382 351808 217410
rect 352392 217382 352728 217410
rect 353312 217382 353556 217410
rect 354048 217382 354384 217410
rect 354876 217382 355212 217410
rect 356040 217382 356100 217410
rect 356532 217410 356560 221342
rect 357360 217410 357388 222090
rect 357728 220386 357756 231676
rect 358004 225078 358032 231676
rect 358372 225282 358400 231676
rect 358740 226982 358768 231676
rect 359122 231662 359412 231690
rect 359096 228744 359148 228750
rect 359096 228686 359148 228692
rect 358728 226976 358780 226982
rect 358728 226918 358780 226924
rect 358360 225276 358412 225282
rect 358360 225218 358412 225224
rect 357992 225072 358044 225078
rect 357992 225014 358044 225020
rect 358268 222012 358320 222018
rect 358268 221954 358320 221960
rect 357716 220380 357768 220386
rect 357716 220322 357768 220328
rect 358280 217410 358308 221954
rect 359108 217410 359136 228686
rect 359384 220454 359412 231662
rect 359476 225010 359504 231676
rect 359844 229770 359872 231676
rect 359832 229764 359884 229770
rect 359832 229706 359884 229712
rect 360212 229702 360240 231676
rect 360200 229696 360252 229702
rect 360200 229638 360252 229644
rect 359464 225004 359516 225010
rect 359464 224946 359516 224952
rect 359924 221468 359976 221474
rect 359924 221410 359976 221416
rect 359372 220448 359424 220454
rect 359372 220390 359424 220396
rect 359936 217410 359964 221410
rect 360580 220250 360608 231676
rect 360856 225894 360884 231676
rect 361224 226710 361252 231676
rect 361592 227050 361620 231676
rect 361580 227044 361632 227050
rect 361580 226986 361632 226992
rect 361212 226704 361264 226710
rect 361212 226646 361264 226652
rect 360844 225888 360896 225894
rect 360844 225830 360896 225836
rect 361764 223576 361816 223582
rect 361764 223518 361816 223524
rect 360752 223508 360804 223514
rect 360752 223450 360804 223456
rect 360568 220244 360620 220250
rect 360568 220186 360620 220192
rect 360764 217410 360792 223450
rect 361776 217410 361804 223518
rect 361960 220318 361988 231676
rect 362328 225826 362356 231676
rect 362408 226840 362460 226846
rect 362408 226782 362460 226788
rect 362316 225820 362368 225826
rect 362316 225762 362368 225768
rect 361948 220312 362000 220318
rect 361948 220254 362000 220260
rect 362420 217410 362448 226782
rect 362696 225758 362724 231676
rect 363064 229022 363092 231676
rect 362960 229016 363012 229022
rect 362960 228958 363012 228964
rect 363052 229016 363104 229022
rect 363052 228958 363104 228964
rect 362972 228478 363000 228958
rect 362960 228472 363012 228478
rect 362960 228414 363012 228420
rect 362684 225752 362736 225758
rect 362684 225694 362736 225700
rect 363236 223372 363288 223378
rect 363236 223314 363288 223320
rect 363248 217410 363276 223314
rect 363432 220114 363460 231676
rect 363708 225690 363736 231676
rect 364076 229498 364104 231676
rect 364444 229634 364472 231676
rect 364432 229628 364484 229634
rect 364432 229570 364484 229576
rect 364064 229492 364116 229498
rect 364064 229434 364116 229440
rect 364340 227384 364392 227390
rect 364340 227326 364392 227332
rect 363696 225684 363748 225690
rect 363696 225626 363748 225632
rect 364352 223582 364380 227326
rect 364340 223576 364392 223582
rect 364340 223518 364392 223524
rect 364340 223440 364392 223446
rect 364340 223382 364392 223388
rect 363420 220108 363472 220114
rect 363420 220050 363472 220056
rect 364352 217410 364380 223382
rect 364812 220182 364840 231676
rect 365180 225622 365208 231676
rect 365548 229566 365576 231676
rect 365930 231662 366220 231690
rect 365536 229560 365588 229566
rect 365536 229502 365588 229508
rect 365904 229016 365956 229022
rect 365904 228958 365956 228964
rect 365916 226334 365944 228958
rect 366192 227118 366220 231662
rect 366180 227112 366232 227118
rect 366180 227054 366232 227060
rect 365916 226306 366036 226334
rect 365168 225616 365220 225622
rect 365168 225558 365220 225564
rect 365904 223576 365956 223582
rect 365904 223518 365956 223524
rect 364984 223304 365036 223310
rect 364984 223246 365036 223252
rect 364800 220176 364852 220182
rect 364800 220118 364852 220124
rect 364996 217410 365024 223246
rect 365916 223038 365944 223518
rect 365812 223032 365864 223038
rect 365812 222974 365864 222980
rect 365904 223032 365956 223038
rect 365904 222974 365956 222980
rect 365824 217410 365852 222974
rect 366008 221338 366036 226306
rect 365996 221332 366048 221338
rect 365996 221274 366048 221280
rect 366284 219910 366312 231676
rect 366560 225486 366588 231676
rect 366928 226846 366956 231676
rect 366916 226840 366968 226846
rect 366916 226782 366968 226788
rect 366548 225480 366600 225486
rect 366548 225422 366600 225428
rect 366640 221536 366692 221542
rect 366640 221478 366692 221484
rect 366272 219904 366324 219910
rect 366272 219846 366324 219852
rect 366652 217410 366680 221478
rect 367296 221406 367324 231676
rect 367468 222828 367520 222834
rect 367468 222770 367520 222776
rect 367284 221400 367336 221406
rect 367284 221342 367336 221348
rect 367480 217410 367508 222770
rect 367664 219978 367692 231676
rect 368032 226370 368060 231676
rect 368020 226364 368072 226370
rect 368020 226306 368072 226312
rect 368204 225548 368256 225554
rect 368204 225490 368256 225496
rect 368216 221202 368244 225490
rect 368296 223236 368348 223242
rect 368296 223178 368348 223184
rect 368204 221196 368256 221202
rect 368204 221138 368256 221144
rect 367652 219972 367704 219978
rect 367652 219914 367704 219920
rect 368308 217410 368336 223178
rect 368400 220046 368428 231676
rect 368768 227322 368796 231676
rect 369150 231662 369348 231690
rect 368756 227316 368808 227322
rect 368756 227258 368808 227264
rect 369124 223100 369176 223106
rect 369124 223042 369176 223048
rect 368388 220040 368440 220046
rect 368388 219982 368440 219988
rect 369136 217410 369164 223042
rect 369320 219774 369348 231662
rect 369412 224641 369440 231676
rect 369780 226334 369808 231676
rect 370148 229430 370176 231676
rect 370136 229424 370188 229430
rect 370136 229366 370188 229372
rect 369688 226306 369808 226334
rect 369952 226364 370004 226370
rect 369952 226306 370004 226312
rect 369688 225418 369716 226306
rect 369964 226250 369992 226306
rect 369780 226222 369992 226250
rect 369780 225554 369808 226222
rect 370228 226024 370280 226030
rect 370228 225966 370280 225972
rect 369768 225548 369820 225554
rect 369768 225490 369820 225496
rect 369584 225412 369636 225418
rect 369584 225354 369636 225360
rect 369676 225412 369728 225418
rect 369676 225354 369728 225360
rect 369398 224632 369454 224641
rect 369398 224567 369454 224576
rect 369596 222834 369624 225354
rect 370240 222902 370268 225966
rect 370044 222896 370096 222902
rect 370044 222838 370096 222844
rect 370228 222896 370280 222902
rect 370228 222838 370280 222844
rect 369584 222828 369636 222834
rect 369584 222770 369636 222776
rect 369308 219768 369360 219774
rect 369308 219710 369360 219716
rect 370056 217410 370084 222838
rect 370516 219842 370544 231676
rect 370884 224505 370912 231676
rect 371252 229362 371280 231676
rect 371240 229356 371292 229362
rect 371240 229298 371292 229304
rect 371620 227254 371648 231676
rect 371608 227248 371660 227254
rect 371608 227190 371660 227196
rect 371988 226642 372016 231676
rect 371976 226636 372028 226642
rect 371976 226578 372028 226584
rect 372264 224777 372292 231676
rect 372250 224768 372306 224777
rect 372250 224703 372306 224712
rect 370870 224496 370926 224505
rect 370870 224431 370926 224440
rect 372632 224369 372660 231676
rect 372618 224360 372674 224369
rect 372618 224295 372674 224304
rect 371700 223168 371752 223174
rect 371700 223110 371752 223116
rect 370872 222964 370924 222970
rect 370872 222906 370924 222912
rect 370504 219836 370556 219842
rect 370504 219778 370556 219784
rect 370884 217410 370912 222906
rect 371712 217410 371740 223110
rect 372620 222488 372672 222494
rect 372620 222430 372672 222436
rect 372632 217410 372660 222430
rect 373000 221474 373028 231676
rect 373368 226438 373396 231676
rect 373356 226432 373408 226438
rect 373356 226374 373408 226380
rect 373736 226273 373764 231676
rect 373908 229084 373960 229090
rect 373908 229026 373960 229032
rect 373722 226264 373778 226273
rect 373722 226199 373778 226208
rect 373920 222494 373948 229026
rect 374104 226574 374132 231676
rect 374472 227390 374500 231676
rect 374840 229294 374868 231676
rect 374828 229288 374880 229294
rect 374828 229230 374880 229236
rect 374460 227384 374512 227390
rect 374460 227326 374512 227332
rect 374092 226568 374144 226574
rect 374092 226510 374144 226516
rect 374184 222760 374236 222766
rect 374184 222702 374236 222708
rect 373908 222488 373960 222494
rect 373908 222430 373960 222436
rect 373356 221672 373408 221678
rect 373356 221614 373408 221620
rect 372988 221468 373040 221474
rect 372988 221410 373040 221416
rect 373368 217410 373396 221614
rect 374196 217410 374224 222702
rect 375116 221542 375144 231676
rect 375484 228682 375512 231676
rect 375472 228676 375524 228682
rect 375472 228618 375524 228624
rect 375380 222624 375432 222630
rect 375380 222566 375432 222572
rect 375104 221536 375156 221542
rect 375104 221478 375156 221484
rect 375392 217410 375420 222566
rect 375852 222057 375880 231676
rect 375932 228540 375984 228546
rect 375932 228482 375984 228488
rect 375838 222048 375894 222057
rect 375838 221983 375894 221992
rect 356532 217382 356868 217410
rect 357360 217382 357696 217410
rect 358280 217382 358616 217410
rect 359108 217382 359444 217410
rect 359936 217382 360272 217410
rect 360764 217382 361100 217410
rect 361776 217382 361928 217410
rect 362420 217382 362756 217410
rect 363248 217382 363584 217410
rect 364352 217382 364504 217410
rect 364996 217382 365332 217410
rect 365824 217382 366160 217410
rect 366652 217382 366988 217410
rect 367480 217382 367816 217410
rect 368308 217382 368644 217410
rect 369136 217382 369472 217410
rect 370056 217382 370392 217410
rect 370884 217382 371220 217410
rect 371712 217382 372048 217410
rect 372632 217382 372876 217410
rect 373368 217382 373704 217410
rect 374196 217382 374532 217410
rect 375360 217382 375420 217410
rect 375944 217410 375972 228482
rect 376220 227186 376248 231676
rect 376588 228750 376616 231676
rect 376576 228744 376628 228750
rect 376576 228686 376628 228692
rect 376668 228608 376720 228614
rect 376668 228550 376720 228556
rect 376208 227180 376260 227186
rect 376208 227122 376260 227128
rect 376576 226772 376628 226778
rect 376576 226714 376628 226720
rect 376588 223990 376616 226714
rect 376576 223984 376628 223990
rect 376576 223926 376628 223932
rect 376680 222630 376708 228550
rect 376852 227656 376904 227662
rect 376852 227598 376904 227604
rect 376668 222624 376720 222630
rect 376668 222566 376720 222572
rect 376864 222426 376892 227598
rect 376956 227361 376984 231676
rect 376942 227352 376998 227361
rect 376942 227287 376998 227296
rect 377324 227225 377352 231676
rect 377310 227216 377366 227225
rect 377310 227151 377366 227160
rect 377588 222692 377640 222698
rect 377588 222634 377640 222640
rect 376760 222420 376812 222426
rect 376760 222362 376812 222368
rect 376852 222420 376904 222426
rect 376852 222362 376904 222368
rect 376772 217410 376800 222362
rect 377600 217410 377628 222634
rect 377692 221678 377720 231676
rect 377968 221814 377996 231676
rect 378232 228472 378284 228478
rect 378232 228414 378284 228420
rect 378140 227588 378192 227594
rect 378140 227530 378192 227536
rect 378152 223922 378180 227530
rect 378244 224058 378272 228414
rect 378232 224052 378284 224058
rect 378232 223994 378284 224000
rect 378140 223916 378192 223922
rect 378140 223858 378192 223864
rect 378336 223553 378364 231676
rect 378322 223544 378378 223553
rect 378322 223479 378378 223488
rect 378704 223417 378732 231676
rect 378690 223408 378746 223417
rect 378690 223343 378746 223352
rect 378416 222556 378468 222562
rect 378416 222498 378468 222504
rect 377956 221808 378008 221814
rect 377956 221750 378008 221756
rect 377680 221672 377732 221678
rect 377680 221614 377732 221620
rect 378428 217410 378456 222498
rect 379072 221610 379100 231676
rect 379440 228614 379468 231676
rect 379428 228608 379480 228614
rect 379428 228550 379480 228556
rect 379808 226778 379836 231676
rect 380176 227497 380204 231676
rect 380162 227488 380218 227497
rect 380162 227423 380218 227432
rect 379796 226772 379848 226778
rect 379796 226714 379848 226720
rect 379244 226500 379296 226506
rect 379244 226442 379296 226448
rect 379060 221604 379112 221610
rect 379060 221546 379112 221552
rect 379256 217410 379284 226442
rect 380072 221944 380124 221950
rect 380072 221886 380124 221892
rect 380084 217410 380112 221886
rect 380544 221882 380572 231676
rect 380532 221876 380584 221882
rect 380532 221818 380584 221824
rect 380820 221746 380848 231676
rect 380992 228948 381044 228954
rect 380992 228890 381044 228896
rect 380900 228880 380952 228886
rect 380900 228822 380952 228828
rect 380912 224670 380940 228822
rect 380900 224664 380952 224670
rect 380900 224606 380952 224612
rect 381004 223854 381032 228890
rect 380992 223848 381044 223854
rect 380992 223790 381044 223796
rect 381188 223281 381216 231676
rect 381174 223272 381230 223281
rect 381174 223207 381230 223216
rect 381556 223145 381584 231676
rect 381542 223136 381598 223145
rect 381542 223071 381598 223080
rect 381082 223000 381138 223009
rect 381082 222935 381138 222944
rect 380808 221740 380860 221746
rect 380808 221682 380860 221688
rect 381096 217410 381124 222935
rect 381820 222284 381872 222290
rect 381820 222226 381872 222232
rect 381832 217410 381860 222226
rect 381924 222018 381952 231676
rect 381912 222012 381964 222018
rect 381912 221954 381964 221960
rect 382292 221950 382320 231676
rect 382660 227089 382688 231676
rect 383028 227526 383056 231676
rect 383016 227520 383068 227526
rect 383016 227462 383068 227468
rect 382646 227080 382702 227089
rect 382646 227015 382702 227024
rect 382648 223032 382700 223038
rect 382648 222974 382700 222980
rect 382280 221944 382332 221950
rect 382280 221886 382332 221892
rect 382660 217410 382688 222974
rect 383396 222086 383424 231676
rect 383686 231662 383976 231690
rect 383752 228812 383804 228818
rect 383752 228754 383804 228760
rect 383660 226704 383712 226710
rect 383660 226646 383712 226652
rect 383672 224126 383700 226646
rect 383660 224120 383712 224126
rect 383660 224062 383712 224068
rect 383658 222864 383714 222873
rect 383658 222799 383714 222808
rect 383384 222080 383436 222086
rect 383384 222022 383436 222028
rect 383672 217410 383700 222799
rect 383764 221134 383792 228754
rect 383948 223009 383976 231662
rect 383934 223000 383990 223009
rect 383934 222935 383990 222944
rect 384040 222154 384068 231676
rect 384408 228546 384436 231676
rect 384776 228993 384804 231676
rect 384762 228984 384818 228993
rect 384762 228919 384818 228928
rect 384396 228540 384448 228546
rect 384396 228482 384448 228488
rect 385144 227594 385172 231676
rect 385132 227588 385184 227594
rect 385132 227530 385184 227536
rect 384302 222592 384358 222601
rect 384302 222527 384358 222536
rect 384028 222148 384080 222154
rect 384028 222090 384080 222096
rect 383752 221128 383804 221134
rect 383752 221070 383804 221076
rect 384316 217410 384344 222527
rect 385132 222352 385184 222358
rect 385132 222294 385184 222300
rect 385144 217410 385172 222294
rect 385512 220998 385540 231676
rect 385880 222873 385908 231676
rect 385960 228404 386012 228410
rect 385960 228346 386012 228352
rect 385866 222864 385922 222873
rect 385866 222799 385922 222808
rect 385500 220992 385552 220998
rect 385500 220934 385552 220940
rect 385972 217410 386000 228346
rect 386248 221066 386276 231676
rect 386524 228478 386552 231676
rect 386892 228857 386920 231676
rect 386878 228848 386934 228857
rect 386878 228783 386934 228792
rect 386512 228472 386564 228478
rect 386512 228414 386564 228420
rect 387260 227662 387288 231676
rect 387248 227656 387300 227662
rect 387248 227598 387300 227604
rect 387628 223514 387656 231676
rect 387616 223508 387668 223514
rect 387616 223450 387668 223456
rect 387996 222737 388024 231676
rect 388364 229226 388392 231676
rect 388352 229220 388404 229226
rect 388352 229162 388404 229168
rect 388732 223378 388760 231676
rect 389008 231662 389114 231690
rect 388720 223372 388772 223378
rect 388720 223314 388772 223320
rect 386786 222728 386842 222737
rect 386786 222663 386842 222672
rect 387982 222728 388038 222737
rect 387982 222663 388038 222672
rect 386236 221060 386288 221066
rect 386236 221002 386288 221008
rect 386800 217410 386828 222663
rect 389008 222601 389036 231662
rect 389088 228336 389140 228342
rect 389088 228278 389140 228284
rect 388994 222592 389050 222601
rect 388994 222527 389050 222536
rect 387706 222456 387762 222465
rect 387706 222391 387762 222400
rect 387720 217410 387748 222391
rect 388534 221912 388590 221921
rect 388534 221847 388590 221856
rect 388548 217410 388576 221847
rect 389100 221082 389128 228278
rect 389376 226370 389404 231676
rect 389744 229090 389772 231676
rect 389732 229084 389784 229090
rect 389732 229026 389784 229032
rect 390112 228721 390140 231676
rect 390098 228712 390154 228721
rect 390098 228647 390154 228656
rect 389916 228132 389968 228138
rect 389916 228074 389968 228080
rect 389364 226364 389416 226370
rect 389364 226306 389416 226312
rect 389928 221270 389956 228074
rect 390480 226001 390508 231676
rect 390466 225992 390522 226001
rect 390466 225927 390522 225936
rect 390848 223310 390876 231676
rect 391020 224936 391072 224942
rect 391020 224878 391072 224884
rect 390836 223304 390888 223310
rect 390836 223246 390888 223252
rect 390190 222320 390246 222329
rect 390190 222255 390246 222264
rect 389916 221264 389968 221270
rect 389916 221206 389968 221212
rect 389100 221054 389312 221082
rect 389284 217410 389312 221054
rect 390204 217410 390232 222255
rect 391032 217410 391060 224878
rect 391216 222465 391244 231676
rect 391584 225729 391612 231676
rect 391952 229022 391980 231676
rect 391940 229016 391992 229022
rect 391940 228958 391992 228964
rect 392228 228585 392256 231676
rect 392214 228576 392270 228585
rect 392214 228511 392270 228520
rect 391940 228268 391992 228274
rect 391940 228210 391992 228216
rect 391756 226772 391808 226778
rect 391756 226714 391808 226720
rect 391570 225720 391626 225729
rect 391570 225655 391626 225664
rect 391202 222456 391258 222465
rect 391202 222391 391258 222400
rect 391768 221921 391796 226714
rect 391754 221912 391810 221921
rect 391754 221847 391810 221856
rect 391952 217410 391980 228210
rect 392596 225865 392624 231676
rect 392582 225856 392638 225865
rect 392582 225791 392638 225800
rect 392964 223242 392992 231676
rect 392952 223236 393004 223242
rect 392952 223178 393004 223184
rect 393332 222329 393360 231676
rect 393700 225593 393728 231676
rect 394068 228818 394096 231676
rect 394056 228812 394108 228818
rect 394056 228754 394108 228760
rect 394436 228449 394464 231676
rect 394422 228440 394478 228449
rect 394422 228375 394478 228384
rect 393780 228200 393832 228206
rect 393780 228142 393832 228148
rect 393686 225584 393742 225593
rect 393686 225519 393742 225528
rect 393318 222320 393374 222329
rect 393318 222255 393374 222264
rect 393596 222216 393648 222222
rect 393596 222158 393648 222164
rect 392676 221264 392728 221270
rect 392676 221206 392728 221212
rect 392688 217410 392716 221206
rect 393608 217410 393636 222158
rect 393792 220930 393820 228142
rect 394804 225457 394832 231676
rect 394790 225448 394846 225457
rect 394790 225383 394846 225392
rect 395080 223174 395108 231676
rect 395252 227996 395304 228002
rect 395252 227938 395304 227944
rect 395068 223168 395120 223174
rect 395068 223110 395120 223116
rect 394700 222624 394752 222630
rect 394700 222566 394752 222572
rect 393780 220924 393832 220930
rect 393780 220866 393832 220872
rect 394712 217410 394740 222566
rect 395264 217410 395292 227938
rect 395448 223106 395476 231676
rect 395816 226506 395844 231676
rect 396184 228886 396212 231676
rect 396172 228880 396224 228886
rect 396172 228822 396224 228828
rect 396552 228313 396580 231676
rect 396920 229158 396948 231676
rect 396908 229152 396960 229158
rect 396908 229094 396960 229100
rect 396538 228304 396594 228313
rect 396538 228239 396594 228248
rect 396172 228064 396224 228070
rect 396172 228006 396224 228012
rect 395804 226500 395856 226506
rect 395804 226442 395856 226448
rect 395436 223100 395488 223106
rect 395436 223042 395488 223048
rect 396184 222290 396212 228006
rect 397288 223038 397316 231676
rect 397552 226636 397604 226642
rect 397552 226578 397604 226584
rect 397460 226432 397512 226438
rect 397460 226374 397512 226380
rect 397472 226030 397500 226374
rect 397460 226024 397512 226030
rect 397460 225966 397512 225972
rect 397276 223032 397328 223038
rect 397276 222974 397328 222980
rect 396172 222284 396224 222290
rect 396172 222226 396224 222232
rect 396906 222184 396962 222193
rect 396906 222119 396962 222128
rect 396080 221128 396132 221134
rect 396080 221070 396132 221076
rect 396092 217410 396120 221070
rect 396920 217410 396948 222119
rect 397564 221270 397592 226578
rect 397656 222193 397684 231676
rect 397932 225321 397960 231676
rect 398300 228954 398328 231676
rect 398288 228948 398340 228954
rect 398288 228890 398340 228896
rect 398668 228177 398696 231676
rect 398654 228168 398710 228177
rect 398654 228103 398710 228112
rect 399036 226710 399064 231676
rect 399024 226704 399076 226710
rect 399024 226646 399076 226652
rect 397918 225312 397974 225321
rect 397918 225247 397974 225256
rect 399404 222970 399432 231676
rect 399772 228041 399800 231676
rect 399758 228032 399814 228041
rect 399758 227967 399814 227976
rect 400036 227928 400088 227934
rect 400036 227870 400088 227876
rect 399392 222964 399444 222970
rect 399392 222906 399444 222912
rect 398564 222828 398616 222834
rect 398564 222770 398616 222776
rect 397736 222488 397788 222494
rect 397736 222430 397788 222436
rect 397642 222184 397698 222193
rect 397642 222119 397698 222128
rect 397552 221264 397604 221270
rect 397552 221206 397604 221212
rect 397748 217410 397776 222430
rect 398576 217410 398604 222770
rect 400048 222222 400076 227870
rect 400140 222834 400168 231676
rect 400508 228410 400536 231676
rect 400496 228404 400548 228410
rect 400496 228346 400548 228352
rect 400784 222902 400812 231676
rect 401152 225185 401180 231676
rect 401138 225176 401194 225185
rect 401138 225111 401194 225120
rect 400404 222896 400456 222902
rect 400404 222838 400456 222844
rect 400772 222896 400824 222902
rect 400772 222838 400824 222844
rect 400128 222828 400180 222834
rect 400128 222770 400180 222776
rect 400036 222216 400088 222222
rect 400036 222158 400088 222164
rect 399484 220924 399536 220930
rect 399484 220866 399536 220872
rect 399496 217410 399524 220866
rect 400416 217410 400444 222838
rect 401520 222766 401548 231676
rect 401888 228342 401916 231676
rect 401876 228336 401928 228342
rect 401876 228278 401928 228284
rect 402256 226778 402284 231676
rect 402624 228274 402652 231676
rect 403006 231662 403296 231690
rect 402612 228268 402664 228274
rect 402612 228210 402664 228216
rect 402796 227860 402848 227866
rect 402796 227802 402848 227808
rect 402244 226772 402296 226778
rect 402244 226714 402296 226720
rect 402808 226334 402836 227802
rect 402980 226568 403032 226574
rect 402980 226510 403032 226516
rect 402808 226306 402928 226334
rect 402796 224664 402848 224670
rect 402796 224606 402848 224612
rect 402808 224466 402836 224606
rect 402796 224460 402848 224466
rect 402796 224402 402848 224408
rect 402612 224392 402664 224398
rect 402612 224334 402664 224340
rect 402624 223786 402652 224334
rect 402612 223780 402664 223786
rect 402612 223722 402664 223728
rect 401508 222760 401560 222766
rect 401508 222702 401560 222708
rect 401140 222420 401192 222426
rect 401140 222362 401192 222368
rect 401152 217410 401180 222362
rect 401968 222284 402020 222290
rect 401968 222226 402020 222232
rect 401980 217410 402008 222226
rect 402900 220946 402928 226306
rect 402992 224670 403020 226510
rect 402980 224664 403032 224670
rect 402980 224606 403032 224612
rect 403268 222630 403296 231662
rect 403360 222698 403388 231676
rect 403636 228206 403664 231676
rect 403624 228200 403676 228206
rect 403624 228142 403676 228148
rect 404004 227905 404032 231676
rect 403990 227896 404046 227905
rect 403990 227831 404046 227840
rect 403716 227792 403768 227798
rect 403716 227734 403768 227740
rect 403348 222692 403400 222698
rect 403348 222634 403400 222640
rect 403256 222624 403308 222630
rect 403256 222566 403308 222572
rect 403624 222216 403676 222222
rect 403624 222158 403676 222164
rect 402900 220918 403020 220946
rect 402992 217410 403020 220918
rect 403636 217410 403664 222158
rect 403728 221202 403756 227734
rect 404372 226642 404400 231676
rect 404360 226636 404412 226642
rect 404360 226578 404412 226584
rect 404452 224460 404504 224466
rect 404452 224402 404504 224408
rect 403716 221196 403768 221202
rect 403716 221138 403768 221144
rect 404464 217410 404492 224402
rect 404740 222562 404768 231676
rect 404728 222556 404780 222562
rect 404728 222498 404780 222504
rect 405108 222426 405136 231676
rect 405096 222420 405148 222426
rect 405096 222362 405148 222368
rect 405476 222358 405504 231676
rect 405740 223848 405792 223854
rect 405740 223790 405792 223796
rect 405464 222352 405516 222358
rect 405464 222294 405516 222300
rect 405752 217410 405780 223790
rect 405844 222494 405872 231676
rect 406212 228070 406240 231676
rect 406200 228064 406252 228070
rect 406200 228006 406252 228012
rect 406488 224942 406516 231676
rect 406856 228138 406884 231676
rect 406844 228132 406896 228138
rect 406844 228074 406896 228080
rect 407224 227934 407252 231676
rect 407212 227928 407264 227934
rect 407212 227870 407264 227876
rect 407592 225049 407620 231676
rect 407578 225040 407634 225049
rect 407578 224975 407634 224984
rect 406476 224936 406528 224942
rect 406476 224878 406528 224884
rect 407856 224052 407908 224058
rect 407856 223994 407908 224000
rect 405832 222488 405884 222494
rect 405832 222430 405884 222436
rect 406200 221196 406252 221202
rect 406200 221138 406252 221144
rect 375944 217382 376280 217410
rect 376772 217382 377108 217410
rect 377600 217382 377936 217410
rect 378428 217382 378764 217410
rect 379256 217382 379592 217410
rect 380084 217382 380420 217410
rect 381096 217382 381248 217410
rect 381832 217382 382168 217410
rect 382660 217382 382996 217410
rect 383672 217382 383824 217410
rect 384316 217382 384652 217410
rect 385144 217382 385480 217410
rect 385972 217382 386308 217410
rect 386800 217382 387136 217410
rect 387720 217382 388056 217410
rect 388548 217382 388884 217410
rect 389284 217382 389712 217410
rect 390204 217382 390540 217410
rect 391032 217382 391368 217410
rect 391952 217382 392196 217410
rect 392688 217382 393024 217410
rect 393608 217382 393944 217410
rect 394712 217382 394772 217410
rect 395264 217382 395600 217410
rect 396092 217382 396428 217410
rect 396920 217382 397256 217410
rect 397748 217382 398084 217410
rect 398576 217382 398912 217410
rect 399496 217382 399832 217410
rect 400416 217382 400660 217410
rect 401152 217382 401488 217410
rect 401980 217382 402316 217410
rect 402992 217382 403144 217410
rect 403636 217382 403972 217410
rect 404464 217382 404800 217410
rect 405720 217382 405780 217410
rect 406212 217410 406240 221138
rect 407028 221128 407080 221134
rect 407028 221070 407080 221076
rect 407040 217410 407068 221070
rect 407868 217410 407896 223994
rect 407960 221134 407988 231676
rect 408328 227866 408356 231676
rect 408316 227860 408368 227866
rect 408316 227802 408368 227808
rect 408696 226914 408724 231676
rect 409064 228002 409092 231676
rect 409052 227996 409104 228002
rect 409052 227938 409104 227944
rect 408316 226908 408368 226914
rect 408316 226850 408368 226856
rect 408684 226908 408736 226914
rect 408684 226850 408736 226856
rect 408328 221202 408356 226850
rect 408408 226840 408460 226846
rect 408408 226782 408460 226788
rect 408420 224058 408448 226782
rect 408684 224256 408736 224262
rect 408684 224198 408736 224204
rect 408408 224052 408460 224058
rect 408408 223994 408460 224000
rect 408316 221196 408368 221202
rect 408316 221138 408368 221144
rect 407948 221128 408000 221134
rect 407948 221070 408000 221076
rect 408696 217410 408724 224198
rect 409340 222290 409368 231676
rect 409708 226846 409736 231676
rect 410076 227769 410104 231676
rect 410444 227798 410472 231676
rect 410432 227792 410484 227798
rect 410062 227760 410118 227769
rect 410432 227734 410484 227740
rect 410062 227695 410118 227704
rect 410340 227724 410392 227730
rect 410340 227666 410392 227672
rect 409696 226840 409748 226846
rect 409696 226782 409748 226788
rect 409328 222284 409380 222290
rect 409328 222226 409380 222232
rect 409512 219088 409564 219094
rect 409512 219030 409564 219036
rect 409524 217410 409552 219030
rect 410352 217410 410380 227666
rect 410812 224913 410840 231676
rect 411180 227633 411208 231676
rect 411548 227730 411576 231676
rect 411536 227724 411588 227730
rect 411536 227666 411588 227672
rect 411166 227624 411222 227633
rect 411166 227559 411222 227568
rect 411076 227452 411128 227458
rect 411076 227394 411128 227400
rect 410798 224904 410854 224913
rect 410798 224839 410854 224848
rect 411088 223650 411116 227394
rect 411914 226414 411942 231698
rect 414020 230104 414072 230110
rect 414020 230046 414072 230052
rect 411996 226976 412048 226982
rect 411996 226918 412048 226924
rect 411902 226408 411954 226414
rect 411168 226364 411220 226370
rect 411902 226350 411954 226356
rect 411168 226306 411220 226312
rect 411180 226137 411208 226306
rect 411166 226128 411222 226137
rect 411166 226063 411222 226072
rect 412008 224262 412036 226918
rect 411996 224256 412048 224262
rect 411996 224198 412048 224204
rect 412088 224188 412140 224194
rect 412088 224130 412140 224136
rect 411260 223916 411312 223922
rect 411260 223858 411312 223864
rect 411076 223644 411128 223650
rect 411076 223586 411128 223592
rect 411272 217410 411300 223858
rect 412100 217410 412128 224130
rect 412916 219156 412968 219162
rect 412916 219098 412968 219104
rect 412928 217410 412956 219098
rect 414032 217410 414060 230046
rect 418080 226334 418108 243063
rect 418158 240000 418214 240009
rect 418158 239935 418214 239944
rect 417896 226306 418108 226334
rect 415400 224324 415452 224330
rect 415400 224266 415452 224272
rect 414572 223984 414624 223990
rect 414572 223926 414624 223932
rect 414584 217410 414612 223926
rect 415412 217410 415440 224266
rect 417148 223644 417200 223650
rect 417148 223586 417200 223592
rect 416228 219224 416280 219230
rect 416228 219166 416280 219172
rect 416240 217410 416268 219166
rect 417160 217410 417188 223586
rect 406212 217382 406548 217410
rect 407040 217382 407376 217410
rect 407868 217382 408204 217410
rect 408696 217382 409032 217410
rect 409524 217382 409860 217410
rect 410352 217382 410688 217410
rect 411272 217382 411608 217410
rect 412100 217382 412436 217410
rect 412928 217382 413264 217410
rect 414032 217382 414092 217410
rect 414584 217382 414920 217410
rect 415412 217382 415748 217410
rect 416240 217382 416576 217410
rect 417160 217382 417496 217410
rect 417896 216850 417924 226306
rect 417976 224392 418028 224398
rect 417976 224334 418028 224340
rect 417988 217410 418016 224334
rect 418172 218006 418200 239935
rect 418434 236736 418490 236745
rect 418434 236671 418490 236680
rect 418160 218000 418212 218006
rect 418160 217942 418212 217948
rect 417988 217382 418324 217410
rect 418448 216918 418476 236671
rect 418526 233608 418582 233617
rect 418526 233543 418582 233552
rect 418540 217054 418568 233543
rect 423864 230240 423916 230246
rect 423864 230182 423916 230188
rect 420460 230172 420512 230178
rect 420460 230114 420512 230120
rect 419540 227112 419592 227118
rect 419540 227054 419592 227060
rect 418896 227044 418948 227050
rect 418896 226986 418948 226992
rect 418908 224330 418936 226986
rect 419552 224534 419580 227054
rect 419540 224528 419592 224534
rect 419540 224470 419592 224476
rect 418896 224324 418948 224330
rect 418896 224266 418948 224272
rect 418804 223780 418856 223786
rect 418804 223722 418856 223728
rect 418620 218000 418672 218006
rect 418620 217942 418672 217948
rect 418528 217048 418580 217054
rect 418528 216990 418580 216996
rect 418632 216986 418660 217942
rect 418816 217410 418844 223722
rect 419724 219360 419776 219366
rect 419724 219302 419776 219308
rect 419736 217410 419764 219302
rect 420472 217410 420500 230114
rect 422300 226500 422352 226506
rect 422300 226442 422352 226448
rect 422312 225214 422340 226442
rect 422208 225208 422260 225214
rect 422208 225150 422260 225156
rect 422300 225208 422352 225214
rect 422300 225150 422352 225156
rect 422220 225026 422248 225150
rect 422220 224998 422340 225026
rect 421288 224392 421340 224398
rect 421288 224334 421340 224340
rect 421300 217410 421328 224334
rect 422312 217410 422340 224998
rect 423036 219292 423088 219298
rect 423036 219234 423088 219240
rect 423048 217410 423076 219234
rect 423876 217410 423904 230182
rect 427176 230036 427228 230042
rect 427176 229978 427228 229984
rect 425704 227316 425756 227322
rect 425704 227258 425756 227264
rect 425716 224806 425744 227258
rect 425060 224800 425112 224806
rect 425060 224742 425112 224748
rect 425704 224800 425756 224806
rect 425704 224742 425756 224748
rect 425072 217410 425100 224742
rect 425520 224596 425572 224602
rect 425520 224538 425572 224544
rect 418816 217382 419152 217410
rect 419736 217382 419980 217410
rect 420472 217382 420808 217410
rect 421300 217382 421636 217410
rect 422312 217382 422464 217410
rect 423048 217382 423384 217410
rect 423876 217382 424212 217410
rect 425040 217382 425100 217410
rect 425532 217410 425560 224538
rect 426348 220788 426400 220794
rect 426348 220730 426400 220736
rect 426360 217410 426388 220730
rect 427188 217410 427216 229978
rect 433892 229968 433944 229974
rect 433892 229910 433944 229916
rect 430580 229900 430632 229906
rect 430580 229842 430632 229848
rect 430488 227248 430540 227254
rect 430488 227190 430540 227196
rect 429108 225276 429160 225282
rect 429108 225218 429160 225224
rect 428004 224868 428056 224874
rect 428004 224810 428056 224816
rect 428016 217410 428044 224810
rect 429120 224738 429148 225218
rect 430500 224874 430528 227190
rect 430488 224868 430540 224874
rect 430488 224810 430540 224816
rect 428924 224732 428976 224738
rect 428924 224674 428976 224680
rect 429108 224732 429160 224738
rect 429108 224674 429160 224680
rect 428936 217410 428964 224674
rect 429752 220720 429804 220726
rect 429752 220662 429804 220668
rect 429764 217410 429792 220662
rect 430592 217410 430620 229842
rect 433248 227384 433300 227390
rect 433248 227326 433300 227332
rect 432236 226296 432288 226302
rect 432236 226238 432288 226244
rect 431408 226160 431460 226166
rect 431408 226102 431460 226108
rect 431420 217410 431448 226102
rect 432248 217410 432276 226238
rect 433260 226166 433288 227326
rect 433248 226160 433300 226166
rect 433248 226102 433300 226108
rect 433340 220652 433392 220658
rect 433340 220594 433392 220600
rect 433352 217410 433380 220594
rect 433904 217410 433932 229910
rect 440700 229832 440752 229838
rect 440700 229774 440752 229780
rect 434628 227180 434680 227186
rect 434628 227122 434680 227128
rect 434640 226098 434668 227122
rect 436100 226704 436152 226710
rect 436100 226646 436152 226652
rect 434812 226296 434864 226302
rect 434812 226238 434864 226244
rect 434628 226092 434680 226098
rect 434628 226034 434680 226040
rect 434824 217410 434852 226238
rect 435640 226228 435692 226234
rect 435640 226170 435692 226176
rect 435652 217410 435680 226170
rect 436112 225350 436140 226646
rect 438860 226636 438912 226642
rect 438860 226578 438912 226584
rect 436100 225344 436152 225350
rect 436100 225286 436152 225292
rect 438124 225276 438176 225282
rect 438124 225218 438176 225224
rect 437296 221196 437348 221202
rect 437296 221138 437348 221144
rect 436468 220584 436520 220590
rect 436468 220526 436520 220532
rect 436480 217410 436508 220526
rect 437308 217410 437336 221138
rect 438136 217410 438164 225218
rect 438872 225146 438900 226578
rect 438768 225140 438820 225146
rect 438768 225082 438820 225088
rect 438860 225140 438912 225146
rect 438860 225082 438912 225088
rect 438780 225026 438808 225082
rect 438780 224998 438900 225026
rect 438872 217410 438900 224998
rect 439780 220516 439832 220522
rect 439780 220458 439832 220464
rect 439792 217410 439820 220458
rect 440712 217410 440740 229774
rect 445668 229764 445720 229770
rect 445668 229706 445720 229712
rect 441620 226772 441672 226778
rect 441620 226714 441672 226720
rect 441632 225282 441660 226714
rect 441712 225956 441764 225962
rect 441712 225898 441764 225904
rect 441620 225276 441672 225282
rect 441620 225218 441672 225224
rect 441724 217410 441752 225898
rect 444840 225072 444892 225078
rect 444840 225014 444892 225020
rect 442356 224732 442408 224738
rect 442356 224674 442408 224680
rect 442368 217410 442396 224674
rect 444380 224256 444432 224262
rect 444380 224198 444432 224204
rect 443184 220380 443236 220386
rect 443184 220322 443236 220328
rect 443196 217410 443224 220322
rect 444392 217410 444420 224198
rect 425532 217382 425868 217410
rect 426360 217382 426696 217410
rect 427188 217382 427524 217410
rect 428016 217382 428352 217410
rect 428936 217382 429272 217410
rect 429764 217382 430100 217410
rect 430592 217382 430928 217410
rect 431420 217382 431756 217410
rect 432248 217382 432584 217410
rect 433352 217382 433412 217410
rect 433904 217382 434240 217410
rect 434824 217382 435160 217410
rect 435652 217382 435988 217410
rect 436480 217382 436816 217410
rect 437308 217382 437644 217410
rect 438136 217382 438472 217410
rect 438872 217382 439300 217410
rect 439792 217382 440128 217410
rect 440712 217382 441048 217410
rect 441724 217382 441876 217410
rect 442368 217382 442704 217410
rect 443196 217382 443532 217410
rect 444360 217382 444420 217410
rect 444852 217410 444880 225014
rect 445680 217410 445708 229706
rect 447416 229696 447468 229702
rect 447416 229638 447468 229644
rect 446588 220448 446640 220454
rect 446588 220390 446640 220396
rect 446600 217410 446628 220390
rect 447428 217410 447456 229638
rect 457444 229628 457496 229634
rect 457444 229570 457496 229576
rect 455788 229492 455840 229498
rect 455788 229434 455840 229440
rect 453856 227520 453908 227526
rect 453856 227462 453908 227468
rect 449716 226908 449768 226914
rect 449716 226850 449768 226856
rect 448796 226840 448848 226846
rect 448796 226782 448848 226788
rect 448808 225010 448836 226782
rect 449728 225078 449756 226850
rect 451556 225888 451608 225894
rect 451556 225830 451608 225836
rect 449716 225072 449768 225078
rect 449716 225014 449768 225020
rect 448244 225004 448296 225010
rect 448244 224946 448296 224952
rect 448796 225004 448848 225010
rect 448796 224946 448848 224952
rect 448256 217410 448284 224946
rect 450728 224324 450780 224330
rect 450728 224266 450780 224272
rect 449072 224120 449124 224126
rect 449072 224062 449124 224068
rect 449084 217410 449112 224062
rect 449900 220244 449952 220250
rect 449900 220186 449952 220192
rect 449912 217410 449940 220186
rect 450740 217410 450768 224266
rect 451568 217410 451596 225830
rect 453868 225758 453896 227462
rect 454960 225820 455012 225826
rect 454960 225762 455012 225768
rect 452660 225752 452712 225758
rect 452660 225694 452712 225700
rect 453856 225752 453908 225758
rect 453856 225694 453908 225700
rect 452672 217410 452700 225694
rect 454132 221332 454184 221338
rect 454132 221274 454184 221280
rect 453304 220312 453356 220318
rect 453304 220254 453356 220260
rect 453316 217410 453344 220254
rect 454144 217410 454172 221274
rect 454972 217410 455000 225762
rect 455800 217410 455828 229434
rect 456616 220108 456668 220114
rect 456616 220050 456668 220056
rect 456628 217410 456656 220050
rect 457456 217410 457484 229570
rect 459192 229560 459244 229566
rect 459192 229502 459244 229508
rect 458180 227588 458232 227594
rect 458180 227530 458232 227536
rect 458192 225826 458220 227530
rect 458180 225820 458232 225826
rect 458180 225762 458232 225768
rect 458456 225684 458508 225690
rect 458456 225626 458508 225632
rect 458468 217410 458496 225626
rect 459204 217410 459232 229502
rect 470968 229424 471020 229430
rect 470968 229366 471020 229372
rect 469128 229084 469180 229090
rect 469128 229026 469180 229032
rect 466368 228744 466420 228750
rect 466368 228686 466420 228692
rect 460940 227656 460992 227662
rect 460940 227598 460992 227604
rect 460952 225690 460980 227598
rect 466380 226234 466408 228686
rect 466368 226228 466420 226234
rect 466368 226170 466420 226176
rect 460940 225684 460992 225690
rect 460940 225626 460992 225632
rect 461676 225616 461728 225622
rect 461676 225558 461728 225564
rect 460940 224528 460992 224534
rect 460940 224470 460992 224476
rect 460020 220176 460072 220182
rect 460020 220118 460072 220124
rect 460032 217410 460060 220118
rect 460952 217410 460980 224470
rect 461688 217410 461716 225558
rect 469140 225554 469168 229026
rect 468392 225548 468444 225554
rect 468392 225490 468444 225496
rect 469128 225548 469180 225554
rect 469128 225490 469180 225496
rect 465080 225480 465132 225486
rect 465080 225422 465132 225428
rect 462504 224052 462556 224058
rect 462504 223994 462556 224000
rect 462516 217410 462544 223994
rect 464252 221400 464304 221406
rect 464252 221342 464304 221348
rect 463700 219904 463752 219910
rect 463700 219846 463752 219852
rect 463712 217410 463740 219846
rect 444852 217382 445188 217410
rect 445680 217382 446016 217410
rect 446600 217382 446936 217410
rect 447428 217382 447764 217410
rect 448256 217382 448592 217410
rect 449084 217382 449420 217410
rect 449912 217382 450248 217410
rect 450740 217382 451076 217410
rect 451568 217382 451904 217410
rect 452672 217382 452824 217410
rect 453316 217382 453652 217410
rect 454144 217382 454480 217410
rect 454972 217382 455308 217410
rect 455800 217382 456136 217410
rect 456628 217382 456964 217410
rect 457456 217382 457792 217410
rect 458468 217382 458712 217410
rect 459204 217382 459540 217410
rect 460032 217382 460368 217410
rect 460952 217382 461196 217410
rect 461688 217382 462024 217410
rect 462516 217382 462852 217410
rect 463680 217382 463740 217410
rect 464264 217410 464292 221342
rect 465092 217410 465120 225422
rect 467564 224800 467616 224806
rect 467564 224742 467616 224748
rect 465908 220040 465960 220046
rect 465908 219982 465960 219988
rect 465920 217410 465948 219982
rect 466736 219972 466788 219978
rect 466736 219914 466788 219920
rect 466748 217410 466776 219914
rect 467576 217410 467604 224742
rect 468404 217410 468432 225490
rect 469220 225412 469272 225418
rect 469220 225354 469272 225360
rect 469232 217410 469260 225354
rect 470140 219768 470192 219774
rect 470140 219710 470192 219716
rect 470152 217410 470180 219710
rect 470980 217410 471008 229366
rect 472624 229356 472676 229362
rect 472624 229298 472676 229304
rect 472072 229016 472124 229022
rect 472072 228958 472124 228964
rect 472084 225894 472112 228958
rect 472072 225888 472124 225894
rect 472072 225830 472124 225836
rect 471978 224632 472034 224641
rect 471978 224567 472034 224576
rect 471992 217410 472020 224567
rect 472636 217410 472664 229298
rect 483020 229288 483072 229294
rect 483020 229230 483072 229236
rect 477500 228948 477552 228954
rect 477500 228890 477552 228896
rect 474832 228880 474884 228886
rect 474832 228822 474884 228828
rect 474740 228812 474792 228818
rect 474740 228754 474792 228760
rect 474752 225622 474780 228754
rect 474740 225616 474792 225622
rect 474740 225558 474792 225564
rect 474844 225486 474872 228822
rect 474832 225480 474884 225486
rect 474832 225422 474884 225428
rect 477512 225418 477540 228890
rect 480258 227080 480314 227089
rect 480258 227015 480314 227024
rect 480272 225962 480300 227015
rect 481914 226264 481970 226273
rect 481914 226199 481970 226208
rect 480996 226160 481048 226166
rect 480996 226102 481048 226108
rect 480352 226024 480404 226030
rect 480352 225966 480404 225972
rect 480260 225956 480312 225962
rect 480260 225898 480312 225904
rect 477500 225412 477552 225418
rect 477500 225354 477552 225360
rect 474280 224868 474332 224874
rect 474280 224810 474332 224816
rect 473452 219836 473504 219842
rect 473452 219778 473504 219784
rect 473464 217410 473492 219778
rect 474292 217410 474320 224810
rect 478510 224768 478566 224777
rect 478510 224703 478566 224712
rect 475106 224496 475162 224505
rect 475106 224431 475162 224440
rect 475120 217410 475148 224431
rect 476026 224360 476082 224369
rect 476026 224295 476082 224304
rect 476040 217410 476068 224295
rect 477776 221468 477828 221474
rect 477776 221410 477828 221416
rect 476856 221264 476908 221270
rect 476856 221206 476908 221212
rect 476868 217410 476896 221206
rect 477788 217410 477816 221410
rect 478524 217410 478552 224703
rect 479340 224664 479392 224670
rect 479340 224606 479392 224612
rect 479352 217410 479380 224606
rect 480364 217410 480392 225966
rect 481008 217410 481036 226102
rect 481928 217410 481956 226199
rect 483032 217410 483060 229230
rect 515496 229220 515548 229226
rect 515496 229162 515548 229168
rect 507398 228984 507454 228993
rect 507398 228919 507454 228928
rect 484400 228676 484452 228682
rect 484400 228618 484452 228624
rect 483572 221536 483624 221542
rect 483572 221478 483624 221484
rect 483584 217410 483612 221478
rect 484412 217410 484440 228618
rect 494520 228608 494572 228614
rect 494520 228550 494572 228556
rect 488906 227352 488962 227361
rect 488906 227287 488962 227296
rect 488446 227216 488502 227225
rect 488446 227151 488502 227160
rect 485552 226406 485604 226412
rect 485552 226348 485604 226354
rect 464264 217382 464600 217410
rect 465092 217382 465428 217410
rect 465920 217382 466256 217410
rect 466748 217382 467084 217410
rect 467576 217382 467912 217410
rect 468404 217382 468740 217410
rect 469232 217382 469568 217410
rect 470152 217382 470488 217410
rect 470980 217382 471316 217410
rect 471992 217382 472144 217410
rect 472636 217382 472972 217410
rect 473464 217382 473800 217410
rect 474292 217382 474628 217410
rect 475120 217382 475456 217410
rect 476040 217382 476376 217410
rect 476868 217382 477204 217410
rect 477788 217382 478032 217410
rect 478524 217382 478860 217410
rect 479352 217382 479688 217410
rect 480364 217382 480516 217410
rect 481008 217382 481344 217410
rect 481928 217382 482264 217410
rect 483032 217382 483092 217410
rect 483584 217382 483920 217410
rect 484412 217382 484748 217410
rect 485564 217388 485592 226348
rect 487804 226228 487856 226234
rect 487804 226170 487856 226176
rect 487160 226092 487212 226098
rect 487160 226034 487212 226040
rect 486330 222048 486386 222057
rect 486330 221983 486386 221992
rect 486344 217410 486372 221983
rect 487172 218074 487200 226034
rect 487160 218068 487212 218074
rect 487160 218010 487212 218016
rect 487172 217410 487200 218010
rect 487816 217410 487844 226170
rect 488460 223650 488488 227151
rect 488448 223644 488500 223650
rect 488448 223586 488500 223592
rect 488920 221241 488948 227287
rect 489736 223644 489788 223650
rect 489736 223586 489788 223592
rect 488906 221232 488962 221241
rect 488906 221167 488962 221176
rect 488920 217410 488948 221167
rect 489748 217410 489776 223586
rect 494060 223576 494112 223582
rect 491942 223544 491998 223553
rect 494060 223518 494112 223524
rect 491942 223479 491998 223488
rect 491300 221808 491352 221814
rect 491300 221750 491352 221756
rect 490288 221672 490340 221678
rect 490288 221614 490340 221620
rect 490300 218142 490328 221614
rect 490288 218136 490340 218142
rect 490288 218078 490340 218084
rect 490300 217410 490328 218078
rect 491312 217410 491340 221750
rect 491956 217410 491984 223479
rect 492770 223408 492826 223417
rect 492770 223343 492826 223352
rect 492266 217592 492318 217598
rect 492266 217534 492318 217540
rect 492278 217410 492306 217534
rect 486344 217382 486740 217410
rect 487172 217382 487232 217410
rect 487816 217382 488152 217410
rect 488920 217382 488980 217410
rect 489748 217382 490144 217410
rect 490300 217382 490636 217410
rect 491312 217382 491464 217410
rect 491956 217396 492306 217410
rect 492784 217410 492812 223343
rect 494072 221610 494100 223518
rect 494060 221604 494112 221610
rect 494060 221546 494112 221552
rect 494072 217410 494100 221546
rect 491956 217382 492292 217396
rect 492784 217382 493272 217410
rect 494040 217382 494100 217410
rect 494532 217410 494560 228550
rect 506296 228540 506348 228546
rect 506296 228482 506348 228488
rect 496174 227488 496230 227497
rect 496174 227423 496230 227432
rect 495622 221912 495678 221921
rect 495622 221847 495678 221856
rect 495636 217410 495664 221847
rect 496188 220969 496216 227423
rect 502340 225956 502392 225962
rect 502340 225898 502392 225904
rect 499488 223440 499540 223446
rect 499488 223382 499540 223388
rect 499302 223272 499358 223281
rect 499302 223207 499358 223216
rect 497372 221876 497424 221882
rect 497372 221818 497424 221824
rect 496174 220960 496230 220969
rect 496174 220895 496230 220904
rect 496188 217410 496216 220895
rect 497384 217410 497412 221818
rect 497832 221740 497884 221746
rect 497832 221682 497884 221688
rect 494532 217382 494868 217410
rect 495636 217382 495696 217410
rect 496188 217382 496524 217410
rect 497352 217382 497412 217410
rect 497844 217410 497872 221682
rect 499316 220862 499344 223207
rect 499500 221882 499528 223382
rect 500222 223136 500278 223145
rect 500222 223071 500278 223080
rect 499488 221876 499540 221882
rect 499488 221818 499540 221824
rect 500236 221105 500264 223071
rect 501052 222012 501104 222018
rect 501052 221954 501104 221960
rect 501064 221338 501092 221954
rect 501236 221944 501288 221950
rect 501236 221886 501288 221892
rect 501052 221332 501104 221338
rect 501052 221274 501104 221280
rect 500222 221096 500278 221105
rect 500222 221031 500278 221040
rect 499304 220856 499356 220862
rect 499304 220798 499356 220804
rect 499316 217410 499344 220798
rect 500236 217410 500264 221031
rect 501064 217410 501092 221274
rect 497844 217382 498180 217410
rect 499008 217382 499344 217410
rect 499928 217382 500264 217410
rect 500756 217382 501092 217410
rect 501248 217410 501276 221886
rect 502352 217410 502380 225898
rect 503168 225752 503220 225758
rect 503168 225694 503220 225700
rect 503180 217410 503208 225694
rect 504822 223000 504878 223009
rect 504822 222935 504878 222944
rect 503720 222080 503772 222086
rect 503720 222022 503772 222028
rect 503732 217410 503760 222022
rect 504836 220930 504864 222935
rect 505744 222148 505796 222154
rect 505744 222090 505796 222096
rect 505756 221406 505784 222090
rect 505744 221400 505796 221406
rect 505744 221342 505796 221348
rect 504824 220924 504876 220930
rect 504824 220866 504876 220872
rect 504836 217410 504864 220866
rect 505756 217410 505784 221342
rect 506308 217410 506336 228482
rect 507412 217410 507440 228919
rect 512182 228848 512238 228857
rect 512182 228783 512238 228792
rect 511356 228472 511408 228478
rect 511356 228414 511408 228420
rect 507952 225820 508004 225826
rect 507952 225762 508004 225768
rect 501248 217382 501584 217410
rect 502352 217382 502748 217410
rect 503180 217382 503576 217410
rect 503732 217382 504068 217410
rect 504836 217382 504896 217410
rect 505756 217382 505816 217410
rect 506308 217382 506644 217410
rect 507412 217382 507808 217410
rect 418620 216980 418672 216986
rect 418620 216922 418672 216928
rect 418436 216912 418488 216918
rect 418436 216854 418488 216860
rect 417884 216844 417936 216850
rect 417884 216786 417936 216792
rect 52276 216776 52328 216782
rect 52276 216718 52328 216724
rect 169668 216776 169720 216782
rect 169668 216718 169720 216724
rect 187608 216776 187660 216782
rect 187608 216718 187660 216724
rect 52184 53916 52236 53922
rect 52184 53858 52236 53864
rect 52288 52426 52316 216718
rect 486712 216442 486740 217382
rect 490116 216442 490144 217382
rect 493244 216442 493272 217382
rect 502720 216510 502748 217382
rect 503548 216578 503576 217382
rect 503536 216572 503588 216578
rect 503536 216514 503588 216520
rect 502708 216504 502760 216510
rect 502708 216446 502760 216452
rect 507780 216442 507808 217382
rect 507964 217138 507992 225762
rect 509606 222864 509662 222873
rect 509606 222799 509662 222808
rect 509620 220998 509648 222799
rect 510620 221536 510672 221542
rect 510620 221478 510672 221484
rect 510632 221066 510660 221478
rect 510620 221060 510672 221066
rect 510620 221002 510672 221008
rect 508780 220992 508832 220998
rect 508780 220934 508832 220940
rect 509608 220992 509660 220998
rect 509608 220934 509660 220940
rect 508792 217410 508820 220934
rect 509620 217410 509648 220934
rect 510632 217410 510660 221002
rect 511368 217410 511396 228414
rect 508792 217382 509128 217410
rect 509620 217382 509956 217410
rect 510632 217382 510784 217410
rect 511368 217382 511704 217410
rect 507964 217122 508636 217138
rect 507964 217116 508648 217122
rect 507964 217110 508596 217116
rect 508596 217058 508648 217064
rect 512196 216458 512224 228783
rect 513472 225684 513524 225690
rect 513472 225626 513524 225632
rect 513378 222728 513434 222737
rect 513378 222663 513434 222672
rect 513392 221202 513420 222663
rect 513380 221196 513432 221202
rect 513380 221138 513432 221144
rect 513484 216458 513512 225626
rect 513840 223508 513892 223514
rect 513840 223450 513892 223456
rect 513852 217410 513880 223450
rect 514944 221196 514996 221202
rect 514944 221138 514996 221144
rect 514956 217410 514984 221138
rect 515508 218210 515536 229162
rect 535460 229152 535512 229158
rect 535460 229094 535512 229100
rect 518990 228712 519046 228721
rect 518990 228647 519046 228656
rect 518622 226128 518678 226137
rect 518622 226063 518678 226072
rect 516416 223372 516468 223378
rect 516416 223314 516468 223320
rect 515496 218204 515548 218210
rect 515496 218146 515548 218152
rect 515508 217410 515536 218146
rect 516428 217410 516456 223314
rect 517242 222592 517298 222601
rect 517242 222527 517298 222536
rect 513852 217382 514188 217410
rect 514956 217382 515016 217410
rect 515508 217382 515844 217410
rect 516428 217382 516672 217410
rect 517256 216458 517284 222527
rect 518636 218278 518664 226063
rect 518900 225548 518952 225554
rect 518900 225490 518952 225496
rect 518624 218272 518676 218278
rect 518624 218214 518676 218220
rect 518636 217410 518664 218214
rect 518420 217382 518664 217410
rect 518912 217410 518940 225490
rect 519004 221270 519032 228647
rect 525062 228576 525118 228585
rect 525062 228511 525118 228520
rect 520830 225992 520886 226001
rect 520830 225927 520886 225936
rect 518992 221264 519044 221270
rect 518992 221206 519044 221212
rect 520004 221264 520056 221270
rect 520004 221206 520056 221212
rect 520016 217410 520044 221206
rect 520844 218346 520872 225927
rect 523960 225888 524012 225894
rect 523960 225830 524012 225836
rect 523406 225720 523462 225729
rect 523406 225655 523462 225664
rect 521660 223304 521712 223310
rect 521660 223246 521712 223252
rect 520832 218340 520884 218346
rect 520832 218282 520884 218288
rect 520844 217410 520872 218282
rect 521672 217410 521700 223246
rect 522210 222456 522266 222465
rect 522210 222391 522266 222400
rect 518912 217382 519248 217410
rect 520016 217382 520076 217410
rect 520844 217382 520904 217410
rect 521672 217382 521732 217410
rect 522224 216458 522252 222391
rect 523420 218414 523448 225655
rect 523408 218408 523460 218414
rect 523408 218350 523460 218356
rect 523420 217410 523448 218350
rect 523972 217410 524000 225830
rect 525076 221474 525104 228511
rect 530122 228440 530178 228449
rect 530122 228375 530178 228384
rect 525798 225856 525854 225865
rect 525798 225791 525854 225800
rect 525064 221468 525116 221474
rect 525064 221410 525116 221416
rect 525076 217410 525104 221410
rect 525812 218482 525840 225791
rect 529020 225616 529072 225622
rect 528098 225584 528154 225593
rect 529020 225558 529072 225564
rect 528098 225519 528154 225528
rect 526444 223236 526496 223242
rect 526444 223178 526496 223184
rect 525800 218476 525852 218482
rect 525800 218418 525852 218424
rect 525812 217410 525840 218418
rect 526456 217410 526484 223178
rect 527270 222320 527326 222329
rect 527270 222255 527326 222264
rect 523420 217382 523480 217410
rect 523972 217382 524308 217410
rect 525076 217382 525136 217410
rect 525812 217382 525964 217410
rect 526456 217382 526792 217410
rect 524052 216572 524104 216578
rect 524052 216514 524104 216520
rect 512196 216442 512868 216458
rect 513360 216442 513696 216458
rect 517256 216442 517928 216458
rect 522224 216442 522896 216458
rect 524064 216442 524092 216514
rect 527284 216458 527312 222255
rect 528112 221882 528140 225519
rect 528100 221876 528152 221882
rect 528100 221818 528152 221824
rect 528112 217410 528140 221818
rect 529032 217410 529060 225558
rect 530136 221610 530164 228375
rect 534906 228304 534962 228313
rect 534906 228239 534962 228248
rect 533988 225480 534040 225486
rect 530674 225448 530730 225457
rect 533988 225422 534040 225428
rect 530674 225383 530730 225392
rect 530688 221950 530716 225383
rect 532792 225208 532844 225214
rect 532792 225150 532844 225156
rect 531504 223168 531556 223174
rect 531504 223110 531556 223116
rect 530676 221944 530728 221950
rect 530676 221886 530728 221892
rect 530124 221604 530176 221610
rect 530124 221546 530176 221552
rect 530136 217410 530164 221546
rect 530688 217410 530716 221886
rect 531516 217410 531544 223110
rect 532700 223100 532752 223106
rect 532700 223042 532752 223048
rect 528112 217382 528448 217410
rect 529032 217382 529368 217410
rect 530136 217382 530196 217410
rect 530688 217382 531024 217410
rect 531516 217382 531852 217410
rect 532712 216594 532740 223042
rect 532804 222154 532832 225150
rect 532792 222148 532844 222154
rect 532792 222090 532844 222096
rect 533436 222148 533488 222154
rect 533436 222090 533488 222096
rect 533448 217410 533476 222090
rect 534000 217410 534028 225422
rect 534920 221678 534948 228239
rect 535472 223514 535500 229094
rect 544108 228404 544160 228410
rect 544108 228346 544160 228352
rect 538310 228168 538366 228177
rect 538310 228103 538366 228112
rect 535460 223508 535512 223514
rect 535460 223450 535512 223456
rect 536104 223508 536156 223514
rect 536104 223450 536156 223456
rect 534908 221672 534960 221678
rect 534908 221614 534960 221620
rect 534920 217410 534948 221614
rect 536116 217410 536144 223450
rect 536564 223032 536616 223038
rect 536564 222974 536616 222980
rect 533448 217382 533508 217410
rect 534000 217382 534336 217410
rect 534920 217382 535256 217410
rect 536084 217382 536144 217410
rect 536576 217410 536604 222974
rect 537390 222184 537446 222193
rect 537390 222119 537446 222128
rect 536576 217382 536912 217410
rect 533068 217116 533120 217122
rect 533068 217058 533120 217064
rect 532680 216578 533016 216594
rect 532680 216572 533028 216578
rect 532680 216566 532976 216572
rect 532976 216514 533028 216520
rect 527284 216442 527956 216458
rect 533080 216442 533108 217058
rect 537404 216458 537432 222119
rect 538324 221746 538352 228103
rect 542726 228032 542782 228041
rect 542726 227967 542782 227976
rect 539048 225412 539100 225418
rect 539048 225354 539100 225360
rect 538864 223304 538916 223310
rect 538864 223246 538916 223252
rect 538312 221740 538364 221746
rect 538312 221682 538364 221688
rect 538876 217410 538904 223246
rect 538568 217382 538904 217410
rect 539060 217410 539088 225354
rect 541440 225344 541492 225350
rect 539322 225312 539378 225321
rect 541440 225286 541492 225292
rect 539322 225247 539378 225256
rect 539336 223310 539364 225247
rect 541452 223378 541480 225286
rect 541440 223372 541492 223378
rect 541440 223314 541492 223320
rect 539324 223304 539376 223310
rect 539324 223246 539376 223252
rect 540152 221740 540204 221746
rect 540152 221682 540204 221688
rect 540164 217410 540192 221682
rect 541452 217410 541480 223314
rect 541624 222964 541676 222970
rect 541624 222906 541676 222912
rect 539060 217382 539396 217410
rect 540164 217382 540224 217410
rect 541144 217382 541480 217410
rect 541636 217410 541664 222906
rect 542740 221814 542768 227967
rect 543648 222828 543700 222834
rect 543648 222770 543700 222776
rect 543660 222222 543688 222770
rect 543648 222216 543700 222222
rect 543648 222158 543700 222164
rect 542728 221808 542780 221814
rect 542728 221750 542780 221756
rect 542740 217410 542768 221750
rect 543660 217410 543688 222158
rect 541636 217382 541972 217410
rect 542740 217382 542800 217410
rect 543628 217382 543688 217410
rect 544120 217410 544148 228346
rect 547788 228336 547840 228342
rect 547788 228278 547840 228284
rect 546500 225276 546552 225282
rect 546500 225218 546552 225224
rect 545762 225176 545818 225185
rect 545762 225111 545818 225120
rect 545120 222896 545172 222902
rect 545120 222838 545172 222844
rect 545132 217410 545160 222838
rect 545776 222834 545804 225111
rect 546512 223242 546540 225218
rect 546500 223236 546552 223242
rect 546500 223178 546552 223184
rect 545764 222828 545816 222834
rect 545764 222770 545816 222776
rect 545776 217410 545804 222770
rect 546684 222760 546736 222766
rect 546684 222702 546736 222708
rect 546696 217410 546724 222702
rect 547800 222018 547828 228278
rect 549260 228268 549312 228274
rect 549260 228210 549312 228216
rect 548616 223236 548668 223242
rect 548616 223178 548668 223184
rect 547788 222012 547840 222018
rect 547788 221954 547840 221960
rect 547800 217410 547828 221954
rect 548628 217410 548656 223178
rect 549272 217410 549300 228210
rect 552020 228200 552072 228206
rect 552020 228142 552072 228148
rect 549352 222692 549404 222698
rect 549352 222634 549404 222640
rect 549364 221066 549392 222634
rect 549996 222624 550048 222630
rect 549996 222566 550048 222572
rect 549352 221060 549404 221066
rect 549352 221002 549404 221008
rect 550008 217410 550036 222566
rect 551100 221060 551152 221066
rect 551100 221002 551152 221008
rect 551112 217410 551140 221002
rect 552032 217410 552060 228142
rect 559288 228132 559340 228138
rect 559288 228074 559340 228080
rect 557632 228064 557684 228070
rect 557632 228006 557684 228012
rect 552570 227896 552626 227905
rect 552570 227831 552626 227840
rect 552584 222086 552612 227831
rect 554320 225140 554372 225146
rect 554320 225082 554372 225088
rect 553768 222624 553820 222630
rect 553768 222566 553820 222572
rect 552572 222080 552624 222086
rect 552572 222022 552624 222028
rect 553216 222080 553268 222086
rect 553216 222022 553268 222028
rect 553228 217410 553256 222022
rect 553780 217410 553808 222566
rect 554332 222562 554360 225082
rect 557448 223168 557500 223174
rect 557448 223110 557500 223116
rect 554228 222556 554280 222562
rect 554228 222498 554280 222504
rect 554320 222556 554372 222562
rect 554320 222498 554372 222504
rect 544120 217382 544456 217410
rect 545132 217382 545620 217410
rect 545776 217382 546112 217410
rect 546696 217382 547032 217410
rect 547800 217382 547860 217410
rect 548628 217382 548688 217410
rect 549272 217382 549516 217410
rect 550008 217382 550496 217410
rect 551112 217382 551172 217410
rect 552000 217382 552060 217410
rect 552920 217382 553256 217410
rect 553748 217382 553808 217410
rect 554240 217410 554268 222498
rect 556712 222488 556764 222494
rect 556712 222430 556764 222436
rect 555056 222420 555108 222426
rect 555056 222362 555108 222368
rect 554240 217382 554576 217410
rect 545592 216578 545620 217382
rect 550468 217122 550496 217382
rect 555068 217138 555096 222362
rect 556252 222352 556304 222358
rect 556252 222294 556304 222300
rect 556264 217410 556292 222294
rect 556232 217382 556292 217410
rect 556724 217410 556752 222430
rect 557460 222358 557488 223110
rect 557644 222358 557672 228006
rect 559104 224936 559156 224942
rect 559104 224878 559156 224884
rect 559116 222494 559144 224878
rect 559104 222488 559156 222494
rect 559104 222430 559156 222436
rect 557448 222352 557500 222358
rect 557448 222294 557500 222300
rect 557632 222352 557684 222358
rect 557632 222294 557684 222300
rect 557644 217410 557672 222294
rect 559116 217410 559144 222430
rect 556724 217382 557060 217410
rect 557644 217382 557888 217410
rect 558808 217382 559144 217410
rect 559300 217410 559328 228074
rect 560392 227928 560444 227934
rect 560392 227870 560444 227876
rect 560404 217682 560432 227870
rect 562876 227860 562928 227866
rect 562876 227802 562928 227808
rect 561218 225040 561274 225049
rect 561218 224975 561274 224984
rect 561232 222630 561260 224975
rect 561220 222624 561272 222630
rect 561220 222566 561272 222572
rect 560404 217654 560478 217682
rect 560450 217410 560478 217654
rect 561232 217410 561260 222566
rect 562888 222426 562916 227802
rect 563704 225072 563756 225078
rect 563704 225014 563756 225020
rect 563716 222698 563744 225014
rect 563704 222692 563756 222698
rect 563704 222634 563756 222640
rect 562876 222420 562928 222426
rect 562876 222362 562928 222368
rect 561772 221128 561824 221134
rect 561772 221070 561824 221076
rect 561784 217410 561812 221070
rect 562888 217410 562916 222362
rect 563716 217410 563744 222634
rect 564360 221513 564388 245618
rect 564440 227996 564492 228002
rect 564440 227938 564492 227944
rect 564346 221504 564402 221513
rect 564346 221439 564402 221448
rect 564452 217410 564480 227938
rect 566830 227760 566886 227769
rect 566830 227695 566886 227704
rect 566004 225004 566056 225010
rect 566004 224946 566056 224952
rect 566016 223106 566044 224946
rect 566004 223100 566056 223106
rect 566004 223042 566056 223048
rect 565176 222284 565228 222290
rect 565176 222226 565228 222232
rect 565188 217410 565216 222226
rect 566016 217410 566044 223042
rect 566844 217410 566872 227695
rect 567120 221785 567148 251194
rect 567292 248464 567344 248470
rect 567292 248406 567344 248412
rect 567304 222193 567332 248406
rect 567936 227792 567988 227798
rect 567936 227734 567988 227740
rect 567290 222184 567346 222193
rect 567290 222119 567346 222128
rect 567106 221776 567162 221785
rect 567106 221711 567162 221720
rect 567948 217410 567976 227734
rect 570236 227724 570288 227730
rect 570236 227666 570288 227672
rect 569314 227624 569370 227633
rect 569314 227559 569370 227568
rect 568578 224904 568634 224913
rect 568578 224839 568634 224848
rect 568592 222902 568620 224839
rect 568580 222896 568632 222902
rect 568580 222838 568632 222844
rect 568592 217410 568620 222838
rect 569328 217410 569356 227559
rect 570248 217410 570276 227666
rect 570880 217456 570932 217462
rect 559300 217382 559636 217410
rect 560450 217396 560524 217410
rect 560464 217382 560524 217396
rect 561232 217382 561292 217410
rect 561784 217382 562120 217410
rect 562888 217382 562948 217410
rect 563716 217382 563776 217410
rect 564452 217382 564696 217410
rect 565188 217382 565676 217410
rect 566016 217382 566352 217410
rect 566844 217382 567180 217410
rect 567948 217394 568344 217410
rect 567948 217388 568356 217394
rect 567948 217382 568304 217388
rect 555700 217184 555752 217190
rect 555068 217132 555700 217138
rect 560496 217138 560524 217382
rect 565648 217326 565676 217382
rect 568592 217382 568836 217410
rect 569328 217382 569664 217410
rect 570248 217404 570880 217410
rect 570248 217398 570932 217404
rect 570248 217382 570920 217398
rect 571410 217348 571438 255852
rect 572234 217352 572262 259115
rect 573060 217364 573088 262251
rect 654140 230988 654192 230994
rect 654140 230930 654192 230936
rect 654152 226334 654180 230930
rect 654152 226306 655192 226334
rect 607588 223576 607640 223582
rect 607588 223518 607640 223524
rect 574374 222184 574430 222193
rect 574374 222119 574430 222128
rect 573546 221504 573602 221513
rect 573546 221439 573602 221448
rect 573560 217410 573588 221439
rect 574388 217410 574416 222119
rect 575202 221776 575258 221785
rect 575202 221711 575258 221720
rect 575216 217410 575244 221711
rect 607128 218136 607180 218142
rect 607128 218078 607180 218084
rect 606668 218068 606720 218074
rect 606668 218010 606720 218016
rect 573560 217382 573896 217410
rect 574388 217382 574724 217410
rect 575216 217382 575552 217410
rect 568304 217330 568356 217336
rect 565636 217320 565688 217326
rect 565636 217262 565688 217268
rect 560760 217252 560812 217258
rect 560760 217194 560812 217200
rect 560772 217138 560800 217194
rect 555068 217126 555752 217132
rect 550456 217116 550508 217122
rect 555068 217110 555740 217126
rect 560464 217110 560800 217138
rect 550456 217058 550508 217064
rect 603448 216776 603500 216782
rect 603448 216718 603500 216724
rect 545580 216572 545632 216578
rect 545580 216514 545632 216520
rect 538036 216504 538088 216510
rect 537404 216452 538036 216458
rect 537404 216446 538088 216452
rect 486700 216436 486752 216442
rect 486700 216378 486752 216384
rect 490104 216436 490156 216442
rect 490104 216378 490156 216384
rect 493232 216436 493284 216442
rect 493232 216378 493284 216384
rect 507768 216436 507820 216442
rect 512196 216436 512880 216442
rect 512196 216430 512828 216436
rect 507768 216378 507820 216384
rect 513360 216436 513708 216442
rect 513360 216430 513656 216436
rect 512828 216378 512880 216384
rect 517256 216436 517940 216442
rect 517256 216430 517888 216436
rect 513656 216378 513708 216384
rect 522224 216436 522908 216442
rect 522224 216430 522856 216436
rect 517888 216378 517940 216384
rect 522856 216378 522908 216384
rect 524052 216436 524104 216442
rect 527284 216436 527968 216442
rect 527284 216430 527916 216436
rect 524052 216378 524104 216384
rect 527916 216378 527968 216384
rect 533068 216436 533120 216442
rect 537404 216430 538076 216446
rect 533068 216378 533120 216384
rect 582286 216200 582342 216209
rect 582286 216135 582342 216144
rect 580908 215756 580960 215762
rect 580908 215698 580960 215704
rect 580446 214704 580502 214713
rect 580446 214639 580502 214648
rect 580170 213208 580226 213217
rect 580170 213143 580226 213152
rect 580184 212634 580212 213143
rect 580172 212628 580224 212634
rect 580172 212570 580224 212576
rect 580460 212566 580488 214639
rect 580448 212560 580500 212566
rect 580448 212502 580500 212508
rect 580078 211712 580134 211721
rect 580078 211647 580134 211656
rect 580092 209846 580120 211647
rect 580080 209840 580132 209846
rect 580080 209782 580132 209788
rect 579802 208720 579858 208729
rect 579802 208655 579858 208664
rect 579816 207058 579844 208655
rect 579804 207052 579856 207058
rect 579804 206994 579856 207000
rect 580630 204232 580686 204241
rect 580630 204167 580686 204176
rect 580644 201550 580672 204167
rect 580632 201544 580684 201550
rect 580632 201486 580684 201492
rect 580722 198248 580778 198257
rect 580722 198183 580778 198192
rect 580736 197334 580764 198183
rect 580724 197328 580776 197334
rect 580724 197270 580776 197276
rect 579804 184884 579856 184890
rect 579804 184826 579856 184832
rect 579816 183161 579844 184826
rect 579802 183152 579858 183161
rect 579802 183087 579858 183096
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 180169 580212 182106
rect 580170 180160 580226 180169
rect 580170 180095 580226 180104
rect 580540 179376 580592 179382
rect 580540 179318 580592 179324
rect 580264 179308 580316 179314
rect 580264 179250 580316 179256
rect 580276 177177 580304 179250
rect 580552 178673 580580 179318
rect 580538 178664 580594 178673
rect 580538 178599 580594 178608
rect 580262 177168 580318 177177
rect 580262 177103 580318 177112
rect 580540 176656 580592 176662
rect 580540 176598 580592 176604
rect 580552 174185 580580 176598
rect 580816 176588 580868 176594
rect 580816 176530 580868 176536
rect 580828 175681 580856 176530
rect 580814 175672 580870 175681
rect 580814 175607 580870 175616
rect 580538 174176 580594 174185
rect 580538 174111 580594 174120
rect 579896 171148 579948 171154
rect 579896 171090 579948 171096
rect 579804 168564 579856 168570
rect 579804 168506 579856 168512
rect 579712 168428 579764 168434
rect 579712 168370 579764 168376
rect 579724 157593 579752 168370
rect 579816 159089 579844 168506
rect 579908 162081 579936 171090
rect 580264 165572 580316 165578
rect 580264 165514 580316 165520
rect 580276 163577 580304 165514
rect 580262 163568 580318 163577
rect 580262 163503 580318 163512
rect 579894 162072 579950 162081
rect 579894 162007 579950 162016
rect 579802 159080 579858 159089
rect 579802 159015 579858 159024
rect 579710 157584 579766 157593
rect 579710 157519 579766 157528
rect 580724 157412 580776 157418
rect 580724 157354 580776 157360
rect 580448 154624 580500 154630
rect 580448 154566 580500 154572
rect 579896 138032 579948 138038
rect 580460 138009 580488 154566
rect 580632 151836 580684 151842
rect 580632 151778 580684 151784
rect 580540 146328 580592 146334
rect 580540 146270 580592 146276
rect 579896 137974 579948 137980
rect 580446 138000 580502 138009
rect 579804 132524 579856 132530
rect 579804 132466 579856 132472
rect 579816 104961 579844 132466
rect 579908 110945 579936 137974
rect 580446 137935 580502 137944
rect 579988 135312 580040 135318
rect 579988 135254 580040 135260
rect 579894 110936 579950 110945
rect 579894 110871 579950 110880
rect 580000 106457 580028 135254
rect 580448 132592 580500 132598
rect 580448 132534 580500 132540
rect 580080 129804 580132 129810
rect 580080 129746 580132 129752
rect 579986 106448 580042 106457
rect 579986 106383 580042 106392
rect 579802 104952 579858 104961
rect 579802 104887 579858 104896
rect 580092 100337 580120 129746
rect 580264 127016 580316 127022
rect 580264 126958 580316 126964
rect 580172 124228 580224 124234
rect 580172 124170 580224 124176
rect 580078 100328 580134 100337
rect 580078 100263 580134 100272
rect 575664 95260 575716 95266
rect 575664 95202 575716 95208
rect 145380 53632 145432 53640
rect 145380 53574 145432 53580
rect 339408 53612 339460 53620
rect 84824 52686 85160 52714
rect 52276 52420 52328 52426
rect 52276 52362 52328 52368
rect 85132 45626 85160 52686
rect 145392 50810 145420 53574
rect 339408 53554 339460 53560
rect 543648 53612 543700 53622
rect 543648 53554 543700 53560
rect 149992 52686 150388 52714
rect 215832 52686 216168 52714
rect 281336 52686 281488 52714
rect 149992 52426 150020 52686
rect 149980 52420 150032 52426
rect 149980 52362 150032 52368
rect 145084 50782 145420 50810
rect 150360 49706 150388 52686
rect 184938 51096 184994 51105
rect 184938 51031 184994 51040
rect 184952 49706 184980 51031
rect 150348 49700 150400 49706
rect 150348 49642 150400 49648
rect 184940 49700 184992 49706
rect 184940 49642 184992 49648
rect 216140 48249 216168 52686
rect 281460 48346 281488 52686
rect 339420 52465 339448 53554
rect 339406 52456 339462 52465
rect 346826 52442 346854 52700
rect 412344 52686 412680 52714
rect 477848 52686 478184 52714
rect 346950 52456 347006 52465
rect 346826 52414 346950 52442
rect 339406 52391 339462 52400
rect 346950 52391 347006 52400
rect 412652 48414 412680 52686
rect 478156 48482 478184 52686
rect 543016 52686 543352 52714
rect 478144 48476 478196 48482
rect 478144 48418 478196 48424
rect 526168 48476 526220 48482
rect 526168 48418 526220 48424
rect 412640 48408 412692 48414
rect 412640 48350 412692 48356
rect 506388 48408 506440 48414
rect 506388 48350 506440 48356
rect 281448 48340 281500 48346
rect 281448 48282 281500 48288
rect 216126 48240 216182 48249
rect 216126 48175 216182 48184
rect 141804 46702 142370 46730
rect 85120 45620 85172 45626
rect 85120 45562 85172 45568
rect 141804 40202 141832 46702
rect 460664 45824 460716 45830
rect 460664 45766 460716 45772
rect 367100 45756 367152 45762
rect 367100 45698 367152 45704
rect 312820 45688 312872 45694
rect 312820 45630 312872 45636
rect 187332 45552 187384 45558
rect 187332 45494 187384 45500
rect 187344 42092 187372 45494
rect 312832 44198 312860 45630
rect 367112 44198 367140 45698
rect 312820 44192 312872 44198
rect 312820 44134 312872 44140
rect 367100 44192 367152 44198
rect 367100 44134 367152 44140
rect 310428 44124 310480 44130
rect 310428 44066 310480 44072
rect 365168 44124 365220 44130
rect 365168 44066 365220 44072
rect 223580 43104 223632 43110
rect 223580 43046 223632 43052
rect 194322 41848 194378 41857
rect 194074 41806 194322 41834
rect 194322 41783 194378 41792
rect 223592 41313 223620 43046
rect 310440 42106 310468 44066
rect 365180 42106 365208 44066
rect 390192 43172 390244 43178
rect 390192 43114 390244 43120
rect 310132 42078 310468 42106
rect 364918 42078 365208 42106
rect 307298 41848 307354 41857
rect 307004 41806 307298 41834
rect 361946 41848 362002 41857
rect 361790 41806 361946 41834
rect 307298 41783 307354 41792
rect 361946 41783 362002 41792
rect 390204 41313 390232 43114
rect 460676 42106 460704 45766
rect 475568 45620 475620 45626
rect 475568 45562 475620 45568
rect 470138 43208 470194 43217
rect 470138 43143 470194 43152
rect 470152 42650 470180 43143
rect 470152 42622 470198 42650
rect 475476 42628 475528 42634
rect 475476 42570 475528 42576
rect 460368 42078 460704 42106
rect 405582 41954 405872 41970
rect 405582 41948 405884 41954
rect 405582 41942 405832 41948
rect 405832 41890 405884 41896
rect 420644 41948 420696 41954
rect 420644 41890 420696 41896
rect 415490 41848 415546 41857
rect 415426 41806 415490 41834
rect 416778 41848 416834 41857
rect 416622 41806 416778 41834
rect 415490 41783 415546 41792
rect 419814 41848 419870 41857
rect 419750 41806 419814 41834
rect 416778 41783 416834 41792
rect 419814 41783 419870 41792
rect 420656 41750 420684 41890
rect 471702 41848 471758 41857
rect 471408 41806 471702 41834
rect 471702 41783 471758 41792
rect 420644 41744 420696 41750
rect 420644 41686 420696 41692
rect 223578 41304 223634 41313
rect 223578 41239 223634 41248
rect 390190 41304 390246 41313
rect 390190 41239 390246 41248
rect 475488 41041 475516 42570
rect 475474 41032 475530 41041
rect 475474 40967 475530 40976
rect 141758 40174 141832 40202
rect 141758 39984 141786 40174
rect 475580 38622 475608 45562
rect 506400 41410 506428 48350
rect 507860 48340 507912 48346
rect 507860 48282 507912 48288
rect 506388 41404 506440 41410
rect 506388 41346 506440 41352
rect 507872 41342 507900 48282
rect 521750 42120 521806 42129
rect 521806 42078 521870 42106
rect 526180 42092 526208 48418
rect 521750 42055 521806 42064
rect 513288 42016 513340 42022
rect 518532 42016 518584 42022
rect 513288 41958 513340 41964
rect 513194 41712 513250 41721
rect 513194 41647 513250 41656
rect 513208 41342 513236 41647
rect 513300 41410 513328 41958
rect 514864 41954 515154 41970
rect 518584 41964 518830 41970
rect 518532 41958 518830 41964
rect 514024 41948 514076 41954
rect 514024 41890 514076 41896
rect 514852 41948 515154 41954
rect 514904 41942 515154 41948
rect 518544 41942 518830 41958
rect 529322 41954 529704 41970
rect 529322 41948 529716 41954
rect 529322 41942 529664 41948
rect 514852 41890 514904 41896
rect 529664 41890 529716 41896
rect 530492 41948 530544 41954
rect 530492 41890 530544 41896
rect 513288 41404 513340 41410
rect 513288 41346 513340 41352
rect 507860 41336 507912 41342
rect 507860 41278 507912 41284
rect 513196 41336 513248 41342
rect 513196 41278 513248 41284
rect 514036 38622 514064 41890
rect 520370 41848 520426 41857
rect 520426 41806 520674 41834
rect 520370 41783 520426 41792
rect 530308 41404 530360 41410
rect 530308 41346 530360 41352
rect 530320 41177 530348 41346
rect 530400 41336 530452 41342
rect 530400 41278 530452 41284
rect 530306 41168 530362 41177
rect 530306 41103 530362 41112
rect 530412 41041 530440 41278
rect 530398 41032 530454 41041
rect 530398 40967 530454 40976
rect 530504 38622 530532 41890
rect 543016 38622 543044 52686
rect 543660 41313 543688 53554
rect 568580 51060 568632 51066
rect 568580 51002 568632 51008
rect 568592 41449 568620 51002
rect 575676 43178 575704 95202
rect 580184 92857 580212 124170
rect 580276 94353 580304 126958
rect 580356 124296 580408 124302
rect 580356 124238 580408 124244
rect 580262 94344 580318 94353
rect 580262 94279 580318 94288
rect 580170 92848 580226 92857
rect 580170 92783 580226 92792
rect 580368 91361 580396 124238
rect 580460 101969 580488 132534
rect 580552 127537 580580 146270
rect 580644 133521 580672 151778
rect 580736 136513 580764 157354
rect 580816 151904 580868 151910
rect 580816 151846 580868 151852
rect 580722 136504 580778 136513
rect 580722 136439 580778 136448
rect 580630 133512 580686 133521
rect 580630 133447 580686 133456
rect 580828 132025 580856 151846
rect 580920 146985 580948 215698
rect 582300 215354 582328 216135
rect 603460 215354 603488 216718
rect 582288 215348 582340 215354
rect 582288 215290 582340 215296
rect 599860 215348 599912 215354
rect 599860 215290 599912 215296
rect 603448 215348 603500 215354
rect 603448 215290 603500 215296
rect 604368 215348 604420 215354
rect 604368 215290 604420 215296
rect 598940 212628 598992 212634
rect 598940 212570 598992 212576
rect 582286 210216 582342 210225
rect 582286 210151 582342 210160
rect 582300 209914 582328 210151
rect 582288 209908 582340 209914
rect 582288 209850 582340 209856
rect 598952 207505 598980 212570
rect 599124 209908 599176 209914
rect 599124 209850 599176 209856
rect 598938 207496 598994 207505
rect 598938 207431 598994 207440
rect 582286 207224 582342 207233
rect 582286 207159 582342 207168
rect 582300 207126 582328 207159
rect 582288 207120 582340 207126
rect 582288 207062 582340 207068
rect 581458 205728 581514 205737
rect 581458 205663 581514 205672
rect 581472 204338 581500 205663
rect 599136 205465 599164 209850
rect 599872 209545 599900 215290
rect 599952 212560 600004 212566
rect 599952 212502 600004 212508
rect 599858 209536 599914 209545
rect 599858 209471 599914 209480
rect 599964 208593 599992 212502
rect 601148 209840 601200 209846
rect 601148 209782 601200 209788
rect 599950 208584 600006 208593
rect 599950 208519 600006 208528
rect 600964 207052 601016 207058
rect 600964 206994 601016 207000
rect 599122 205456 599178 205465
rect 599122 205391 599178 205400
rect 600976 204513 601004 206994
rect 601160 206553 601188 209782
rect 601516 207120 601568 207126
rect 601516 207062 601568 207068
rect 601146 206544 601202 206553
rect 601146 206479 601202 206488
rect 600962 204504 601018 204513
rect 600962 204439 601018 204448
rect 581460 204332 581512 204338
rect 581460 204274 581512 204280
rect 599952 204332 600004 204338
rect 599952 204274 600004 204280
rect 582286 202736 582342 202745
rect 582286 202671 582342 202680
rect 582300 201618 582328 202671
rect 599964 202473 599992 204274
rect 601528 203425 601556 207062
rect 601514 203416 601570 203425
rect 601514 203351 601570 203360
rect 599950 202464 600006 202473
rect 599950 202399 600006 202408
rect 582288 201612 582340 201618
rect 582288 201554 582340 201560
rect 599952 201612 600004 201618
rect 599952 201554 600004 201560
rect 598940 201544 598992 201550
rect 598940 201486 598992 201492
rect 598952 201385 598980 201486
rect 598938 201376 598994 201385
rect 598938 201311 598994 201320
rect 582286 201240 582342 201249
rect 582286 201175 582342 201184
rect 582300 200122 582328 201175
rect 599964 200433 599992 201554
rect 599950 200424 600006 200433
rect 599950 200359 600006 200368
rect 582288 200116 582340 200122
rect 582288 200058 582340 200064
rect 599952 200116 600004 200122
rect 599952 200058 600004 200064
rect 581090 199744 581146 199753
rect 581090 199679 581146 199688
rect 581104 198762 581132 199679
rect 599964 199345 599992 200058
rect 599950 199336 600006 199345
rect 599950 199271 600006 199280
rect 581092 198756 581144 198762
rect 581092 198698 581144 198704
rect 599124 198756 599176 198762
rect 599124 198698 599176 198704
rect 599136 198393 599164 198698
rect 599122 198384 599178 198393
rect 599122 198319 599178 198328
rect 582288 197396 582340 197402
rect 582288 197338 582340 197344
rect 599308 197396 599360 197402
rect 599308 197338 599360 197344
rect 582300 196761 582328 197338
rect 599320 197305 599348 197338
rect 599952 197328 600004 197334
rect 599306 197296 599362 197305
rect 599952 197270 600004 197276
rect 599306 197231 599362 197240
rect 582286 196752 582342 196761
rect 582286 196687 582342 196696
rect 599964 196353 599992 197270
rect 599950 196344 600006 196353
rect 599950 196279 600006 196288
rect 582286 195256 582342 195265
rect 582286 195191 582342 195200
rect 599950 195256 600006 195265
rect 599950 195191 600006 195200
rect 582196 194676 582248 194682
rect 582196 194618 582248 194624
rect 582208 193633 582236 194618
rect 582300 194614 582328 195191
rect 599124 194676 599176 194682
rect 599124 194618 599176 194624
rect 582288 194608 582340 194614
rect 582288 194550 582340 194556
rect 599136 194313 599164 194618
rect 599964 194614 599992 195191
rect 599952 194608 600004 194614
rect 599952 194550 600004 194556
rect 599122 194304 599178 194313
rect 599122 194239 599178 194248
rect 582194 193624 582250 193633
rect 582194 193559 582250 193568
rect 599950 193216 600006 193225
rect 599950 193151 600006 193160
rect 599122 192264 599178 192273
rect 599122 192199 599178 192208
rect 582286 192128 582342 192137
rect 582286 192063 582342 192072
rect 582196 191888 582248 191894
rect 582196 191830 582248 191836
rect 582208 190641 582236 191830
rect 582300 191826 582328 192063
rect 599136 191894 599164 192199
rect 599124 191888 599176 191894
rect 599124 191830 599176 191836
rect 599964 191826 599992 193151
rect 582288 191820 582340 191826
rect 582288 191762 582340 191768
rect 599952 191820 600004 191826
rect 599952 191762 600004 191768
rect 599858 191176 599914 191185
rect 599858 191111 599914 191120
rect 582194 190632 582250 190641
rect 582194 190567 582250 190576
rect 599872 190466 599900 191111
rect 581368 190460 581420 190466
rect 581368 190402 581420 190408
rect 599860 190460 599912 190466
rect 599860 190402 599912 190408
rect 581380 189145 581408 190402
rect 600962 190224 601018 190233
rect 600962 190159 601018 190168
rect 581366 189136 581422 189145
rect 581366 189071 581422 189080
rect 582196 187672 582248 187678
rect 582196 187614 582248 187620
rect 582286 187640 582342 187649
rect 582208 186153 582236 187614
rect 600976 187610 601004 190159
rect 601606 189136 601662 189145
rect 601606 189071 601662 189080
rect 601514 188184 601570 188193
rect 601514 188119 601570 188128
rect 582286 187575 582288 187584
rect 582340 187575 582342 187584
rect 600964 187604 601016 187610
rect 582288 187546 582340 187552
rect 600964 187546 601016 187552
rect 599950 187096 600006 187105
rect 599950 187031 600006 187040
rect 582194 186144 582250 186153
rect 582194 186079 582250 186088
rect 599858 185056 599914 185065
rect 599858 184991 599914 185000
rect 582288 184816 582340 184822
rect 582288 184758 582340 184764
rect 582300 184657 582328 184758
rect 582286 184648 582342 184657
rect 582286 184583 582342 184592
rect 599766 184104 599822 184113
rect 599766 184039 599822 184048
rect 582288 182096 582340 182102
rect 582288 182038 582340 182044
rect 582300 181665 582328 182038
rect 582286 181656 582342 181665
rect 582286 181591 582342 181600
rect 599674 180024 599730 180033
rect 599674 179959 599730 179968
rect 598938 176896 598994 176905
rect 598938 176831 598994 176840
rect 598952 176730 598980 176831
rect 581276 176724 581328 176730
rect 581276 176666 581328 176672
rect 598940 176724 598992 176730
rect 598940 176666 598992 176672
rect 581000 173936 581052 173942
rect 581000 173878 581052 173884
rect 581012 165073 581040 173878
rect 581288 168065 581316 176666
rect 599688 173874 599716 179959
rect 599780 179382 599808 184039
rect 599872 182170 599900 184991
rect 599964 184890 599992 187031
rect 600042 186144 600098 186153
rect 600042 186079 600098 186088
rect 599952 184884 600004 184890
rect 599952 184826 600004 184832
rect 599950 183016 600006 183025
rect 599950 182951 600006 182960
rect 599860 182164 599912 182170
rect 599860 182106 599912 182112
rect 599858 180976 599914 180985
rect 599858 180911 599914 180920
rect 599768 179376 599820 179382
rect 599768 179318 599820 179324
rect 599766 177984 599822 177993
rect 599766 177919 599822 177928
rect 582288 173868 582340 173874
rect 582288 173810 582340 173816
rect 599676 173868 599728 173874
rect 599676 173810 599728 173816
rect 582196 173800 582248 173806
rect 582196 173742 582248 173748
rect 582012 171216 582064 171222
rect 582208 171193 582236 173742
rect 582300 172689 582328 173810
rect 582286 172680 582342 172689
rect 582286 172615 582342 172624
rect 582012 171158 582064 171164
rect 582194 171184 582250 171193
rect 581736 168496 581788 168502
rect 581736 168438 581788 168444
rect 581460 168360 581512 168366
rect 581460 168302 581512 168308
rect 581274 168056 581330 168065
rect 581274 167991 581330 168000
rect 581472 166569 581500 168302
rect 581458 166560 581514 166569
rect 581458 166495 581514 166504
rect 580998 165064 581054 165073
rect 580998 164999 581054 165008
rect 581460 162920 581512 162926
rect 581460 162862 581512 162868
rect 581276 160268 581328 160274
rect 581276 160210 581328 160216
rect 581000 160200 581052 160206
rect 581000 160142 581052 160148
rect 580906 146976 580962 146985
rect 580906 146911 580962 146920
rect 581012 143993 581040 160142
rect 581092 157480 581144 157486
rect 581092 157422 581144 157428
rect 580998 143984 581054 143993
rect 580998 143919 581054 143928
rect 581104 141001 581132 157422
rect 581184 154692 581236 154698
rect 581184 154634 581236 154640
rect 581090 140992 581146 141001
rect 581090 140927 581146 140936
rect 581000 140820 581052 140826
rect 581000 140762 581052 140768
rect 580908 132660 580960 132666
rect 580908 132602 580960 132608
rect 580814 132016 580870 132025
rect 580814 131951 580870 131960
rect 580632 129872 580684 129878
rect 580632 129814 580684 129820
rect 580538 127528 580594 127537
rect 580538 127463 580594 127472
rect 580540 121508 580592 121514
rect 580540 121450 580592 121456
rect 580446 101960 580502 101969
rect 580446 101895 580502 101904
rect 580354 91352 580410 91361
rect 580354 91287 580410 91296
rect 580552 88369 580580 121450
rect 580644 98841 580672 129814
rect 580724 124364 580776 124370
rect 580724 124306 580776 124312
rect 580630 98832 580686 98841
rect 580630 98767 580686 98776
rect 580736 89865 580764 124306
rect 580816 121576 580868 121582
rect 580816 121518 580868 121524
rect 580722 89856 580778 89865
rect 580722 89791 580778 89800
rect 580538 88360 580594 88369
rect 580538 88295 580594 88304
rect 580828 86873 580856 121518
rect 580920 103465 580948 132602
rect 581012 113937 581040 140762
rect 581092 138100 581144 138106
rect 581092 138042 581144 138048
rect 580998 113928 581054 113937
rect 580998 113863 581054 113872
rect 581104 109449 581132 138042
rect 581196 135017 581224 154634
rect 581288 145489 581316 160210
rect 581368 160132 581420 160138
rect 581368 160074 581420 160080
rect 581274 145480 581330 145489
rect 581274 145415 581330 145424
rect 581276 140888 581328 140894
rect 581276 140830 581328 140836
rect 581182 135008 581238 135017
rect 581182 134943 581238 134952
rect 581184 129940 581236 129946
rect 581184 129882 581236 129888
rect 581090 109440 581146 109449
rect 581090 109375 581146 109384
rect 581000 107704 581052 107710
rect 581000 107646 581052 107652
rect 580906 103456 580962 103465
rect 580906 103391 580962 103400
rect 580908 99408 580960 99414
rect 580908 99350 580960 99356
rect 580814 86864 580870 86873
rect 580814 86799 580870 86808
rect 580816 84312 580868 84318
rect 580816 84254 580868 84260
rect 580724 84244 580776 84250
rect 580724 84186 580776 84192
rect 580632 84176 580684 84182
rect 580632 84118 580684 84124
rect 579988 82816 580040 82822
rect 579988 82758 580040 82764
rect 580000 82385 580028 82758
rect 579986 82376 580042 82385
rect 579620 82340 579672 82346
rect 579986 82311 580042 82320
rect 579620 82282 579672 82288
rect 579632 80889 579660 82282
rect 579618 80880 579674 80889
rect 579618 80815 579674 80824
rect 575756 80164 575808 80170
rect 575756 80106 575808 80112
rect 575664 43172 575716 43178
rect 575664 43114 575716 43120
rect 568578 41440 568634 41449
rect 568578 41375 568634 41384
rect 575768 41342 575796 80106
rect 578148 74792 578200 74798
rect 578148 74734 578200 74740
rect 578160 45558 578188 74734
rect 579620 60444 579672 60450
rect 579620 60386 579672 60392
rect 579632 59809 579660 60386
rect 579618 59800 579674 59809
rect 579618 59735 579674 59744
rect 579620 58336 579672 58342
rect 579618 58304 579620 58313
rect 579672 58304 579674 58313
rect 579618 58239 579674 58248
rect 580644 55321 580672 84118
rect 580736 61305 580764 84186
rect 580722 61296 580778 61305
rect 580722 61231 580778 61240
rect 580828 56817 580856 84254
rect 580814 56808 580870 56817
rect 580814 56743 580870 56752
rect 580630 55312 580686 55321
rect 580630 55247 580686 55256
rect 580920 53825 580948 99350
rect 581012 65793 581040 107646
rect 581092 104916 581144 104922
rect 581092 104858 581144 104864
rect 580998 65784 581054 65793
rect 580998 65719 581054 65728
rect 581104 62801 581132 104858
rect 581196 97345 581224 129882
rect 581288 115433 581316 140830
rect 581380 139505 581408 160074
rect 581472 148617 581500 162862
rect 581552 157548 581604 157554
rect 581552 157490 581604 157496
rect 581458 148608 581514 148617
rect 581458 148543 581514 148552
rect 581460 143608 581512 143614
rect 581460 143550 581512 143556
rect 581366 139496 581422 139505
rect 581366 139431 581422 139440
rect 581368 135380 581420 135386
rect 581368 135322 581420 135328
rect 581274 115424 581330 115433
rect 581274 115359 581330 115368
rect 581276 110560 581328 110566
rect 581276 110502 581328 110508
rect 581182 97336 581238 97345
rect 581182 97271 581238 97280
rect 581184 95328 581236 95334
rect 581184 95270 581236 95276
rect 581090 62792 581146 62801
rect 581090 62727 581146 62736
rect 580906 53816 580962 53825
rect 580906 53751 580962 53760
rect 581196 51066 581224 95270
rect 581288 70281 581316 110502
rect 581380 107953 581408 135322
rect 581472 118425 581500 143550
rect 581564 142497 581592 157490
rect 581748 156097 581776 168438
rect 581920 165708 581972 165714
rect 581920 165650 581972 165656
rect 581828 165640 581880 165646
rect 581828 165582 581880 165588
rect 581734 156088 581790 156097
rect 581734 156023 581790 156032
rect 581840 151609 581868 165582
rect 581932 153105 581960 165650
rect 582024 160585 582052 171158
rect 582194 171119 582250 171128
rect 599780 171086 599808 177919
rect 599872 176662 599900 180911
rect 599964 179314 599992 182951
rect 600056 182102 600084 186079
rect 601528 184822 601556 188119
rect 601620 187678 601648 189071
rect 601608 187672 601660 187678
rect 601608 187614 601660 187620
rect 601516 184816 601568 184822
rect 601516 184758 601568 184764
rect 600044 182096 600096 182102
rect 600044 182038 600096 182044
rect 600134 182064 600190 182073
rect 600134 181999 600190 182008
rect 599952 179308 600004 179314
rect 599952 179250 600004 179256
rect 600042 178936 600098 178945
rect 600042 178871 600098 178880
rect 599860 176656 599912 176662
rect 599860 176598 599912 176604
rect 599950 174856 600006 174865
rect 599950 174791 600006 174800
rect 599964 173942 599992 174791
rect 599952 173936 600004 173942
rect 599952 173878 600004 173884
rect 600056 173806 600084 178871
rect 600148 176594 600176 181999
rect 600136 176588 600188 176594
rect 600136 176530 600188 176536
rect 600318 175944 600374 175953
rect 600318 175879 600374 175888
rect 600134 173904 600190 173913
rect 600134 173839 600190 173848
rect 600044 173800 600096 173806
rect 600044 173742 600096 173748
rect 599858 172816 599914 172825
rect 599858 172751 599914 172760
rect 599872 171154 599900 172751
rect 599950 171864 600006 171873
rect 599950 171799 600006 171808
rect 599964 171222 599992 171799
rect 599952 171216 600004 171222
rect 599952 171158 600004 171164
rect 599860 171148 599912 171154
rect 599860 171090 599912 171096
rect 582288 171080 582340 171086
rect 582288 171022 582340 171028
rect 599768 171080 599820 171086
rect 599768 171022 599820 171028
rect 582300 169561 582328 171022
rect 599950 170776 600006 170785
rect 599950 170711 600006 170720
rect 599858 169824 599914 169833
rect 599858 169759 599914 169768
rect 582286 169552 582342 169561
rect 582286 169487 582342 169496
rect 599030 168736 599086 168745
rect 599030 168671 599086 168680
rect 599044 168502 599072 168671
rect 599032 168496 599084 168502
rect 599032 168438 599084 168444
rect 599872 168434 599900 169759
rect 599964 168570 599992 170711
rect 599952 168564 600004 168570
rect 599952 168506 600004 168512
rect 599860 168428 599912 168434
rect 599860 168370 599912 168376
rect 599858 167784 599914 167793
rect 599858 167719 599914 167728
rect 599872 165782 599900 167719
rect 600042 166696 600098 166705
rect 600042 166631 600098 166640
rect 582288 165776 582340 165782
rect 582288 165718 582340 165724
rect 599860 165776 599912 165782
rect 599860 165718 599912 165724
rect 599950 165744 600006 165753
rect 582104 162988 582156 162994
rect 582104 162930 582156 162936
rect 582010 160576 582066 160585
rect 582010 160511 582066 160520
rect 581918 153096 581974 153105
rect 581918 153031 581974 153040
rect 581826 151600 581882 151609
rect 581826 151535 581882 151544
rect 582116 150113 582144 162930
rect 582300 154601 582328 165718
rect 600056 165714 600084 166631
rect 599950 165679 600006 165688
rect 600044 165708 600096 165714
rect 599964 165646 599992 165679
rect 600044 165650 600096 165656
rect 599952 165640 600004 165646
rect 599952 165582 600004 165588
rect 600148 165578 600176 173839
rect 600332 168366 600360 175879
rect 600320 168360 600372 168366
rect 600320 168302 600372 168308
rect 600136 165572 600188 165578
rect 600136 165514 600188 165520
rect 599858 164656 599914 164665
rect 599858 164591 599914 164600
rect 599872 162994 599900 164591
rect 599950 163704 600006 163713
rect 599950 163639 600006 163648
rect 599860 162988 599912 162994
rect 599860 162930 599912 162936
rect 599964 162926 599992 163639
rect 599952 162920 600004 162926
rect 599952 162862 600004 162868
rect 599858 162616 599914 162625
rect 599858 162551 599914 162560
rect 599306 160576 599362 160585
rect 599306 160511 599362 160520
rect 599320 160138 599348 160511
rect 599872 160274 599900 162551
rect 599950 161664 600006 161673
rect 599950 161599 600006 161608
rect 599860 160268 599912 160274
rect 599860 160210 599912 160216
rect 599964 160206 599992 161599
rect 599952 160200 600004 160206
rect 599952 160142 600004 160148
rect 599308 160132 599360 160138
rect 599308 160074 599360 160080
rect 600042 159624 600098 159633
rect 600042 159559 600098 159568
rect 599950 158536 600006 158545
rect 599950 158471 600006 158480
rect 599858 157584 599914 157593
rect 599964 157554 599992 158471
rect 599858 157519 599914 157528
rect 599952 157548 600004 157554
rect 599872 157418 599900 157519
rect 599952 157490 600004 157496
rect 600056 157486 600084 159559
rect 600044 157480 600096 157486
rect 600044 157422 600096 157428
rect 599860 157412 599912 157418
rect 599860 157354 599912 157360
rect 599858 156496 599914 156505
rect 599858 156431 599914 156440
rect 599872 154630 599900 156431
rect 599950 155544 600006 155553
rect 599950 155479 600006 155488
rect 599964 154698 599992 155479
rect 599952 154692 600004 154698
rect 599952 154634 600004 154640
rect 599860 154624 599912 154630
rect 582286 154592 582342 154601
rect 599860 154566 599912 154572
rect 582286 154527 582342 154536
rect 599858 154456 599914 154465
rect 599858 154391 599914 154400
rect 599306 152416 599362 152425
rect 599306 152351 599362 152360
rect 599320 151978 599348 152351
rect 582196 151972 582248 151978
rect 582196 151914 582248 151920
rect 599308 151972 599360 151978
rect 599308 151914 599360 151920
rect 582102 150104 582158 150113
rect 582102 150039 582158 150048
rect 582012 149252 582064 149258
rect 582012 149194 582064 149200
rect 581828 149116 581880 149122
rect 581828 149058 581880 149064
rect 581644 146396 581696 146402
rect 581644 146338 581696 146344
rect 581550 142488 581606 142497
rect 581550 142423 581606 142432
rect 581552 138168 581604 138174
rect 581552 138110 581604 138116
rect 581458 118416 581514 118425
rect 581458 118351 581514 118360
rect 581564 112441 581592 138110
rect 581656 122913 581684 146338
rect 581736 143676 581788 143682
rect 581736 143618 581788 143624
rect 581642 122904 581698 122913
rect 581642 122839 581698 122848
rect 581748 119921 581776 143618
rect 581840 126041 581868 149058
rect 581920 140956 581972 140962
rect 581920 140898 581972 140904
rect 581826 126032 581882 126041
rect 581826 125967 581882 125976
rect 581734 119912 581790 119921
rect 581734 119847 581790 119856
rect 581932 116929 581960 140898
rect 582024 124545 582052 149194
rect 582104 143744 582156 143750
rect 582104 143686 582156 143692
rect 582010 124536 582066 124545
rect 582010 124471 582066 124480
rect 582012 121644 582064 121650
rect 582012 121586 582064 121592
rect 581918 116920 581974 116929
rect 581918 116855 581974 116864
rect 581828 116000 581880 116006
rect 581828 115942 581880 115948
rect 581644 113280 581696 113286
rect 581644 113222 581696 113228
rect 581550 112432 581606 112441
rect 581550 112367 581606 112376
rect 581460 110492 581512 110498
rect 581460 110434 581512 110440
rect 581366 107944 581422 107953
rect 581366 107879 581422 107888
rect 581368 104984 581420 104990
rect 581368 104926 581420 104932
rect 581274 70272 581330 70281
rect 581274 70207 581330 70216
rect 581380 64297 581408 104926
rect 581472 71777 581500 110434
rect 581552 107772 581604 107778
rect 581552 107714 581604 107720
rect 581458 71768 581514 71777
rect 581458 71703 581514 71712
rect 581564 67289 581592 107714
rect 581656 73273 581684 113222
rect 581736 113212 581788 113218
rect 581736 113154 581788 113160
rect 581748 76265 581776 113154
rect 581840 77897 581868 115942
rect 581920 113348 581972 113354
rect 581920 113290 581972 113296
rect 581826 77888 581882 77897
rect 581826 77823 581882 77832
rect 581734 76256 581790 76265
rect 581734 76191 581790 76200
rect 581932 74769 581960 113290
rect 582024 85377 582052 121586
rect 582116 121417 582144 143686
rect 582208 130529 582236 151914
rect 599872 151842 599900 154391
rect 599950 153504 600006 153513
rect 599950 153439 600006 153448
rect 599964 151910 599992 153439
rect 599952 151904 600004 151910
rect 599952 151846 600004 151852
rect 599860 151836 599912 151842
rect 599860 151778 599912 151784
rect 598938 151464 598994 151473
rect 598938 151399 598994 151408
rect 598952 149190 598980 151399
rect 599766 150376 599822 150385
rect 599766 150311 599822 150320
rect 599780 149258 599808 150311
rect 599950 149424 600006 149433
rect 599950 149359 600006 149368
rect 599768 149252 599820 149258
rect 599768 149194 599820 149200
rect 582288 149184 582340 149190
rect 582288 149126 582340 149132
rect 598940 149184 598992 149190
rect 598940 149126 598992 149132
rect 582194 130520 582250 130529
rect 582194 130455 582250 130464
rect 582300 129033 582328 149126
rect 599964 149122 599992 149359
rect 599952 149116 600004 149122
rect 599952 149058 600004 149064
rect 599858 148336 599914 148345
rect 599858 148271 599914 148280
rect 599872 146334 599900 148271
rect 599950 147384 600006 147393
rect 599950 147319 600006 147328
rect 599964 146402 599992 147319
rect 599952 146396 600004 146402
rect 599952 146338 600004 146344
rect 599860 146328 599912 146334
rect 599860 146270 599912 146276
rect 600042 146296 600098 146305
rect 600042 146231 600098 146240
rect 599858 145344 599914 145353
rect 599858 145279 599914 145288
rect 599872 143682 599900 145279
rect 599950 144256 600006 144265
rect 599950 144191 600006 144200
rect 599860 143676 599912 143682
rect 599860 143618 599912 143624
rect 599964 143614 599992 144191
rect 600056 143750 600084 146231
rect 600044 143744 600096 143750
rect 600044 143686 600096 143692
rect 599952 143608 600004 143614
rect 599952 143550 600004 143556
rect 599858 143304 599914 143313
rect 599858 143239 599914 143248
rect 599306 141264 599362 141273
rect 599306 141199 599362 141208
rect 599320 140826 599348 141199
rect 599872 140962 599900 143239
rect 599950 142216 600006 142225
rect 599950 142151 600006 142160
rect 599860 140956 599912 140962
rect 599860 140898 599912 140904
rect 599964 140894 599992 142151
rect 599952 140888 600004 140894
rect 599952 140830 600004 140836
rect 599308 140820 599360 140826
rect 599308 140762 599360 140768
rect 599858 140176 599914 140185
rect 599858 140111 599914 140120
rect 599872 138174 599900 140111
rect 600042 139224 600098 139233
rect 600042 139159 600098 139168
rect 599860 138168 599912 138174
rect 599860 138110 599912 138116
rect 599950 138136 600006 138145
rect 599950 138071 599952 138080
rect 600004 138071 600006 138080
rect 599952 138042 600004 138048
rect 600056 138038 600084 139159
rect 600044 138032 600096 138038
rect 600044 137974 600096 137980
rect 599858 137184 599914 137193
rect 599858 137119 599914 137128
rect 599872 135386 599900 137119
rect 599950 136096 600006 136105
rect 599950 136031 600006 136040
rect 599860 135380 599912 135386
rect 599860 135322 599912 135328
rect 599964 135318 599992 136031
rect 599952 135312 600004 135318
rect 599952 135254 600004 135260
rect 600042 135144 600098 135153
rect 600042 135079 600098 135088
rect 599858 134056 599914 134065
rect 599858 133991 599914 134000
rect 599872 132666 599900 133991
rect 599950 133104 600006 133113
rect 599950 133039 600006 133048
rect 599860 132660 599912 132666
rect 599860 132602 599912 132608
rect 599964 132598 599992 133039
rect 599952 132592 600004 132598
rect 599952 132534 600004 132540
rect 600056 132530 600084 135079
rect 600044 132524 600096 132530
rect 600044 132466 600096 132472
rect 598938 132016 598994 132025
rect 598938 131951 598994 131960
rect 598952 129810 598980 131951
rect 599766 131064 599822 131073
rect 599766 130999 599822 131008
rect 599780 129878 599808 130999
rect 599950 129976 600006 129985
rect 599950 129911 599952 129920
rect 600004 129911 600006 129920
rect 599952 129882 600004 129888
rect 599768 129872 599820 129878
rect 599768 129814 599820 129820
rect 598940 129804 598992 129810
rect 598940 129746 598992 129752
rect 582286 129024 582342 129033
rect 582286 128959 582342 128968
rect 599858 129024 599914 129033
rect 599858 128959 599914 128968
rect 599872 127090 599900 128959
rect 599950 127936 600006 127945
rect 599950 127871 600006 127880
rect 582196 127084 582248 127090
rect 582196 127026 582248 127032
rect 599860 127084 599912 127090
rect 599860 127026 599912 127032
rect 582102 121408 582158 121417
rect 582102 121343 582158 121352
rect 582104 116068 582156 116074
rect 582104 116010 582156 116016
rect 582010 85368 582066 85377
rect 582010 85303 582066 85312
rect 582116 79393 582144 116010
rect 582208 95849 582236 127026
rect 599964 127022 599992 127871
rect 599952 127016 600004 127022
rect 599952 126958 600004 126964
rect 600042 126984 600098 126993
rect 600042 126919 600098 126928
rect 599858 125896 599914 125905
rect 599858 125831 599914 125840
rect 599872 124302 599900 125831
rect 599950 124944 600006 124953
rect 599950 124879 600006 124888
rect 599964 124370 599992 124879
rect 599952 124364 600004 124370
rect 599952 124306 600004 124312
rect 599860 124296 599912 124302
rect 599860 124238 599912 124244
rect 600056 124234 600084 126919
rect 600044 124228 600096 124234
rect 600044 124170 600096 124176
rect 599858 123856 599914 123865
rect 599858 123791 599914 123800
rect 599582 121816 599638 121825
rect 599582 121751 599638 121760
rect 599596 121650 599624 121751
rect 599584 121644 599636 121650
rect 599584 121586 599636 121592
rect 599872 121514 599900 123791
rect 599950 122904 600006 122913
rect 599950 122839 600006 122848
rect 599964 121582 599992 122839
rect 599952 121576 600004 121582
rect 599952 121518 600004 121524
rect 599860 121508 599912 121514
rect 599860 121450 599912 121456
rect 600042 120864 600098 120873
rect 600042 120799 600098 120808
rect 599858 119776 599914 119785
rect 599858 119711 599914 119720
rect 599872 118862 599900 119711
rect 586428 118856 586480 118862
rect 586428 118798 586480 118804
rect 599860 118856 599912 118862
rect 599860 118798 599912 118804
rect 599950 118824 600006 118833
rect 583668 118788 583720 118794
rect 583668 118730 583720 118736
rect 582288 118720 582340 118726
rect 582288 118662 582340 118668
rect 582194 95840 582250 95849
rect 582194 95775 582250 95784
rect 582196 88392 582248 88398
rect 582196 88334 582248 88340
rect 582102 79384 582158 79393
rect 582102 79319 582158 79328
rect 581918 74760 581974 74769
rect 581918 74695 581974 74704
rect 581642 73264 581698 73273
rect 581642 73199 581698 73208
rect 581550 67280 581606 67289
rect 581550 67215 581606 67224
rect 581366 64288 581422 64297
rect 581366 64223 581422 64232
rect 582208 53922 582236 88334
rect 582300 83881 582328 118662
rect 582286 83872 582342 83881
rect 582286 83807 582342 83816
rect 583680 82346 583708 118730
rect 585140 89684 585192 89690
rect 585140 89626 585192 89632
rect 583760 84448 583812 84454
rect 583760 84390 583812 84396
rect 583668 82340 583720 82346
rect 583668 82282 583720 82288
rect 583772 60450 583800 84390
rect 583852 84380 583904 84386
rect 583852 84322 583904 84328
rect 583760 60444 583812 60450
rect 583760 60386 583812 60392
rect 583864 58342 583892 84322
rect 585152 80170 585180 89626
rect 586440 82822 586468 118798
rect 599950 118759 599952 118768
rect 600004 118759 600006 118768
rect 599952 118730 600004 118736
rect 600056 118726 600084 120799
rect 600044 118720 600096 118726
rect 600044 118662 600096 118668
rect 599858 117736 599914 117745
rect 599858 117671 599914 117680
rect 599872 116074 599900 117671
rect 599950 116784 600006 116793
rect 599950 116719 600006 116728
rect 599860 116068 599912 116074
rect 599860 116010 599912 116016
rect 599964 116006 599992 116719
rect 599952 116000 600004 116006
rect 599952 115942 600004 115948
rect 599858 115696 599914 115705
rect 599858 115631 599914 115640
rect 599872 113218 599900 115631
rect 600042 114744 600098 114753
rect 600042 114679 600098 114688
rect 599950 113656 600006 113665
rect 599950 113591 600006 113600
rect 599964 113286 599992 113591
rect 600056 113354 600084 114679
rect 600044 113348 600096 113354
rect 600044 113290 600096 113296
rect 599952 113280 600004 113286
rect 599952 113222 600004 113228
rect 599860 113212 599912 113218
rect 599860 113154 599912 113160
rect 598938 112704 598994 112713
rect 598938 112639 598994 112648
rect 598952 110498 598980 112639
rect 599950 111616 600006 111625
rect 599950 111551 600006 111560
rect 599964 110566 599992 111551
rect 599952 110560 600004 110566
rect 599952 110502 600004 110508
rect 598940 110492 598992 110498
rect 598940 110434 598992 110440
rect 599858 109576 599914 109585
rect 599858 109511 599914 109520
rect 599872 107778 599900 109511
rect 599950 108624 600006 108633
rect 599950 108559 600006 108568
rect 599860 107772 599912 107778
rect 599860 107714 599912 107720
rect 599964 107710 599992 108559
rect 599952 107704 600004 107710
rect 599952 107646 600004 107652
rect 599858 107536 599914 107545
rect 599858 107471 599914 107480
rect 599872 104990 599900 107471
rect 599950 106584 600006 106593
rect 599950 106519 600006 106528
rect 599860 104984 599912 104990
rect 599860 104926 599912 104932
rect 599964 104922 599992 106519
rect 600226 105496 600282 105505
rect 600226 105431 600282 105440
rect 599952 104916 600004 104922
rect 599952 104858 600004 104864
rect 599950 100464 600006 100473
rect 599950 100399 600006 100408
rect 599964 99414 599992 100399
rect 599952 99408 600004 99414
rect 599952 99350 600004 99356
rect 596180 95668 596232 95674
rect 596180 95610 596232 95616
rect 588084 95396 588136 95402
rect 588084 95338 588136 95344
rect 588096 88398 588124 95338
rect 588084 88392 588136 88398
rect 588084 88334 588136 88340
rect 596192 86018 596220 95610
rect 591948 86012 592000 86018
rect 591948 85954 592000 85960
rect 596180 86012 596232 86018
rect 596180 85954 596232 85960
rect 586428 82816 586480 82822
rect 586428 82758 586480 82764
rect 585140 80164 585192 80170
rect 585140 80106 585192 80112
rect 591960 69465 591988 85954
rect 600240 84250 600268 105431
rect 600502 104544 600558 104553
rect 600502 104479 600558 104488
rect 600318 102504 600374 102513
rect 600318 102439 600374 102448
rect 600332 84318 600360 102439
rect 600410 101416 600466 101425
rect 600410 101351 600466 101360
rect 600320 84312 600372 84318
rect 600320 84254 600372 84260
rect 600228 84244 600280 84250
rect 600228 84186 600280 84192
rect 600424 84182 600452 101351
rect 600516 84454 600544 104479
rect 600686 103456 600742 103465
rect 600686 103391 600742 103400
rect 600504 84448 600556 84454
rect 600504 84390 600556 84396
rect 600700 84386 600728 103391
rect 600688 84380 600740 84386
rect 600688 84322 600740 84328
rect 600412 84176 600464 84182
rect 600412 84118 600464 84124
rect 602988 82884 603040 82890
rect 602988 82826 603040 82832
rect 591946 69456 592002 69465
rect 591946 69391 592002 69400
rect 598940 66496 598992 66502
rect 598940 66438 598992 66444
rect 597468 58404 597520 58410
rect 597468 58346 597520 58352
rect 583852 58336 583904 58342
rect 583852 58278 583904 58284
rect 594800 57996 594852 58002
rect 594800 57938 594852 57944
rect 582196 53916 582248 53922
rect 582196 53858 582248 53864
rect 594812 53854 594840 57938
rect 594800 53848 594852 53854
rect 594800 53790 594852 53796
rect 581184 51060 581236 51066
rect 581184 51002 581236 51008
rect 597480 49745 597508 58346
rect 598952 58002 598980 66438
rect 603000 58410 603028 82826
rect 604380 81326 604408 215290
rect 606680 210202 606708 218010
rect 607140 210202 607168 218078
rect 607600 210202 607628 223518
rect 615040 223508 615092 223514
rect 615040 223450 615092 223456
rect 608048 223440 608100 223446
rect 608048 223382 608100 223388
rect 608060 210202 608088 223382
rect 614580 222148 614632 222154
rect 614580 222090 614632 222096
rect 614028 221944 614080 221950
rect 614028 221886 614080 221892
rect 613568 221876 613620 221882
rect 613568 221818 613620 221824
rect 610348 221536 610400 221542
rect 610348 221478 610400 221484
rect 609428 221400 609480 221406
rect 609428 221342 609480 221348
rect 608508 221332 608560 221338
rect 608508 221274 608560 221280
rect 608520 210202 608548 221274
rect 608968 216164 609020 216170
rect 608968 216106 609020 216112
rect 608980 210202 609008 216106
rect 609440 210202 609468 221342
rect 609888 216300 609940 216306
rect 609888 216242 609940 216248
rect 609900 210202 609928 216242
rect 610360 210202 610388 221478
rect 613108 218476 613160 218482
rect 613108 218418 613160 218424
rect 612648 218408 612700 218414
rect 612648 218350 612700 218356
rect 612188 218340 612240 218346
rect 612188 218282 612240 218288
rect 611728 218272 611780 218278
rect 611728 218214 611780 218220
rect 611268 218204 611320 218210
rect 611268 218146 611320 218152
rect 610808 216368 610860 216374
rect 610808 216310 610860 216316
rect 610820 210202 610848 216310
rect 611280 210202 611308 218146
rect 611740 210202 611768 218214
rect 612200 210202 612228 218282
rect 612660 210202 612688 218350
rect 613120 210202 613148 218418
rect 613580 210202 613608 221818
rect 614040 210202 614068 221886
rect 614592 210202 614620 222090
rect 615052 210202 615080 223450
rect 615960 223372 616012 223378
rect 615960 223314 616012 223320
rect 615500 223304 615552 223310
rect 615500 223246 615552 223252
rect 615512 210202 615540 223246
rect 615972 210202 616000 223314
rect 617340 223236 617392 223242
rect 617340 223178 617392 223184
rect 616880 222828 616932 222834
rect 616880 222770 616932 222776
rect 616420 222216 616472 222222
rect 616420 222158 616472 222164
rect 616432 210202 616460 222158
rect 616892 210202 616920 222770
rect 617352 210202 617380 223178
rect 618720 223168 618772 223174
rect 618720 223110 618772 223116
rect 618260 222556 618312 222562
rect 618260 222498 618312 222504
rect 617800 221060 617852 221066
rect 617800 221002 617852 221008
rect 617812 210202 617840 221002
rect 618272 210202 618300 222498
rect 618732 210202 618760 223110
rect 620560 223100 620612 223106
rect 620560 223042 620612 223048
rect 620100 222692 620152 222698
rect 620100 222634 620152 222640
rect 619640 222624 619692 222630
rect 619640 222566 619692 222572
rect 619180 222488 619232 222494
rect 619180 222430 619232 222436
rect 619192 210202 619220 222430
rect 619652 210202 619680 222566
rect 620112 210202 620140 222634
rect 620572 210202 620600 223042
rect 621020 222896 621072 222902
rect 621020 222838 621072 222844
rect 621032 210202 621060 222838
rect 634544 222420 634596 222426
rect 634544 222362 634596 222368
rect 633624 222352 633676 222358
rect 633624 222294 633676 222300
rect 632704 222080 632756 222086
rect 632704 222022 632756 222028
rect 631784 222012 631836 222018
rect 631784 221954 631836 221960
rect 630864 221808 630916 221814
rect 630864 221750 630916 221756
rect 630404 221740 630456 221746
rect 630404 221682 630456 221688
rect 629484 221672 629536 221678
rect 629484 221614 629536 221620
rect 628472 221604 628524 221610
rect 628472 221546 628524 221552
rect 627552 221468 627604 221474
rect 627552 221410 627604 221416
rect 622490 221368 622546 221377
rect 622490 221303 622546 221312
rect 621478 221232 621534 221241
rect 621478 221167 621534 221176
rect 621492 210202 621520 221167
rect 622032 217592 622084 217598
rect 622032 217534 622084 217540
rect 622044 210202 622072 217534
rect 622504 210202 622532 221303
rect 626632 221264 626684 221270
rect 626632 221206 626684 221212
rect 625712 221196 625764 221202
rect 625712 221138 625764 221144
rect 624792 220992 624844 220998
rect 624792 220934 624844 220940
rect 623872 220924 623924 220930
rect 623872 220866 623924 220872
rect 622952 220856 623004 220862
rect 622952 220798 623004 220804
rect 622964 210202 622992 220798
rect 623412 215892 623464 215898
rect 623412 215834 623464 215840
rect 623424 210202 623452 215834
rect 623884 210202 623912 220866
rect 624332 215824 624384 215830
rect 624332 215766 624384 215772
rect 624344 210202 624372 215766
rect 624804 210202 624832 220934
rect 625252 215960 625304 215966
rect 625252 215902 625304 215908
rect 625264 210202 625292 215902
rect 625724 210202 625752 221138
rect 626172 216028 626224 216034
rect 626172 215970 626224 215976
rect 626184 210202 626212 215970
rect 626644 210202 626672 221206
rect 627092 216096 627144 216102
rect 627092 216038 627144 216044
rect 627104 210202 627132 216038
rect 627564 210202 627592 221410
rect 628012 216232 628064 216238
rect 628012 216174 628064 216180
rect 628024 210202 628052 216174
rect 628484 210202 628512 221546
rect 628932 216436 628984 216442
rect 628932 216378 628984 216384
rect 628944 210202 628972 216378
rect 629496 210202 629524 221614
rect 629944 216504 629996 216510
rect 629944 216446 629996 216452
rect 629956 210202 629984 216446
rect 630416 210202 630444 221682
rect 630876 210202 630904 221750
rect 631324 216572 631376 216578
rect 631324 216514 631376 216520
rect 631336 210202 631364 216514
rect 631796 210202 631824 221954
rect 632244 217116 632296 217122
rect 632244 217058 632296 217064
rect 632256 210202 632284 217058
rect 632716 210202 632744 222022
rect 633164 217184 633216 217190
rect 633164 217126 633216 217132
rect 633176 210202 633204 217126
rect 633636 210202 633664 222294
rect 634084 217252 634136 217258
rect 634084 217194 634136 217200
rect 634096 210202 634124 217194
rect 634556 210202 634584 222362
rect 637854 221096 637910 221105
rect 637854 221031 637910 221040
rect 637394 220960 637450 220969
rect 637394 220895 637450 220904
rect 635924 217456 635976 217462
rect 635924 217398 635976 217404
rect 635464 217388 635516 217394
rect 635464 217330 635516 217336
rect 635004 217320 635056 217326
rect 635004 217262 635056 217268
rect 635016 210202 635044 217262
rect 635476 210202 635504 217330
rect 635936 210202 635964 217398
rect 636936 215688 636988 215694
rect 636936 215630 636988 215636
rect 636384 215620 636436 215626
rect 636384 215562 636436 215568
rect 636396 210202 636424 215562
rect 636948 210202 636976 215630
rect 637408 210202 637436 220895
rect 637868 210202 637896 221031
rect 648528 219700 648580 219706
rect 648528 219642 648580 219648
rect 639696 217048 639748 217054
rect 639696 216990 639748 216996
rect 638776 215756 638828 215762
rect 638776 215698 638828 215704
rect 638316 215552 638368 215558
rect 638316 215494 638368 215500
rect 638328 210202 638356 215494
rect 638788 210202 638816 215698
rect 639236 215348 639288 215354
rect 639236 215290 639288 215296
rect 639248 210202 639276 215290
rect 639708 210202 639736 216990
rect 640156 216980 640208 216986
rect 640156 216922 640208 216928
rect 640168 210202 640196 216922
rect 640616 216912 640668 216918
rect 640616 216854 640668 216860
rect 640628 210202 640656 216854
rect 641076 216844 641128 216850
rect 641076 216786 641128 216792
rect 641088 210202 641116 216786
rect 643204 210310 643508 210338
rect 643204 210202 643232 210310
rect 606648 210174 606708 210202
rect 607108 210174 607168 210202
rect 607568 210174 607628 210202
rect 608028 210174 608088 210202
rect 608488 210174 608548 210202
rect 608948 210174 609008 210202
rect 609408 210174 609468 210202
rect 609868 210174 609928 210202
rect 610328 210174 610388 210202
rect 610788 210174 610848 210202
rect 611248 210174 611308 210202
rect 611708 210174 611768 210202
rect 612168 210174 612228 210202
rect 612628 210174 612688 210202
rect 613088 210174 613148 210202
rect 613548 210174 613608 210202
rect 614008 210174 614068 210202
rect 614560 210174 614620 210202
rect 615020 210174 615080 210202
rect 615480 210174 615540 210202
rect 615940 210174 616000 210202
rect 616400 210174 616460 210202
rect 616860 210174 616920 210202
rect 617320 210174 617380 210202
rect 617780 210174 617840 210202
rect 618240 210174 618300 210202
rect 618700 210174 618760 210202
rect 619160 210174 619220 210202
rect 619620 210174 619680 210202
rect 620080 210174 620140 210202
rect 620540 210174 620600 210202
rect 621000 210174 621060 210202
rect 621460 210174 621520 210202
rect 622012 210174 622072 210202
rect 622472 210174 622532 210202
rect 622932 210174 622992 210202
rect 623392 210174 623452 210202
rect 623852 210174 623912 210202
rect 624312 210174 624372 210202
rect 624772 210174 624832 210202
rect 625232 210174 625292 210202
rect 625692 210174 625752 210202
rect 626152 210174 626212 210202
rect 626612 210174 626672 210202
rect 627072 210174 627132 210202
rect 627532 210174 627592 210202
rect 627992 210174 628052 210202
rect 628452 210174 628512 210202
rect 628912 210174 628972 210202
rect 629464 210174 629524 210202
rect 629924 210174 629984 210202
rect 630384 210174 630444 210202
rect 630844 210174 630904 210202
rect 631304 210174 631364 210202
rect 631764 210174 631824 210202
rect 632224 210174 632284 210202
rect 632684 210174 632744 210202
rect 633144 210174 633204 210202
rect 633604 210174 633664 210202
rect 634064 210174 634124 210202
rect 634524 210174 634584 210202
rect 634984 210174 635044 210202
rect 635444 210174 635504 210202
rect 635904 210174 635964 210202
rect 636364 210174 636424 210202
rect 636916 210174 636976 210202
rect 637376 210174 637436 210202
rect 637836 210174 637896 210202
rect 638296 210174 638356 210202
rect 638756 210174 638816 210202
rect 639216 210174 639276 210202
rect 639676 210174 639736 210202
rect 640136 210174 640196 210202
rect 640596 210174 640656 210202
rect 641056 210174 641116 210202
rect 642896 210174 643232 210202
rect 643480 210066 643508 210310
rect 646056 210310 646360 210338
rect 646056 210202 646084 210310
rect 645748 210174 646084 210202
rect 646332 210066 646360 210310
rect 648540 210202 648568 219642
rect 649908 219632 649960 219638
rect 649908 219574 649960 219580
rect 648816 210310 649120 210338
rect 648816 210202 648844 210310
rect 648508 210174 648844 210202
rect 649092 210066 649120 210310
rect 649920 210202 649948 219574
rect 651288 219564 651340 219570
rect 651288 219506 651340 219512
rect 650196 210310 650500 210338
rect 650196 210202 650224 210310
rect 649888 210174 650224 210202
rect 650472 210066 650500 210310
rect 651300 210202 651328 219506
rect 652760 219496 652812 219502
rect 652760 219438 652812 219444
rect 651668 210310 651972 210338
rect 651668 210202 651696 210310
rect 651268 210174 651696 210202
rect 651944 210066 651972 210310
rect 652772 210202 652800 219438
rect 654140 219428 654192 219434
rect 654140 219370 654192 219376
rect 653048 210310 653352 210338
rect 653048 210202 653076 210310
rect 652740 210174 653076 210202
rect 653324 210066 653352 210310
rect 654152 210202 654180 219370
rect 654428 210310 654732 210338
rect 654428 210202 654456 210310
rect 654120 210174 654456 210202
rect 654704 210066 654732 210310
rect 655164 210066 655192 226306
rect 655440 212498 655468 283183
rect 655532 220862 655560 292703
rect 655610 290456 655666 290465
rect 655610 290391 655666 290400
rect 655624 221066 655652 290391
rect 655716 245614 655744 293927
rect 655794 291544 655850 291553
rect 655794 291479 655850 291488
rect 655704 245608 655756 245614
rect 655704 245550 655756 245556
rect 655808 221202 655836 291479
rect 655900 267782 655928 296239
rect 656084 267986 656112 297463
rect 656254 295352 656310 295361
rect 656254 295287 656310 295296
rect 656268 268122 656296 295287
rect 666836 288584 666888 288590
rect 666836 288526 666888 288532
rect 656806 287328 656862 287337
rect 656806 287263 656862 287272
rect 656820 287162 656848 287263
rect 656808 287156 656860 287162
rect 656808 287098 656860 287104
rect 666744 284708 666796 284714
rect 666744 284650 666796 284656
rect 656806 282160 656862 282169
rect 656806 282095 656862 282104
rect 656820 281654 656848 282095
rect 656808 281648 656860 281654
rect 656808 281590 656860 281596
rect 666652 278996 666704 279002
rect 666652 278938 666704 278944
rect 666560 277364 666612 277370
rect 666560 277306 666612 277312
rect 656256 268116 656308 268122
rect 656256 268058 656308 268064
rect 656072 267980 656124 267986
rect 656072 267922 656124 267928
rect 655888 267776 655940 267782
rect 655888 267718 655940 267724
rect 656992 230920 657044 230926
rect 656992 230862 657044 230868
rect 656900 230852 656952 230858
rect 656900 230794 656952 230800
rect 655796 221196 655848 221202
rect 655796 221138 655848 221144
rect 655612 221060 655664 221066
rect 655612 221002 655664 221008
rect 655520 220856 655572 220862
rect 655520 220798 655572 220804
rect 655428 212492 655480 212498
rect 655428 212434 655480 212440
rect 655808 210310 656112 210338
rect 655808 210066 655836 210310
rect 643480 210038 643816 210066
rect 646332 210038 646668 210066
rect 649092 210038 649428 210066
rect 650472 210038 650808 210066
rect 651944 210038 652280 210066
rect 653324 210038 653660 210066
rect 654704 210038 655040 210066
rect 655164 210038 655836 210066
rect 656084 210066 656112 210310
rect 656912 210202 656940 230794
rect 657004 226334 657032 230862
rect 659660 230784 659712 230790
rect 659660 230726 659712 230732
rect 657004 226306 657952 226334
rect 657188 210310 657492 210338
rect 657188 210202 657216 210310
rect 656880 210174 657216 210202
rect 657464 210066 657492 210310
rect 657924 210066 657952 226306
rect 659672 215150 659700 230726
rect 662788 230716 662840 230722
rect 662788 230658 662840 230664
rect 659752 230580 659804 230586
rect 659752 230522 659804 230528
rect 659660 215144 659712 215150
rect 659660 215086 659712 215092
rect 658568 210310 658872 210338
rect 658568 210066 658596 210310
rect 656084 210038 656420 210066
rect 657464 210038 657800 210066
rect 657924 210038 658596 210066
rect 658844 210066 658872 210310
rect 659764 210202 659792 230522
rect 662604 230512 662656 230518
rect 662604 230454 662656 230460
rect 660764 215144 660816 215150
rect 660764 215086 660816 215092
rect 660040 210310 660344 210338
rect 660040 210202 660068 210310
rect 659732 210174 660068 210202
rect 660316 210066 660344 210310
rect 660776 210066 660804 215086
rect 661420 210310 661724 210338
rect 661420 210066 661448 210310
rect 658844 210038 659272 210066
rect 660316 210038 660652 210066
rect 660776 210038 661448 210066
rect 661696 210066 661724 210310
rect 662616 210202 662644 230454
rect 662696 230444 662748 230450
rect 662696 230386 662748 230392
rect 662492 210174 662644 210202
rect 662708 210118 662736 230386
rect 662696 210112 662748 210118
rect 661696 210038 662032 210066
rect 662696 210054 662748 210060
rect 662800 210066 662828 230658
rect 662880 230648 662932 230654
rect 662880 230590 662932 230596
rect 662892 226334 662920 230590
rect 662892 226306 663104 226334
rect 663076 210066 663104 226306
rect 666572 218618 666600 277306
rect 666560 218612 666612 218618
rect 666560 218554 666612 218560
rect 665732 217524 665784 217530
rect 665732 217466 665784 217472
rect 664812 216708 664864 216714
rect 664812 216650 664864 216656
rect 664352 216640 664404 216646
rect 664352 216582 664404 216588
rect 664364 210202 664392 216582
rect 664824 210202 664852 216650
rect 665272 215416 665324 215422
rect 665272 215358 665324 215364
rect 665284 210202 665312 215358
rect 665744 210202 665772 217466
rect 666192 215484 666244 215490
rect 666192 215426 666244 215432
rect 666204 210202 666232 215426
rect 664332 210174 664392 210202
rect 664792 210174 664852 210202
rect 665252 210174 665312 210202
rect 665712 210174 665772 210202
rect 666172 210174 666232 210202
rect 663524 210112 663576 210118
rect 662800 210038 662952 210066
rect 663076 210038 663412 210066
rect 663576 210060 663872 210066
rect 663524 210054 663872 210060
rect 663536 210038 663872 210054
rect 641812 209840 641864 209846
rect 641516 209788 641812 209794
rect 641516 209782 641864 209788
rect 642088 209840 642140 209846
rect 644664 209840 644716 209846
rect 642140 209788 642436 209794
rect 642088 209782 642436 209788
rect 641516 209766 641852 209782
rect 642100 209766 642436 209782
rect 644368 209788 644664 209794
rect 644368 209782 644716 209788
rect 644940 209840 644992 209846
rect 647424 209840 647476 209846
rect 644992 209788 645288 209794
rect 644940 209782 645288 209788
rect 644368 209766 644704 209782
rect 644952 209766 645288 209782
rect 647128 209788 647424 209794
rect 647128 209782 647476 209788
rect 647700 209840 647752 209846
rect 647752 209788 648048 209794
rect 647700 209782 648048 209788
rect 647128 209766 647464 209782
rect 647712 209766 648048 209782
rect 666558 209264 666614 209273
rect 666558 209199 666614 209208
rect 666572 205873 666600 209199
rect 666558 205864 666614 205873
rect 666558 205799 666614 205808
rect 666558 204232 666614 204241
rect 666558 204167 666614 204176
rect 666572 200841 666600 204167
rect 666558 200832 666614 200841
rect 666558 200767 666614 200776
rect 666558 199064 666614 199073
rect 666558 198999 666614 199008
rect 666572 195673 666600 198999
rect 666558 195664 666614 195673
rect 666558 195599 666614 195608
rect 666558 189000 666614 189009
rect 666558 188935 666614 188944
rect 666572 185609 666600 188935
rect 666558 185600 666614 185609
rect 666558 185535 666614 185544
rect 666558 183832 666614 183841
rect 666558 183767 666614 183776
rect 666572 180441 666600 183767
rect 666558 180432 666614 180441
rect 666558 180367 666614 180376
rect 666558 178800 666614 178809
rect 666558 178735 666614 178744
rect 666572 175409 666600 178735
rect 666558 175400 666614 175409
rect 666558 175335 666614 175344
rect 666558 173632 666614 173641
rect 666558 173567 666614 173576
rect 666572 170241 666600 173567
rect 666558 170232 666614 170241
rect 666558 170167 666614 170176
rect 666560 165980 666612 165986
rect 666560 165922 666612 165928
rect 606404 100014 606740 100042
rect 607384 100014 607444 100042
rect 606404 95266 606432 100014
rect 606392 95260 606444 95266
rect 606392 95202 606444 95208
rect 607220 93900 607272 93906
rect 607220 93842 607272 93848
rect 607232 89690 607260 93842
rect 607220 89684 607272 89690
rect 607220 89626 607272 89632
rect 604368 81320 604420 81326
rect 604368 81262 604420 81268
rect 602988 58404 603040 58410
rect 602988 58346 603040 58352
rect 598940 57996 598992 58002
rect 598940 57938 598992 57944
rect 600044 52488 600096 52494
rect 600044 52430 600096 52436
rect 597466 49736 597522 49745
rect 597466 49671 597522 49680
rect 578148 45552 578200 45558
rect 578148 45494 578200 45500
rect 600056 43217 600084 52430
rect 607416 45762 607444 100014
rect 607692 100014 608028 100042
rect 608152 100014 608672 100042
rect 608980 100014 609316 100042
rect 609960 100014 610204 100042
rect 607692 95674 607720 100014
rect 607680 95668 607732 95674
rect 607680 95610 607732 95616
rect 607496 95600 607548 95606
rect 607496 95542 607548 95548
rect 607404 45756 607456 45762
rect 607404 45698 607456 45704
rect 600042 43208 600098 43217
rect 600042 43143 600098 43152
rect 607508 41478 607536 95542
rect 608152 91094 608180 100014
rect 608980 95606 609008 100014
rect 608968 95600 609020 95606
rect 608968 95542 609020 95548
rect 607600 91066 608180 91094
rect 607600 45694 607628 91066
rect 610176 82890 610204 100014
rect 610268 100014 610604 100042
rect 610912 100014 611248 100042
rect 611556 100014 611892 100042
rect 612200 100014 612536 100042
rect 613028 100014 613180 100042
rect 613580 100014 613916 100042
rect 614560 100014 614896 100042
rect 615204 100014 615356 100042
rect 615848 100014 616184 100042
rect 616492 100014 616828 100042
rect 617136 100014 617472 100042
rect 617780 100014 618116 100042
rect 618424 100014 618760 100042
rect 619068 100014 619404 100042
rect 619712 100014 620048 100042
rect 620448 100014 620784 100042
rect 621092 100014 621428 100042
rect 621736 100014 622072 100042
rect 622380 100014 622716 100042
rect 623024 100014 623544 100042
rect 623668 100014 623728 100042
rect 610164 82884 610216 82890
rect 610164 82826 610216 82832
rect 607588 45688 607640 45694
rect 607588 45630 607640 45636
rect 607496 41472 607548 41478
rect 607496 41414 607548 41420
rect 610268 41410 610296 100014
rect 610348 95600 610400 95606
rect 610348 95542 610400 95548
rect 610360 45830 610388 95542
rect 610912 95402 610940 100014
rect 611556 95606 611584 100014
rect 611544 95600 611596 95606
rect 611544 95542 611596 95548
rect 610900 95396 610952 95402
rect 610900 95338 610952 95344
rect 612200 95334 612228 100014
rect 612188 95328 612240 95334
rect 612188 95270 612240 95276
rect 612740 75812 612792 75818
rect 612740 75754 612792 75760
rect 612752 66502 612780 75754
rect 612740 66496 612792 66502
rect 612740 66438 612792 66444
rect 613028 52494 613056 100014
rect 613580 93906 613608 100014
rect 614868 94994 614896 100014
rect 614856 94988 614908 94994
rect 614856 94930 614908 94936
rect 613568 93900 613620 93906
rect 613568 93842 613620 93848
rect 615328 77246 615356 100014
rect 616156 95606 616184 100014
rect 616144 95600 616196 95606
rect 616144 95542 616196 95548
rect 615408 94988 615460 94994
rect 615408 94930 615460 94936
rect 615316 77240 615368 77246
rect 615316 77182 615368 77188
rect 613016 52488 613068 52494
rect 613016 52430 613068 52436
rect 615420 49570 615448 94930
rect 616800 94926 616828 100014
rect 617444 95130 617472 100014
rect 617432 95124 617484 95130
rect 617432 95066 617484 95072
rect 616788 94920 616840 94926
rect 616788 94862 616840 94868
rect 618088 94586 618116 100014
rect 618732 94994 618760 100014
rect 619376 95538 619404 100014
rect 619364 95532 619416 95538
rect 619364 95474 619416 95480
rect 620020 95470 620048 100014
rect 620008 95464 620060 95470
rect 620008 95406 620060 95412
rect 620756 95334 620784 100014
rect 621400 95810 621428 100014
rect 622044 96150 622072 100014
rect 622032 96144 622084 96150
rect 622032 96086 622084 96092
rect 621388 95804 621440 95810
rect 621388 95746 621440 95752
rect 621204 95532 621256 95538
rect 621204 95474 621256 95480
rect 620744 95328 620796 95334
rect 620744 95270 620796 95276
rect 618720 94988 618772 94994
rect 618720 94930 618772 94936
rect 618076 94580 618128 94586
rect 618076 94522 618128 94528
rect 621216 86057 621244 95474
rect 622688 95266 622716 100014
rect 623228 95600 623280 95606
rect 623228 95542 623280 95548
rect 623516 95554 623544 100014
rect 623700 95878 623728 100014
rect 623976 100014 624312 100042
rect 624620 100014 624956 100042
rect 625600 100014 625936 100042
rect 626244 100014 626488 100042
rect 626980 100014 627316 100042
rect 627624 100014 627960 100042
rect 628268 100014 628328 100042
rect 623688 95872 623740 95878
rect 623688 95814 623740 95820
rect 623780 95600 623832 95606
rect 622676 95260 622728 95266
rect 622676 95202 622728 95208
rect 621940 95124 621992 95130
rect 621940 95066 621992 95072
rect 621202 86048 621258 86057
rect 621202 85983 621258 85992
rect 621952 83201 621980 95066
rect 622492 94920 622544 94926
rect 622492 94862 622544 94868
rect 622504 88913 622532 94862
rect 623136 94580 623188 94586
rect 623136 94522 623188 94528
rect 622490 88904 622546 88913
rect 622490 88839 622546 88848
rect 623148 84153 623176 94522
rect 623240 87961 623268 95542
rect 623516 95526 623636 95554
rect 623780 95542 623832 95548
rect 623504 95464 623556 95470
rect 623504 95406 623556 95412
rect 623320 94988 623372 94994
rect 623320 94930 623372 94936
rect 623226 87952 623282 87961
rect 623226 87887 623282 87896
rect 623332 85105 623360 94930
rect 623516 87009 623544 95406
rect 623502 87000 623558 87009
rect 623502 86935 623558 86944
rect 623318 85096 623374 85105
rect 623318 85031 623374 85040
rect 623134 84144 623190 84153
rect 623134 84079 623190 84088
rect 621938 83192 621994 83201
rect 621938 83127 621994 83136
rect 623608 75886 623636 95526
rect 623688 95260 623740 95266
rect 623688 95202 623740 95208
rect 623700 76022 623728 95202
rect 623792 90681 623820 95542
rect 623778 90672 623834 90681
rect 623778 90607 623834 90616
rect 623976 89729 624004 100014
rect 624620 95606 624648 100014
rect 624608 95600 624660 95606
rect 624608 95542 624660 95548
rect 625908 91633 625936 100014
rect 626460 92585 626488 100014
rect 626540 95736 626592 95742
rect 626540 95678 626592 95684
rect 626446 92576 626502 92585
rect 626446 92511 626502 92520
rect 625894 91624 625950 91633
rect 625894 91559 625950 91568
rect 623962 89720 624018 89729
rect 623962 89655 624018 89664
rect 626552 80209 626580 95678
rect 627288 93537 627316 100014
rect 627932 94489 627960 100014
rect 628300 95985 628328 100014
rect 628760 100014 628912 100042
rect 629556 100014 629708 100042
rect 630200 100014 630628 100042
rect 630844 100014 631180 100042
rect 631488 100014 631824 100042
rect 632132 100014 632468 100042
rect 632776 100014 633112 100042
rect 633512 100014 633848 100042
rect 634156 100014 634492 100042
rect 634800 100014 635136 100042
rect 635444 100014 635780 100042
rect 636088 100014 636332 100042
rect 636732 100014 637068 100042
rect 637376 100014 637528 100042
rect 638020 100014 638356 100042
rect 638664 100014 639000 100042
rect 639308 100014 639644 100042
rect 639952 100014 640104 100042
rect 640688 100014 640932 100042
rect 641332 100014 641668 100042
rect 628286 95976 628342 95985
rect 628286 95911 628342 95920
rect 628760 95826 628788 100014
rect 628728 95798 628788 95826
rect 629680 95826 629708 100014
rect 630600 95826 630628 100014
rect 631152 96082 631180 100014
rect 631140 96076 631192 96082
rect 631140 96018 631192 96024
rect 631796 95946 631824 100014
rect 632440 96082 632468 100014
rect 633084 96354 633112 100014
rect 633820 96626 633848 100014
rect 633808 96620 633860 96626
rect 633808 96562 633860 96568
rect 634464 96558 634492 100014
rect 634452 96552 634504 96558
rect 634452 96494 634504 96500
rect 633072 96348 633124 96354
rect 633072 96290 633124 96296
rect 635108 96082 635136 100014
rect 635752 96490 635780 100014
rect 635740 96484 635792 96490
rect 635740 96426 635792 96432
rect 636304 96422 636332 100014
rect 637040 96626 637068 100014
rect 636384 96620 636436 96626
rect 636384 96562 636436 96568
rect 637028 96620 637080 96626
rect 637028 96562 637080 96568
rect 636292 96416 636344 96422
rect 636292 96358 636344 96364
rect 635280 96348 635332 96354
rect 635280 96290 635332 96296
rect 632106 96076 632158 96082
rect 632106 96018 632158 96024
rect 632428 96076 632480 96082
rect 632428 96018 632480 96024
rect 634406 96076 634458 96082
rect 634406 96018 634458 96024
rect 635096 96076 635148 96082
rect 635096 96018 635148 96024
rect 631784 95940 631836 95946
rect 631784 95882 631836 95888
rect 629680 95798 629832 95826
rect 630600 95798 631028 95826
rect 632118 95812 632146 96018
rect 632980 95940 633032 95946
rect 632980 95882 633032 95888
rect 632992 95826 633020 95882
rect 632992 95798 633328 95826
rect 634418 95812 634446 96018
rect 635292 95826 635320 96290
rect 636396 95826 636424 96562
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637500 95606 637528 100014
rect 637580 96552 637632 96558
rect 637580 96494 637632 96500
rect 637592 95826 637620 96494
rect 637592 95798 637928 95826
rect 638328 95674 638356 100014
rect 638972 96218 639000 100014
rect 638960 96212 639012 96218
rect 638960 96154 639012 96160
rect 639006 96076 639058 96082
rect 639006 96018 639058 96024
rect 639018 95812 639046 96018
rect 639616 95946 639644 100014
rect 639880 96484 639932 96490
rect 639880 96426 639932 96432
rect 639604 95940 639656 95946
rect 639604 95882 639656 95888
rect 639892 95826 639920 96426
rect 640076 96014 640104 100014
rect 640340 96280 640392 96286
rect 640340 96222 640392 96228
rect 640064 96008 640116 96014
rect 640064 95950 640116 95956
rect 639892 95798 640228 95826
rect 640352 95742 640380 96222
rect 640904 95742 640932 100014
rect 640984 96416 641036 96422
rect 640984 96358 641036 96364
rect 640996 95826 641024 96358
rect 640996 95798 641332 95826
rect 640340 95736 640392 95742
rect 640340 95678 640392 95684
rect 640892 95736 640944 95742
rect 640892 95678 640944 95684
rect 638316 95668 638368 95674
rect 638316 95610 638368 95616
rect 641640 95606 641668 100014
rect 641732 100014 641976 100042
rect 642284 100014 642620 100042
rect 643264 100014 643600 100042
rect 643908 100014 644244 100042
rect 644552 100014 644796 100042
rect 641732 96286 641760 100014
rect 642180 96620 642232 96626
rect 642180 96562 642232 96568
rect 641720 96280 641772 96286
rect 641720 96222 641772 96228
rect 642192 95826 642220 96562
rect 642284 95985 642312 100014
rect 642824 96144 642876 96150
rect 642824 96086 642876 96092
rect 642270 95976 642326 95985
rect 642270 95911 642326 95920
rect 642192 95798 642528 95826
rect 642640 95668 642692 95674
rect 642640 95610 642692 95616
rect 637488 95600 637540 95606
rect 637488 95542 637540 95548
rect 641628 95600 641680 95606
rect 641628 95542 641680 95548
rect 627918 94480 627974 94489
rect 627918 94415 627974 94424
rect 627274 93528 627330 93537
rect 627274 93463 627330 93472
rect 642652 92721 642680 95610
rect 642732 95532 642784 95538
rect 642732 95474 642784 95480
rect 642744 95169 642772 95474
rect 642836 95470 642864 96086
rect 642916 95872 642968 95878
rect 642916 95814 642968 95820
rect 642824 95464 642876 95470
rect 642824 95406 642876 95412
rect 642824 95328 642876 95334
rect 642824 95270 642876 95276
rect 642730 95160 642786 95169
rect 642730 95095 642786 95104
rect 642836 95010 642864 95270
rect 642744 94982 642864 95010
rect 642638 92712 642694 92721
rect 642638 92647 642694 92656
rect 642744 91094 642772 94982
rect 642928 94874 642956 95814
rect 643008 95804 643060 95810
rect 643008 95746 643060 95752
rect 642652 91066 642772 91094
rect 642836 94846 642956 94874
rect 628562 81696 628618 81705
rect 628562 81631 628618 81640
rect 628576 81258 628604 81631
rect 631324 81320 631376 81326
rect 631324 81262 631376 81268
rect 628564 81252 628616 81258
rect 628564 81194 628616 81200
rect 629206 80880 629262 80889
rect 629206 80815 629262 80824
rect 626538 80200 626594 80209
rect 626538 80135 626594 80144
rect 628470 80200 628526 80209
rect 628470 80135 628526 80144
rect 623688 76016 623740 76022
rect 623688 75958 623740 75964
rect 623596 75880 623648 75886
rect 623596 75822 623648 75828
rect 623090 75812 623142 75818
rect 623090 75754 623142 75760
rect 623102 75548 623130 75754
rect 628484 75585 628512 80135
rect 629220 80102 629248 80815
rect 629208 80096 629260 80102
rect 629208 80038 629260 80044
rect 628470 75576 628526 75585
rect 631336 75562 631364 81262
rect 637028 81252 637080 81258
rect 637028 81194 637080 81200
rect 631520 80974 631856 81002
rect 631520 75818 631548 80974
rect 634174 80200 634230 80209
rect 634174 80135 634230 80144
rect 631508 75812 631560 75818
rect 631508 75754 631560 75760
rect 634188 75585 634216 80135
rect 634174 75576 634230 75585
rect 628526 75534 628820 75562
rect 631336 75534 631672 75562
rect 628470 75511 628526 75520
rect 637040 75562 637068 81194
rect 638972 80974 639308 81002
rect 634230 75534 634524 75562
rect 637040 75534 637376 75562
rect 634174 75511 634230 75520
rect 628484 75451 628512 75511
rect 634188 75451 634216 75511
rect 625632 75002 625968 75018
rect 638972 75002 639000 80974
rect 639880 80096 639932 80102
rect 639880 80038 639932 80044
rect 639892 75562 639920 80038
rect 640340 77240 640392 77246
rect 640340 77182 640392 77188
rect 639892 75534 640228 75562
rect 640352 75449 640380 77182
rect 641076 76016 641128 76022
rect 641076 75958 641128 75964
rect 640984 75880 641036 75886
rect 640984 75822 641036 75828
rect 640338 75440 640394 75449
rect 640338 75375 640394 75384
rect 625620 74996 625968 75002
rect 625672 74990 625968 74996
rect 638960 74996 639012 75002
rect 625620 74938 625672 74944
rect 638960 74938 639012 74944
rect 640996 72457 641024 75822
rect 640982 72448 641038 72457
rect 640982 72383 641038 72392
rect 641088 70961 641116 75958
rect 641074 70952 641130 70961
rect 641074 70887 641130 70896
rect 642652 65929 642680 91066
rect 642836 73409 642864 94846
rect 642916 94784 642968 94790
rect 642916 94726 642968 94732
rect 642822 73400 642878 73409
rect 642822 73335 642878 73344
rect 642928 68921 642956 94726
rect 642914 68912 642970 68921
rect 642914 68847 642970 68856
rect 643020 67425 643048 95746
rect 643100 95600 643152 95606
rect 643100 95542 643152 95548
rect 643006 67416 643062 67425
rect 643006 67351 643062 67360
rect 642638 65920 642694 65929
rect 642638 65855 642694 65864
rect 643112 64433 643140 95542
rect 643468 95124 643520 95130
rect 643468 95066 643520 95072
rect 643480 85270 643508 95066
rect 643572 94246 643600 100014
rect 643560 94240 643612 94246
rect 643560 94182 643612 94188
rect 644216 94110 644244 100014
rect 644768 94178 644796 100014
rect 644860 100014 645196 100042
rect 645840 100014 646176 100042
rect 646484 100014 646820 100042
rect 647220 100014 647556 100042
rect 647864 100014 648108 100042
rect 644860 95130 644888 100014
rect 646044 96008 646096 96014
rect 646044 95950 646096 95956
rect 645952 95940 646004 95946
rect 645952 95882 646004 95888
rect 645860 95736 645912 95742
rect 645860 95678 645912 95684
rect 644848 95124 644900 95130
rect 644848 95066 644900 95072
rect 644756 94172 644808 94178
rect 644756 94114 644808 94120
rect 644204 94104 644256 94110
rect 644204 94046 644256 94052
rect 643468 85264 643520 85270
rect 643468 85206 643520 85212
rect 645872 82249 645900 95678
rect 645964 87145 645992 95882
rect 646056 95010 646084 95950
rect 646148 95198 646176 100014
rect 646228 96212 646280 96218
rect 646228 96154 646280 96160
rect 646136 95192 646188 95198
rect 646136 95134 646188 95140
rect 646056 94982 646176 95010
rect 646044 94920 646096 94926
rect 646044 94862 646096 94868
rect 646056 89729 646084 94862
rect 646042 89720 646098 89729
rect 646042 89655 646098 89664
rect 645950 87136 646006 87145
rect 645950 87071 646006 87080
rect 646148 84697 646176 94982
rect 646240 94926 646268 96154
rect 646792 95334 646820 100014
rect 647528 95878 647556 100014
rect 647516 95872 647568 95878
rect 647516 95814 647568 95820
rect 646780 95328 646832 95334
rect 646780 95270 646832 95276
rect 646228 94920 646280 94926
rect 646228 94862 646280 94868
rect 647516 94716 647568 94722
rect 647516 94658 647568 94664
rect 647528 85202 647556 94658
rect 648080 94518 648108 100014
rect 648172 100014 648508 100042
rect 649152 100014 649396 100042
rect 648172 94722 648200 100014
rect 648620 94988 648672 94994
rect 648620 94930 648672 94936
rect 648160 94716 648212 94722
rect 648160 94658 648212 94664
rect 648068 94512 648120 94518
rect 648068 94454 648120 94460
rect 648632 85338 648660 94930
rect 648712 94852 648764 94858
rect 648712 94794 648764 94800
rect 648724 85406 648752 94794
rect 648804 94580 648856 94586
rect 648804 94522 648856 94528
rect 648816 85542 648844 94522
rect 649368 93906 649396 100014
rect 649460 100014 649796 100042
rect 650104 100014 650440 100042
rect 650748 100014 651084 100042
rect 651728 100014 652064 100042
rect 652372 100014 652708 100042
rect 653016 100014 653352 100042
rect 649460 94858 649488 100014
rect 649448 94852 649500 94858
rect 649448 94794 649500 94800
rect 650104 94586 650132 100014
rect 650748 94994 650776 100014
rect 652036 96490 652064 100014
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 651564 95872 651616 95878
rect 651564 95814 651616 95820
rect 650736 94988 650788 94994
rect 650736 94930 650788 94936
rect 650092 94580 650144 94586
rect 650092 94522 650144 94528
rect 649356 93900 649408 93906
rect 649356 93842 649408 93848
rect 651576 92585 651604 95814
rect 652680 95674 652708 100014
rect 652668 95668 652720 95674
rect 652668 95610 652720 95616
rect 653324 94790 653352 100014
rect 653416 100014 653752 100042
rect 654396 100014 654732 100042
rect 655040 100014 655376 100042
rect 655684 100014 656020 100042
rect 656328 100014 656664 100042
rect 656972 100014 657308 100042
rect 653312 94784 653364 94790
rect 653312 94726 653364 94732
rect 653416 94722 653444 100014
rect 654704 96558 654732 100014
rect 654692 96552 654744 96558
rect 654692 96494 654744 96500
rect 651840 94716 651892 94722
rect 651840 94658 651892 94664
rect 653404 94716 653456 94722
rect 653404 94658 653456 94664
rect 651562 92576 651618 92585
rect 651562 92511 651618 92520
rect 648804 85536 648856 85542
rect 648804 85478 648856 85484
rect 651852 85474 651880 94658
rect 652760 94172 652812 94178
rect 652760 94114 652812 94120
rect 652772 90681 652800 94114
rect 654048 94104 654100 94110
rect 654048 94046 654100 94052
rect 654060 91497 654088 94046
rect 655348 93401 655376 100014
rect 655992 96626 656020 100014
rect 655980 96620 656032 96626
rect 655980 96562 656032 96568
rect 656636 94722 656664 100014
rect 656992 95600 657044 95606
rect 656992 95542 657044 95548
rect 656624 94716 656676 94722
rect 656624 94658 656676 94664
rect 656900 94580 656952 94586
rect 656900 94522 656952 94528
rect 656912 93906 656940 94522
rect 656900 93900 656952 93906
rect 656900 93842 656952 93848
rect 655334 93392 655390 93401
rect 655334 93327 655390 93336
rect 654046 91488 654102 91497
rect 654046 91423 654102 91432
rect 657004 91094 657032 95542
rect 657084 95260 657136 95266
rect 657084 95202 657136 95208
rect 656912 91066 657032 91094
rect 652758 90672 652814 90681
rect 652758 90607 652814 90616
rect 656912 90409 656940 91066
rect 656898 90400 656954 90409
rect 656898 90335 656954 90344
rect 657096 88874 657124 95202
rect 657280 94654 657308 100014
rect 657372 100014 657616 100042
rect 657924 100014 658260 100042
rect 658904 100014 659148 100042
rect 657372 94761 657400 100014
rect 657728 99816 657780 99822
rect 657728 99758 657780 99764
rect 657740 95132 657768 99758
rect 657924 95266 657952 100014
rect 659120 96558 659148 100014
rect 659212 100014 659548 100042
rect 660284 100014 660620 100042
rect 658280 96552 658332 96558
rect 658280 96494 658332 96500
rect 659108 96552 659160 96558
rect 659108 96494 659160 96500
rect 657912 95260 657964 95266
rect 657912 95202 657964 95208
rect 658292 95132 658320 96494
rect 659212 95606 659240 100014
rect 659568 96620 659620 96626
rect 659568 96562 659620 96568
rect 659200 95600 659252 95606
rect 659200 95542 659252 95548
rect 659580 95132 659608 96562
rect 660592 95538 660620 100014
rect 660914 99822 660942 100028
rect 661572 100014 661908 100042
rect 662216 100014 662276 100042
rect 662860 100014 663288 100042
rect 663504 100014 663656 100042
rect 660902 99816 660954 99822
rect 660902 99758 660954 99764
rect 661880 96626 661908 100014
rect 661868 96620 661920 96626
rect 661868 96562 661920 96568
rect 661960 96484 662012 96490
rect 661960 96426 662012 96432
rect 660580 95532 660632 95538
rect 660580 95474 660632 95480
rect 661408 95532 661460 95538
rect 661408 95474 661460 95480
rect 661420 95132 661448 95474
rect 661972 95132 662000 96426
rect 662248 95577 662276 100014
rect 663064 96620 663116 96626
rect 663064 96562 663116 96568
rect 662512 96552 662564 96558
rect 662512 96494 662564 96500
rect 662234 95568 662290 95577
rect 662234 95503 662290 95512
rect 662524 95132 662552 96494
rect 663076 95132 663104 96562
rect 657358 94752 657414 94761
rect 657358 94687 657414 94696
rect 657268 94648 657320 94654
rect 657268 94590 657320 94596
rect 658568 94586 658858 94602
rect 658556 94580 658858 94586
rect 658608 94574 658858 94580
rect 658556 94522 658608 94528
rect 659844 94512 659896 94518
rect 660396 94512 660448 94518
rect 659896 94460 660146 94466
rect 659844 94454 660146 94460
rect 660448 94460 660698 94466
rect 660396 94454 660698 94460
rect 659856 94438 660146 94454
rect 660408 94438 660698 94454
rect 663260 93809 663288 100014
rect 663340 95328 663392 95334
rect 663340 95270 663392 95276
rect 663246 93800 663302 93809
rect 663246 93735 663302 93744
rect 663352 93129 663380 95270
rect 663432 95192 663484 95198
rect 663432 95134 663484 95140
rect 663338 93120 663394 93129
rect 663338 93055 663394 93064
rect 663444 92313 663472 95134
rect 663524 94648 663576 94654
rect 663524 94590 663576 94596
rect 663430 92304 663486 92313
rect 663430 92239 663486 92248
rect 663536 89593 663564 94590
rect 663522 89584 663578 89593
rect 663522 89519 663578 89528
rect 658016 88874 658306 88890
rect 659488 88874 659594 88890
rect 663628 88874 663656 100014
rect 663800 95668 663852 95674
rect 663800 95610 663852 95616
rect 663708 94784 663760 94790
rect 663708 94726 663760 94732
rect 663720 90409 663748 94726
rect 663706 90400 663762 90409
rect 663706 90335 663762 90344
rect 657084 88868 657136 88874
rect 657084 88810 657136 88816
rect 658004 88868 658306 88874
rect 658056 88862 658306 88868
rect 659476 88868 659594 88874
rect 658004 88810 658056 88816
rect 659528 88862 659594 88868
rect 663616 88868 663668 88874
rect 659476 88810 659528 88816
rect 663616 88810 663668 88816
rect 662142 88768 662198 88777
rect 661986 88726 662142 88754
rect 663812 88754 663840 95610
rect 663892 94716 663944 94722
rect 663892 94658 663944 94664
rect 663904 91089 663932 94658
rect 663890 91080 663946 91089
rect 663890 91015 663946 91024
rect 662538 88726 663840 88754
rect 662142 88703 662198 88712
rect 651840 85468 651892 85474
rect 651840 85410 651892 85416
rect 648712 85400 648764 85406
rect 648712 85342 648764 85348
rect 657188 85338 657216 88196
rect 657740 85542 657768 88196
rect 657728 85536 657780 85542
rect 657728 85478 657780 85484
rect 658844 85474 658872 88196
rect 658832 85468 658884 85474
rect 658832 85410 658884 85416
rect 648620 85332 648672 85338
rect 648620 85274 648672 85280
rect 657176 85332 657228 85338
rect 657176 85274 657228 85280
rect 660132 85270 660160 88196
rect 660684 85406 660712 88196
rect 660672 85400 660724 85406
rect 660672 85342 660724 85348
rect 660120 85264 660172 85270
rect 660120 85206 660172 85212
rect 661420 85202 661448 88196
rect 647516 85196 647568 85202
rect 647516 85138 647568 85144
rect 661408 85196 661460 85202
rect 661408 85138 661460 85144
rect 646134 84688 646190 84697
rect 646134 84623 646190 84632
rect 645858 82240 645914 82249
rect 645858 82175 645914 82184
rect 643098 64424 643154 64433
rect 643098 64359 643154 64368
rect 650000 49632 650052 49638
rect 650000 49574 650052 49580
rect 615408 49564 615460 49570
rect 615408 49506 615460 49512
rect 650012 46986 650040 49574
rect 666572 49065 666600 165922
rect 666664 128058 666692 278938
rect 666756 179414 666784 284650
rect 666848 226334 666876 288526
rect 669412 287156 669464 287162
rect 669412 287098 669464 287104
rect 669228 281648 669280 281654
rect 669228 281590 669280 281596
rect 666848 226306 666968 226334
rect 666836 218612 666888 218618
rect 666836 218554 666888 218560
rect 666848 187694 666876 218554
rect 666940 206990 666968 226306
rect 666928 206984 666980 206990
rect 666928 206926 666980 206932
rect 666848 187666 666968 187694
rect 666756 179386 666876 179414
rect 666742 168600 666798 168609
rect 666742 168535 666798 168544
rect 666756 165209 666784 168535
rect 666742 165200 666798 165209
rect 666742 165135 666798 165144
rect 666742 163568 666798 163577
rect 666742 163503 666798 163512
rect 666756 160177 666784 163503
rect 666742 160168 666798 160177
rect 666742 160103 666798 160112
rect 666742 158400 666798 158409
rect 666742 158335 666798 158344
rect 666756 155009 666784 158335
rect 666848 157350 666876 179386
rect 666940 165986 666968 187666
rect 666928 165980 666980 165986
rect 666928 165922 666980 165928
rect 666836 157344 666888 157350
rect 666836 157286 666888 157292
rect 666742 155000 666798 155009
rect 666742 154935 666798 154944
rect 666742 153368 666798 153377
rect 666742 153303 666798 153312
rect 666756 149977 666784 153303
rect 666742 149968 666798 149977
rect 666742 149903 666798 149912
rect 666742 148200 666798 148209
rect 666742 148135 666798 148144
rect 666756 144945 666784 148135
rect 666742 144936 666798 144945
rect 666742 144871 666798 144880
rect 666742 143168 666798 143177
rect 666742 143103 666798 143112
rect 666756 139777 666784 143103
rect 666742 139768 666798 139777
rect 666742 139703 666798 139712
rect 666742 132968 666798 132977
rect 666742 132903 666798 132912
rect 666756 129577 666784 132903
rect 669240 132666 669268 281590
rect 669320 280220 669372 280226
rect 669320 280162 669372 280168
rect 669332 132802 669360 280162
rect 669424 178838 669452 287098
rect 669504 287088 669556 287094
rect 669504 287030 669556 287036
rect 669412 178832 669464 178838
rect 669412 178774 669464 178780
rect 669516 178158 669544 287030
rect 669596 284980 669648 284986
rect 669596 284922 669648 284928
rect 669504 178152 669556 178158
rect 669504 178094 669556 178100
rect 669608 177750 669636 284922
rect 670884 213648 670936 213654
rect 670884 213590 670936 213596
rect 669688 212492 669740 212498
rect 669688 212434 669740 212440
rect 669596 177744 669648 177750
rect 669596 177686 669648 177692
rect 669700 132938 669728 212434
rect 670698 194032 670754 194041
rect 670698 193967 670754 193976
rect 670712 190641 670740 193967
rect 670698 190632 670754 190641
rect 670698 190567 670754 190576
rect 670340 168342 670400 168351
rect 670340 168273 670400 168282
rect 669688 132932 669740 132938
rect 669688 132874 669740 132880
rect 669320 132796 669372 132802
rect 669320 132738 669372 132744
rect 669228 132660 669280 132666
rect 669228 132602 669280 132608
rect 666742 129568 666798 129577
rect 666742 129503 666798 129512
rect 666664 128030 666784 128058
rect 666650 127936 666706 127945
rect 666650 127871 666706 127880
rect 666664 124545 666692 127871
rect 666650 124536 666706 124545
rect 666650 124471 666706 124480
rect 666650 122904 666706 122913
rect 666650 122839 666706 122848
rect 666664 119513 666692 122839
rect 666650 119504 666706 119513
rect 666650 119439 666706 119448
rect 666756 115938 666784 128030
rect 670356 117793 670384 168273
rect 670506 167932 670566 167941
rect 670506 167863 670566 167872
rect 670346 117784 670402 117793
rect 670346 117719 670402 117728
rect 670522 116163 670550 167863
rect 670698 138136 670754 138145
rect 670698 138071 670754 138080
rect 670712 134745 670740 138071
rect 670698 134736 670754 134745
rect 670698 134671 670754 134680
rect 670502 116154 670558 116163
rect 670502 116089 670558 116098
rect 666744 115932 666796 115938
rect 666744 115874 666796 115880
rect 670896 107545 670924 213590
rect 671804 213580 671856 213586
rect 671804 213522 671856 213528
rect 671712 176860 671764 176866
rect 671712 176802 671764 176808
rect 671724 132326 671752 176802
rect 671712 132320 671764 132326
rect 671712 132262 671764 132268
rect 671816 130082 671844 213522
rect 671896 213444 671948 213450
rect 671896 213386 671948 213392
rect 671908 131714 671936 213386
rect 672000 178809 672028 884954
rect 673288 747974 673316 892978
rect 673196 747946 673316 747974
rect 673196 723246 673224 747946
rect 673276 732488 673328 732494
rect 673276 732430 673328 732436
rect 673288 728822 673316 732430
rect 673276 728816 673328 728822
rect 673276 728758 673328 728764
rect 673184 723240 673236 723246
rect 673184 723182 673236 723188
rect 673380 723178 673408 894610
rect 676048 894402 676076 896679
rect 676126 896064 676182 896073
rect 676126 895999 676182 896008
rect 676036 894396 676088 894402
rect 676036 894338 676088 894344
rect 676140 894334 676168 895999
rect 676128 894328 676180 894334
rect 676128 894270 676180 894276
rect 676034 893072 676090 893081
rect 676034 893007 676036 893016
rect 676088 893007 676090 893016
rect 676036 892978 676088 892984
rect 679162 892664 679218 892673
rect 679162 892599 679218 892608
rect 676034 892256 676090 892265
rect 676034 892191 676090 892200
rect 676048 891546 676076 892191
rect 674748 891540 674800 891546
rect 674748 891482 674800 891488
rect 676036 891540 676088 891546
rect 676036 891482 676088 891488
rect 673736 887868 673788 887874
rect 673736 887810 673788 887816
rect 673748 874206 673776 887810
rect 674288 887460 674340 887466
rect 674288 887402 674340 887408
rect 674196 886032 674248 886038
rect 674196 885974 674248 885980
rect 673736 874200 673788 874206
rect 673736 874142 673788 874148
rect 674208 869446 674236 885974
rect 674300 869990 674328 887402
rect 674760 883214 674788 891482
rect 676034 891032 676090 891041
rect 676034 890967 676090 890976
rect 676048 890730 676076 890967
rect 674932 890724 674984 890730
rect 674932 890666 674984 890672
rect 676036 890724 676088 890730
rect 676036 890666 676088 890672
rect 674392 883186 674788 883214
rect 674392 875906 674420 883186
rect 674944 880818 674972 890666
rect 676034 890624 676090 890633
rect 676034 890559 676090 890568
rect 676048 889098 676076 890559
rect 675024 889092 675076 889098
rect 675024 889034 675076 889040
rect 676036 889092 676088 889098
rect 676036 889034 676088 889040
rect 674760 880790 674972 880818
rect 674472 880728 674524 880734
rect 674472 880670 674524 880676
rect 674380 875900 674432 875906
rect 674380 875842 674432 875848
rect 674288 869984 674340 869990
rect 674288 869926 674340 869932
rect 674196 869440 674248 869446
rect 674196 869382 674248 869388
rect 674484 867610 674512 880670
rect 674564 878688 674616 878694
rect 674564 878630 674616 878636
rect 674576 873798 674604 878630
rect 674656 878620 674708 878626
rect 674656 878562 674708 878568
rect 674668 874342 674696 878562
rect 674656 874336 674708 874342
rect 674656 874278 674708 874284
rect 674656 874200 674708 874206
rect 674656 874142 674708 874148
rect 674564 873792 674616 873798
rect 674564 873734 674616 873740
rect 674668 869378 674696 874142
rect 674760 872506 674788 880790
rect 674840 880660 674892 880666
rect 674840 880602 674892 880608
rect 674852 877266 674880 880602
rect 674932 878552 674984 878558
rect 674932 878494 674984 878500
rect 674840 877260 674892 877266
rect 674840 877202 674892 877208
rect 674840 875900 674892 875906
rect 674840 875842 674892 875848
rect 674748 872500 674800 872506
rect 674748 872442 674800 872448
rect 674852 872386 674880 875842
rect 674944 872658 674972 878494
rect 675036 872778 675064 889034
rect 676034 888992 676090 889001
rect 676034 888927 676090 888936
rect 676048 888758 676076 888927
rect 675208 888752 675260 888758
rect 675208 888694 675260 888700
rect 676036 888752 676088 888758
rect 676036 888694 676088 888700
rect 675220 880734 675248 888694
rect 676034 888584 676090 888593
rect 676034 888519 676090 888528
rect 676048 887874 676076 888519
rect 679070 888176 679126 888185
rect 679070 888111 679126 888120
rect 676036 887868 676088 887874
rect 676036 887810 676088 887816
rect 676034 887768 676090 887777
rect 676034 887703 676090 887712
rect 676048 887466 676076 887703
rect 676036 887460 676088 887466
rect 676036 887402 676088 887408
rect 676034 887360 676090 887369
rect 676034 887295 676090 887304
rect 676048 886038 676076 887295
rect 676036 886032 676088 886038
rect 676036 885974 676088 885980
rect 678978 885048 679034 885057
rect 678978 884983 678980 884992
rect 679032 884983 679034 884992
rect 678980 884954 679032 884960
rect 675392 883312 675444 883318
rect 675392 883254 675444 883260
rect 675208 880728 675260 880734
rect 675208 880670 675260 880676
rect 675208 880592 675260 880598
rect 675208 880534 675260 880540
rect 675116 878824 675168 878830
rect 675116 878766 675168 878772
rect 675128 874426 675156 878766
rect 675220 876262 675248 880534
rect 675300 880524 675352 880530
rect 675300 880466 675352 880472
rect 675312 877418 675340 880466
rect 675404 878084 675432 883254
rect 679084 878558 679112 888111
rect 679176 880598 679204 892599
rect 679438 891848 679494 891857
rect 679438 891783 679494 891792
rect 679254 891440 679310 891449
rect 679254 891375 679310 891384
rect 679164 880592 679216 880598
rect 679164 880534 679216 880540
rect 679268 878830 679296 891375
rect 679452 880530 679480 891783
rect 680266 890216 680322 890225
rect 680266 890151 680322 890160
rect 679714 889808 679770 889817
rect 679714 889743 679770 889752
rect 679530 889400 679586 889409
rect 679530 889335 679586 889344
rect 679440 880524 679492 880530
rect 679440 880466 679492 880472
rect 679256 878824 679308 878830
rect 679256 878766 679308 878772
rect 679544 878694 679572 889335
rect 679532 878688 679584 878694
rect 679532 878630 679584 878636
rect 679728 878626 679756 889743
rect 680280 880666 680308 890151
rect 680268 880660 680320 880666
rect 680268 880602 680320 880608
rect 679716 878620 679768 878626
rect 679716 878562 679768 878568
rect 679072 878552 679124 878558
rect 679072 878494 679124 878500
rect 675404 877418 675432 877540
rect 675312 877390 675432 877418
rect 675392 877260 675444 877266
rect 675392 877202 675444 877208
rect 675404 876860 675432 877202
rect 675220 876234 675418 876262
rect 675128 874398 675340 874426
rect 675116 874336 675168 874342
rect 675116 874278 675168 874284
rect 675312 874290 675340 874398
rect 675404 874290 675432 874412
rect 675128 873882 675156 874278
rect 675312 874262 675432 874290
rect 675128 873854 675340 873882
rect 675116 873792 675168 873798
rect 675116 873734 675168 873740
rect 675312 873746 675340 873854
rect 675404 873746 675432 873868
rect 675128 873202 675156 873734
rect 675312 873718 675432 873746
rect 675128 873174 675418 873202
rect 675024 872772 675076 872778
rect 675024 872714 675076 872720
rect 674944 872630 675156 872658
rect 675128 872590 675156 872630
rect 675024 872568 675076 872574
rect 675128 872562 675340 872590
rect 675024 872510 675076 872516
rect 675312 872522 675340 872562
rect 675404 872522 675432 872576
rect 674760 872358 674880 872386
rect 674656 869372 674708 869378
rect 674656 869314 674708 869320
rect 674472 867604 674524 867610
rect 674472 867546 674524 867552
rect 674760 865774 674788 872358
rect 674748 865768 674800 865774
rect 674748 865710 674800 865716
rect 675036 863342 675064 872510
rect 675208 872500 675260 872506
rect 675312 872494 675432 872522
rect 675208 872442 675260 872448
rect 675116 872228 675168 872234
rect 675116 872170 675168 872176
rect 675128 867694 675156 872170
rect 675220 870074 675248 872442
rect 675220 870046 675418 870074
rect 675208 869984 675260 869990
rect 675208 869926 675260 869932
rect 675220 869530 675248 869926
rect 675220 869502 675418 869530
rect 675208 869440 675260 869446
rect 675208 869382 675260 869388
rect 675220 868238 675248 869382
rect 675300 869372 675352 869378
rect 675300 869314 675352 869320
rect 675312 868889 675340 869314
rect 675312 868861 675418 868889
rect 675220 868210 675418 868238
rect 675128 867666 675418 867694
rect 675116 867604 675168 867610
rect 675116 867546 675168 867552
rect 675128 867049 675156 867546
rect 675128 867021 675418 867049
rect 675128 865830 675418 865858
rect 675128 863870 675156 865830
rect 675208 865768 675260 865774
rect 675208 865710 675260 865716
rect 675220 865209 675248 865710
rect 675220 865181 675418 865209
rect 675116 863864 675168 863870
rect 675116 863806 675168 863812
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675036 863314 675340 863342
rect 675404 863328 675432 863382
rect 675392 792192 675444 792198
rect 675392 792134 675444 792140
rect 675404 788868 675432 792134
rect 675114 788352 675170 788361
rect 675170 788310 675418 788338
rect 675114 788287 675170 788296
rect 675220 787665 675418 787693
rect 675220 787137 675248 787665
rect 675206 787128 675262 787137
rect 675206 787063 675262 787072
rect 675312 787018 675418 787046
rect 675312 786865 675340 787018
rect 675298 786856 675354 786865
rect 675298 786791 675354 786800
rect 675128 785182 675418 785210
rect 675128 784786 675156 785182
rect 673828 784780 673880 784786
rect 673828 784722 673880 784728
rect 675116 784780 675168 784786
rect 675116 784722 675168 784728
rect 673644 779816 673696 779822
rect 673644 779758 673696 779764
rect 673460 744252 673512 744258
rect 673460 744194 673512 744200
rect 673472 732494 673500 744194
rect 673552 744184 673604 744190
rect 673552 744126 673604 744132
rect 673460 732488 673512 732494
rect 673460 732430 673512 732436
rect 673460 732352 673512 732358
rect 673460 732294 673512 732300
rect 673472 728770 673500 732294
rect 673564 728890 673592 744126
rect 673552 728884 673604 728890
rect 673552 728826 673604 728832
rect 673472 728742 673592 728770
rect 673460 728612 673512 728618
rect 673460 728554 673512 728560
rect 673368 723172 673420 723178
rect 673368 723114 673420 723120
rect 673276 714944 673328 714950
rect 673276 714886 673328 714892
rect 673184 714060 673236 714066
rect 673184 714002 673236 714008
rect 673092 712428 673144 712434
rect 673092 712370 673144 712376
rect 672080 705152 672132 705158
rect 672080 705094 672132 705100
rect 671986 178800 672042 178809
rect 671986 178735 672042 178744
rect 672092 173641 672120 705094
rect 673104 680882 673132 712370
rect 673092 680876 673144 680882
rect 673092 680818 673144 680824
rect 673196 680814 673224 714002
rect 673288 681494 673316 714886
rect 673472 714610 673500 728554
rect 673460 714604 673512 714610
rect 673460 714546 673512 714552
rect 673368 713244 673420 713250
rect 673368 713186 673420 713192
rect 673276 681488 673328 681494
rect 673276 681430 673328 681436
rect 673184 680808 673236 680814
rect 673184 680750 673236 680756
rect 673380 668710 673408 713186
rect 673564 710734 673592 728742
rect 673552 710728 673604 710734
rect 673552 710670 673604 710676
rect 673656 708694 673684 779758
rect 673736 778796 673788 778802
rect 673736 778738 673788 778744
rect 673748 742801 673776 778738
rect 673734 742792 673790 742801
rect 673734 742727 673790 742736
rect 673736 738404 673788 738410
rect 673736 738346 673788 738352
rect 673748 728618 673776 738346
rect 673736 728612 673788 728618
rect 673736 728554 673788 728560
rect 673734 728512 673790 728521
rect 673734 728447 673790 728456
rect 673644 708688 673696 708694
rect 673644 708630 673696 708636
rect 673552 669044 673604 669050
rect 673552 668986 673604 668992
rect 673368 668704 673420 668710
rect 673368 668646 673420 668652
rect 672172 659728 672224 659734
rect 672172 659670 672224 659676
rect 672078 173632 672134 173641
rect 672078 173567 672134 173576
rect 672184 168609 672212 659670
rect 673460 646196 673512 646202
rect 673460 646138 673512 646144
rect 673184 644292 673236 644298
rect 673184 644234 673236 644240
rect 673196 637362 673224 644234
rect 673276 642252 673328 642258
rect 673276 642194 673328 642200
rect 673288 637430 673316 642194
rect 673472 640370 673500 646138
rect 673564 644298 673592 668986
rect 673748 662386 673776 728447
rect 673840 714678 673868 784722
rect 674760 784638 675418 784666
rect 674564 780496 674616 780502
rect 674564 780438 674616 780444
rect 674288 780020 674340 780026
rect 674288 779962 674340 779968
rect 674300 742665 674328 779962
rect 674472 778592 674524 778598
rect 674472 778534 674524 778540
rect 674286 742656 674342 742665
rect 674286 742591 674342 742600
rect 674288 734188 674340 734194
rect 674288 734130 674340 734136
rect 673828 714672 673880 714678
rect 673828 714614 673880 714620
rect 673828 689376 673880 689382
rect 673828 689318 673880 689324
rect 673736 662380 673788 662386
rect 673736 662322 673788 662328
rect 673736 645244 673788 645250
rect 673736 645186 673788 645192
rect 673644 644632 673696 644638
rect 673644 644574 673696 644580
rect 673552 644292 673604 644298
rect 673552 644234 673604 644240
rect 673552 644156 673604 644162
rect 673552 644098 673604 644104
rect 673380 640342 673500 640370
rect 673380 637498 673408 640342
rect 673458 640248 673514 640257
rect 673458 640183 673514 640192
rect 673368 637492 673420 637498
rect 673368 637434 673420 637440
rect 673276 637424 673328 637430
rect 673276 637366 673328 637372
rect 673184 637356 673236 637362
rect 673184 637298 673236 637304
rect 673368 623960 673420 623966
rect 673368 623902 673420 623908
rect 673276 621988 673328 621994
rect 673276 621930 673328 621936
rect 672264 614644 672316 614650
rect 672264 614586 672316 614592
rect 672170 168600 672226 168609
rect 672170 168535 672226 168544
rect 671988 167068 672040 167074
rect 671988 167010 672040 167016
rect 671896 131708 671948 131714
rect 671896 131650 671948 131656
rect 671804 130076 671856 130082
rect 671804 130018 671856 130024
rect 672000 114345 672028 167010
rect 672276 163577 672304 614586
rect 673184 597304 673236 597310
rect 673184 597246 673236 597252
rect 673196 593434 673224 597246
rect 673184 593428 673236 593434
rect 673184 593370 673236 593376
rect 673288 587994 673316 621930
rect 673276 587988 673328 587994
rect 673276 587930 673328 587936
rect 673380 587926 673408 623902
rect 673472 621382 673500 640183
rect 673564 637786 673592 644098
rect 673656 637922 673684 644574
rect 673748 638042 673776 645186
rect 673736 638036 673788 638042
rect 673736 637978 673788 637984
rect 673656 637894 673776 637922
rect 673564 637758 673684 637786
rect 673550 637664 673606 637673
rect 673550 637599 673606 637608
rect 673564 629377 673592 637599
rect 673550 629368 673606 629377
rect 673550 629303 673606 629312
rect 673460 621376 673512 621382
rect 673460 621318 673512 621324
rect 673552 599820 673604 599826
rect 673552 599762 673604 599768
rect 673460 598596 673512 598602
rect 673460 598538 673512 598544
rect 673368 587920 673420 587926
rect 673368 587862 673420 587868
rect 673472 583778 673500 598538
rect 673564 593570 673592 599762
rect 673552 593564 673604 593570
rect 673552 593506 673604 593512
rect 673552 593428 673604 593434
rect 673552 593370 673604 593376
rect 673460 583772 673512 583778
rect 673460 583714 673512 583720
rect 673564 582350 673592 593370
rect 673552 582344 673604 582350
rect 673552 582286 673604 582292
rect 673656 572830 673684 637758
rect 673748 609249 673776 637894
rect 673840 618186 673868 689318
rect 674300 663134 674328 734130
rect 674484 724810 674512 778534
rect 674472 724804 674524 724810
rect 674472 724746 674524 724752
rect 674470 724704 674526 724713
rect 674470 724639 674526 724648
rect 674484 721585 674512 724639
rect 674470 721576 674526 721585
rect 674470 721511 674526 721520
rect 674576 714746 674604 780438
rect 674656 777368 674708 777374
rect 674656 777310 674708 777316
rect 674668 767378 674696 777310
rect 674760 773362 674788 784638
rect 675312 784094 675432 784122
rect 675312 783986 675340 784094
rect 674944 783958 675340 783986
rect 675404 783972 675432 784094
rect 674944 776914 674972 783958
rect 675116 783896 675168 783902
rect 675116 783838 675168 783844
rect 675128 778478 675156 783838
rect 675220 783346 675418 783374
rect 675220 779822 675248 783346
rect 675496 780502 675524 780844
rect 675484 780496 675536 780502
rect 675484 780438 675536 780444
rect 675496 780026 675524 780300
rect 675484 780020 675536 780026
rect 675484 779962 675536 779968
rect 675208 779816 675260 779822
rect 675208 779758 675260 779764
rect 675220 779674 675418 779702
rect 675220 778598 675248 779674
rect 675496 778802 675524 779008
rect 675484 778796 675536 778802
rect 675484 778738 675536 778744
rect 675208 778592 675260 778598
rect 675208 778534 675260 778540
rect 675128 778450 675418 778478
rect 675404 777374 675432 777852
rect 675392 777368 675444 777374
rect 675392 777310 675444 777316
rect 674944 776898 675064 776914
rect 674944 776892 675076 776898
rect 674944 776886 675024 776892
rect 675024 776834 675076 776840
rect 675024 776688 675076 776694
rect 675024 776630 675076 776636
rect 675036 773430 675064 776630
rect 675128 776614 675418 776642
rect 675128 775538 675156 776614
rect 675220 776002 675340 776030
rect 675116 775532 675168 775538
rect 675116 775474 675168 775480
rect 675024 773424 675076 773430
rect 675024 773366 675076 773372
rect 674748 773356 674800 773362
rect 674748 773298 674800 773304
rect 675220 771610 675248 776002
rect 675312 775962 675340 776002
rect 675404 775962 675432 776016
rect 675312 775934 675432 775962
rect 675404 773650 675432 774180
rect 674852 771582 675248 771610
rect 675312 773622 675432 773650
rect 674656 767372 674708 767378
rect 674656 767314 674708 767320
rect 674656 757648 674708 757654
rect 674656 757590 674708 757596
rect 674668 738410 674696 757590
rect 674852 747974 674880 771582
rect 674932 767372 674984 767378
rect 674932 767314 674984 767320
rect 674760 747946 674880 747974
rect 674656 738404 674708 738410
rect 674656 738346 674708 738352
rect 674760 738290 674788 747946
rect 674668 738262 674788 738290
rect 674668 714814 674696 738262
rect 674748 735684 674800 735690
rect 674748 735626 674800 735632
rect 674656 714808 674708 714814
rect 674656 714750 674708 714756
rect 674564 714740 674616 714746
rect 674564 714682 674616 714688
rect 674656 710728 674708 710734
rect 674656 710670 674708 710676
rect 674564 687336 674616 687342
rect 674564 687278 674616 687284
rect 674470 681184 674526 681193
rect 674470 681119 674526 681128
rect 674484 674121 674512 681119
rect 674470 674112 674526 674121
rect 674470 674047 674526 674056
rect 674576 673962 674604 687278
rect 674484 673934 674604 673962
rect 674288 663128 674340 663134
rect 674288 663070 674340 663076
rect 674288 647896 674340 647902
rect 674288 647838 674340 647844
rect 674300 642258 674328 647838
rect 674288 642252 674340 642258
rect 674288 642194 674340 642200
rect 674288 642116 674340 642122
rect 674288 642058 674340 642064
rect 673828 618180 673880 618186
rect 673828 618122 673880 618128
rect 673734 609240 673790 609249
rect 673734 609175 673790 609184
rect 673736 609068 673788 609074
rect 673736 609010 673788 609016
rect 673748 593609 673776 609010
rect 673828 606960 673880 606966
rect 673828 606902 673880 606908
rect 673840 597310 673868 606902
rect 673828 597304 673880 597310
rect 673828 597246 673880 597252
rect 673828 597168 673880 597174
rect 673828 597110 673880 597116
rect 673734 593600 673790 593609
rect 673734 593535 673790 593544
rect 673736 593496 673788 593502
rect 673736 593438 673788 593444
rect 673644 572824 673696 572830
rect 673644 572766 673696 572772
rect 672356 568608 672408 568614
rect 672356 568550 672408 568556
rect 672262 163568 672318 163577
rect 672262 163503 672318 163512
rect 672368 158409 672396 568550
rect 673644 559564 673696 559570
rect 673644 559506 673696 559512
rect 673460 558272 673512 558278
rect 673460 558214 673512 558220
rect 673368 553580 673420 553586
rect 673368 553522 673420 553528
rect 673380 547210 673408 553522
rect 673472 547346 673500 558214
rect 673552 557524 673604 557530
rect 673552 557466 673604 557472
rect 673564 547482 673592 557466
rect 673656 553586 673684 559506
rect 673644 553580 673696 553586
rect 673644 553522 673696 553528
rect 673644 553444 673696 553450
rect 673644 553386 673696 553392
rect 673656 547618 673684 553386
rect 673748 547738 673776 593438
rect 673840 576706 673868 597110
rect 673828 576700 673880 576706
rect 673828 576642 673880 576648
rect 674300 573646 674328 642058
rect 674484 618254 674512 673934
rect 674564 673872 674616 673878
rect 674564 673814 674616 673820
rect 674472 618248 674524 618254
rect 674472 618190 674524 618196
rect 674576 618118 674604 673814
rect 674668 664766 674696 710670
rect 674760 667894 674788 735626
rect 674840 735004 674892 735010
rect 674840 734946 674892 734952
rect 674852 732018 674880 734946
rect 674840 732012 674892 732018
rect 674840 731954 674892 731960
rect 674840 731876 674892 731882
rect 674840 731818 674892 731824
rect 674852 728793 674880 731818
rect 674838 728784 674894 728793
rect 674838 728719 674894 728728
rect 674840 728680 674892 728686
rect 674944 728657 674972 767314
rect 675312 757654 675340 773622
rect 675668 773424 675720 773430
rect 675668 773366 675720 773372
rect 675300 757648 675352 757654
rect 675300 757590 675352 757596
rect 675392 747992 675444 747998
rect 675392 747934 675444 747940
rect 675404 743852 675432 747934
rect 675680 744190 675708 773366
rect 675760 773356 675812 773362
rect 675760 773298 675812 773304
rect 675772 744258 675800 773298
rect 675760 744252 675812 744258
rect 675760 744194 675812 744200
rect 675668 744184 675720 744190
rect 675668 744126 675720 744132
rect 675404 742937 675432 743308
rect 675390 742928 675446 742937
rect 675390 742863 675446 742872
rect 675680 742529 675708 742696
rect 675666 742520 675722 742529
rect 675666 742455 675722 742464
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 675128 742002 675340 742030
rect 675404 742016 675432 742070
rect 675128 740353 675156 742002
rect 675114 740344 675170 740353
rect 675114 740279 675170 740288
rect 675114 740208 675170 740217
rect 675170 740166 675418 740194
rect 675114 740143 675170 740152
rect 675114 739664 675170 739673
rect 675170 739622 675418 739650
rect 675114 739599 675170 739608
rect 675404 738721 675432 739024
rect 675390 738712 675446 738721
rect 675390 738647 675446 738656
rect 675772 738041 675800 738344
rect 675758 738032 675814 738041
rect 675758 737967 675814 737976
rect 675208 737044 675260 737050
rect 675208 736986 675260 736992
rect 675220 733666 675248 736986
rect 675300 736976 675352 736982
rect 675300 736918 675352 736924
rect 675312 733786 675340 736918
rect 675404 735690 675432 735896
rect 675392 735684 675444 735690
rect 675392 735626 675444 735632
rect 675404 735010 675432 735319
rect 675392 735004 675444 735010
rect 675392 734946 675444 734952
rect 675404 734194 675432 734672
rect 675392 734188 675444 734194
rect 675392 734130 675444 734136
rect 675404 733786 675432 734031
rect 675300 733780 675352 733786
rect 675300 733722 675352 733728
rect 675392 733780 675444 733786
rect 675392 733722 675444 733728
rect 675220 733638 675432 733666
rect 675404 733479 675432 733638
rect 675300 733440 675352 733446
rect 675300 733382 675352 733388
rect 675208 733372 675260 733378
rect 675208 733314 675260 733320
rect 675220 732154 675248 733314
rect 675208 732148 675260 732154
rect 675208 732090 675260 732096
rect 675312 732034 675340 733382
rect 675404 732358 675432 732836
rect 675392 732352 675444 732358
rect 675392 732294 675444 732300
rect 675208 732012 675260 732018
rect 675312 732006 675432 732034
rect 675208 731954 675260 731960
rect 675220 728906 675248 731954
rect 675404 731612 675432 732006
rect 675312 730986 675418 731014
rect 675312 729065 675340 730986
rect 675298 729056 675354 729065
rect 675298 728991 675354 729000
rect 675220 728878 675340 728906
rect 675208 728816 675260 728822
rect 675208 728758 675260 728764
rect 674840 728622 674892 728628
rect 674930 728648 674986 728657
rect 674852 709238 674880 728622
rect 674930 728583 674986 728592
rect 674932 728544 674984 728550
rect 674932 728486 674984 728492
rect 674840 709232 674892 709238
rect 674840 709174 674892 709180
rect 674944 701054 674972 728486
rect 675022 728376 675078 728385
rect 675022 728311 675078 728320
rect 675036 712026 675064 728311
rect 675116 724804 675168 724810
rect 675116 724746 675168 724752
rect 675128 712094 675156 724746
rect 675116 712088 675168 712094
rect 675116 712030 675168 712036
rect 675024 712020 675076 712026
rect 675024 711962 675076 711968
rect 675220 709306 675248 728758
rect 675312 728362 675340 728878
rect 675404 728686 675432 729164
rect 675392 728680 675444 728686
rect 675392 728622 675444 728628
rect 675312 728334 675432 728362
rect 675298 728240 675354 728249
rect 675298 728175 675354 728184
rect 675208 709300 675260 709306
rect 675208 709242 675260 709248
rect 674944 701026 675248 701054
rect 675024 692912 675076 692918
rect 675024 692854 675076 692860
rect 675036 688974 675064 692854
rect 675116 690056 675168 690062
rect 675116 689998 675168 690004
rect 675024 688968 675076 688974
rect 675024 688910 675076 688916
rect 675024 688628 675076 688634
rect 675024 688570 675076 688576
rect 675036 683754 675064 688570
rect 675128 687070 675156 689998
rect 675116 687064 675168 687070
rect 675116 687006 675168 687012
rect 675116 685500 675168 685506
rect 675116 685442 675168 685448
rect 674944 683726 675064 683754
rect 674944 673878 674972 683726
rect 675024 683664 675076 683670
rect 675024 683606 675076 683612
rect 674932 673872 674984 673878
rect 674932 673814 674984 673820
rect 674932 668024 674984 668030
rect 674932 667966 674984 667972
rect 674748 667888 674800 667894
rect 674748 667830 674800 667836
rect 674656 664760 674708 664766
rect 674656 664702 674708 664708
rect 674656 649596 674708 649602
rect 674656 649538 674708 649544
rect 674668 638178 674696 649538
rect 674748 648644 674800 648650
rect 674748 648586 674800 648592
rect 674760 643550 674788 648586
rect 674944 647902 674972 667966
rect 674932 647896 674984 647902
rect 674932 647838 674984 647844
rect 674932 647760 674984 647766
rect 674932 647702 674984 647708
rect 674748 643544 674800 643550
rect 674748 643486 674800 643492
rect 674748 643408 674800 643414
rect 674748 643350 674800 643356
rect 674760 639266 674788 643350
rect 674748 639260 674800 639266
rect 674748 639202 674800 639208
rect 674748 639124 674800 639130
rect 674748 639066 674800 639072
rect 674656 638172 674708 638178
rect 674656 638114 674708 638120
rect 674656 638036 674708 638042
rect 674656 637978 674708 637984
rect 674564 618112 674616 618118
rect 674564 618054 674616 618060
rect 674564 609136 674616 609142
rect 674564 609078 674616 609084
rect 674472 609000 674524 609006
rect 674472 608942 674524 608948
rect 674484 596358 674512 608942
rect 674576 598534 674604 609078
rect 674564 598528 674616 598534
rect 674564 598470 674616 598476
rect 674564 598392 674616 598398
rect 674564 598334 674616 598340
rect 674472 596352 674524 596358
rect 674472 596294 674524 596300
rect 674472 595332 674524 595338
rect 674472 595274 674524 595280
rect 674484 583914 674512 595274
rect 674472 583908 674524 583914
rect 674472 583850 674524 583856
rect 674472 583772 674524 583778
rect 674472 583714 674524 583720
rect 674288 573640 674340 573646
rect 674288 573582 674340 573588
rect 674288 568812 674340 568818
rect 674288 568754 674340 568760
rect 673828 554940 673880 554946
rect 673828 554882 673880 554888
rect 673840 547738 673868 554882
rect 674300 553897 674328 568754
rect 674286 553888 674342 553897
rect 674286 553823 674342 553832
rect 674288 553784 674340 553790
rect 674288 553726 674340 553732
rect 674300 547874 674328 553726
rect 674288 547868 674340 547874
rect 674288 547810 674340 547816
rect 673736 547732 673788 547738
rect 673736 547674 673788 547680
rect 673828 547732 673880 547738
rect 673828 547674 673880 547680
rect 674288 547732 674340 547738
rect 674288 547674 674340 547680
rect 673656 547590 673868 547618
rect 673736 547528 673788 547534
rect 673564 547454 673684 547482
rect 673736 547470 673788 547476
rect 673472 547318 673592 547346
rect 673380 547182 673500 547210
rect 673472 537130 673500 547182
rect 673460 537124 673512 537130
rect 673460 537066 673512 537072
rect 673564 537010 673592 547318
rect 673472 536982 673592 537010
rect 673472 536790 673500 536982
rect 673656 536874 673684 547454
rect 673564 536846 673684 536874
rect 673460 536784 673512 536790
rect 673460 536726 673512 536732
rect 673460 536648 673512 536654
rect 673460 536590 673512 536596
rect 672448 524476 672500 524482
rect 672448 524418 672500 524424
rect 672354 158400 672410 158409
rect 672354 158335 672410 158344
rect 672460 153377 672488 524418
rect 673472 488374 673500 536590
rect 673460 488368 673512 488374
rect 673460 488310 673512 488316
rect 673564 483478 673592 536846
rect 673644 536784 673696 536790
rect 673644 536726 673696 536732
rect 673656 485722 673684 536726
rect 673748 527066 673776 547470
rect 673736 527060 673788 527066
rect 673736 527002 673788 527008
rect 673644 485716 673696 485722
rect 673644 485658 673696 485664
rect 673552 483472 673604 483478
rect 673552 483414 673604 483420
rect 673840 483002 673868 547590
rect 674300 539510 674328 547674
rect 674288 539504 674340 539510
rect 674288 539446 674340 539452
rect 674288 537124 674340 537130
rect 674288 537066 674340 537072
rect 674300 488442 674328 537066
rect 674484 527134 674512 583714
rect 674576 527882 674604 598334
rect 674668 575278 674696 637978
rect 674760 576774 674788 639066
rect 674944 638246 674972 647702
rect 674840 638240 674892 638246
rect 674840 638182 674892 638188
rect 674932 638240 674984 638246
rect 674932 638182 674984 638188
rect 674852 637566 674880 638182
rect 674840 637560 674892 637566
rect 674840 637502 674892 637508
rect 675036 635474 675064 683606
rect 674852 635446 675064 635474
rect 675128 635458 675156 685442
rect 675220 665174 675248 701026
rect 675312 666505 675340 728175
rect 675404 720374 675432 728334
rect 679072 723240 679124 723246
rect 679072 723182 679124 723188
rect 678980 723172 679032 723178
rect 678980 723114 679032 723120
rect 675404 720346 675616 720374
rect 675392 703928 675444 703934
rect 675392 703870 675444 703876
rect 675404 698875 675432 703870
rect 675588 699689 675616 720346
rect 675942 716544 675998 716553
rect 675942 716479 675998 716488
rect 675850 716136 675906 716145
rect 675850 716071 675906 716080
rect 675864 715018 675892 716071
rect 675956 715290 675984 716479
rect 676034 715728 676090 715737
rect 676034 715663 676090 715672
rect 675944 715284 675996 715290
rect 675944 715226 675996 715232
rect 676048 715154 676076 715663
rect 676036 715148 676088 715154
rect 676036 715090 676088 715096
rect 675852 715012 675904 715018
rect 675852 714954 675904 714960
rect 676036 714944 676088 714950
rect 676034 714912 676036 714921
rect 676088 714912 676090 714921
rect 676034 714847 676090 714856
rect 676036 714808 676088 714814
rect 676036 714750 676088 714756
rect 675760 714740 675812 714746
rect 675760 714682 675812 714688
rect 675668 714672 675720 714678
rect 675668 714614 675720 714620
rect 675680 710841 675708 714614
rect 675666 710832 675722 710841
rect 675666 710767 675722 710776
rect 675772 710433 675800 714682
rect 675942 714096 675998 714105
rect 675942 714031 675944 714040
rect 675996 714031 675998 714040
rect 675944 714002 675996 714008
rect 675942 713280 675998 713289
rect 675942 713215 675944 713224
rect 675996 713215 675998 713224
rect 675944 713186 675996 713192
rect 675942 712464 675998 712473
rect 675942 712399 675944 712408
rect 675996 712399 675998 712408
rect 675944 712370 675996 712376
rect 675944 712088 675996 712094
rect 675944 712030 675996 712036
rect 675852 712020 675904 712026
rect 675852 711962 675904 711968
rect 675758 710424 675814 710433
rect 675758 710359 675814 710368
rect 675760 709232 675812 709238
rect 675758 709200 675760 709209
rect 675812 709200 675814 709209
rect 675758 709135 675814 709144
rect 675864 708393 675892 711962
rect 675850 708384 675906 708393
rect 675850 708319 675906 708328
rect 675956 707985 675984 712030
rect 676048 711657 676076 714750
rect 676128 714604 676180 714610
rect 676128 714546 676180 714552
rect 676034 711648 676090 711657
rect 676034 711583 676090 711592
rect 676034 710016 676090 710025
rect 676140 710002 676168 714546
rect 678992 714513 679020 723114
rect 678978 714504 679034 714513
rect 678978 714439 679034 714448
rect 679084 712881 679112 723182
rect 703694 717196 703722 717332
rect 704154 717196 704182 717332
rect 704614 717196 704642 717332
rect 705074 717196 705102 717332
rect 705534 717196 705562 717332
rect 705994 717196 706022 717332
rect 706454 717196 706482 717332
rect 706914 717196 706942 717332
rect 707374 717196 707402 717332
rect 707834 717196 707862 717332
rect 708294 717196 708322 717332
rect 708754 717196 708782 717332
rect 709214 717196 709242 717332
rect 679070 712872 679126 712881
rect 679070 712807 679126 712816
rect 676090 709974 676168 710002
rect 676034 709951 676090 709960
rect 676036 709300 676088 709306
rect 676036 709242 676088 709248
rect 676048 708801 676076 709242
rect 676034 708792 676090 708801
rect 676034 708727 676090 708736
rect 676036 708688 676088 708694
rect 676036 708630 676088 708636
rect 675942 707976 675998 707985
rect 675942 707911 675998 707920
rect 676048 707577 676076 708630
rect 676034 707568 676090 707577
rect 676034 707503 676090 707512
rect 676034 706344 676090 706353
rect 676034 706279 676090 706288
rect 676048 705158 676076 706279
rect 676036 705152 676088 705158
rect 676034 705120 676036 705129
rect 676088 705120 676090 705129
rect 676034 705055 676090 705064
rect 676048 705029 676076 705055
rect 675574 699680 675630 699689
rect 675574 699615 675630 699624
rect 675404 698193 675432 698323
rect 675390 698184 675446 698193
rect 675390 698119 675446 698128
rect 675772 697241 675800 697680
rect 675758 697232 675814 697241
rect 675758 697167 675814 697176
rect 675772 696697 675800 697035
rect 675758 696688 675814 696697
rect 675758 696623 675814 696632
rect 675772 694793 675800 695195
rect 675758 694784 675814 694793
rect 675758 694719 675814 694728
rect 675496 694385 675524 694620
rect 675482 694376 675538 694385
rect 675482 694311 675538 694320
rect 675772 693569 675800 694008
rect 675758 693560 675814 693569
rect 675758 693495 675814 693504
rect 675772 693025 675800 693328
rect 675758 693016 675814 693025
rect 675758 692951 675814 692960
rect 675404 690577 675432 690880
rect 675390 690568 675446 690577
rect 675390 690503 675446 690512
rect 675404 690169 675432 690336
rect 675390 690160 675446 690169
rect 675390 690095 675446 690104
rect 675496 689382 675524 689656
rect 675484 689376 675536 689382
rect 675484 689318 675536 689324
rect 675404 688634 675432 689044
rect 675484 688968 675536 688974
rect 675484 688910 675536 688916
rect 675392 688628 675444 688634
rect 675392 688570 675444 688576
rect 675496 688500 675524 688910
rect 675404 687342 675432 687820
rect 675392 687336 675444 687342
rect 675392 687278 675444 687284
rect 675484 687064 675536 687070
rect 675484 687006 675536 687012
rect 675496 686664 675524 687006
rect 675404 685506 675432 685984
rect 675392 685500 675444 685506
rect 675392 685442 675444 685448
rect 675404 683670 675432 684148
rect 675392 683664 675444 683670
rect 675392 683606 675444 683612
rect 679164 681488 679216 681494
rect 679164 681430 679216 681436
rect 679072 680808 679124 680814
rect 679072 680750 679124 680756
rect 675942 678464 675998 678473
rect 675942 678399 675998 678408
rect 675956 674801 675984 678399
rect 675942 674792 675998 674801
rect 675942 674727 675998 674736
rect 676218 671120 676274 671129
rect 676218 671055 676274 671064
rect 676034 670984 676090 670993
rect 676232 670954 676260 671055
rect 676034 670919 676090 670928
rect 676220 670948 676272 670954
rect 676048 670818 676076 670919
rect 676220 670890 676272 670896
rect 676036 670812 676088 670818
rect 676036 670754 676088 670760
rect 678978 670304 679034 670313
rect 678978 670239 679034 670248
rect 676034 669760 676090 669769
rect 676034 669695 676090 669704
rect 676048 669050 676076 669695
rect 676036 669044 676088 669050
rect 676036 668986 676088 668992
rect 676034 668944 676090 668953
rect 676034 668879 676090 668888
rect 675482 668128 675538 668137
rect 675482 668063 675538 668072
rect 675390 667312 675446 667321
rect 675390 667247 675446 667256
rect 675298 666496 675354 666505
rect 675298 666431 675354 666440
rect 675208 665168 675260 665174
rect 675208 665110 675260 665116
rect 675404 659274 675432 667247
rect 675220 659246 675432 659274
rect 675220 646202 675248 659246
rect 675496 659138 675524 668063
rect 676048 668030 676076 668879
rect 676220 668704 676272 668710
rect 676218 668672 676220 668681
rect 676272 668672 676274 668681
rect 676218 668607 676274 668616
rect 678992 668098 679020 670239
rect 679084 669497 679112 680750
rect 679176 670313 679204 681430
rect 679256 680876 679308 680882
rect 679256 680818 679308 680824
rect 679162 670304 679218 670313
rect 679162 670239 679218 670248
rect 679070 669488 679126 669497
rect 679070 669423 679126 669432
rect 678980 668092 679032 668098
rect 678980 668034 679032 668040
rect 676036 668024 676088 668030
rect 676036 667966 676088 667972
rect 676036 667888 676088 667894
rect 679268 667865 679296 680818
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 676036 667830 676088 667836
rect 679254 667856 679310 667865
rect 676048 665281 676076 667830
rect 679254 667791 679310 667800
rect 676034 665272 676090 665281
rect 676034 665207 676090 665216
rect 676036 665168 676088 665174
rect 676036 665110 676088 665116
rect 676048 664873 676076 665110
rect 676034 664864 676090 664873
rect 676034 664799 676090 664808
rect 676036 664760 676088 664766
rect 676036 664702 676088 664708
rect 676048 663241 676076 664702
rect 676034 663232 676090 663241
rect 676034 663167 676090 663176
rect 676036 663128 676088 663134
rect 676036 663070 676088 663076
rect 676048 662833 676076 663070
rect 676034 662824 676090 662833
rect 676034 662759 676090 662768
rect 676036 662380 676088 662386
rect 676036 662322 676088 662328
rect 676048 661609 676076 662322
rect 676034 661600 676090 661609
rect 676034 661535 676090 661544
rect 678978 660920 679034 660929
rect 678978 660855 679034 660864
rect 678992 660113 679020 660855
rect 678978 660104 679034 660113
rect 678978 660039 679034 660048
rect 678992 659734 679020 660039
rect 678980 659728 679032 659734
rect 678980 659670 679032 659676
rect 675312 659110 675524 659138
rect 675208 646196 675260 646202
rect 675208 646138 675260 646144
rect 675312 646082 675340 659110
rect 675392 656940 675444 656946
rect 675392 656882 675444 656888
rect 675404 653684 675432 656882
rect 675680 652633 675708 653140
rect 675666 652624 675722 652633
rect 675666 652559 675722 652568
rect 675496 652225 675524 652460
rect 675482 652216 675538 652225
rect 675482 652151 675538 652160
rect 675404 651681 675432 651848
rect 675390 651672 675446 651681
rect 675390 651607 675446 651616
rect 675404 649602 675432 650012
rect 675392 649596 675444 649602
rect 675392 649538 675444 649544
rect 675404 648961 675432 649468
rect 675390 648952 675446 648961
rect 675390 648887 675446 648896
rect 675404 648689 675432 648788
rect 675390 648680 675446 648689
rect 675390 648615 675446 648624
rect 675404 647766 675432 648176
rect 675392 647760 675444 647766
rect 675392 647702 675444 647708
rect 675220 646054 675340 646082
rect 675220 643958 675248 646054
rect 675300 645924 675352 645930
rect 675300 645866 675352 645872
rect 675208 643952 675260 643958
rect 675208 643894 675260 643900
rect 675312 643890 675340 645866
rect 675404 645250 675432 645660
rect 675392 645244 675444 645250
rect 675392 645186 675444 645192
rect 675404 644638 675432 645116
rect 675392 644632 675444 644638
rect 675392 644574 675444 644580
rect 675404 644162 675432 644475
rect 675392 644156 675444 644162
rect 675392 644098 675444 644104
rect 675300 643884 675352 643890
rect 675300 643826 675352 643832
rect 675404 643770 675432 643824
rect 675220 643742 675432 643770
rect 675220 639010 675248 643742
rect 675300 643476 675352 643482
rect 675300 643418 675352 643424
rect 675312 641458 675340 643418
rect 675392 643408 675444 643414
rect 675392 643350 675444 643356
rect 675404 643280 675432 643350
rect 675404 642122 675432 642635
rect 675392 642116 675444 642122
rect 675392 642058 675444 642064
rect 675312 641430 675418 641458
rect 675312 640781 675418 640809
rect 675312 639130 675340 640781
rect 675300 639124 675352 639130
rect 675300 639066 675352 639072
rect 675220 638982 675340 639010
rect 675312 638722 675340 638982
rect 675300 638716 675352 638722
rect 675300 638658 675352 638664
rect 675496 638602 675524 638928
rect 675220 638574 675524 638602
rect 675116 635452 675168 635458
rect 674852 620974 674880 635446
rect 675116 635394 675168 635400
rect 675220 635338 675248 638574
rect 675300 638444 675352 638450
rect 675300 638386 675352 638392
rect 674944 635310 675248 635338
rect 674840 620968 674892 620974
rect 674840 620910 674892 620916
rect 674840 576972 674892 576978
rect 674840 576914 674892 576920
rect 674748 576768 674800 576774
rect 674748 576710 674800 576716
rect 674656 575272 674708 575278
rect 674656 575214 674708 575220
rect 674852 574094 674880 576914
rect 674944 574870 674972 635310
rect 675116 635112 675168 635118
rect 675116 635054 675168 635060
rect 675128 623762 675156 635054
rect 675312 632054 675340 638386
rect 675576 638240 675628 638246
rect 675576 638182 675628 638188
rect 675758 638208 675814 638217
rect 675484 638172 675536 638178
rect 675484 638114 675536 638120
rect 675220 632026 675340 632054
rect 675116 623756 675168 623762
rect 675116 623698 675168 623704
rect 675220 617137 675248 632026
rect 675298 624744 675354 624753
rect 675298 624679 675354 624688
rect 675206 617128 675262 617137
rect 675206 617063 675262 617072
rect 675312 606966 675340 624679
rect 675496 609074 675524 638114
rect 675484 609068 675536 609074
rect 675484 609010 675536 609016
rect 675588 609006 675616 638182
rect 675758 638143 675814 638152
rect 675668 612876 675720 612882
rect 675668 612818 675720 612824
rect 675576 609000 675628 609006
rect 675576 608942 675628 608948
rect 675680 608668 675708 612818
rect 675772 609142 675800 638143
rect 679256 637560 679308 637566
rect 679256 637502 679308 637508
rect 679164 637424 679216 637430
rect 679164 637366 679216 637372
rect 679072 637356 679124 637362
rect 679072 637298 679124 637304
rect 678978 626104 679034 626113
rect 678978 626039 679034 626048
rect 676218 625696 676274 625705
rect 676218 625631 676274 625640
rect 676126 625288 676182 625297
rect 676126 625223 676182 625232
rect 676036 623960 676088 623966
rect 676034 623928 676036 623937
rect 676088 623928 676090 623937
rect 676140 623898 676168 625223
rect 676232 624170 676260 625631
rect 676220 624164 676272 624170
rect 676220 624106 676272 624112
rect 678992 624034 679020 626039
rect 679084 625297 679112 637298
rect 679070 625288 679126 625297
rect 679070 625223 679126 625232
rect 679176 624481 679204 637366
rect 679162 624472 679218 624481
rect 679162 624407 679218 624416
rect 678980 624028 679032 624034
rect 678980 623970 679032 623976
rect 676034 623863 676090 623872
rect 676128 623892 676180 623898
rect 676128 623834 676180 623840
rect 676036 623756 676088 623762
rect 676036 623698 676088 623704
rect 676048 621489 676076 623698
rect 679268 623665 679296 637502
rect 679348 637492 679400 637498
rect 679348 637434 679400 637440
rect 679254 623656 679310 623665
rect 679254 623591 679310 623600
rect 679360 622849 679388 637434
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 679346 622840 679402 622849
rect 679346 622775 679402 622784
rect 676218 622024 676274 622033
rect 676218 621959 676220 621968
rect 676272 621959 676274 621968
rect 676220 621930 676272 621936
rect 676034 621480 676090 621489
rect 676034 621415 676090 621424
rect 676036 621376 676088 621382
rect 676036 621318 676088 621324
rect 676048 621081 676076 621318
rect 676034 621072 676090 621081
rect 676034 621007 676090 621016
rect 676036 620968 676088 620974
rect 676036 620910 676088 620916
rect 676048 619857 676076 620910
rect 676034 619848 676090 619857
rect 676034 619783 676090 619792
rect 676036 618248 676088 618254
rect 676034 618216 676036 618225
rect 676088 618216 676090 618225
rect 676034 618151 676090 618160
rect 676128 618180 676180 618186
rect 676128 618122 676180 618128
rect 676036 618112 676088 618118
rect 676036 618054 676088 618060
rect 676048 616593 676076 618054
rect 676140 617953 676168 618122
rect 676126 617944 676182 617953
rect 676126 617879 676182 617888
rect 676034 616584 676090 616593
rect 676034 616519 676090 616528
rect 678978 615904 679034 615913
rect 678978 615839 679034 615848
rect 678992 615097 679020 615839
rect 678978 615088 679034 615097
rect 678978 615023 679034 615032
rect 678992 614650 679020 615023
rect 678980 614644 679032 614650
rect 678980 614586 679032 614592
rect 675760 609136 675812 609142
rect 675760 609078 675812 609084
rect 675404 607889 675432 608124
rect 675390 607880 675446 607889
rect 675390 607815 675446 607824
rect 675772 607345 675800 607479
rect 675758 607336 675814 607345
rect 675758 607271 675814 607280
rect 675300 606960 675352 606966
rect 675300 606902 675352 606908
rect 675128 606818 675418 606846
rect 675128 604489 675156 606818
rect 675206 605024 675262 605033
rect 675262 604982 675418 605010
rect 675206 604959 675262 604968
rect 675114 604480 675170 604489
rect 675114 604415 675170 604424
rect 675298 604480 675354 604489
rect 675354 604438 675418 604466
rect 675298 604415 675354 604424
rect 675312 603894 675432 603922
rect 675114 603800 675170 603809
rect 675312 603786 675340 603894
rect 675170 603758 675340 603786
rect 675404 603772 675432 603894
rect 675114 603735 675170 603744
rect 675128 603146 675418 603174
rect 675128 601905 675156 603146
rect 675114 601896 675170 601905
rect 675114 601831 675170 601840
rect 675116 601792 675168 601798
rect 675116 601734 675168 601740
rect 675024 601724 675076 601730
rect 675024 601666 675076 601672
rect 675036 598126 675064 601666
rect 675128 598738 675156 601734
rect 675312 600766 675432 600794
rect 675312 600658 675340 600766
rect 675220 600630 675340 600658
rect 675404 600644 675432 600766
rect 675116 598732 675168 598738
rect 675116 598674 675168 598680
rect 675116 598528 675168 598534
rect 675116 598470 675168 598476
rect 675024 598120 675076 598126
rect 675024 598062 675076 598068
rect 675128 597106 675156 598470
rect 675116 597100 675168 597106
rect 675116 597042 675168 597048
rect 675220 596986 675248 600630
rect 675496 599826 675524 600100
rect 675484 599820 675536 599826
rect 675484 599762 675536 599768
rect 675312 599474 675418 599502
rect 675312 598398 675340 599474
rect 675392 598732 675444 598738
rect 675392 598674 675444 598680
rect 675300 598392 675352 598398
rect 675300 598334 675352 598340
rect 675404 598264 675432 598674
rect 675496 598602 675524 598808
rect 675484 598596 675536 598602
rect 675484 598538 675536 598544
rect 675300 598120 675352 598126
rect 675300 598062 675352 598068
rect 675036 596958 675248 596986
rect 674932 574864 674984 574870
rect 674932 574806 674984 574812
rect 674760 574066 674880 574094
rect 674760 565814 674788 574066
rect 674760 565786 674972 565814
rect 674748 557592 674800 557598
rect 674748 557534 674800 557540
rect 674656 555076 674708 555082
rect 674656 555018 674708 555024
rect 674668 548010 674696 555018
rect 674760 553518 674788 557534
rect 674748 553512 674800 553518
rect 674748 553454 674800 553460
rect 674748 551948 674800 551954
rect 674748 551890 674800 551896
rect 674656 548004 674708 548010
rect 674656 547946 674708 547952
rect 674656 547868 674708 547874
rect 674656 547810 674708 547816
rect 674564 527876 674616 527882
rect 674564 527818 674616 527824
rect 674472 527128 674524 527134
rect 674472 527070 674524 527076
rect 674288 488436 674340 488442
rect 674288 488378 674340 488384
rect 674668 483886 674696 547810
rect 674760 485518 674788 551890
rect 674840 548004 674892 548010
rect 674840 547946 674892 547952
rect 674852 536874 674880 547946
rect 674944 543794 674972 565786
rect 674932 543788 674984 543794
rect 674932 543730 674984 543736
rect 674852 536846 674972 536874
rect 674840 536784 674892 536790
rect 674840 536726 674892 536732
rect 674852 485790 674880 536726
rect 674944 488510 674972 536846
rect 675036 532710 675064 596958
rect 675208 596896 675260 596902
rect 675208 596838 675260 596844
rect 675220 593314 675248 596838
rect 675312 596442 675340 598062
rect 675404 597174 675432 597652
rect 675392 597168 675444 597174
rect 675392 597110 675444 597116
rect 675312 596414 675418 596442
rect 675300 596352 675352 596358
rect 675300 596294 675352 596300
rect 675128 593286 675248 593314
rect 675128 576842 675156 593286
rect 675208 593224 675260 593230
rect 675208 593166 675260 593172
rect 675116 576836 675168 576842
rect 675116 576778 675168 576784
rect 675116 576700 675168 576706
rect 675116 576642 675168 576648
rect 675024 532704 675076 532710
rect 675024 532646 675076 532652
rect 675128 529514 675156 576642
rect 675220 529922 675248 593166
rect 675312 583794 675340 596294
rect 675404 595338 675432 595816
rect 675392 595332 675444 595338
rect 675392 595274 675444 595280
rect 675680 593434 675708 593980
rect 675668 593428 675720 593434
rect 675668 593370 675720 593376
rect 675574 593192 675630 593201
rect 675574 593127 675630 593136
rect 675312 583766 675524 583794
rect 675392 583704 675444 583710
rect 675392 583646 675444 583652
rect 675404 568818 675432 583646
rect 675496 572121 675524 583766
rect 675588 575385 675616 593127
rect 679072 587988 679124 587994
rect 679072 587930 679124 587936
rect 678980 587920 679032 587926
rect 678980 587862 679032 587868
rect 676034 587752 676090 587761
rect 676034 587687 676090 587696
rect 676048 586265 676076 587687
rect 676034 586256 676090 586265
rect 676034 586191 676090 586200
rect 676036 582344 676088 582350
rect 676036 582286 676088 582292
rect 676048 579873 676076 582286
rect 676126 580952 676182 580961
rect 676126 580887 676182 580896
rect 676140 579970 676168 580887
rect 676310 580544 676366 580553
rect 676310 580479 676366 580488
rect 676218 580136 676274 580145
rect 676218 580071 676220 580080
rect 676272 580071 676274 580080
rect 676220 580042 676272 580048
rect 676128 579964 676180 579970
rect 676128 579906 676180 579912
rect 676034 579864 676090 579873
rect 676324 579834 676352 580479
rect 676034 579799 676090 579808
rect 676312 579828 676364 579834
rect 676312 579770 676364 579776
rect 678992 579329 679020 587862
rect 678978 579320 679034 579329
rect 678978 579255 679034 579264
rect 676034 578640 676090 578649
rect 676034 578575 676090 578584
rect 676048 576978 676076 578575
rect 679084 577697 679112 587930
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 679070 577688 679126 577697
rect 679070 577623 679126 577632
rect 676036 576972 676088 576978
rect 676036 576914 676088 576920
rect 676036 576836 676088 576842
rect 676036 576778 676088 576784
rect 675944 576768 675996 576774
rect 675944 576710 675996 576716
rect 675956 576201 675984 576710
rect 675942 576192 675998 576201
rect 675942 576127 675998 576136
rect 676048 575793 676076 576778
rect 676034 575784 676090 575793
rect 676034 575719 676090 575728
rect 675574 575376 675630 575385
rect 675574 575311 675630 575320
rect 676036 575272 676088 575278
rect 676036 575214 676088 575220
rect 676048 574977 676076 575214
rect 676034 574968 676090 574977
rect 676034 574903 676090 574912
rect 676036 574864 676088 574870
rect 676036 574806 676088 574812
rect 676048 574569 676076 574806
rect 676034 574560 676090 574569
rect 676034 574495 676090 574504
rect 676036 573640 676088 573646
rect 676036 573582 676088 573588
rect 676048 572937 676076 573582
rect 676034 572928 676090 572937
rect 676034 572863 676090 572872
rect 676036 572824 676088 572830
rect 676036 572766 676088 572772
rect 676048 572529 676076 572766
rect 676034 572520 676090 572529
rect 676034 572455 676090 572464
rect 675482 572112 675538 572121
rect 675482 572047 675538 572056
rect 678978 570752 679034 570761
rect 678978 570687 679034 570696
rect 678992 569945 679020 570687
rect 678978 569936 679034 569945
rect 678978 569871 679034 569880
rect 675392 568812 675444 568818
rect 675392 568754 675444 568760
rect 675392 568676 675444 568682
rect 675392 568618 675444 568624
rect 675404 563448 675432 568618
rect 678992 568614 679020 569871
rect 678980 568608 679032 568614
rect 678980 568550 679032 568556
rect 675496 562465 675524 562904
rect 675482 562456 675538 562465
rect 675482 562391 675538 562400
rect 675298 562320 675354 562329
rect 675354 562278 675418 562306
rect 675298 562255 675354 562264
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675496 559570 675524 559776
rect 675484 559564 675536 559570
rect 675484 559506 675536 559512
rect 675312 559218 675418 559246
rect 675312 557569 675340 559218
rect 675404 558278 675432 558620
rect 675392 558272 675444 558278
rect 675392 558214 675444 558220
rect 675298 557560 675354 557569
rect 675404 557530 675432 557940
rect 675298 557495 675354 557504
rect 675392 557524 675444 557530
rect 675392 557466 675444 557472
rect 675404 555082 675432 555492
rect 675392 555076 675444 555082
rect 675392 555018 675444 555024
rect 675300 554940 675352 554946
rect 675352 554905 675418 554933
rect 675300 554882 675352 554888
rect 675300 554804 675352 554810
rect 675300 554746 675352 554752
rect 675312 551253 675340 554746
rect 675404 553790 675432 554268
rect 675392 553784 675444 553790
rect 675392 553726 675444 553732
rect 675392 553512 675444 553518
rect 675392 553454 675444 553460
rect 675404 553079 675432 553454
rect 675496 553450 675524 553656
rect 675484 553444 675536 553450
rect 675484 553386 675536 553392
rect 675404 551954 675432 552432
rect 675392 551948 675444 551954
rect 675392 551890 675444 551896
rect 675312 551225 675418 551253
rect 675312 550582 675418 550610
rect 675312 548026 675340 550582
rect 675680 548282 675708 548760
rect 675668 548276 675720 548282
rect 675668 548218 675720 548224
rect 675482 548040 675538 548049
rect 675312 547998 675432 548026
rect 675300 547936 675352 547942
rect 675300 547878 675352 547884
rect 675312 536790 675340 547878
rect 675300 536784 675352 536790
rect 675300 536726 675352 536732
rect 675404 536654 675432 547998
rect 675482 547975 675538 547984
rect 675392 536648 675444 536654
rect 675392 536590 675444 536596
rect 675496 531321 675524 547975
rect 679254 544096 679310 544105
rect 679254 544031 679310 544040
rect 679070 543960 679126 543969
rect 679070 543895 679126 543904
rect 678978 543824 679034 543833
rect 678978 543759 679034 543768
rect 676126 542736 676182 542745
rect 676126 542671 676182 542680
rect 676140 541249 676168 542671
rect 676126 541240 676182 541249
rect 676126 541175 676182 541184
rect 675576 539504 675628 539510
rect 675576 539446 675628 539452
rect 675482 531312 675538 531321
rect 675482 531247 675538 531256
rect 675208 529916 675260 529922
rect 675208 529858 675260 529864
rect 675116 529508 675168 529514
rect 675116 529450 675168 529456
rect 675390 488880 675446 488889
rect 675390 488815 675446 488824
rect 674932 488504 674984 488510
rect 674932 488446 674984 488452
rect 674840 485784 674892 485790
rect 674840 485726 674892 485732
rect 674748 485512 674800 485518
rect 674748 485454 674800 485460
rect 674656 483880 674708 483886
rect 674656 483822 674708 483828
rect 673828 482996 673880 483002
rect 673828 482938 673880 482944
rect 672540 480752 672592 480758
rect 672540 480694 672592 480700
rect 672446 153368 672502 153377
rect 672446 153303 672502 153312
rect 672552 148209 672580 480694
rect 675404 477578 675432 488815
rect 675484 488368 675536 488374
rect 675484 488310 675536 488316
rect 675496 487257 675524 488310
rect 675482 487248 675538 487257
rect 675482 487183 675538 487192
rect 675588 482769 675616 539446
rect 676218 535936 676274 535945
rect 676218 535871 676274 535880
rect 676036 535764 676088 535770
rect 676034 535732 676036 535741
rect 676088 535732 676090 535741
rect 676034 535667 676090 535676
rect 676232 535634 676260 535871
rect 676220 535628 676272 535634
rect 676220 535570 676272 535576
rect 678992 535129 679020 543759
rect 678978 535120 679034 535129
rect 678978 535055 679034 535064
rect 676036 532704 676088 532710
rect 679084 532681 679112 543895
rect 679162 535120 679218 535129
rect 679162 535055 679218 535064
rect 679176 532914 679204 535055
rect 679268 533497 679296 544031
rect 679348 543788 679400 543794
rect 679348 543730 679400 543736
rect 679360 534313 679388 543730
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 679346 534304 679402 534313
rect 679346 534239 679402 534248
rect 679530 534304 679586 534313
rect 679530 534239 679586 534248
rect 679254 533488 679310 533497
rect 679438 533488 679494 533497
rect 679254 533423 679310 533432
rect 679360 533446 679438 533474
rect 679164 532908 679216 532914
rect 679164 532850 679216 532856
rect 676036 532646 676088 532652
rect 679070 532672 679126 532681
rect 676048 530029 676076 532646
rect 679254 532672 679310 532681
rect 679070 532607 679126 532616
rect 679176 532630 679254 532658
rect 678978 531856 679034 531865
rect 678978 531791 679034 531800
rect 676034 530020 676090 530029
rect 676034 529955 676090 529964
rect 676036 529916 676088 529922
rect 676036 529858 676088 529864
rect 676048 529621 676076 529858
rect 676034 529612 676090 529621
rect 676034 529547 676090 529556
rect 676036 529508 676088 529514
rect 676036 529450 676088 529456
rect 676048 527989 676076 529450
rect 676034 527980 676090 527989
rect 676034 527915 676090 527924
rect 676036 527876 676088 527882
rect 676036 527818 676088 527824
rect 676048 527581 676076 527818
rect 676034 527572 676090 527581
rect 676034 527507 676090 527516
rect 676036 527128 676088 527134
rect 676036 527070 676088 527076
rect 675944 527060 675996 527066
rect 675944 527002 675996 527008
rect 675956 526765 675984 527002
rect 675942 526756 675998 526765
rect 675942 526691 675998 526700
rect 676048 526357 676076 527070
rect 676034 526348 676090 526357
rect 676034 526283 676090 526292
rect 678992 521626 679020 531791
rect 679070 525736 679126 525745
rect 679070 525671 679126 525680
rect 679084 524929 679112 525671
rect 679070 524920 679126 524929
rect 679070 524855 679126 524864
rect 679084 524482 679112 524855
rect 679072 524476 679124 524482
rect 679072 524418 679124 524424
rect 676128 521620 676180 521626
rect 676128 521562 676180 521568
rect 678980 521620 679032 521626
rect 678980 521562 679032 521568
rect 676034 492144 676090 492153
rect 676034 492079 676090 492088
rect 675942 491736 675998 491745
rect 676048 491706 676076 492079
rect 675942 491671 675998 491680
rect 676036 491700 676088 491706
rect 675956 491434 675984 491671
rect 676036 491642 676088 491648
rect 676036 491564 676088 491570
rect 676036 491506 676088 491512
rect 675944 491428 675996 491434
rect 675944 491370 675996 491376
rect 676048 491337 676076 491506
rect 676034 491328 676090 491337
rect 676034 491263 676090 491272
rect 676140 491178 676168 521562
rect 679176 521558 679204 532630
rect 679254 532607 679310 532616
rect 679360 530414 679388 533446
rect 679438 533423 679494 533432
rect 679268 530386 679388 530414
rect 677396 521552 677448 521558
rect 677396 521494 677448 521500
rect 679164 521552 679216 521558
rect 679164 521494 679216 521500
rect 677304 521484 677356 521490
rect 677304 521426 677356 521432
rect 677316 491298 677344 521426
rect 676220 491292 676272 491298
rect 676220 491234 676272 491240
rect 677304 491292 677356 491298
rect 677304 491234 677356 491240
rect 675956 491150 676168 491178
rect 675758 490512 675814 490521
rect 675758 490447 675814 490456
rect 675772 484106 675800 490447
rect 675956 488481 675984 491150
rect 676034 490920 676090 490929
rect 676232 490906 676260 491234
rect 676090 490878 676260 490906
rect 676034 490855 676090 490864
rect 676220 490816 676272 490822
rect 676220 490758 676272 490764
rect 676034 490104 676090 490113
rect 676232 490090 676260 490758
rect 676090 490062 676260 490090
rect 676034 490039 676090 490048
rect 677408 490006 677436 521494
rect 679268 521422 679296 530386
rect 679544 527174 679572 534239
rect 679360 527146 679572 527174
rect 679360 521490 679388 527146
rect 679348 521484 679400 521490
rect 679348 521426 679400 521432
rect 677488 521416 677540 521422
rect 677488 521358 677540 521364
rect 679256 521416 679308 521422
rect 679256 521358 679308 521364
rect 677500 490822 677528 521358
rect 703694 492796 703722 492932
rect 704154 492796 704182 492932
rect 704614 492796 704642 492932
rect 705074 492796 705102 492932
rect 705534 492796 705562 492932
rect 705994 492796 706022 492932
rect 706454 492796 706482 492932
rect 706914 492796 706942 492932
rect 707374 492796 707402 492932
rect 707834 492796 707862 492932
rect 708294 492796 708322 492932
rect 708754 492796 708782 492932
rect 709214 492796 709242 492932
rect 677488 490816 677540 490822
rect 677488 490758 677540 490764
rect 676220 490000 676272 490006
rect 676220 489942 676272 489948
rect 677396 490000 677448 490006
rect 677396 489942 677448 489948
rect 676034 489696 676090 489705
rect 676034 489631 676090 489640
rect 676048 489394 676076 489631
rect 676036 489388 676088 489394
rect 676036 489330 676088 489336
rect 676034 489288 676090 489297
rect 676232 489274 676260 489942
rect 676090 489246 676260 489274
rect 676034 489223 676090 489232
rect 676128 489184 676180 489190
rect 676128 489126 676180 489132
rect 676036 488504 676088 488510
rect 675942 488472 675998 488481
rect 675852 488436 675904 488442
rect 676036 488446 676088 488452
rect 675942 488407 675998 488416
rect 675852 488378 675904 488384
rect 675864 486441 675892 488378
rect 675942 488064 675998 488073
rect 675942 487999 675998 488008
rect 675850 486432 675906 486441
rect 675850 486367 675906 486376
rect 675852 485716 675904 485722
rect 675852 485658 675904 485664
rect 675864 484401 675892 485658
rect 675850 484392 675906 484401
rect 675850 484327 675906 484336
rect 675772 484078 675892 484106
rect 675574 482760 675630 482769
rect 675574 482695 675630 482704
rect 675404 477550 675800 477578
rect 675772 402506 675800 477550
rect 675864 402665 675892 484078
rect 675850 402656 675906 402665
rect 675850 402591 675906 402600
rect 675772 402478 675892 402506
rect 675298 402248 675354 402257
rect 675298 402183 675354 402192
rect 674288 399492 674340 399498
rect 674288 399434 674340 399440
rect 673644 397588 673696 397594
rect 673644 397530 673696 397536
rect 673460 395412 673512 395418
rect 673460 395354 673512 395360
rect 672632 392080 672684 392086
rect 672632 392022 672684 392028
rect 672538 148200 672594 148209
rect 672538 148135 672594 148144
rect 672644 143177 672672 392022
rect 673472 375766 673500 395354
rect 673552 394936 673604 394942
rect 673552 394878 673604 394884
rect 673564 377466 673592 394878
rect 673656 381070 673684 397530
rect 673736 394188 673788 394194
rect 673736 394130 673788 394136
rect 673644 381064 673696 381070
rect 673644 381006 673696 381012
rect 673644 380928 673696 380934
rect 673644 380870 673696 380876
rect 673656 378826 673684 380870
rect 673644 378820 673696 378826
rect 673644 378762 673696 378768
rect 673748 378010 673776 394130
rect 673828 392012 673880 392018
rect 673828 391954 673880 391960
rect 673736 378004 673788 378010
rect 673736 377946 673788 377952
rect 673552 377460 673604 377466
rect 673552 377402 673604 377408
rect 673840 376990 673868 391954
rect 674300 385014 674328 399434
rect 674564 398268 674616 398274
rect 674564 398210 674616 398216
rect 674472 397044 674524 397050
rect 674472 396986 674524 396992
rect 674288 385008 674340 385014
rect 674288 384950 674340 384956
rect 674288 384872 674340 384878
rect 674288 384814 674340 384820
rect 674300 380934 674328 384814
rect 674484 381018 674512 396986
rect 674576 384810 674604 398210
rect 675024 397656 675076 397662
rect 675024 397598 675076 397604
rect 674656 397520 674708 397526
rect 674656 397462 674708 397468
rect 674564 384804 674616 384810
rect 674564 384746 674616 384752
rect 674668 383178 674696 397462
rect 674748 395004 674800 395010
rect 674748 394946 674800 394952
rect 674656 383172 674708 383178
rect 674656 383114 674708 383120
rect 674760 381954 674788 394946
rect 674840 394868 674892 394874
rect 674840 394810 674892 394816
rect 674852 382498 674880 394810
rect 674932 390584 674984 390590
rect 674932 390526 674984 390532
rect 674840 382492 674892 382498
rect 674840 382434 674892 382440
rect 674748 381948 674800 381954
rect 674748 381890 674800 381896
rect 674944 381138 674972 390526
rect 675036 386170 675064 397598
rect 675116 394800 675168 394806
rect 675116 394742 675168 394748
rect 675024 386164 675076 386170
rect 675024 386106 675076 386112
rect 675024 386028 675076 386034
rect 675024 385970 675076 385976
rect 674932 381132 674984 381138
rect 674932 381074 674984 381080
rect 674484 380990 674972 381018
rect 674288 380928 674340 380934
rect 674288 380870 674340 380876
rect 674472 380928 674524 380934
rect 674472 380870 674524 380876
rect 673828 376984 673880 376990
rect 673828 376926 673880 376932
rect 673460 375760 673512 375766
rect 673460 375702 673512 375708
rect 674484 373930 674512 380870
rect 674944 379250 674972 380990
rect 674668 379222 674972 379250
rect 674472 373924 674524 373930
rect 674472 373866 674524 373872
rect 674668 372094 674696 379222
rect 675036 372570 675064 385970
rect 675128 381274 675156 394742
rect 675208 394732 675260 394738
rect 675208 394674 675260 394680
rect 675220 385626 675248 394674
rect 675208 385620 675260 385626
rect 675208 385562 675260 385568
rect 675208 385008 675260 385014
rect 675208 384950 675260 384956
rect 675116 381268 675168 381274
rect 675116 381210 675168 381216
rect 675116 381132 675168 381138
rect 675116 381074 675168 381080
rect 675024 372564 675076 372570
rect 675024 372506 675076 372512
rect 674656 372088 674708 372094
rect 674656 372030 674708 372036
rect 675128 370734 675156 381074
rect 675220 370802 675248 384950
rect 675208 370796 675260 370802
rect 675208 370738 675260 370744
rect 675116 370728 675168 370734
rect 675116 370670 675168 370676
rect 675312 357513 675340 402183
rect 675758 401432 675814 401441
rect 675758 401367 675814 401376
rect 675666 395720 675722 395729
rect 675666 395655 675722 395664
rect 675680 395418 675708 395655
rect 675668 395412 675720 395418
rect 675668 395354 675720 395360
rect 675666 395312 675722 395321
rect 675666 395247 675722 395256
rect 675680 394942 675708 395247
rect 675668 394936 675720 394942
rect 675668 394878 675720 394884
rect 675772 390590 675800 401367
rect 675864 401033 675892 402478
rect 675850 401024 675906 401033
rect 675850 400959 675906 400968
rect 675956 400217 675984 487999
rect 676048 486033 676076 488446
rect 676034 486024 676090 486033
rect 676034 485959 676090 485968
rect 676036 485784 676088 485790
rect 676036 485726 676088 485732
rect 676048 485625 676076 485726
rect 676034 485616 676090 485625
rect 676034 485551 676090 485560
rect 676036 485512 676088 485518
rect 676036 485454 676088 485460
rect 676048 483993 676076 485454
rect 676034 483984 676090 483993
rect 676034 483919 676090 483928
rect 676036 483880 676088 483886
rect 676036 483822 676088 483828
rect 676048 483585 676076 483822
rect 676034 483576 676090 483585
rect 676034 483511 676090 483520
rect 676036 483472 676088 483478
rect 676036 483414 676088 483420
rect 676048 483177 676076 483414
rect 676034 483168 676090 483177
rect 676034 483103 676090 483112
rect 676036 482996 676088 483002
rect 676036 482938 676088 482944
rect 676048 482361 676076 482938
rect 676034 482352 676090 482361
rect 676034 482287 676090 482296
rect 676034 481944 676090 481953
rect 676034 481879 676090 481888
rect 676048 480758 676076 481879
rect 676036 480752 676088 480758
rect 676034 480720 676036 480729
rect 676088 480720 676090 480729
rect 676034 480655 676090 480664
rect 676048 480629 676076 480655
rect 676140 477494 676168 489126
rect 676048 477466 676168 477494
rect 676048 401849 676076 477466
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 676126 403744 676182 403753
rect 676126 403679 676182 403688
rect 676140 403170 676168 403679
rect 676218 403336 676274 403345
rect 676218 403271 676274 403280
rect 676128 403164 676180 403170
rect 676128 403106 676180 403112
rect 676232 403102 676260 403271
rect 676220 403096 676272 403102
rect 676220 403038 676272 403044
rect 676128 403028 676180 403034
rect 676128 402970 676180 402976
rect 676140 402937 676168 402970
rect 676126 402928 676182 402937
rect 676126 402863 676182 402872
rect 676034 401840 676090 401849
rect 676034 401775 676090 401784
rect 675942 400208 675998 400217
rect 675942 400143 675998 400152
rect 676034 399800 676090 399809
rect 676034 399735 676090 399744
rect 676048 399498 676076 399735
rect 676036 399492 676088 399498
rect 676036 399434 676088 399440
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675850 398576 675906 398585
rect 675850 398511 675906 398520
rect 675760 390584 675812 390590
rect 675760 390526 675812 390532
rect 675864 390402 675892 398511
rect 676048 398274 676076 399327
rect 676126 398848 676182 398857
rect 676126 398783 676182 398792
rect 676036 398268 676088 398274
rect 676036 398210 676088 398216
rect 676034 398168 676090 398177
rect 676034 398103 676090 398112
rect 675942 397760 675998 397769
rect 675942 397695 675998 397704
rect 675956 397662 675984 397695
rect 675944 397656 675996 397662
rect 675944 397598 675996 397604
rect 676048 397526 676076 398103
rect 676140 397594 676168 398783
rect 676128 397588 676180 397594
rect 676128 397530 676180 397536
rect 676036 397520 676088 397526
rect 676036 397462 676088 397468
rect 676034 397352 676090 397361
rect 676034 397287 676090 397296
rect 676048 397050 676076 397287
rect 676036 397044 676088 397050
rect 676036 396986 676088 396992
rect 676034 396944 676090 396953
rect 676034 396879 676090 396888
rect 675942 396128 675998 396137
rect 675942 396063 675998 396072
rect 675956 395010 675984 396063
rect 675944 395004 675996 395010
rect 675944 394946 675996 394952
rect 675942 394904 675998 394913
rect 675942 394839 675998 394848
rect 675956 394806 675984 394839
rect 675944 394800 675996 394806
rect 675944 394742 675996 394748
rect 676048 394738 676076 396879
rect 676126 396400 676182 396409
rect 676126 396335 676182 396344
rect 676140 394874 676168 396335
rect 676128 394868 676180 394874
rect 676128 394810 676180 394816
rect 676036 394732 676088 394738
rect 676036 394674 676088 394680
rect 676034 394496 676090 394505
rect 676034 394431 676090 394440
rect 676048 394194 676076 394431
rect 676036 394188 676088 394194
rect 676036 394130 676088 394136
rect 676034 394088 676090 394097
rect 676034 394023 676090 394032
rect 676048 392018 676076 394023
rect 678978 393544 679034 393553
rect 678978 393479 679034 393488
rect 678992 392737 679020 393479
rect 678978 392728 679034 392737
rect 678978 392663 679034 392672
rect 678992 392086 679020 392663
rect 678980 392080 679032 392086
rect 678980 392022 679032 392028
rect 676036 392012 676088 392018
rect 676036 391954 676088 391960
rect 675772 390374 675892 390402
rect 675772 386646 675800 390374
rect 675760 386640 675812 386646
rect 675760 386582 675812 386588
rect 675404 386034 675432 386275
rect 675392 386028 675444 386034
rect 675392 385970 675444 385976
rect 675760 386028 675812 386034
rect 675760 385970 675812 385976
rect 675772 385696 675800 385970
rect 675392 385620 675444 385626
rect 675392 385562 675444 385568
rect 675404 385084 675432 385562
rect 675392 384804 675444 384810
rect 675392 384746 675444 384752
rect 675404 384435 675432 384746
rect 675392 383172 675444 383178
rect 675392 383114 675444 383120
rect 675404 382568 675432 383114
rect 675392 382492 675444 382498
rect 675392 382434 675444 382440
rect 675404 382024 675432 382434
rect 675392 381948 675444 381954
rect 675392 381890 675444 381896
rect 675404 381412 675432 381890
rect 675392 381132 675444 381138
rect 675392 381074 675444 381080
rect 675404 380732 675432 381074
rect 675392 378820 675444 378826
rect 675392 378762 675444 378768
rect 675404 378284 675432 378762
rect 675484 378004 675536 378010
rect 675484 377946 675536 377952
rect 675496 377740 675524 377946
rect 675392 377460 675444 377466
rect 675392 377402 675444 377408
rect 675404 377060 675432 377402
rect 675484 376984 675536 376990
rect 675484 376926 675536 376932
rect 675496 376448 675524 376926
rect 675392 375760 675444 375766
rect 675392 375702 675444 375708
rect 675404 375224 675432 375702
rect 675392 373924 675444 373930
rect 675392 373866 675444 373872
rect 675404 373388 675432 373866
rect 675392 372088 675444 372094
rect 675392 372030 675444 372036
rect 675404 371552 675432 372030
rect 675668 370796 675720 370802
rect 675668 370738 675720 370744
rect 675298 357504 675354 357513
rect 675298 357439 675354 357448
rect 675206 357096 675262 357105
rect 675206 357031 675262 357040
rect 673368 356176 673420 356182
rect 673368 356118 673420 356124
rect 672724 347268 672776 347274
rect 672724 347210 672776 347216
rect 672630 143168 672686 143177
rect 672630 143103 672686 143112
rect 672736 138417 672764 347210
rect 673276 342576 673328 342582
rect 673276 342518 673328 342524
rect 673288 340134 673316 342518
rect 673276 340128 673328 340134
rect 673276 340070 673328 340076
rect 673000 311908 673052 311914
rect 673000 311850 673052 311856
rect 672816 300892 672868 300898
rect 672816 300834 672868 300840
rect 672722 138408 672778 138417
rect 672722 138343 672778 138352
rect 672828 132977 672856 300834
rect 673012 267510 673040 311850
rect 673380 311710 673408 356118
rect 674656 353524 674708 353530
rect 674656 353466 674708 353472
rect 674564 352300 674616 352306
rect 674564 352242 674616 352248
rect 673644 351484 673696 351490
rect 673644 351426 673696 351432
rect 673552 350804 673604 350810
rect 673552 350746 673604 350752
rect 673460 347948 673512 347954
rect 673460 347890 673512 347896
rect 673472 342514 673500 347890
rect 673564 342582 673592 350746
rect 673552 342576 673604 342582
rect 673552 342518 673604 342524
rect 673460 342508 673512 342514
rect 673460 342450 673512 342456
rect 673656 342394 673684 351426
rect 674288 350736 674340 350742
rect 674288 350678 674340 350684
rect 673828 349852 673880 349858
rect 673828 349794 673880 349800
rect 673736 347880 673788 347886
rect 673736 347822 673788 347828
rect 673564 342366 673684 342394
rect 673460 342304 673512 342310
rect 673460 342246 673512 342252
rect 673472 331634 673500 342246
rect 673460 331628 673512 331634
rect 673460 331570 673512 331576
rect 673564 326942 673592 342366
rect 673644 342304 673696 342310
rect 673644 342246 673696 342252
rect 673656 333606 673684 342246
rect 673644 333600 673696 333606
rect 673644 333542 673696 333548
rect 673748 332790 673776 347822
rect 673736 332784 673788 332790
rect 673736 332726 673788 332732
rect 673840 332246 673868 349794
rect 674300 336598 674328 350678
rect 674472 347812 674524 347818
rect 674472 347754 674524 347760
rect 674288 336592 674340 336598
rect 674288 336534 674340 336540
rect 674484 336122 674512 347754
rect 674576 342310 674604 352242
rect 674564 342304 674616 342310
rect 674564 342246 674616 342252
rect 674564 341488 674616 341494
rect 674564 341430 674616 341436
rect 674472 336116 674524 336122
rect 674472 336058 674524 336064
rect 674576 332450 674604 341430
rect 674668 339590 674696 353466
rect 674932 353320 674984 353326
rect 674932 353262 674984 353268
rect 674840 351892 674892 351898
rect 674840 351834 674892 351840
rect 674748 350668 674800 350674
rect 674748 350610 674800 350616
rect 674656 339584 674708 339590
rect 674656 339526 674708 339532
rect 674760 337142 674788 350610
rect 674852 337958 674880 351834
rect 674944 341018 674972 353262
rect 675024 350600 675076 350606
rect 675024 350542 675076 350548
rect 674932 341012 674984 341018
rect 674932 340954 674984 340960
rect 675036 340950 675064 350542
rect 675116 341420 675168 341426
rect 675116 341362 675168 341368
rect 675024 340944 675076 340950
rect 675024 340886 675076 340892
rect 675128 340762 675156 341362
rect 674944 340734 675156 340762
rect 674840 337952 674892 337958
rect 674840 337894 674892 337900
rect 674748 337136 674800 337142
rect 674748 337078 674800 337084
rect 674564 332444 674616 332450
rect 674564 332386 674616 332392
rect 673828 332240 673880 332246
rect 673828 332182 673880 332188
rect 674944 328778 674972 340734
rect 675024 340672 675076 340678
rect 675024 340614 675076 340620
rect 675116 340672 675168 340678
rect 675116 340614 675168 340620
rect 675036 340270 675064 340614
rect 675024 340264 675076 340270
rect 675024 340206 675076 340212
rect 675024 340128 675076 340134
rect 675024 340070 675076 340076
rect 675036 330614 675064 340070
rect 675128 335374 675156 340614
rect 675116 335368 675168 335374
rect 675116 335310 675168 335316
rect 675116 332580 675168 332586
rect 675116 332522 675168 332528
rect 675024 330608 675076 330614
rect 675024 330550 675076 330556
rect 674932 328772 674984 328778
rect 674932 328714 674984 328720
rect 673552 326936 673604 326942
rect 673552 326878 673604 326884
rect 673368 311704 673420 311710
rect 673368 311646 673420 311652
rect 675128 311574 675156 332522
rect 675220 314634 675248 357031
rect 675680 355065 675708 370738
rect 675760 370728 675812 370734
rect 675760 370670 675812 370676
rect 675772 356697 675800 370670
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675850 358728 675906 358737
rect 675850 358663 675906 358672
rect 675758 356688 675814 356697
rect 675758 356623 675814 356632
rect 675864 356318 675892 358663
rect 676034 358320 676090 358329
rect 676034 358255 676090 358264
rect 675942 357912 675998 357921
rect 675942 357847 675998 357856
rect 675852 356312 675904 356318
rect 675852 356254 675904 356260
rect 675956 356250 675984 357847
rect 676048 356454 676076 358255
rect 676036 356448 676088 356454
rect 676036 356390 676088 356396
rect 676034 356280 676090 356289
rect 675944 356244 675996 356250
rect 676034 356215 676090 356224
rect 675944 356186 675996 356192
rect 676048 356182 676076 356215
rect 676036 356176 676088 356182
rect 676036 356118 676088 356124
rect 675758 355464 675814 355473
rect 675758 355399 675814 355408
rect 675666 355056 675722 355065
rect 675666 354991 675722 355000
rect 675298 354648 675354 354657
rect 675298 354583 675354 354592
rect 675312 332586 675340 354583
rect 675390 353832 675446 353841
rect 675390 353767 675446 353776
rect 675404 341426 675432 353767
rect 675668 350804 675720 350810
rect 675668 350746 675720 350752
rect 675680 350577 675708 350746
rect 675666 350568 675722 350577
rect 675666 350503 675722 350512
rect 675772 341494 675800 355399
rect 676034 354240 676090 354249
rect 676034 354175 676090 354184
rect 676048 353530 676076 354175
rect 676036 353524 676088 353530
rect 676036 353466 676088 353472
rect 676034 353424 676090 353433
rect 676034 353359 676090 353368
rect 676048 353326 676076 353359
rect 676036 353320 676088 353326
rect 676036 353262 676088 353268
rect 676034 353016 676090 353025
rect 676034 352951 676090 352960
rect 675942 352608 675998 352617
rect 675942 352543 675998 352552
rect 675956 352306 675984 352543
rect 675944 352300 675996 352306
rect 675944 352242 675996 352248
rect 675942 352200 675998 352209
rect 675942 352135 675998 352144
rect 675956 351490 675984 352135
rect 676048 351898 676076 352951
rect 676036 351892 676088 351898
rect 676036 351834 676088 351840
rect 676034 351792 676090 351801
rect 676034 351727 676090 351736
rect 675944 351484 675996 351490
rect 675944 351426 675996 351432
rect 675942 351384 675998 351393
rect 675942 351319 675998 351328
rect 675850 350976 675906 350985
rect 675850 350911 675906 350920
rect 675864 350742 675892 350911
rect 675852 350736 675904 350742
rect 675852 350678 675904 350684
rect 675956 350674 675984 351319
rect 675944 350668 675996 350674
rect 675944 350610 675996 350616
rect 676048 350606 676076 351727
rect 676036 350600 676088 350606
rect 676036 350542 676088 350548
rect 676034 350160 676090 350169
rect 676034 350095 676090 350104
rect 676048 349858 676076 350095
rect 676036 349852 676088 349858
rect 676036 349794 676088 349800
rect 676034 349752 676090 349761
rect 676034 349687 676090 349696
rect 675942 349344 675998 349353
rect 675942 349279 675998 349288
rect 675850 348936 675906 348945
rect 675850 348871 675906 348880
rect 675864 347954 675892 348871
rect 675852 347948 675904 347954
rect 675852 347890 675904 347896
rect 675956 347886 675984 349279
rect 675944 347880 675996 347886
rect 675944 347822 675996 347828
rect 676048 347818 676076 349687
rect 676036 347812 676088 347818
rect 676036 347754 676088 347760
rect 676034 347304 676090 347313
rect 676034 347239 676036 347248
rect 676088 347239 676090 347248
rect 676036 347210 676088 347216
rect 675760 341488 675812 341494
rect 675760 341430 675812 341436
rect 675392 341420 675444 341426
rect 675392 341362 675444 341368
rect 675404 340678 675432 341088
rect 675484 341012 675536 341018
rect 675484 340954 675536 340960
rect 675392 340672 675444 340678
rect 675392 340614 675444 340620
rect 675496 340544 675524 340954
rect 675392 340264 675444 340270
rect 675392 340206 675444 340212
rect 675404 339864 675432 340206
rect 675484 339584 675536 339590
rect 675484 339526 675536 339532
rect 675496 339252 675524 339526
rect 675484 337952 675536 337958
rect 675484 337894 675536 337900
rect 675496 337416 675524 337894
rect 675392 337136 675444 337142
rect 675392 337078 675444 337084
rect 675404 336843 675432 337078
rect 675392 336592 675444 336598
rect 675392 336534 675444 336540
rect 675404 336192 675432 336534
rect 675484 336116 675536 336122
rect 675484 336058 675536 336064
rect 675496 335580 675524 336058
rect 675392 333600 675444 333606
rect 675392 333542 675444 333548
rect 675404 333064 675432 333542
rect 675392 332784 675444 332790
rect 675392 332726 675444 332732
rect 675300 332580 675352 332586
rect 675300 332522 675352 332528
rect 675404 332520 675432 332726
rect 675300 332444 675352 332450
rect 675300 332386 675352 332392
rect 675208 314628 675260 314634
rect 675208 314570 675260 314576
rect 675116 311568 675168 311574
rect 675116 311510 675168 311516
rect 673276 311092 673328 311098
rect 673276 311034 673328 311040
rect 673184 310276 673236 310282
rect 673184 310218 673236 310224
rect 673092 309460 673144 309466
rect 673092 309402 673144 309408
rect 673000 267504 673052 267510
rect 673000 267446 673052 267452
rect 673104 264994 673132 309402
rect 673196 265878 673224 310218
rect 673288 266694 673316 311034
rect 675312 310865 675340 332386
rect 675392 332240 675444 332246
rect 675392 332182 675444 332188
rect 675404 331875 675432 332182
rect 675392 331628 675444 331634
rect 675392 331570 675444 331576
rect 675404 331228 675432 331570
rect 675392 330608 675444 330614
rect 675392 330550 675444 330556
rect 675404 330035 675432 330550
rect 675392 328772 675444 328778
rect 675392 328714 675444 328720
rect 675404 328168 675432 328714
rect 675392 326936 675444 326942
rect 675392 326878 675444 326884
rect 675404 326332 675432 326878
rect 676036 314628 676088 314634
rect 676036 314570 676088 314576
rect 676048 312497 676076 314570
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676310 313576 676366 313585
rect 676310 313511 676366 313520
rect 676126 313168 676182 313177
rect 676126 313103 676182 313112
rect 676034 312488 676090 312497
rect 676034 312423 676090 312432
rect 676140 311982 676168 313103
rect 676218 312760 676274 312769
rect 676218 312695 676274 312704
rect 676232 312118 676260 312695
rect 676220 312112 676272 312118
rect 676220 312054 676272 312060
rect 676324 312050 676352 313511
rect 676312 312044 676364 312050
rect 676312 311986 676364 311992
rect 676128 311976 676180 311982
rect 676128 311918 676180 311924
rect 676218 311944 676274 311953
rect 676218 311879 676220 311888
rect 676272 311879 676274 311888
rect 676220 311850 676272 311856
rect 676036 311704 676088 311710
rect 676034 311672 676036 311681
rect 676088 311672 676090 311681
rect 676034 311607 676090 311616
rect 676036 311568 676088 311574
rect 676036 311510 676088 311516
rect 675298 310856 675354 310865
rect 675298 310791 675354 310800
rect 676048 310049 676076 311510
rect 676218 311128 676274 311137
rect 676218 311063 676220 311072
rect 676272 311063 676274 311072
rect 676220 311034 676272 311040
rect 676218 310312 676274 310321
rect 676218 310247 676220 310256
rect 676272 310247 676274 310256
rect 676220 310218 676272 310224
rect 676034 310040 676090 310049
rect 676034 309975 676090 309984
rect 676218 309496 676274 309505
rect 676218 309431 676220 309440
rect 676272 309431 676274 309440
rect 676220 309402 676272 309408
rect 676034 309224 676090 309233
rect 674656 309188 674708 309194
rect 676034 309159 676036 309168
rect 674656 309130 674708 309136
rect 676088 309159 676090 309168
rect 676036 309130 676088 309136
rect 673552 308100 673604 308106
rect 673552 308042 673604 308048
rect 673564 283762 673592 308042
rect 674288 306468 674340 306474
rect 674288 306410 674340 306416
rect 673828 305108 673880 305114
rect 673828 305050 673880 305056
rect 673736 304360 673788 304366
rect 673736 304302 673788 304308
rect 673644 303748 673696 303754
rect 673644 303690 673696 303696
rect 673656 286618 673684 303690
rect 673748 287434 673776 304302
rect 673736 287428 673788 287434
rect 673736 287370 673788 287376
rect 673840 286822 673868 305050
rect 674300 288658 674328 306410
rect 674472 303952 674524 303958
rect 674472 303894 674524 303900
rect 674484 290494 674512 303894
rect 674668 294574 674696 309130
rect 676034 308816 676090 308825
rect 676034 308751 676090 308760
rect 675758 308408 675814 308417
rect 675758 308343 675814 308352
rect 674932 307284 674984 307290
rect 674932 307226 674984 307232
rect 674840 306876 674892 306882
rect 674840 306818 674892 306824
rect 674852 300218 674880 306818
rect 674840 300212 674892 300218
rect 674840 300154 674892 300160
rect 674944 300098 674972 307226
rect 675024 306400 675076 306406
rect 675024 306342 675076 306348
rect 675298 306368 675354 306377
rect 674760 300070 674972 300098
rect 675036 300082 675064 306342
rect 675298 306303 675354 306312
rect 675116 304836 675168 304842
rect 675116 304778 675168 304784
rect 675024 300076 675076 300082
rect 674760 294778 674788 300070
rect 675024 300018 675076 300024
rect 674840 300008 674892 300014
rect 675128 299962 675156 304778
rect 675208 304224 675260 304230
rect 675208 304166 675260 304172
rect 674840 299950 674892 299956
rect 674748 294772 674800 294778
rect 674748 294714 674800 294720
rect 674656 294568 674708 294574
rect 674656 294510 674708 294516
rect 674472 290488 674524 290494
rect 674472 290430 674524 290436
rect 674288 288652 674340 288658
rect 674288 288594 674340 288600
rect 673828 286816 673880 286822
rect 673828 286758 673880 286764
rect 673644 286612 673696 286618
rect 673644 286554 673696 286560
rect 674852 284294 674880 299950
rect 674944 299934 675156 299962
rect 674944 291582 674972 299934
rect 675024 299872 675076 299878
rect 675220 299826 675248 304166
rect 675024 299814 675076 299820
rect 675036 295458 675064 299814
rect 675128 299798 675248 299826
rect 675024 295452 675076 295458
rect 675024 295394 675076 295400
rect 675128 295338 675156 299798
rect 675312 299690 675340 306303
rect 675036 295310 675156 295338
rect 675220 299662 675340 299690
rect 675036 291802 675064 295310
rect 675220 291870 675248 299662
rect 675772 299554 675800 308343
rect 676048 308106 676076 308751
rect 676036 308100 676088 308106
rect 676036 308042 676088 308048
rect 676034 308000 676090 308009
rect 676034 307935 676090 307944
rect 676048 307290 676076 307935
rect 676126 307456 676182 307465
rect 676126 307391 676182 307400
rect 676036 307284 676088 307290
rect 676036 307226 676088 307232
rect 676034 307184 676090 307193
rect 676034 307119 676090 307128
rect 676048 306882 676076 307119
rect 676036 306876 676088 306882
rect 676036 306818 676088 306824
rect 676034 306776 676090 306785
rect 676034 306711 676090 306720
rect 676048 306406 676076 306711
rect 676140 306474 676168 307391
rect 676128 306468 676180 306474
rect 676128 306410 676180 306416
rect 676036 306400 676088 306406
rect 676036 306342 676088 306348
rect 676034 305960 676090 305969
rect 676034 305895 676090 305904
rect 676048 304842 676076 305895
rect 676126 305416 676182 305425
rect 676126 305351 676182 305360
rect 676140 305114 676168 305351
rect 676128 305108 676180 305114
rect 676128 305050 676180 305056
rect 676126 305008 676182 305017
rect 676126 304943 676182 304952
rect 676036 304836 676088 304842
rect 676036 304778 676088 304784
rect 676034 304736 676090 304745
rect 676034 304671 676090 304680
rect 676048 304230 676076 304671
rect 676140 304366 676168 304943
rect 676128 304360 676180 304366
rect 676128 304302 676180 304308
rect 676036 304224 676088 304230
rect 676036 304166 676088 304172
rect 676126 304192 676182 304201
rect 676126 304127 676182 304136
rect 676140 303958 676168 304127
rect 676128 303952 676180 303958
rect 676034 303920 676090 303929
rect 676128 303894 676180 303900
rect 676034 303855 676090 303864
rect 676048 303754 676076 303855
rect 676036 303748 676088 303754
rect 676036 303690 676088 303696
rect 678978 303376 679034 303385
rect 678978 303311 679034 303320
rect 678992 302569 679020 303311
rect 678978 302560 679034 302569
rect 678978 302495 679034 302504
rect 678992 300898 679020 302495
rect 678980 300892 679032 300898
rect 678980 300834 679032 300840
rect 675312 299526 675800 299554
rect 675312 295542 675340 299526
rect 675392 298172 675444 298178
rect 675392 298114 675444 298120
rect 675404 296072 675432 298114
rect 675312 295514 675418 295542
rect 675300 295452 675352 295458
rect 675300 295394 675352 295400
rect 675312 294893 675340 295394
rect 675312 294865 675418 294893
rect 675300 294772 675352 294778
rect 675300 294714 675352 294720
rect 675312 292414 675340 294714
rect 675392 294568 675444 294574
rect 675392 294510 675444 294516
rect 675404 294236 675432 294510
rect 675312 292386 675418 292414
rect 675220 291842 675418 291870
rect 675036 291774 675248 291802
rect 674932 291576 674984 291582
rect 674932 291518 674984 291524
rect 675220 290578 675248 291774
rect 675392 291576 675444 291582
rect 675392 291518 675444 291524
rect 675404 291176 675432 291518
rect 675220 290550 675418 290578
rect 675116 290488 675168 290494
rect 675116 290430 675168 290436
rect 675128 287518 675156 290430
rect 675392 288652 675444 288658
rect 675392 288594 675444 288600
rect 675404 288048 675432 288594
rect 675128 287490 675418 287518
rect 675116 287428 675168 287434
rect 675116 287370 675168 287376
rect 675128 286906 675156 287370
rect 675128 286878 675340 286906
rect 675116 286816 675168 286822
rect 675116 286758 675168 286764
rect 675312 286770 675340 286878
rect 675404 286770 675432 286892
rect 675128 285070 675156 286758
rect 675312 286742 675432 286770
rect 675392 286612 675444 286618
rect 675392 286554 675444 286560
rect 675404 286212 675432 286554
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 674852 284266 675248 284294
rect 673552 283756 673604 283762
rect 673552 283698 673604 283704
rect 675220 281369 675248 284266
rect 675484 283756 675536 283762
rect 675484 283698 675536 283704
rect 675496 283220 675524 283698
rect 675220 281341 675418 281369
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 676126 268560 676182 268569
rect 676126 268495 676182 268504
rect 676034 268288 676090 268297
rect 676034 268223 676090 268232
rect 676048 267986 676076 268223
rect 676036 267980 676088 267986
rect 676036 267922 676088 267928
rect 676140 267782 676168 268495
rect 676218 268152 676274 268161
rect 676218 268087 676220 268096
rect 676272 268087 676274 268096
rect 676220 268058 676272 268064
rect 676128 267776 676180 267782
rect 676128 267718 676180 267724
rect 676036 267504 676088 267510
rect 676034 267472 676036 267481
rect 676088 267472 676090 267481
rect 676034 267407 676090 267416
rect 675666 267064 675722 267073
rect 675666 266999 675722 267008
rect 673276 266688 673328 266694
rect 673276 266630 673328 266636
rect 673184 265872 673236 265878
rect 673184 265814 673236 265820
rect 673092 264988 673144 264994
rect 675680 264974 675708 266999
rect 676036 266688 676088 266694
rect 676034 266656 676036 266665
rect 676088 266656 676090 266665
rect 676034 266591 676090 266600
rect 675758 266248 675814 266257
rect 675758 266183 675814 266192
rect 673092 264930 673144 264936
rect 675312 264946 675708 264974
rect 674288 264308 674340 264314
rect 674288 264250 674340 264256
rect 673644 262336 673696 262342
rect 673644 262278 673696 262284
rect 673460 260228 673512 260234
rect 673460 260170 673512 260176
rect 672908 256896 672960 256902
rect 672908 256838 672960 256844
rect 672814 132968 672870 132977
rect 672814 132903 672870 132912
rect 672172 131708 672224 131714
rect 672172 131650 672224 131656
rect 672080 130076 672132 130082
rect 672080 130018 672132 130024
rect 671986 114336 672042 114345
rect 671986 114271 672042 114280
rect 670882 107536 670938 107545
rect 670882 107471 670938 107480
rect 672092 100881 672120 130018
rect 672184 104145 672212 131650
rect 672264 130892 672316 130898
rect 672264 130834 672316 130840
rect 672276 105913 672304 130834
rect 672356 129464 672408 129470
rect 672356 129406 672408 129412
rect 672262 105904 672318 105913
rect 672262 105839 672318 105848
rect 672170 104136 672226 104145
rect 672170 104071 672226 104080
rect 672368 102513 672396 129406
rect 672920 127945 672948 256838
rect 673368 250980 673420 250986
rect 673368 250922 673420 250928
rect 673380 249354 673408 250922
rect 673368 249348 673420 249354
rect 673368 249290 673420 249296
rect 673472 240582 673500 260170
rect 673552 259616 673604 259622
rect 673552 259558 673604 259564
rect 673564 242214 673592 259558
rect 673656 246430 673684 262278
rect 673828 261452 673880 261458
rect 673828 261394 673880 261400
rect 673736 256828 673788 256834
rect 673736 256770 673788 256776
rect 673644 246424 673696 246430
rect 673644 246366 673696 246372
rect 673644 246288 673696 246294
rect 673644 246230 673696 246236
rect 673656 243642 673684 246230
rect 673644 243636 673696 243642
rect 673644 243578 673696 243584
rect 673552 242208 673604 242214
rect 673552 242150 673604 242156
rect 673748 241806 673776 256770
rect 673840 249490 673868 261394
rect 673828 249484 673880 249490
rect 673828 249426 673880 249432
rect 673828 249348 673880 249354
rect 673828 249290 673880 249296
rect 673840 246294 673868 249290
rect 673828 246288 673880 246294
rect 673828 246230 673880 246236
rect 674300 246158 674328 264250
rect 674472 263084 674524 263090
rect 674472 263026 674524 263032
rect 674484 249626 674512 263026
rect 674932 262404 674984 262410
rect 674932 262346 674984 262352
rect 674564 262268 674616 262274
rect 674564 262210 674616 262216
rect 674472 249620 674524 249626
rect 674472 249562 674524 249568
rect 674472 249484 674524 249490
rect 674472 249426 674524 249432
rect 674288 246152 674340 246158
rect 674288 246094 674340 246100
rect 673736 241800 673788 241806
rect 673736 241742 673788 241748
rect 673460 240576 673512 240582
rect 673460 240518 673512 240524
rect 674484 236910 674512 249426
rect 674576 247926 674604 262210
rect 674748 259548 674800 259554
rect 674748 259490 674800 259496
rect 674656 256760 674708 256766
rect 674656 256702 674708 256708
rect 674564 247920 674616 247926
rect 674564 247862 674616 247868
rect 674668 247178 674696 256702
rect 674656 247172 674708 247178
rect 674656 247114 674708 247120
rect 674760 246566 674788 259490
rect 674840 259480 674892 259486
rect 674840 259422 674892 259428
rect 674748 246560 674800 246566
rect 674748 246502 674800 246508
rect 674748 246424 674800 246430
rect 674748 246366 674800 246372
rect 674760 238746 674788 246366
rect 674852 246090 674880 259422
rect 674944 250986 674972 262346
rect 675024 259820 675076 259826
rect 675024 259762 675076 259768
rect 674932 250980 674984 250986
rect 674932 250922 674984 250928
rect 674932 250844 674984 250850
rect 674932 250786 674984 250792
rect 674840 246084 674892 246090
rect 674840 246026 674892 246032
rect 674944 245614 674972 250786
rect 675036 247314 675064 259762
rect 675116 255332 675168 255338
rect 675116 255274 675168 255280
rect 675024 247308 675076 247314
rect 675024 247250 675076 247256
rect 675024 247172 675076 247178
rect 675024 247114 675076 247120
rect 674932 245608 674984 245614
rect 674932 245550 674984 245556
rect 675036 242826 675064 247114
rect 675024 242820 675076 242826
rect 675024 242762 675076 242768
rect 675128 242706 675156 255274
rect 675206 250200 675262 250209
rect 675206 250135 675262 250144
rect 675220 246265 675248 250135
rect 675206 246256 675262 246265
rect 675206 246191 675262 246200
rect 675208 246152 675260 246158
rect 675208 246094 675260 246100
rect 675036 242678 675156 242706
rect 674748 238740 674800 238746
rect 674748 238682 674800 238688
rect 674472 236904 674524 236910
rect 674472 236846 674524 236852
rect 675036 235618 675064 242678
rect 675024 235612 675076 235618
rect 675024 235554 675076 235560
rect 675220 220794 675248 246094
rect 675312 235634 675340 264946
rect 675482 263392 675538 263401
rect 675482 263327 675538 263336
rect 675496 251394 675524 263327
rect 675772 255338 675800 266183
rect 676036 265872 676088 265878
rect 676034 265840 676036 265849
rect 676088 265840 676090 265849
rect 676034 265775 676090 265784
rect 676220 264988 676272 264994
rect 676220 264930 676272 264936
rect 676232 264897 676260 264930
rect 676218 264888 676274 264897
rect 676218 264823 676274 264832
rect 676034 264616 676090 264625
rect 676034 264551 676090 264560
rect 676048 264314 676076 264551
rect 676036 264308 676088 264314
rect 676036 264250 676088 264256
rect 676034 264208 676090 264217
rect 676034 264143 676090 264152
rect 676048 263090 676076 264143
rect 676126 263664 676182 263673
rect 676126 263599 676182 263608
rect 676036 263084 676088 263090
rect 676036 263026 676088 263032
rect 676034 262984 676090 262993
rect 676034 262919 676090 262928
rect 675942 262576 675998 262585
rect 675942 262511 675998 262520
rect 675956 262410 675984 262511
rect 675944 262404 675996 262410
rect 675944 262346 675996 262352
rect 676048 262274 676076 262919
rect 676140 262342 676168 263599
rect 676128 262336 676180 262342
rect 676128 262278 676180 262284
rect 676036 262268 676088 262274
rect 676036 262210 676088 262216
rect 676034 262168 676090 262177
rect 676034 262103 676090 262112
rect 675850 261760 675906 261769
rect 675850 261695 675906 261704
rect 675760 255332 675812 255338
rect 675760 255274 675812 255280
rect 675864 255218 675892 261695
rect 676048 261458 676076 262103
rect 676036 261452 676088 261458
rect 676036 261394 676088 261400
rect 676034 261352 676090 261361
rect 676034 261287 676090 261296
rect 675942 260536 675998 260545
rect 675942 260471 675998 260480
rect 675956 260234 675984 260471
rect 675944 260228 675996 260234
rect 675944 260170 675996 260176
rect 675942 260128 675998 260137
rect 675942 260063 675998 260072
rect 675956 259622 675984 260063
rect 676048 259826 676076 261287
rect 676126 260808 676182 260817
rect 676126 260743 676182 260752
rect 676036 259820 676088 259826
rect 676036 259762 676088 259768
rect 676034 259720 676090 259729
rect 676034 259655 676090 259664
rect 675944 259616 675996 259622
rect 675944 259558 675996 259564
rect 676048 259486 676076 259655
rect 676140 259554 676168 260743
rect 676128 259548 676180 259554
rect 676128 259490 676180 259496
rect 676036 259480 676088 259486
rect 676036 259422 676088 259428
rect 676034 259312 676090 259321
rect 676034 259247 676090 259256
rect 676048 256766 676076 259247
rect 676126 258768 676182 258777
rect 676126 258703 676182 258712
rect 676140 256834 676168 258703
rect 678978 258360 679034 258369
rect 678978 258295 679034 258304
rect 678992 257553 679020 258295
rect 678978 257544 679034 257553
rect 678978 257479 679034 257488
rect 678992 256902 679020 257479
rect 678980 256896 679032 256902
rect 678980 256838 679032 256844
rect 676128 256828 676180 256834
rect 676128 256770 676180 256776
rect 676036 256760 676088 256766
rect 676036 256702 676088 256708
rect 675772 255190 675892 255218
rect 675772 251394 675800 255190
rect 675484 251388 675536 251394
rect 675484 251330 675536 251336
rect 675760 251388 675812 251394
rect 675760 251330 675812 251336
rect 675392 250980 675444 250986
rect 675392 250922 675444 250928
rect 675404 250512 675432 250922
rect 675496 250850 675524 251056
rect 675484 250844 675536 250850
rect 675484 250786 675536 250792
rect 675760 250232 675812 250238
rect 675760 250174 675812 250180
rect 675772 249900 675800 250174
rect 675392 249620 675444 249626
rect 675392 249562 675444 249568
rect 675404 249220 675432 249562
rect 675392 247920 675444 247926
rect 675392 247862 675444 247868
rect 675404 247384 675432 247862
rect 675392 247104 675444 247110
rect 675392 247046 675444 247052
rect 675404 246840 675432 247046
rect 675392 246560 675444 246566
rect 675392 246502 675444 246508
rect 675404 246199 675432 246502
rect 675392 246084 675444 246090
rect 675392 246026 675444 246032
rect 675404 245548 675432 246026
rect 675392 243636 675444 243642
rect 675392 243578 675444 243584
rect 675404 243071 675432 243578
rect 675392 242820 675444 242826
rect 675392 242762 675444 242768
rect 675404 242519 675432 242762
rect 675392 242208 675444 242214
rect 675392 242150 675444 242156
rect 675404 241876 675432 242150
rect 675392 241800 675444 241806
rect 675392 241742 675444 241748
rect 675404 241231 675432 241742
rect 675392 240576 675444 240582
rect 675392 240518 675444 240524
rect 675404 240040 675432 240518
rect 675392 238740 675444 238746
rect 675392 238682 675444 238688
rect 675404 238204 675432 238682
rect 675392 236904 675444 236910
rect 675392 236846 675444 236852
rect 675404 236368 675432 236846
rect 675312 235606 675708 235634
rect 675680 222329 675708 235606
rect 675760 235612 675812 235618
rect 675760 235554 675812 235560
rect 675666 222320 675722 222329
rect 675666 222255 675722 222264
rect 675298 221912 675354 221921
rect 675298 221847 675354 221856
rect 675208 220788 675260 220794
rect 675208 220730 675260 220736
rect 675312 219586 675340 221847
rect 675772 221513 675800 235554
rect 703694 224196 703722 224332
rect 704154 224196 704182 224332
rect 704614 224196 704642 224332
rect 705074 224196 705102 224332
rect 705534 224196 705562 224332
rect 705994 224196 706022 224332
rect 706454 224196 706482 224332
rect 706914 224196 706942 224332
rect 707374 224196 707402 224332
rect 707834 224196 707862 224332
rect 708294 224196 708322 224332
rect 708754 224196 708782 224332
rect 709214 224196 709242 224332
rect 675942 223544 675998 223553
rect 675942 223479 675998 223488
rect 675850 223136 675906 223145
rect 675850 223071 675906 223080
rect 675758 221504 675814 221513
rect 675758 221439 675814 221448
rect 675758 221096 675814 221105
rect 675758 221031 675814 221040
rect 675666 220280 675722 220289
rect 675666 220215 675722 220224
rect 675220 219558 675340 219586
rect 674564 218340 674616 218346
rect 674564 218282 674616 218288
rect 673828 216708 673880 216714
rect 673828 216650 673880 216656
rect 673552 216300 673604 216306
rect 673552 216242 673604 216248
rect 673460 215552 673512 215558
rect 673460 215494 673512 215500
rect 673092 213512 673144 213518
rect 673092 213454 673144 213460
rect 673000 212084 673052 212090
rect 673000 212026 673052 212032
rect 672906 127936 672962 127945
rect 672906 127871 672962 127880
rect 673012 122913 673040 212026
rect 673104 129470 673132 213454
rect 673368 206236 673420 206242
rect 673368 206178 673420 206184
rect 673380 200546 673408 206178
rect 673472 200682 673500 215494
rect 673564 200802 673592 216242
rect 673736 214668 673788 214674
rect 673736 214610 673788 214616
rect 673644 213852 673696 213858
rect 673644 213794 673696 213800
rect 673552 200796 673604 200802
rect 673552 200738 673604 200744
rect 673472 200654 673592 200682
rect 673380 200518 673500 200546
rect 673472 198422 673500 200518
rect 673460 198416 673512 198422
rect 673460 198358 673512 198364
rect 673564 195362 673592 200654
rect 673656 197810 673684 213794
rect 673644 197804 673696 197810
rect 673644 197746 673696 197752
rect 673748 197062 673776 214610
rect 673840 202774 673868 216650
rect 674472 215484 674524 215490
rect 674472 215426 674524 215432
rect 674288 212628 674340 212634
rect 674288 212570 674340 212576
rect 674300 203726 674328 212570
rect 674288 203720 674340 203726
rect 674288 203662 674340 203668
rect 673828 202768 673880 202774
rect 673828 202710 673880 202716
rect 674484 201550 674512 215426
rect 674576 205222 674604 218282
rect 674840 218068 674892 218074
rect 674840 218010 674892 218016
rect 674656 215416 674708 215422
rect 674656 215358 674708 215364
rect 674564 205216 674616 205222
rect 674564 205158 674616 205164
rect 674564 205080 674616 205086
rect 674564 205022 674616 205028
rect 674472 201544 674524 201550
rect 674472 201486 674524 201492
rect 674576 198734 674604 205022
rect 674668 202094 674696 215358
rect 674748 212560 674800 212566
rect 674748 212502 674800 212508
rect 674656 202088 674708 202094
rect 674656 202030 674708 202036
rect 674760 200938 674788 212502
rect 674852 208282 674880 218010
rect 674932 215348 674984 215354
rect 674932 215290 674984 215296
rect 674840 208276 674892 208282
rect 674840 208218 674892 208224
rect 674840 206304 674892 206310
rect 674840 206246 674892 206252
rect 674852 203862 674880 206246
rect 674944 205018 674972 215290
rect 675024 208412 675076 208418
rect 675024 208354 675076 208360
rect 674932 205012 674984 205018
rect 674932 204954 674984 204960
rect 674840 203856 674892 203862
rect 675036 203833 675064 208354
rect 675116 208344 675168 208350
rect 675116 208286 675168 208292
rect 675128 203930 675156 208286
rect 675116 203924 675168 203930
rect 675116 203866 675168 203872
rect 674840 203798 674892 203804
rect 675022 203824 675078 203833
rect 675022 203759 675078 203768
rect 675116 203788 675168 203794
rect 675116 203730 675168 203736
rect 674840 203720 674892 203726
rect 674840 203662 674892 203668
rect 674748 200932 674800 200938
rect 674748 200874 674800 200880
rect 674748 200796 674800 200802
rect 674748 200738 674800 200744
rect 674484 198706 674604 198734
rect 673736 197056 673788 197062
rect 673736 196998 673788 197004
rect 673552 195356 673604 195362
rect 673552 195298 673604 195304
rect 674484 192846 674512 198706
rect 674472 192840 674524 192846
rect 674472 192782 674524 192788
rect 674760 191690 674788 200738
rect 674852 196586 674880 203662
rect 675022 203552 675078 203561
rect 675022 203487 675078 203496
rect 674840 196580 674892 196586
rect 674840 196522 674892 196528
rect 674748 191684 674800 191690
rect 674748 191626 674800 191632
rect 675036 176390 675064 203487
rect 675128 176662 675156 203730
rect 675220 178634 675248 219558
rect 675298 219464 675354 219473
rect 675298 219399 675354 219408
rect 675312 208418 675340 219399
rect 675390 218648 675446 218657
rect 675390 218583 675446 218592
rect 675300 208412 675352 208418
rect 675300 208354 675352 208360
rect 675404 208350 675432 218583
rect 675482 217424 675538 217433
rect 675482 217359 675538 217368
rect 675392 208344 675444 208350
rect 675392 208286 675444 208292
rect 675300 208276 675352 208282
rect 675300 208218 675352 208224
rect 675312 205337 675340 208218
rect 675392 206984 675444 206990
rect 675392 206926 675444 206932
rect 675404 205875 675432 206926
rect 675496 206242 675524 217359
rect 675576 215552 675628 215558
rect 675576 215494 675628 215500
rect 675588 215393 675616 215494
rect 675574 215384 675630 215393
rect 675574 215319 675630 215328
rect 675680 206242 675708 220215
rect 675772 206310 675800 221031
rect 675864 220862 675892 223071
rect 675956 221202 675984 223479
rect 676034 222728 676090 222737
rect 676034 222663 676090 222672
rect 675944 221196 675996 221202
rect 675944 221138 675996 221144
rect 676048 221066 676076 222663
rect 676036 221060 676088 221066
rect 676036 221002 676088 221008
rect 675852 220856 675904 220862
rect 675852 220798 675904 220804
rect 676036 220788 676088 220794
rect 676036 220730 676088 220736
rect 676048 219881 676076 220730
rect 676034 219872 676090 219881
rect 676034 219807 676090 219816
rect 676034 219056 676090 219065
rect 676034 218991 676090 219000
rect 676048 218346 676076 218991
rect 676036 218340 676088 218346
rect 676036 218282 676088 218288
rect 676034 218240 676090 218249
rect 676034 218175 676090 218184
rect 676048 218074 676076 218175
rect 676036 218068 676088 218074
rect 676036 218010 676088 218016
rect 676034 217832 676090 217841
rect 676034 217767 676090 217776
rect 675942 217016 675998 217025
rect 675942 216951 675998 216960
rect 675956 216306 675984 216951
rect 676048 216714 676076 217767
rect 676036 216708 676088 216714
rect 676036 216650 676088 216656
rect 676034 216608 676090 216617
rect 676034 216543 676090 216552
rect 675944 216300 675996 216306
rect 675944 216242 675996 216248
rect 675942 216200 675998 216209
rect 675942 216135 675998 216144
rect 675850 215792 675906 215801
rect 675850 215727 675906 215736
rect 675864 215490 675892 215727
rect 675852 215484 675904 215490
rect 675852 215426 675904 215432
rect 675956 215422 675984 216135
rect 675944 215416 675996 215422
rect 675944 215358 675996 215364
rect 676048 215354 676076 216543
rect 676036 215348 676088 215354
rect 676036 215290 676088 215296
rect 676034 214976 676090 214985
rect 676034 214911 676090 214920
rect 676048 214674 676076 214911
rect 676036 214668 676088 214674
rect 676036 214610 676088 214616
rect 676034 214568 676090 214577
rect 676034 214503 676090 214512
rect 675942 214160 675998 214169
rect 675942 214095 675998 214104
rect 675956 213858 675984 214095
rect 675944 213852 675996 213858
rect 675944 213794 675996 213800
rect 675942 213752 675998 213761
rect 675942 213687 675998 213696
rect 675956 212634 675984 213687
rect 675944 212628 675996 212634
rect 675944 212570 675996 212576
rect 676048 212566 676076 214503
rect 676036 212560 676088 212566
rect 676036 212502 676088 212508
rect 676034 212120 676090 212129
rect 676034 212055 676036 212064
rect 676088 212055 676090 212064
rect 676036 212026 676088 212032
rect 675760 206304 675812 206310
rect 675760 206246 675812 206252
rect 675484 206236 675536 206242
rect 675484 206178 675536 206184
rect 675668 206236 675720 206242
rect 675668 206178 675720 206184
rect 675312 205309 675418 205337
rect 675300 205216 675352 205222
rect 675300 205158 675352 205164
rect 675312 204049 675340 205158
rect 675392 205012 675444 205018
rect 675392 204954 675444 204960
rect 675404 204680 675432 204954
rect 675312 204021 675418 204049
rect 675300 203924 675352 203930
rect 675300 203866 675352 203872
rect 675312 192998 675340 203866
rect 675392 202768 675444 202774
rect 675392 202710 675444 202716
rect 675404 202195 675432 202710
rect 675392 202088 675444 202094
rect 675392 202030 675444 202036
rect 675404 201620 675432 202030
rect 675392 201544 675444 201550
rect 675392 201486 675444 201492
rect 675404 201008 675432 201486
rect 675392 200932 675444 200938
rect 675392 200874 675444 200880
rect 675404 200328 675432 200874
rect 675392 198416 675444 198422
rect 675392 198358 675444 198364
rect 675404 197880 675432 198358
rect 675484 197804 675536 197810
rect 675484 197746 675536 197752
rect 675496 197336 675524 197746
rect 675392 197056 675444 197062
rect 675392 196998 675444 197004
rect 675404 196656 675432 196998
rect 675392 196580 675444 196586
rect 675392 196522 675444 196528
rect 675404 196044 675432 196522
rect 675392 195356 675444 195362
rect 675392 195298 675444 195304
rect 675404 194820 675432 195298
rect 675312 192970 675418 192998
rect 675300 192840 675352 192846
rect 675300 192782 675352 192788
rect 675208 178628 675260 178634
rect 675208 178570 675260 178576
rect 675116 176656 675168 176662
rect 675116 176598 675168 176604
rect 675024 176384 675076 176390
rect 675024 176326 675076 176332
rect 673184 176044 673236 176050
rect 673184 175986 673236 175992
rect 673196 131510 673224 175986
rect 675312 175681 675340 192782
rect 675392 191684 675444 191690
rect 675392 191626 675444 191632
rect 675404 191148 675432 191626
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 676220 178832 676272 178838
rect 676218 178800 676220 178809
rect 676272 178800 676274 178809
rect 676218 178735 676274 178744
rect 676036 178628 676088 178634
rect 676036 178570 676088 178576
rect 675944 178152 675996 178158
rect 675942 178120 675944 178129
rect 675996 178120 675998 178129
rect 675942 178055 675998 178064
rect 675944 177744 675996 177750
rect 675942 177712 675944 177721
rect 675996 177712 675998 177721
rect 675942 177647 675998 177656
rect 676048 177313 676076 178570
rect 676034 177304 676090 177313
rect 676034 177239 676090 177248
rect 676034 176896 676090 176905
rect 676034 176831 676036 176840
rect 676088 176831 676090 176840
rect 676036 176802 676088 176808
rect 676036 176656 676088 176662
rect 676036 176598 676088 176604
rect 676048 176497 676076 176598
rect 676034 176488 676090 176497
rect 676034 176423 676090 176432
rect 676036 176384 676088 176390
rect 676036 176326 676088 176332
rect 675942 176080 675998 176089
rect 675942 176015 675944 176024
rect 675996 176015 675998 176024
rect 675944 175986 675996 175992
rect 675298 175672 675354 175681
rect 675298 175607 675354 175616
rect 675942 175264 675998 175273
rect 673276 175228 673328 175234
rect 675942 175199 675944 175208
rect 673276 175170 673328 175176
rect 675996 175199 675998 175208
rect 675944 175170 675996 175176
rect 673184 131504 673236 131510
rect 673184 131446 673236 131452
rect 673288 130694 673316 175170
rect 676048 174865 676076 176326
rect 676034 174856 676090 174865
rect 676034 174791 676090 174800
rect 676034 174448 676090 174457
rect 673368 174412 673420 174418
rect 676034 174383 676036 174392
rect 673368 174354 673420 174360
rect 676088 174383 676090 174392
rect 676036 174354 676088 174360
rect 673276 130688 673328 130694
rect 673276 130630 673328 130636
rect 673380 129742 673408 174354
rect 676034 174040 676090 174049
rect 676034 173975 676090 173984
rect 676048 173942 676076 173975
rect 674564 173936 674616 173942
rect 674564 173878 674616 173884
rect 676036 173936 676088 173942
rect 676036 173878 676088 173884
rect 673552 172916 673604 172922
rect 673552 172858 673604 172864
rect 673564 148510 673592 172858
rect 673736 172100 673788 172106
rect 673736 172042 673788 172048
rect 673644 169244 673696 169250
rect 673644 169186 673696 169192
rect 673656 152114 673684 169186
rect 673748 155242 673776 172042
rect 674288 169652 674340 169658
rect 674288 169594 674340 169600
rect 673828 168632 673880 168638
rect 673828 168574 673880 168580
rect 673736 155236 673788 155242
rect 673736 155178 673788 155184
rect 673840 152182 673868 168574
rect 674300 152250 674328 169594
rect 674472 168564 674524 168570
rect 674472 168506 674524 168512
rect 674484 155310 674512 168506
rect 674576 159594 674604 173878
rect 676034 173632 676090 173641
rect 676034 173567 676090 173576
rect 675298 173224 675354 173233
rect 675298 173159 675354 173168
rect 674748 171692 674800 171698
rect 674748 171634 674800 171640
rect 674760 160206 674788 171634
rect 674932 171216 674984 171222
rect 674932 171158 674984 171164
rect 674840 168496 674892 168502
rect 674840 168438 674892 168444
rect 674748 160200 674800 160206
rect 674748 160142 674800 160148
rect 674852 159882 674880 168438
rect 674944 160290 674972 171158
rect 675024 171148 675076 171154
rect 675024 171090 675076 171096
rect 675036 160410 675064 171090
rect 675208 168428 675260 168434
rect 675208 168370 675260 168376
rect 675116 160540 675168 160546
rect 675116 160482 675168 160488
rect 675024 160404 675076 160410
rect 675024 160346 675076 160352
rect 674944 160262 675064 160290
rect 674932 160132 674984 160138
rect 674932 160074 674984 160080
rect 674944 160002 674972 160074
rect 675036 160070 675064 160262
rect 675024 160064 675076 160070
rect 675024 160006 675076 160012
rect 674932 159996 674984 160002
rect 674932 159938 674984 159944
rect 674852 159854 675064 159882
rect 674840 159792 674892 159798
rect 674840 159734 674892 159740
rect 674564 159588 674616 159594
rect 674564 159530 674616 159536
rect 674472 155304 674524 155310
rect 674472 155246 674524 155252
rect 674288 152244 674340 152250
rect 674288 152186 674340 152192
rect 673828 152176 673880 152182
rect 673828 152118 673880 152124
rect 673644 152108 673696 152114
rect 673644 152050 673696 152056
rect 673552 148504 673604 148510
rect 673552 148446 673604 148452
rect 674852 146146 674880 159734
rect 675036 155394 675064 159854
rect 675128 157350 675156 160482
rect 675116 157344 675168 157350
rect 675116 157286 675168 157292
rect 675220 156006 675248 168370
rect 675312 160290 675340 173159
rect 676048 172922 676076 173567
rect 676036 172916 676088 172922
rect 676036 172858 676088 172864
rect 676034 172816 676090 172825
rect 676034 172751 676090 172760
rect 675942 172408 675998 172417
rect 675942 172343 675998 172352
rect 675956 172106 675984 172343
rect 675944 172100 675996 172106
rect 675944 172042 675996 172048
rect 675942 172000 675998 172009
rect 675942 171935 675998 171944
rect 675956 171698 675984 171935
rect 675944 171692 675996 171698
rect 675944 171634 675996 171640
rect 675942 171592 675998 171601
rect 675942 171527 675998 171536
rect 675956 171222 675984 171527
rect 675944 171216 675996 171222
rect 675944 171158 675996 171164
rect 676048 171154 676076 172751
rect 676036 171148 676088 171154
rect 676036 171090 676088 171096
rect 676034 170776 676090 170785
rect 676034 170711 676090 170720
rect 675942 170368 675998 170377
rect 675942 170303 675998 170312
rect 675850 169960 675906 169969
rect 675850 169895 675906 169904
rect 675864 169250 675892 169895
rect 675956 169658 675984 170303
rect 675944 169652 675996 169658
rect 675944 169594 675996 169600
rect 675942 169552 675998 169561
rect 675942 169487 675998 169496
rect 675852 169244 675904 169250
rect 675852 169186 675904 169192
rect 675850 169144 675906 169153
rect 675850 169079 675906 169088
rect 675758 168736 675814 168745
rect 675758 168671 675814 168680
rect 675772 168638 675800 168671
rect 675760 168632 675812 168638
rect 675760 168574 675812 168580
rect 675864 168570 675892 169079
rect 675852 168564 675904 168570
rect 675852 168506 675904 168512
rect 675956 168502 675984 169487
rect 675944 168496 675996 168502
rect 675944 168438 675996 168444
rect 676048 168434 676076 170711
rect 676036 168428 676088 168434
rect 676036 168370 676088 168376
rect 676034 167104 676090 167113
rect 676034 167039 676036 167048
rect 676088 167039 676090 167048
rect 676036 167010 676088 167016
rect 675404 160546 675432 160888
rect 675392 160540 675444 160546
rect 675392 160482 675444 160488
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675300 160200 675352 160206
rect 675300 160142 675352 160148
rect 675312 157162 675340 160142
rect 675392 160064 675444 160070
rect 675392 160006 675444 160012
rect 675404 159664 675432 160006
rect 675484 159588 675536 159594
rect 675484 159530 675536 159536
rect 675496 159052 675524 159530
rect 675404 157162 675432 157216
rect 675312 157134 675432 157162
rect 675758 157040 675814 157049
rect 675758 156975 675814 156984
rect 675772 156643 675800 156975
rect 675220 155978 675418 156006
rect 675036 155366 675340 155394
rect 675116 155304 675168 155310
rect 675116 155246 675168 155252
rect 675312 155258 675340 155366
rect 675404 155258 675432 155380
rect 675128 152334 675156 155246
rect 675208 155236 675260 155242
rect 675312 155230 675432 155258
rect 675208 155178 675260 155184
rect 675220 152878 675248 155178
rect 675220 152850 675418 152878
rect 675128 152306 675418 152334
rect 675116 152244 675168 152250
rect 675116 152186 675168 152192
rect 675128 149849 675156 152186
rect 675208 152176 675260 152182
rect 675208 152118 675260 152124
rect 675220 151042 675248 152118
rect 675300 152108 675352 152114
rect 675300 152050 675352 152056
rect 675312 151689 675340 152050
rect 675312 151661 675418 151689
rect 675220 151014 675418 151042
rect 675128 149821 675418 149849
rect 675392 148504 675444 148510
rect 675392 148446 675444 148452
rect 675404 147968 675432 148446
rect 675312 146254 675432 146282
rect 675312 146146 675340 146254
rect 674852 146118 675340 146146
rect 675404 146132 675432 146254
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676126 133104 676182 133113
rect 676126 133039 676182 133048
rect 676034 132968 676090 132977
rect 676034 132903 676036 132912
rect 676088 132903 676090 132912
rect 676036 132874 676088 132880
rect 676140 132666 676168 133039
rect 676220 132796 676272 132802
rect 676220 132738 676272 132744
rect 676232 132705 676260 132738
rect 676218 132696 676274 132705
rect 676128 132660 676180 132666
rect 676218 132631 676274 132640
rect 676128 132602 676180 132608
rect 676220 132320 676272 132326
rect 676218 132288 676220 132297
rect 676272 132288 676274 132297
rect 676218 132223 676274 132232
rect 676034 131744 676090 131753
rect 676034 131679 676036 131688
rect 676088 131679 676090 131688
rect 676036 131650 676088 131656
rect 676220 131504 676272 131510
rect 676218 131472 676220 131481
rect 676272 131472 676274 131481
rect 676218 131407 676274 131416
rect 676034 130928 676090 130937
rect 676034 130863 676036 130872
rect 676088 130863 676090 130872
rect 676036 130834 676088 130840
rect 676220 130688 676272 130694
rect 676218 130656 676220 130665
rect 676272 130656 676274 130665
rect 676218 130591 676274 130600
rect 676034 130112 676090 130121
rect 676034 130047 676036 130056
rect 676088 130047 676090 130056
rect 676036 130018 676088 130024
rect 673368 129736 673420 129742
rect 676036 129736 676088 129742
rect 673368 129678 673420 129684
rect 676034 129704 676036 129713
rect 676088 129704 676090 129713
rect 676034 129639 676090 129648
rect 673092 129464 673144 129470
rect 676220 129464 676272 129470
rect 673092 129406 673144 129412
rect 676218 129432 676220 129441
rect 676272 129432 676274 129441
rect 676218 129367 676274 129376
rect 676034 128888 676090 128897
rect 676034 128823 676090 128832
rect 675942 128480 675998 128489
rect 675942 128415 675998 128424
rect 675574 128072 675630 128081
rect 675574 128007 675630 128016
rect 674656 127764 674708 127770
rect 674656 127706 674708 127712
rect 673552 127356 673604 127362
rect 673552 127298 673604 127304
rect 673294 123141 673322 123142
rect 673278 123132 673338 123141
rect 673278 123063 673338 123072
rect 672998 122904 673054 122913
rect 672998 122839 673054 122848
rect 672448 121644 672500 121650
rect 672448 121586 672500 121592
rect 672460 109313 672488 121586
rect 673294 112755 673322 123063
rect 673442 122739 673470 122740
rect 673426 122730 673486 122739
rect 673426 122661 673486 122670
rect 673284 112746 673340 112755
rect 673284 112681 673340 112690
rect 673442 110991 673470 122661
rect 673418 110982 673474 110991
rect 673418 110917 673474 110926
rect 672446 109304 672502 109313
rect 672446 109239 672502 109248
rect 673564 104582 673592 127298
rect 673828 127084 673880 127090
rect 673828 127026 673880 127032
rect 673644 124636 673696 124642
rect 673644 124578 673696 124584
rect 673656 105738 673684 124578
rect 673736 124364 673788 124370
rect 673736 124306 673788 124312
rect 673748 110090 673776 124306
rect 673736 110084 673788 110090
rect 673736 110026 673788 110032
rect 673840 108254 673868 127026
rect 674564 126132 674616 126138
rect 674564 126074 674616 126080
rect 674288 123684 674340 123690
rect 674288 123626 674340 123632
rect 673828 108248 673880 108254
rect 673828 108190 673880 108196
rect 674300 107574 674328 123626
rect 674576 111738 674604 126074
rect 674668 114374 674696 127706
rect 674748 127016 674800 127022
rect 674748 126958 674800 126964
rect 674656 114368 674708 114374
rect 674656 114310 674708 114316
rect 674760 113762 674788 126958
rect 675298 126440 675354 126449
rect 675298 126375 675354 126384
rect 674932 124500 674984 124506
rect 674932 124442 674984 124448
rect 674840 124296 674892 124302
rect 674840 124238 674892 124244
rect 674748 113756 674800 113762
rect 674748 113698 674800 113704
rect 674576 111710 674788 111738
rect 674288 107568 674340 107574
rect 674288 107510 674340 107516
rect 673644 105732 673696 105738
rect 673644 105674 673696 105680
rect 673552 104576 673604 104582
rect 673552 104518 673604 104524
rect 672354 102504 672410 102513
rect 672354 102439 672410 102448
rect 674760 100994 674788 111710
rect 674852 111178 674880 124238
rect 674944 111926 674972 124442
rect 675208 124228 675260 124234
rect 675208 124170 675260 124176
rect 675024 121508 675076 121514
rect 675024 121450 675076 121456
rect 675220 121454 675248 124170
rect 674932 111920 674984 111926
rect 674932 111862 674984 111868
rect 675036 111738 675064 121450
rect 674944 111710 675064 111738
rect 675128 121426 675248 121454
rect 674840 111172 674892 111178
rect 674840 111114 674892 111120
rect 674944 105822 674972 111710
rect 675128 110174 675156 121426
rect 675312 118402 675340 126375
rect 675220 118374 675340 118402
rect 675220 114493 675248 118374
rect 675588 118266 675616 128007
rect 675956 127362 675984 128415
rect 676048 127770 676076 128823
rect 676036 127764 676088 127770
rect 676036 127706 676088 127712
rect 676034 127664 676090 127673
rect 676034 127599 676090 127608
rect 675944 127356 675996 127362
rect 675944 127298 675996 127304
rect 675942 127256 675998 127265
rect 675942 127191 675998 127200
rect 675956 127090 675984 127191
rect 675944 127084 675996 127090
rect 675944 127026 675996 127032
rect 676048 127022 676076 127599
rect 676036 127016 676088 127022
rect 676036 126958 676088 126964
rect 676034 126848 676090 126857
rect 676034 126783 676090 126792
rect 676048 126138 676076 126783
rect 676036 126132 676088 126138
rect 676036 126074 676088 126080
rect 676034 126032 676090 126041
rect 676034 125967 676090 125976
rect 675942 125624 675998 125633
rect 675942 125559 675998 125568
rect 675956 124302 675984 125559
rect 676048 124506 676076 125967
rect 676126 124944 676182 124953
rect 676126 124879 676182 124888
rect 676140 124642 676168 124879
rect 676128 124636 676180 124642
rect 676128 124578 676180 124584
rect 676126 124536 676182 124545
rect 676036 124500 676088 124506
rect 676126 124471 676182 124480
rect 676036 124442 676088 124448
rect 676034 124400 676090 124409
rect 676140 124370 676168 124471
rect 676034 124335 676090 124344
rect 676128 124364 676180 124370
rect 675944 124296 675996 124302
rect 675944 124238 675996 124244
rect 676048 124234 676076 124335
rect 676128 124306 676180 124312
rect 676036 124228 676088 124234
rect 676036 124170 676088 124176
rect 676034 123992 676090 124001
rect 676034 123927 676090 123936
rect 676048 123690 676076 123927
rect 676036 123684 676088 123690
rect 676036 123626 676088 123632
rect 676034 123584 676090 123593
rect 676034 123519 676090 123528
rect 676048 121514 676076 123519
rect 676218 121680 676274 121689
rect 676218 121615 676220 121624
rect 676272 121615 676274 121624
rect 676220 121586 676272 121592
rect 676036 121508 676088 121514
rect 676036 121450 676088 121456
rect 675312 118238 675616 118266
rect 675312 115138 675340 118238
rect 675392 115932 675444 115938
rect 675392 115874 675444 115880
rect 675404 115668 675432 115874
rect 675312 115110 675418 115138
rect 675220 114465 675418 114493
rect 675208 114368 675260 114374
rect 675208 114310 675260 114316
rect 675220 113846 675248 114310
rect 675220 113818 675418 113846
rect 675208 113756 675260 113762
rect 675208 113698 675260 113704
rect 675220 112010 675248 113698
rect 675220 111982 675418 112010
rect 675208 111920 675260 111926
rect 675208 111862 675260 111868
rect 675220 111466 675248 111862
rect 675220 111438 675418 111466
rect 675392 111172 675444 111178
rect 675392 111114 675444 111120
rect 675404 110772 675432 111114
rect 675128 110146 675418 110174
rect 675116 110084 675168 110090
rect 675116 110026 675168 110032
rect 675128 106502 675156 110026
rect 675392 108248 675444 108254
rect 675392 108190 675444 108196
rect 675404 107644 675432 108190
rect 675392 107568 675444 107574
rect 675392 107510 675444 107516
rect 675404 107100 675432 107510
rect 675128 106474 675418 106502
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 674944 105794 675340 105822
rect 675404 105808 675432 105862
rect 675116 105732 675168 105738
rect 675116 105674 675168 105680
rect 675128 104666 675156 105674
rect 675128 104638 675340 104666
rect 675116 104576 675168 104582
rect 675116 104518 675168 104524
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675128 102830 675156 104518
rect 675312 104502 675432 104530
rect 675128 102802 675340 102830
rect 675312 102762 675340 102802
rect 675404 102762 675432 102816
rect 675312 102734 675432 102762
rect 674760 100966 675340 100994
rect 672078 100872 672134 100881
rect 675312 100858 675340 100966
rect 675404 100858 675432 100980
rect 675312 100830 675432 100858
rect 672078 100807 672134 100816
rect 666558 49056 666614 49065
rect 666558 48991 666614 49000
rect 661040 47388 661092 47394
rect 661040 47330 661092 47336
rect 650000 46980 650052 46986
rect 650000 46922 650052 46928
rect 661052 46912 661080 47330
rect 661052 46884 661500 46912
rect 610348 45824 610400 45830
rect 610348 45766 610400 45772
rect 661472 43110 661500 46884
rect 661460 43104 661512 43110
rect 661460 43046 661512 43052
rect 610256 41404 610308 41410
rect 610256 41346 610308 41352
rect 575756 41336 575808 41342
rect 543646 41304 543702 41313
rect 575756 41278 575808 41284
rect 543646 41239 543702 41248
rect 475568 38616 475620 38622
rect 475568 38558 475620 38564
rect 514024 38616 514076 38622
rect 514024 38558 514076 38564
rect 530492 38616 530544 38622
rect 530492 38558 530544 38564
rect 543004 38616 543056 38622
rect 543004 38558 543056 38564
<< via2 >>
rect 676034 897096 676090 897152
rect 676034 896688 676090 896744
rect 675942 894668 675998 894704
rect 675942 894648 675944 894668
rect 675944 894648 675996 894668
rect 675996 894648 675998 894668
rect 655426 867584 655482 867640
rect 655610 868808 655666 868864
rect 655518 866496 655574 866552
rect 655702 865272 655758 865328
rect 655794 863776 655850 863832
rect 656806 862552 656862 862608
rect 41786 817692 41842 817728
rect 41786 817672 41788 817692
rect 41788 817672 41840 817692
rect 41840 817672 41842 817692
rect 41786 817284 41842 817320
rect 41786 817264 41788 817284
rect 41788 817264 41840 817284
rect 41840 817264 41842 817284
rect 41786 816876 41842 816912
rect 41786 816856 41788 816876
rect 41788 816856 41840 816876
rect 41840 816856 41842 816876
rect 41786 816040 41842 816096
rect 41786 815224 41842 815280
rect 41786 814428 41842 814464
rect 41786 814408 41788 814428
rect 41788 814408 41840 814428
rect 41840 814408 41842 814428
rect 41786 813592 41842 813648
rect 41786 813184 41842 813240
rect 41786 812796 41842 812832
rect 41786 812776 41788 812796
rect 41788 812776 41840 812796
rect 41840 812776 41842 812796
rect 41786 812368 41842 812424
rect 41970 811552 42026 811608
rect 41786 810736 41842 810792
rect 41878 810328 41934 810384
rect 41786 809512 41842 809568
rect 41878 808696 41934 808752
rect 41786 808288 41842 808344
rect 41786 807880 41842 807936
rect 42246 811144 42302 811200
rect 42062 807472 42118 807528
rect 42062 806248 42118 806304
rect 42614 809920 42670 809976
rect 41878 794416 41934 794472
rect 41786 774444 41842 774480
rect 41786 774424 41788 774444
rect 41788 774424 41840 774444
rect 41840 774424 41842 774444
rect 41418 773900 41474 773936
rect 41418 773880 41420 773900
rect 41420 773880 41472 773900
rect 41472 773880 41474 773900
rect 41786 773628 41842 773664
rect 41786 773608 41788 773628
rect 41788 773608 41840 773628
rect 41840 773608 41842 773628
rect 41510 773472 41566 773528
rect 41878 772828 41880 772848
rect 41880 772828 41932 772848
rect 41932 772828 41934 772848
rect 41878 772792 41934 772828
rect 41510 772692 41512 772712
rect 41512 772692 41564 772712
rect 41564 772692 41566 772712
rect 41510 772656 41566 772692
rect 41510 771840 41566 771896
rect 41418 771044 41474 771080
rect 41418 771024 41420 771044
rect 41420 771024 41472 771044
rect 41472 771024 41474 771044
rect 41786 771568 41842 771624
rect 43718 811824 43774 811880
rect 41786 770752 41842 770808
rect 42154 770344 42210 770400
rect 41510 769800 41566 769856
rect 41510 769412 41566 769448
rect 41510 769392 41512 769412
rect 41512 769392 41564 769412
rect 41564 769392 41566 769412
rect 41510 769004 41566 769040
rect 41510 768984 41512 769004
rect 41512 768984 41564 769004
rect 41564 768984 41566 769004
rect 41510 768576 41566 768632
rect 41510 768188 41566 768224
rect 41510 768168 41512 768188
rect 41512 768168 41564 768188
rect 41564 768168 41566 768188
rect 41786 767896 41842 767952
rect 41510 767388 41512 767408
rect 41512 767388 41564 767408
rect 41564 767388 41566 767408
rect 41510 767352 41566 767388
rect 41694 766944 41750 767000
rect 41418 766536 41474 766592
rect 41510 766148 41566 766184
rect 41510 766128 41512 766148
rect 41512 766128 41564 766148
rect 41564 766128 41566 766148
rect 41510 765740 41566 765776
rect 41510 765720 41512 765740
rect 41512 765720 41564 765740
rect 41564 765720 41566 765740
rect 41602 765312 41658 765368
rect 41510 764924 41566 764960
rect 41510 764904 41512 764924
rect 41512 764904 41564 764924
rect 41564 764904 41566 764924
rect 41510 764532 41512 764552
rect 41512 764532 41564 764552
rect 41564 764532 41566 764552
rect 41510 764496 41566 764532
rect 41510 764088 41566 764144
rect 41510 762884 41566 762920
rect 41510 762864 41512 762884
rect 41512 762864 41564 762884
rect 41564 762864 41566 762884
rect 41786 757016 41842 757072
rect 42154 757016 42210 757072
rect 43074 752936 43130 752992
rect 42430 748720 42486 748776
rect 41510 731060 41566 731096
rect 41510 731040 41512 731060
rect 41512 731040 41564 731060
rect 41564 731040 41566 731060
rect 41510 730652 41566 730688
rect 41510 730632 41512 730652
rect 41512 730632 41564 730652
rect 41564 730632 41566 730652
rect 41510 730244 41566 730280
rect 41510 730224 41512 730244
rect 41512 730224 41564 730244
rect 41564 730224 41566 730244
rect 41510 729408 41566 729464
rect 41878 730088 41934 730144
rect 41786 729272 41842 729328
rect 42430 728864 42486 728920
rect 41510 728612 41566 728648
rect 41510 728592 41512 728612
rect 41512 728592 41564 728612
rect 41564 728592 41566 728612
rect 41786 728048 41842 728104
rect 41510 727776 41566 727832
rect 41510 726572 41566 726608
rect 41510 726552 41512 726572
rect 41512 726552 41564 726572
rect 41564 726552 41566 726572
rect 41970 727232 42026 727288
rect 41510 726164 41566 726200
rect 41510 726144 41512 726164
rect 41512 726144 41564 726164
rect 41564 726144 41566 726164
rect 41786 726028 41842 726064
rect 41786 726008 41788 726028
rect 41788 726008 41840 726028
rect 41840 726008 41842 726028
rect 41510 725328 41566 725384
rect 41786 725192 41842 725248
rect 41510 724104 41566 724160
rect 30286 723696 30342 723752
rect 41694 723288 41750 723344
rect 41510 722084 41566 722120
rect 41510 722064 41512 722084
rect 41512 722064 41564 722084
rect 41564 722064 41566 722084
rect 41510 721656 41566 721712
rect 41418 720840 41474 720896
rect 41602 721248 41658 721304
rect 41510 719636 41566 719672
rect 41510 719616 41512 719636
rect 41512 719616 41564 719636
rect 41564 719616 41566 719636
rect 41786 723172 41842 723208
rect 41786 723152 41788 723172
rect 41788 723152 41840 723172
rect 41840 723152 41842 723172
rect 41878 722744 41934 722800
rect 42246 724784 42302 724840
rect 42246 708872 42302 708928
rect 41786 688084 41842 688120
rect 41786 688064 41788 688084
rect 41788 688064 41840 688084
rect 41840 688064 41842 688084
rect 41786 687676 41842 687712
rect 41786 687656 41788 687676
rect 41788 687656 41840 687676
rect 41840 687656 41842 687676
rect 41786 687284 41788 687304
rect 41788 687284 41840 687304
rect 41840 687284 41842 687304
rect 41786 687248 41842 687284
rect 41786 686840 41842 686896
rect 41786 686432 41842 686488
rect 43074 714312 43130 714368
rect 43166 714176 43222 714232
rect 43442 711456 43498 711512
rect 42430 686024 42486 686080
rect 43718 709416 43774 709472
rect 43810 708464 43866 708520
rect 42062 685616 42118 685672
rect 41786 685208 41842 685264
rect 41786 684428 41788 684448
rect 41788 684428 41840 684448
rect 41840 684428 41842 684448
rect 41786 684392 41842 684428
rect 41786 683984 41842 684040
rect 41786 683576 41842 683632
rect 41694 682624 41750 682680
rect 41694 682236 41750 682272
rect 41694 682216 41696 682236
rect 41696 682216 41748 682236
rect 41748 682216 41750 682236
rect 30286 681944 30342 682000
rect 27434 680312 27490 680368
rect 27526 679088 27582 679144
rect 41786 681128 41842 681184
rect 41970 680720 42026 680776
rect 41786 679924 41842 679960
rect 41786 679904 41788 679924
rect 41788 679904 41840 679924
rect 41840 679904 41842 679924
rect 41694 679380 41750 679416
rect 41694 679360 41696 679380
rect 41696 679360 41748 679380
rect 41748 679360 41750 679380
rect 41786 678680 41842 678736
rect 41694 678136 41750 678192
rect 41694 676524 41750 676560
rect 41694 676504 41696 676524
rect 41696 676504 41748 676524
rect 41748 676504 41750 676524
rect 42430 684800 42486 684856
rect 42246 683168 42302 683224
rect 41970 670656 42026 670712
rect 42338 681536 42394 681592
rect 42430 670928 42486 670984
rect 43258 670656 43314 670712
rect 43074 665216 43130 665272
rect 43258 670520 43314 670576
rect 43442 671064 43498 671120
rect 41510 644700 41566 644736
rect 41510 644680 41512 644700
rect 41512 644680 41564 644700
rect 41564 644680 41566 644700
rect 41510 644292 41566 644328
rect 41510 644272 41512 644292
rect 41512 644272 41564 644292
rect 41564 644272 41566 644292
rect 41786 644088 41842 644124
rect 41786 644068 41788 644088
rect 41788 644068 41840 644088
rect 41840 644068 41842 644088
rect 41510 643864 41566 643920
rect 41786 643272 41842 643308
rect 41786 643252 41788 643272
rect 41788 643252 41840 643272
rect 41840 643252 41842 643272
rect 41510 643068 41566 643104
rect 41510 643048 41512 643068
rect 41512 643048 41564 643068
rect 41564 643048 41566 643068
rect 43626 670792 43682 670848
rect 43718 670520 43774 670576
rect 43902 670384 43958 670440
rect 44086 670656 44142 670712
rect 41602 642232 41658 642288
rect 41510 641416 41566 641472
rect 41510 640620 41566 640656
rect 41510 640600 41512 640620
rect 41512 640600 41564 640620
rect 41564 640600 41566 640620
rect 41786 642028 41842 642084
rect 41786 641620 41842 641676
rect 41786 640416 41842 640452
rect 41786 640396 41788 640416
rect 41788 640396 41840 640416
rect 41840 640396 41842 640416
rect 42338 639920 42394 639976
rect 41510 639376 41566 639432
rect 41510 638968 41566 639024
rect 41786 638764 41842 638820
rect 41786 638356 41842 638412
rect 41510 637764 41566 637800
rect 41510 637744 41512 637764
rect 41512 637744 41564 637764
rect 41564 637744 41566 637764
rect 38106 636928 38162 636984
rect 41510 636520 41566 636576
rect 38198 635704 38254 635760
rect 41602 636112 41658 636168
rect 41602 635296 41658 635352
rect 41602 634888 41658 634944
rect 41510 634480 41566 634536
rect 41510 633276 41566 633312
rect 41510 633256 41512 633276
rect 41512 633256 41564 633276
rect 41564 633256 41566 633276
rect 41694 631896 41750 631952
rect 41878 637540 41934 637596
rect 41786 627408 41842 627464
rect 42430 627408 42486 627464
rect 42062 621968 42118 622024
rect 41878 621424 41934 621480
rect 41786 601724 41842 601760
rect 41786 601704 41788 601724
rect 41788 601704 41840 601724
rect 41840 601704 41842 601724
rect 41786 601316 41842 601352
rect 41786 601296 41788 601316
rect 41788 601296 41840 601316
rect 41840 601296 41842 601316
rect 41786 600908 41842 600944
rect 41786 600888 41788 600908
rect 41788 600888 41840 600908
rect 41840 600888 41842 600908
rect 41510 600616 41566 600672
rect 41786 600072 41842 600128
rect 41510 599800 41566 599856
rect 41510 599004 41566 599040
rect 41510 598984 41512 599004
rect 41512 598984 41564 599004
rect 41564 598984 41566 599004
rect 41786 598884 41788 598904
rect 41788 598884 41840 598904
rect 41840 598884 41842 598904
rect 41786 598848 41842 598884
rect 42430 598440 42486 598496
rect 41510 598168 41566 598224
rect 41510 597352 41566 597408
rect 41510 596944 41566 597000
rect 41510 596536 41566 596592
rect 42154 596400 42210 596456
rect 41510 595720 41566 595776
rect 41510 595312 41566 595368
rect 41878 595176 41934 595232
rect 41510 594496 41566 594552
rect 38014 594088 38070 594144
rect 38106 593680 38162 593736
rect 41786 593564 41842 593600
rect 41786 593544 41788 593564
rect 41788 593544 41840 593564
rect 41840 593544 41842 593564
rect 41510 592864 41566 592920
rect 41694 592456 41750 592512
rect 41510 592048 41566 592104
rect 41510 591640 41566 591696
rect 41418 591232 41474 591288
rect 41510 590028 41566 590064
rect 41510 590008 41512 590028
rect 41512 590008 41564 590028
rect 41564 590008 41566 590028
rect 41786 584160 41842 584216
rect 42338 585248 42394 585304
rect 42706 583888 42762 583944
rect 42246 580624 42302 580680
rect 42154 576952 42210 577008
rect 43166 581848 43222 581904
rect 41510 558340 41566 558376
rect 41510 558320 41512 558340
rect 41512 558320 41564 558340
rect 41564 558320 41566 558340
rect 41510 557932 41566 557968
rect 41510 557912 41512 557932
rect 41512 557912 41564 557932
rect 41564 557912 41566 557932
rect 41510 557540 41512 557560
rect 41512 557540 41564 557560
rect 41564 557540 41566 557560
rect 41510 557504 41566 557540
rect 41786 557268 41788 557288
rect 41788 557268 41840 557288
rect 41840 557268 41842 557288
rect 41786 557232 41842 557268
rect 43902 632032 43958 632088
rect 43902 583752 43958 583808
rect 41786 556416 41842 556472
rect 41510 555872 41566 555928
rect 44086 583752 44142 583808
rect 38566 554648 38622 554704
rect 41510 553424 41566 553480
rect 41786 551928 41842 551984
rect 41510 550160 41566 550216
rect 41418 549772 41474 549808
rect 41418 549752 41420 549772
rect 41420 549752 41472 549772
rect 41472 549752 41474 549772
rect 41510 549364 41566 549400
rect 41510 549344 41512 549364
rect 41512 549344 41564 549364
rect 41564 549344 41566 549364
rect 41510 548936 41566 548992
rect 41510 548528 41566 548584
rect 41418 548120 41474 548176
rect 41510 546916 41566 546952
rect 41510 546896 41512 546916
rect 41512 546896 41564 546916
rect 41564 546896 41566 546916
rect 43074 538328 43130 538384
rect 42706 538056 42762 538112
rect 42246 535336 42302 535392
rect 42430 532752 42486 532808
rect 42338 532616 42394 532672
rect 43166 535336 43222 535392
rect 43074 532616 43130 532672
rect 43626 538464 43682 538520
rect 43718 538192 43774 538248
rect 41878 435920 41934 435976
rect 41786 430908 41842 430944
rect 41786 430888 41788 430908
rect 41788 430888 41840 430908
rect 41840 430888 41842 430908
rect 41786 430500 41842 430536
rect 41786 430480 41788 430500
rect 41788 430480 41840 430500
rect 41840 430480 41842 430500
rect 41786 430092 41842 430128
rect 41786 430072 41788 430092
rect 41788 430072 41840 430092
rect 41840 430072 41842 430092
rect 41786 429664 41842 429720
rect 41786 429256 41842 429312
rect 41786 428884 41788 428904
rect 41788 428884 41840 428904
rect 41840 428884 41842 428904
rect 41786 428848 41842 428884
rect 42430 428440 42486 428496
rect 42062 427624 42118 427680
rect 41878 427216 41934 427272
rect 41786 426808 41842 426864
rect 41786 426420 41842 426456
rect 41786 426400 41788 426420
rect 41788 426400 41840 426420
rect 41840 426400 41842 426420
rect 41970 425992 42026 426048
rect 41786 425584 41842 425640
rect 41786 425196 41842 425232
rect 41786 425176 41788 425196
rect 41788 425176 41840 425196
rect 41840 425176 41842 425196
rect 41786 424768 41842 424824
rect 41878 423952 41934 424008
rect 41878 423564 41934 423600
rect 41878 423544 41880 423564
rect 41880 423544 41932 423564
rect 41932 423544 41934 423564
rect 41878 423136 41934 423192
rect 41878 422728 41934 422784
rect 41786 422340 41842 422376
rect 41786 422320 41788 422340
rect 41788 422320 41840 422340
rect 41840 422320 41842 422340
rect 41786 421912 41842 421968
rect 41878 421504 41934 421560
rect 41786 420688 41842 420744
rect 41786 419484 41842 419520
rect 41786 419464 41788 419484
rect 41788 419464 41840 419484
rect 41840 419464 41842 419484
rect 42246 424360 42302 424416
rect 42338 421096 42394 421152
rect 43258 411440 43314 411496
rect 43166 406816 43222 406872
rect 41418 387524 41474 387560
rect 41418 387504 41420 387524
rect 41420 387504 41472 387524
rect 41472 387504 41474 387524
rect 41418 387116 41474 387152
rect 41418 387096 41420 387116
rect 41420 387096 41472 387116
rect 41472 387096 41474 387116
rect 41786 386844 41842 386880
rect 41786 386824 41788 386844
rect 41788 386824 41840 386844
rect 41840 386824 41842 386844
rect 41510 386688 41566 386744
rect 41510 385872 41566 385928
rect 41510 385056 41566 385112
rect 41510 384240 41566 384296
rect 42430 386008 42486 386064
rect 41878 385192 41934 385248
rect 41786 383968 41842 384024
rect 41510 383424 41566 383480
rect 41510 382608 41566 382664
rect 41510 381812 41566 381848
rect 41510 381792 41512 381812
rect 41512 381792 41564 381812
rect 41564 381792 41566 381812
rect 41510 381384 41566 381440
rect 42338 381112 42394 381168
rect 41970 380704 42026 380760
rect 41510 380180 41566 380216
rect 41510 380160 41512 380180
rect 41512 380160 41564 380180
rect 41564 380160 41566 380180
rect 41510 379752 41566 379808
rect 41510 379344 41566 379400
rect 41418 378956 41474 378992
rect 41418 378936 41420 378956
rect 41420 378936 41472 378956
rect 41472 378936 41474 378956
rect 41602 378528 41658 378584
rect 41510 378120 41566 378176
rect 41326 377712 41382 377768
rect 41418 377304 41474 377360
rect 41418 376100 41474 376136
rect 41418 376080 41420 376100
rect 41420 376080 41472 376100
rect 41472 376080 41474 376100
rect 41786 356904 41842 356960
rect 41786 355680 41842 355736
rect 41510 344276 41566 344312
rect 41510 344256 41512 344276
rect 41512 344256 41564 344276
rect 41564 344256 41566 344276
rect 41510 343868 41566 343904
rect 41510 343848 41512 343868
rect 41512 343848 41564 343868
rect 41564 343848 41566 343868
rect 41510 343460 41566 343496
rect 41510 343440 41512 343460
rect 41512 343440 41564 343460
rect 41564 343440 41566 343460
rect 41510 342644 41566 342680
rect 41510 342624 41512 342644
rect 41512 342624 41564 342644
rect 41564 342624 41566 342644
rect 41878 343304 41934 343360
rect 41786 342488 41842 342544
rect 41786 342080 41842 342136
rect 41510 341844 41512 341864
rect 41512 341844 41564 341864
rect 41564 341844 41566 341864
rect 41510 341808 41566 341844
rect 41786 341264 41842 341320
rect 41510 340992 41566 341048
rect 29918 339768 29974 339824
rect 33046 339768 33102 339824
rect 30102 338952 30158 339008
rect 30010 338544 30066 338600
rect 29918 329976 29974 330032
rect 30194 338136 30250 338192
rect 30102 330112 30158 330168
rect 30286 337728 30342 337784
rect 41510 336096 41566 336152
rect 41418 334872 41474 334928
rect 41786 335960 41842 336016
rect 41602 335280 41658 335336
rect 30010 329840 30066 329896
rect 41694 334464 41750 334520
rect 41878 334328 41934 334384
rect 41878 333124 41934 333160
rect 41878 333104 41880 333124
rect 41880 333104 41932 333124
rect 41932 333104 41934 333124
rect 42430 316376 42486 316432
rect 41786 316240 41842 316296
rect 42154 315424 42210 315480
rect 41970 313792 42026 313848
rect 41786 312976 41842 313032
rect 42154 312296 42210 312352
rect 41970 301280 42026 301336
rect 27526 300872 27582 300928
rect 41878 300464 41934 300520
rect 41786 300092 41788 300112
rect 41788 300092 41840 300112
rect 41840 300092 41842 300112
rect 41786 300056 41842 300092
rect 41786 299240 41842 299296
rect 41786 298424 41842 298480
rect 41786 298016 41842 298072
rect 41786 297200 41842 297256
rect 35806 296384 35862 296440
rect 41694 295024 41750 295080
rect 41786 294752 41842 294808
rect 42062 299648 42118 299704
rect 42430 298832 42486 298888
rect 42062 293936 42118 293992
rect 42062 293528 42118 293584
rect 42062 293120 42118 293176
rect 41878 292324 41934 292360
rect 41878 292304 41880 292324
rect 41880 292304 41932 292324
rect 41932 292304 41934 292324
rect 41786 291100 41842 291136
rect 41786 291080 41788 291100
rect 41788 291080 41840 291100
rect 41840 291080 41842 291100
rect 41786 290692 41842 290728
rect 41786 290672 41788 290692
rect 41788 290672 41840 290692
rect 41840 290672 41842 290692
rect 41786 289876 41842 289912
rect 41786 289856 41788 289876
rect 41788 289856 41840 289876
rect 41840 289856 41842 289876
rect 41970 291896 42026 291952
rect 42154 292712 42210 292768
rect 42706 291488 42762 291544
rect 41786 272312 41842 272368
rect 41786 270408 41842 270464
rect 41970 269728 42026 269784
rect 41786 269320 41842 269376
rect 41510 257896 41566 257952
rect 41602 257524 41604 257544
rect 41604 257524 41656 257544
rect 41656 257524 41658 257544
rect 41602 257488 41658 257524
rect 41878 257660 41880 257680
rect 41880 257660 41932 257680
rect 41932 257660 41934 257680
rect 41878 257624 41934 257660
rect 41786 256808 41842 256864
rect 41878 256400 41934 256456
rect 41510 256300 41512 256320
rect 41512 256300 41564 256320
rect 41564 256300 41566 256320
rect 41510 256264 41566 256300
rect 41510 255448 41566 255504
rect 41786 254768 41842 254824
rect 41510 254632 41566 254688
rect 41878 253988 41880 254008
rect 41880 253988 41932 254008
rect 41932 253988 41934 254008
rect 41878 253952 41934 253988
rect 42062 253544 42118 253600
rect 41694 253000 41750 253056
rect 41142 251368 41198 251424
rect 35806 250960 35862 251016
rect 38474 250552 38530 250608
rect 38566 250144 38622 250200
rect 41234 249736 41290 249792
rect 41602 248920 41658 248976
rect 41418 248512 41474 248568
rect 41326 248104 41382 248160
rect 41510 247716 41566 247752
rect 41510 247696 41512 247716
rect 41512 247696 41564 247716
rect 41564 247696 41566 247716
rect 41510 247308 41566 247344
rect 41510 247288 41512 247308
rect 41512 247288 41564 247308
rect 41564 247288 41566 247308
rect 41510 246492 41566 246528
rect 41510 246472 41512 246492
rect 41512 246472 41564 246492
rect 41564 246472 41566 246492
rect 41878 252728 41934 252784
rect 41786 251912 41842 251968
rect 41970 252320 42026 252376
rect 41970 242256 42026 242312
rect 42338 249464 42394 249520
rect 42062 242120 42118 242176
rect 42430 228792 42486 228848
rect 42430 228656 42486 228712
rect 42430 225664 42486 225720
rect 41510 215092 41512 215112
rect 41512 215092 41564 215112
rect 41564 215092 41566 215112
rect 41510 215056 41566 215092
rect 41510 214684 41512 214704
rect 41512 214684 41564 214704
rect 41564 214684 41566 214704
rect 41510 214648 41566 214684
rect 41510 214276 41512 214296
rect 41512 214276 41564 214296
rect 41564 214276 41566 214296
rect 41510 214240 41566 214276
rect 41510 213832 41566 213888
rect 41510 213444 41566 213480
rect 41510 213424 41512 213444
rect 41512 213424 41564 213444
rect 41564 213424 41566 213444
rect 33046 212608 33102 212664
rect 43534 238040 43590 238096
rect 41510 212236 41512 212256
rect 41512 212236 41564 212256
rect 41564 212236 41566 212256
rect 41510 212200 41566 212236
rect 58254 790880 58310 790936
rect 58530 789284 58532 789304
rect 58532 789284 58584 789304
rect 58584 789284 58586 789304
rect 58530 789248 58586 789284
rect 58162 788432 58218 788488
rect 58438 787344 58494 787400
rect 58530 786120 58586 786176
rect 58438 784896 58494 784952
rect 655426 778368 655482 778424
rect 654966 773472 655022 773528
rect 58438 747632 58494 747688
rect 59266 746408 59322 746464
rect 58438 744912 58494 744968
rect 58530 744096 58586 744152
rect 57978 742348 58034 742384
rect 57978 742328 57980 742348
rect 57980 742328 58032 742348
rect 58032 742328 58034 742348
rect 58438 741784 58494 741840
rect 654322 730224 654378 730280
rect 655794 777008 655850 777064
rect 655610 775920 655666 775976
rect 655518 775512 655574 775568
rect 655518 734304 655574 734360
rect 59358 704384 59414 704440
rect 59266 703296 59322 703352
rect 58530 702072 58586 702128
rect 58254 700712 58310 700768
rect 58530 699624 58586 699680
rect 58530 698128 58586 698184
rect 655426 687248 655482 687304
rect 654230 685752 654286 685808
rect 654138 684392 654194 684448
rect 60646 661136 60702 661192
rect 58530 659504 58586 659560
rect 58438 658824 58494 658880
rect 58622 657600 58678 657656
rect 58438 656512 58494 656568
rect 58070 655288 58126 655344
rect 654414 639376 654470 639432
rect 58162 617752 58218 617808
rect 655702 731448 655758 731504
rect 655610 688200 655666 688256
rect 655518 643184 655574 643240
rect 58530 616800 58586 616856
rect 58530 615476 58532 615496
rect 58532 615476 58584 615496
rect 58584 615476 58586 615496
rect 58530 615440 58586 615476
rect 58162 614488 58218 614544
rect 58530 612620 58532 612640
rect 58532 612620 58584 612640
rect 58584 612620 58586 612640
rect 58530 612584 58586 612620
rect 58346 612040 58402 612096
rect 655426 595312 655482 595368
rect 655242 594224 655298 594280
rect 58530 574776 58586 574832
rect 656530 774696 656586 774752
rect 655886 732672 655942 732728
rect 655794 689424 655850 689480
rect 655702 640192 655758 640248
rect 655978 731312 656034 731368
rect 656070 728592 656126 728648
rect 655978 686976 656034 687032
rect 655886 641824 655942 641880
rect 655702 596536 655758 596592
rect 655610 593000 655666 593056
rect 59266 573552 59322 573608
rect 60646 572328 60702 572384
rect 58070 570968 58126 571024
rect 58346 570016 58402 570072
rect 58254 568248 58310 568304
rect 655426 553288 655482 553344
rect 654230 549208 654286 549264
rect 654138 548528 654194 548584
rect 59450 531664 59506 531720
rect 59266 530576 59322 530632
rect 58530 529352 58586 529408
rect 58346 528128 58402 528184
rect 57978 526904 58034 526960
rect 58070 525816 58126 525872
rect 655610 552064 655666 552120
rect 655518 550976 655574 551032
rect 655794 595448 655850 595504
rect 656070 640600 656126 640656
rect 655978 597760 656034 597816
rect 655886 550840 655942 550896
rect 656438 638152 656494 638208
rect 58438 404096 58494 404152
rect 58530 402908 58532 402928
rect 58532 402908 58584 402928
rect 58584 402908 58586 402928
rect 58530 402872 58586 402908
rect 60370 400696 60426 400752
rect 58438 400016 58494 400072
rect 58530 399336 58586 399392
rect 58346 398248 58402 398304
rect 655518 374448 655574 374504
rect 655702 373224 655758 373280
rect 655426 372136 655482 372192
rect 654506 370912 654562 370968
rect 58162 360848 58218 360904
rect 58530 359760 58586 359816
rect 57978 357448 58034 357504
rect 58530 357312 58586 357368
rect 58530 355816 58586 355872
rect 58438 355000 58494 355056
rect 32954 211792 33010 211848
rect 41510 211384 41566 211440
rect 32862 210976 32918 211032
rect 30010 210160 30066 210216
rect 25134 204856 25190 204912
rect 24950 204448 25006 204504
rect 24858 203632 24914 203688
rect 30194 209752 30250 209808
rect 30102 209344 30158 209400
rect 41510 208936 41566 208992
rect 38014 208528 38070 208584
rect 30286 208120 30342 208176
rect 38106 207712 38162 207768
rect 41510 207324 41566 207360
rect 41510 207304 41512 207324
rect 41512 207304 41564 207324
rect 41564 207304 41566 207324
rect 41786 207188 41842 207224
rect 41786 207168 41788 207188
rect 41788 207168 41840 207188
rect 41840 207168 41842 207188
rect 41418 206488 41474 206544
rect 41694 206080 41750 206136
rect 41602 205264 41658 205320
rect 41510 204856 41566 204912
rect 38106 201320 38162 201376
rect 30102 200232 30158 200288
rect 30010 200096 30066 200152
rect 41786 205944 41842 206000
rect 41878 184184 41934 184240
rect 41786 183368 41842 183424
rect 41786 182960 41842 183016
rect 655518 329840 655574 329896
rect 655426 328208 655482 328264
rect 655610 327392 655666 327448
rect 655978 325624 656034 325680
rect 58530 317328 58586 317384
rect 58070 316512 58126 316568
rect 58346 314744 58402 314800
rect 58162 312976 58218 313032
rect 58530 314064 58586 314120
rect 58530 311788 58532 311808
rect 58532 311788 58584 311808
rect 58584 311788 58586 311808
rect 58530 311752 58586 311788
rect 655518 303320 655574 303376
rect 655702 302096 655758 302152
rect 655426 300736 655482 300792
rect 655058 298696 655114 298752
rect 656070 297472 656126 297528
rect 655886 296248 655942 296304
rect 58530 295432 58586 295488
rect 58438 293936 58494 293992
rect 655702 293936 655758 293992
rect 59266 292712 59322 292768
rect 655518 292712 655574 292768
rect 58530 292304 58586 292360
rect 57978 291488 58034 291544
rect 57978 289756 57980 289776
rect 57980 289756 58032 289776
rect 58032 289756 58034 289776
rect 57978 289720 58034 289756
rect 58162 287952 58218 288008
rect 58530 287136 58586 287192
rect 57978 285640 58034 285696
rect 58530 284416 58586 284472
rect 58530 283192 58586 283248
rect 58254 282104 58310 282160
rect 58162 280880 58218 280936
rect 58254 279656 58310 279712
rect 654506 289176 654562 289232
rect 654874 287952 654930 288008
rect 655426 285640 655482 285696
rect 654874 284708 654930 284744
rect 654874 284688 654876 284708
rect 654876 284688 654928 284708
rect 654928 284688 654930 284708
rect 655426 283192 655482 283248
rect 654690 280880 654746 280936
rect 654874 279928 654930 279984
rect 69386 271768 69442 271824
rect 70582 269048 70638 269104
rect 81254 272176 81310 272232
rect 80058 272040 80114 272096
rect 78862 269320 78918 269376
rect 84750 272312 84806 272368
rect 83646 271904 83702 271960
rect 85946 269592 86002 269648
rect 90730 272448 90786 272504
rect 87142 269456 87198 269512
rect 93030 269728 93086 269784
rect 95422 272584 95478 272640
rect 99010 269864 99066 269920
rect 104898 272856 104954 272912
rect 103702 272720 103758 272776
rect 110786 273128 110842 273184
rect 109590 272992 109646 273048
rect 108394 270272 108450 270328
rect 107198 270136 107254 270192
rect 106094 270000 106150 270056
rect 76470 269184 76526 269240
rect 114374 270408 114430 270464
rect 120262 271632 120318 271688
rect 121458 268912 121514 268968
rect 124954 271496 125010 271552
rect 132038 271224 132094 271280
rect 134430 271360 134486 271416
rect 133234 271088 133290 271144
rect 184938 268776 184994 268832
rect 193678 271768 193734 271824
rect 194138 269048 194194 269104
rect 196898 272040 196954 272096
rect 195978 269184 196034 269240
rect 198094 272176 198150 272232
rect 197726 269320 197782 269376
rect 199106 272312 199162 272368
rect 198738 269320 198794 269376
rect 199382 271904 199438 271960
rect 199934 269592 199990 269648
rect 200394 269456 200450 269512
rect 201222 268776 201278 268832
rect 201958 272448 202014 272504
rect 203522 272584 203578 272640
rect 203062 269728 203118 269784
rect 206466 272856 206522 272912
rect 204810 269864 204866 269920
rect 204350 269320 204406 269376
rect 206742 272992 206798 273048
rect 207386 272720 207442 272776
rect 207478 270000 207534 270056
rect 207938 270272 207994 270328
rect 208398 270136 208454 270192
rect 209410 273128 209466 273184
rect 212354 271632 212410 271688
rect 210698 270408 210754 270464
rect 215022 271496 215078 271552
rect 213734 268912 213790 268968
rect 217690 271224 217746 271280
rect 217322 271088 217378 271144
rect 218150 271360 218206 271416
rect 355322 271088 355378 271144
rect 356610 268640 356666 268696
rect 357530 271224 357586 271280
rect 357990 271360 358046 271416
rect 359370 268776 359426 268832
rect 360658 271496 360714 271552
rect 362038 268912 362094 268968
rect 363326 271632 363382 271688
rect 364246 270408 364302 270464
rect 365994 273128 366050 273184
rect 365534 272992 365590 273048
rect 366914 270272 366970 270328
rect 368662 272856 368718 272912
rect 370870 272720 370926 272776
rect 369582 270136 369638 270192
rect 371330 272584 371386 272640
rect 373998 272448 374054 272504
rect 372250 270000 372306 270056
rect 380714 269864 380770 269920
rect 385590 274080 385646 274136
rect 383382 269728 383438 269784
rect 388258 274216 388314 274272
rect 387430 272312 387486 272368
rect 386970 267008 387026 267064
rect 387798 267144 387854 267200
rect 389638 266872 389694 266928
rect 391018 274352 391074 274408
rect 390466 266736 390522 266792
rect 391846 266600 391902 266656
rect 393134 266464 393190 266520
rect 394974 275848 395030 275904
rect 393594 267280 393650 267336
rect 394514 266328 394570 266384
rect 395434 272176 395490 272232
rect 396262 267416 396318 267472
rect 397366 275712 397422 275768
rect 398470 275576 398526 275632
rect 399850 275168 399906 275224
rect 399390 269592 399446 269648
rect 398930 267552 398986 267608
rect 400402 275440 400458 275496
rect 401138 275304 401194 275360
rect 402610 275032 402666 275088
rect 403438 272040 403494 272096
rect 403990 274896 404046 274952
rect 405186 274760 405242 274816
rect 404726 269456 404782 269512
rect 405462 267688 405518 267744
rect 406934 274624 406990 274680
rect 408130 274488 408186 274544
rect 407394 269320 407450 269376
rect 408774 271904 408830 271960
rect 408314 266192 408370 266248
rect 410522 271768 410578 271824
rect 410798 269184 410854 269240
rect 411902 269048 411958 269104
rect 436098 266192 436154 266248
rect 477314 267688 477370 267744
rect 471978 267552 472034 267608
rect 485686 267416 485742 267472
rect 498474 271088 498530 271144
rect 497922 267280 497978 267336
rect 505558 271360 505614 271416
rect 504362 271224 504418 271280
rect 509054 268776 509110 268832
rect 501970 268640 502026 268696
rect 512642 271496 512698 271552
rect 516230 268912 516286 268968
rect 519726 271632 519782 271688
rect 522118 270408 522174 270464
rect 526810 273128 526866 273184
rect 525614 272992 525670 273048
rect 529202 270272 529258 270328
rect 533894 272856 533950 272912
rect 536286 270136 536342 270192
rect 539874 272720 539930 272776
rect 540978 272584 541034 272640
rect 543370 270000 543426 270056
rect 548062 272448 548118 272504
rect 565818 269864 565874 269920
rect 572902 269728 572958 269784
rect 578882 274080 578938 274136
rect 583574 272312 583630 272368
rect 585966 274216 586022 274272
rect 584770 267144 584826 267200
rect 582378 267008 582434 267064
rect 589462 266872 589518 266928
rect 593050 274352 593106 274408
rect 591854 266736 591910 266792
rect 595350 266600 595406 266656
rect 598938 266464 598994 266520
rect 603630 275848 603686 275904
rect 604826 272176 604882 272232
rect 602434 266328 602490 266384
rect 609610 275712 609666 275768
rect 613106 275576 613162 275632
rect 617798 275440 617854 275496
rect 616694 275168 616750 275224
rect 620190 275304 620246 275360
rect 615498 269592 615554 269648
rect 623778 275032 623834 275088
rect 627274 274896 627330 274952
rect 626078 272040 626134 272096
rect 630862 274760 630918 274816
rect 635554 274624 635610 274680
rect 629666 269456 629722 269512
rect 637946 274488 638002 274544
rect 640338 271904 640394 271960
rect 636750 269320 636806 269376
rect 645030 271768 645086 271824
rect 646226 269184 646282 269240
rect 648618 269048 648674 269104
rect 573044 262260 573104 262320
rect 572218 259124 572278 259184
rect 184938 258576 184994 258632
rect 571394 255852 571454 255912
rect 416778 252728 416834 252784
rect 416778 249464 416834 249520
rect 187606 247968 187662 248024
rect 62762 227840 62818 227896
rect 57610 227704 57666 227760
rect 56046 227568 56102 227624
rect 55126 224848 55182 224904
rect 54390 222128 54446 222184
rect 56874 224984 56930 225040
rect 61106 222264 61162 222320
rect 63406 225120 63462 225176
rect 93030 228928 93086 228984
rect 84658 228792 84714 228848
rect 82726 228384 82782 228440
rect 76286 228248 76342 228304
rect 69478 228112 69534 228168
rect 66994 225256 67050 225312
rect 66166 222400 66222 222456
rect 67822 222536 67878 222592
rect 71226 227976 71282 228032
rect 70398 225392 70454 225448
rect 74446 222672 74502 222728
rect 77114 225528 77170 225584
rect 80426 225664 80482 225720
rect 79598 222808 79654 222864
rect 81254 222944 81310 223000
rect 83830 225800 83886 225856
rect 88062 228656 88118 228712
rect 86314 228520 86370 228576
rect 92202 225936 92258 225992
rect 89718 223080 89774 223136
rect 94778 227432 94834 227488
rect 99838 227296 99894 227352
rect 98918 226208 98974 226264
rect 97262 226072 97318 226128
rect 96434 223216 96490 223272
rect 98090 223352 98146 223408
rect 101494 227160 101550 227216
rect 106554 227024 106610 227080
rect 102046 224712 102102 224768
rect 103150 221992 103206 222048
rect 104806 223488 104862 223544
rect 113086 226888 113142 226944
rect 109038 224576 109094 224632
rect 110694 224440 110750 224496
rect 109866 221856 109922 221912
rect 112442 224168 112498 224224
rect 111614 221720 111670 221776
rect 114926 226752 114982 226808
rect 115754 224304 115810 224360
rect 118330 221584 118386 221640
rect 120814 224032 120870 224088
rect 121366 221448 121422 221504
rect 184938 237396 184940 237416
rect 184940 237396 184992 237416
rect 184992 237396 184994 237416
rect 184938 237360 184994 237396
rect 416778 246336 416834 246392
rect 418066 243072 418122 243128
rect 192574 224848 192630 224904
rect 193678 224984 193734 225040
rect 193310 222128 193366 222184
rect 194782 227704 194838 227760
rect 194414 227568 194470 227624
rect 197266 227840 197322 227896
rect 196530 225120 196586 225176
rect 196162 222264 196218 222320
rect 198002 225256 198058 225312
rect 198738 222536 198794 222592
rect 198646 222400 198702 222456
rect 200118 228112 200174 228168
rect 200486 227976 200542 228032
rect 199382 225392 199438 225448
rect 202970 228248 203026 228304
rect 202234 225528 202290 225584
rect 201866 222672 201922 222728
rect 203706 225664 203762 225720
rect 205086 225800 205142 225856
rect 204718 222944 204774 223000
rect 204442 222808 204498 222864
rect 206190 228792 206246 228848
rect 205822 228384 205878 228440
rect 207570 228656 207626 228712
rect 207202 228520 207258 228576
rect 208306 225936 208362 225992
rect 208674 223080 208730 223136
rect 210054 228928 210110 228984
rect 210698 227568 210754 227624
rect 210422 227432 210478 227488
rect 211158 226208 211214 226264
rect 210790 226072 210846 226128
rect 211526 223216 211582 223272
rect 212354 227704 212410 227760
rect 211894 223352 211950 223408
rect 212906 227296 212962 227352
rect 213274 227160 213330 227216
rect 212538 224712 212594 224768
rect 214746 223488 214802 223544
rect 214378 221992 214434 222048
rect 215758 227024 215814 227080
rect 215390 224576 215446 224632
rect 216494 224440 216550 224496
rect 216862 224168 216918 224224
rect 217230 221856 217286 221912
rect 217598 227840 217654 227896
rect 217322 221720 217378 221776
rect 218610 226888 218666 226944
rect 219254 228112 219310 228168
rect 218978 226752 219034 226808
rect 218242 224304 218298 224360
rect 220726 227976 220782 228032
rect 220450 221584 220506 221640
rect 220818 224032 220874 224088
rect 222106 223524 222108 223544
rect 222108 223524 222160 223544
rect 222160 223524 222162 223544
rect 222106 223488 222162 223524
rect 221830 221448 221886 221504
rect 225970 228248 226026 228304
rect 227810 223488 227866 223544
rect 234802 228520 234858 228576
rect 234618 228384 234674 228440
rect 245842 228792 245898 228848
rect 256698 228928 256754 228984
rect 259642 228520 259698 228576
rect 260378 227704 260434 227760
rect 260010 227568 260066 227624
rect 261758 228928 261814 228984
rect 261390 228792 261446 228848
rect 262494 228384 262550 228440
rect 263230 228112 263286 228168
rect 262862 227840 262918 227896
rect 264242 227976 264298 228032
rect 266082 228248 266138 228304
rect 330942 222944 330998 223000
rect 332322 222536 332378 222592
rect 333058 222808 333114 222864
rect 333794 222400 333850 222456
rect 334530 222672 334586 222728
rect 335910 222264 335966 222320
rect 335818 221856 335874 221912
rect 338762 222128 338818 222184
rect 369398 224576 369454 224632
rect 372250 224712 372306 224768
rect 370870 224440 370926 224496
rect 372618 224304 372674 224360
rect 373722 226208 373778 226264
rect 375838 221992 375894 222048
rect 376942 227296 376998 227352
rect 377310 227160 377366 227216
rect 378322 223488 378378 223544
rect 378690 223352 378746 223408
rect 380162 227432 380218 227488
rect 381174 223216 381230 223272
rect 381542 223080 381598 223136
rect 381082 222944 381138 223000
rect 382646 227024 382702 227080
rect 383658 222808 383714 222864
rect 383934 222944 383990 223000
rect 384762 228928 384818 228984
rect 384302 222536 384358 222592
rect 385866 222808 385922 222864
rect 386878 228792 386934 228848
rect 386786 222672 386842 222728
rect 387982 222672 388038 222728
rect 388994 222536 389050 222592
rect 387706 222400 387762 222456
rect 388534 221856 388590 221912
rect 390098 228656 390154 228712
rect 390466 225936 390522 225992
rect 390190 222264 390246 222320
rect 392214 228520 392270 228576
rect 391570 225664 391626 225720
rect 391202 222400 391258 222456
rect 391754 221856 391810 221912
rect 392582 225800 392638 225856
rect 394422 228384 394478 228440
rect 393686 225528 393742 225584
rect 393318 222264 393374 222320
rect 394790 225392 394846 225448
rect 396538 228248 396594 228304
rect 396906 222128 396962 222184
rect 398654 228112 398710 228168
rect 397918 225256 397974 225312
rect 399758 227976 399814 228032
rect 397642 222128 397698 222184
rect 401138 225120 401194 225176
rect 403990 227840 404046 227896
rect 407578 224984 407634 225040
rect 410062 227704 410118 227760
rect 411166 227568 411222 227624
rect 410798 224848 410854 224904
rect 411166 226072 411222 226128
rect 418158 239944 418214 240000
rect 418434 236680 418490 236736
rect 418526 233552 418582 233608
rect 471978 224576 472034 224632
rect 480258 227024 480314 227080
rect 481914 226208 481970 226264
rect 478510 224712 478566 224768
rect 475106 224440 475162 224496
rect 476026 224304 476082 224360
rect 507398 228928 507454 228984
rect 488906 227296 488962 227352
rect 488446 227160 488502 227216
rect 486330 221992 486386 222048
rect 488906 221176 488962 221232
rect 491942 223488 491998 223544
rect 492770 223352 492826 223408
rect 496174 227432 496230 227488
rect 495622 221856 495678 221912
rect 499302 223216 499358 223272
rect 496174 220904 496230 220960
rect 500222 223080 500278 223136
rect 500222 221040 500278 221096
rect 504822 222944 504878 223000
rect 512182 228792 512238 228848
rect 509606 222808 509662 222864
rect 513378 222672 513434 222728
rect 518990 228656 519046 228712
rect 518622 226072 518678 226128
rect 517242 222536 517298 222592
rect 525062 228520 525118 228576
rect 520830 225936 520886 225992
rect 523406 225664 523462 225720
rect 522210 222400 522266 222456
rect 530122 228384 530178 228440
rect 525798 225800 525854 225856
rect 528098 225528 528154 225584
rect 527270 222264 527326 222320
rect 534906 228248 534962 228304
rect 530674 225392 530730 225448
rect 538310 228112 538366 228168
rect 537390 222128 537446 222184
rect 542726 227976 542782 228032
rect 539322 225256 539378 225312
rect 545762 225120 545818 225176
rect 552570 227840 552626 227896
rect 561218 224984 561274 225040
rect 564346 221448 564402 221504
rect 566830 227704 566886 227760
rect 567290 222128 567346 222184
rect 567106 221720 567162 221776
rect 569314 227568 569370 227624
rect 568578 224848 568634 224904
rect 574374 222128 574430 222184
rect 573546 221448 573602 221504
rect 575202 221720 575258 221776
rect 582286 216144 582342 216200
rect 580446 214648 580502 214704
rect 580170 213152 580226 213208
rect 580078 211656 580134 211712
rect 579802 208664 579858 208720
rect 580630 204176 580686 204232
rect 580722 198192 580778 198248
rect 579802 183096 579858 183152
rect 580170 180104 580226 180160
rect 580538 178608 580594 178664
rect 580262 177112 580318 177168
rect 580814 175616 580870 175672
rect 580538 174120 580594 174176
rect 580262 163512 580318 163568
rect 579894 162016 579950 162072
rect 579802 159024 579858 159080
rect 579710 157528 579766 157584
rect 580446 137944 580502 138000
rect 579894 110880 579950 110936
rect 579986 106392 580042 106448
rect 579802 104896 579858 104952
rect 580078 100272 580134 100328
rect 184938 51040 184994 51096
rect 339406 52400 339462 52456
rect 346950 52400 347006 52456
rect 216126 48184 216182 48240
rect 194322 41792 194378 41848
rect 307298 41792 307354 41848
rect 361946 41792 362002 41848
rect 470138 43152 470194 43208
rect 415490 41792 415546 41848
rect 416778 41792 416834 41848
rect 419814 41792 419870 41848
rect 471702 41792 471758 41848
rect 223578 41248 223634 41304
rect 390190 41248 390246 41304
rect 475474 40976 475530 41032
rect 521750 42064 521806 42120
rect 513194 41656 513250 41712
rect 520370 41792 520426 41848
rect 530306 41112 530362 41168
rect 530398 40976 530454 41032
rect 580262 94288 580318 94344
rect 580170 92792 580226 92848
rect 580722 136448 580778 136504
rect 580630 133456 580686 133512
rect 582286 210160 582342 210216
rect 598938 207440 598994 207496
rect 582286 207168 582342 207224
rect 581458 205672 581514 205728
rect 599858 209480 599914 209536
rect 599950 208528 600006 208584
rect 599122 205400 599178 205456
rect 601146 206488 601202 206544
rect 600962 204448 601018 204504
rect 582286 202680 582342 202736
rect 601514 203360 601570 203416
rect 599950 202408 600006 202464
rect 598938 201320 598994 201376
rect 582286 201184 582342 201240
rect 599950 200368 600006 200424
rect 581090 199688 581146 199744
rect 599950 199280 600006 199336
rect 599122 198328 599178 198384
rect 599306 197240 599362 197296
rect 582286 196696 582342 196752
rect 599950 196288 600006 196344
rect 582286 195200 582342 195256
rect 599950 195200 600006 195256
rect 599122 194248 599178 194304
rect 582194 193568 582250 193624
rect 599950 193160 600006 193216
rect 599122 192208 599178 192264
rect 582286 192072 582342 192128
rect 599858 191120 599914 191176
rect 582194 190576 582250 190632
rect 600962 190168 601018 190224
rect 581366 189080 581422 189136
rect 582286 187604 582342 187640
rect 601606 189080 601662 189136
rect 601514 188128 601570 188184
rect 582286 187584 582288 187604
rect 582288 187584 582340 187604
rect 582340 187584 582342 187604
rect 599950 187040 600006 187096
rect 582194 186088 582250 186144
rect 599858 185000 599914 185056
rect 582286 184592 582342 184648
rect 599766 184048 599822 184104
rect 582286 181600 582342 181656
rect 599674 179968 599730 180024
rect 598938 176840 598994 176896
rect 600042 186088 600098 186144
rect 599950 182960 600006 183016
rect 599858 180920 599914 180976
rect 599766 177928 599822 177984
rect 582286 172624 582342 172680
rect 581274 168000 581330 168056
rect 581458 166504 581514 166560
rect 580998 165008 581054 165064
rect 580906 146920 580962 146976
rect 580998 143928 581054 143984
rect 581090 140936 581146 140992
rect 580814 131960 580870 132016
rect 580538 127472 580594 127528
rect 580446 101904 580502 101960
rect 580354 91296 580410 91352
rect 580630 98776 580686 98832
rect 580722 89800 580778 89856
rect 580538 88304 580594 88360
rect 580998 113872 581054 113928
rect 581274 145424 581330 145480
rect 581182 134952 581238 135008
rect 581090 109384 581146 109440
rect 580906 103400 580962 103456
rect 580814 86808 580870 86864
rect 579986 82320 580042 82376
rect 579618 80824 579674 80880
rect 568578 41384 568634 41440
rect 579618 59744 579674 59800
rect 579618 58284 579620 58304
rect 579620 58284 579672 58304
rect 579672 58284 579674 58304
rect 579618 58248 579674 58284
rect 580722 61240 580778 61296
rect 580814 56752 580870 56808
rect 580630 55256 580686 55312
rect 580998 65728 581054 65784
rect 581458 148552 581514 148608
rect 581366 139440 581422 139496
rect 581274 115368 581330 115424
rect 581182 97280 581238 97336
rect 581090 62736 581146 62792
rect 580906 53760 580962 53816
rect 581734 156032 581790 156088
rect 582194 171128 582250 171184
rect 600134 182008 600190 182064
rect 600042 178880 600098 178936
rect 599950 174800 600006 174856
rect 600318 175888 600374 175944
rect 600134 173848 600190 173904
rect 599858 172760 599914 172816
rect 599950 171808 600006 171864
rect 599950 170720 600006 170776
rect 599858 169768 599914 169824
rect 582286 169496 582342 169552
rect 599030 168680 599086 168736
rect 599858 167728 599914 167784
rect 600042 166640 600098 166696
rect 582010 160520 582066 160576
rect 581918 153040 581974 153096
rect 581826 151544 581882 151600
rect 599950 165688 600006 165744
rect 599858 164600 599914 164656
rect 599950 163648 600006 163704
rect 599858 162560 599914 162616
rect 599306 160520 599362 160576
rect 599950 161608 600006 161664
rect 600042 159568 600098 159624
rect 599950 158480 600006 158536
rect 599858 157528 599914 157584
rect 599858 156440 599914 156496
rect 599950 155488 600006 155544
rect 582286 154536 582342 154592
rect 599858 154400 599914 154456
rect 599306 152360 599362 152416
rect 582102 150048 582158 150104
rect 581550 142432 581606 142488
rect 581458 118360 581514 118416
rect 581642 122848 581698 122904
rect 581826 125976 581882 126032
rect 581734 119856 581790 119912
rect 582010 124480 582066 124536
rect 581918 116864 581974 116920
rect 581550 112376 581606 112432
rect 581366 107888 581422 107944
rect 581274 70216 581330 70272
rect 581458 71712 581514 71768
rect 581826 77832 581882 77888
rect 581734 76200 581790 76256
rect 599950 153448 600006 153504
rect 598938 151408 598994 151464
rect 599766 150320 599822 150376
rect 599950 149368 600006 149424
rect 582194 130464 582250 130520
rect 599858 148280 599914 148336
rect 599950 147328 600006 147384
rect 600042 146240 600098 146296
rect 599858 145288 599914 145344
rect 599950 144200 600006 144256
rect 599858 143248 599914 143304
rect 599306 141208 599362 141264
rect 599950 142160 600006 142216
rect 599858 140120 599914 140176
rect 600042 139168 600098 139224
rect 599950 138100 600006 138136
rect 599950 138080 599952 138100
rect 599952 138080 600004 138100
rect 600004 138080 600006 138100
rect 599858 137128 599914 137184
rect 599950 136040 600006 136096
rect 600042 135088 600098 135144
rect 599858 134000 599914 134056
rect 599950 133048 600006 133104
rect 598938 131960 598994 132016
rect 599766 131008 599822 131064
rect 599950 129940 600006 129976
rect 599950 129920 599952 129940
rect 599952 129920 600004 129940
rect 600004 129920 600006 129940
rect 582286 128968 582342 129024
rect 599858 128968 599914 129024
rect 599950 127880 600006 127936
rect 582102 121352 582158 121408
rect 582010 85312 582066 85368
rect 600042 126928 600098 126984
rect 599858 125840 599914 125896
rect 599950 124888 600006 124944
rect 599858 123800 599914 123856
rect 599582 121760 599638 121816
rect 599950 122848 600006 122904
rect 600042 120808 600098 120864
rect 599858 119720 599914 119776
rect 582194 95784 582250 95840
rect 582102 79328 582158 79384
rect 581918 74704 581974 74760
rect 581642 73208 581698 73264
rect 581550 67224 581606 67280
rect 581366 64232 581422 64288
rect 582286 83816 582342 83872
rect 599950 118788 600006 118824
rect 599950 118768 599952 118788
rect 599952 118768 600004 118788
rect 600004 118768 600006 118788
rect 599858 117680 599914 117736
rect 599950 116728 600006 116784
rect 599858 115640 599914 115696
rect 600042 114688 600098 114744
rect 599950 113600 600006 113656
rect 598938 112648 598994 112704
rect 599950 111560 600006 111616
rect 599858 109520 599914 109576
rect 599950 108568 600006 108624
rect 599858 107480 599914 107536
rect 599950 106528 600006 106584
rect 600226 105440 600282 105496
rect 599950 100408 600006 100464
rect 600502 104488 600558 104544
rect 600318 102448 600374 102504
rect 600410 101360 600466 101416
rect 600686 103400 600742 103456
rect 591946 69400 592002 69456
rect 622490 221312 622546 221368
rect 621478 221176 621534 221232
rect 637854 221040 637910 221096
rect 637394 220904 637450 220960
rect 655610 290400 655666 290456
rect 655794 291488 655850 291544
rect 656254 295296 656310 295352
rect 656806 287272 656862 287328
rect 656806 282104 656862 282160
rect 666558 209208 666614 209264
rect 666558 205808 666614 205864
rect 666558 204176 666614 204232
rect 666558 200776 666614 200832
rect 666558 199008 666614 199064
rect 666558 195608 666614 195664
rect 666558 188944 666614 189000
rect 666558 185544 666614 185600
rect 666558 183776 666614 183832
rect 666558 180376 666614 180432
rect 666558 178744 666614 178800
rect 666558 175344 666614 175400
rect 666558 173576 666614 173632
rect 666558 170176 666614 170232
rect 597466 49680 597522 49736
rect 600042 43152 600098 43208
rect 621202 85992 621258 86048
rect 622490 88848 622546 88904
rect 623226 87896 623282 87952
rect 623502 86944 623558 87000
rect 623318 85040 623374 85096
rect 623134 84088 623190 84144
rect 621938 83136 621994 83192
rect 623778 90616 623834 90672
rect 626446 92520 626502 92576
rect 625894 91568 625950 91624
rect 623962 89664 624018 89720
rect 628286 95920 628342 95976
rect 642270 95920 642326 95976
rect 627918 94424 627974 94480
rect 627274 93472 627330 93528
rect 642730 95104 642786 95160
rect 642638 92656 642694 92712
rect 628562 81640 628618 81696
rect 629206 80824 629262 80880
rect 626538 80144 626594 80200
rect 628470 80144 628526 80200
rect 628470 75520 628526 75576
rect 634174 80144 634230 80200
rect 634174 75520 634230 75576
rect 640338 75384 640394 75440
rect 640982 72392 641038 72448
rect 641074 70896 641130 70952
rect 642822 73344 642878 73400
rect 642914 68856 642970 68912
rect 643006 67360 643062 67416
rect 642638 65864 642694 65920
rect 646042 89664 646098 89720
rect 645950 87080 646006 87136
rect 651562 92520 651618 92576
rect 655334 93336 655390 93392
rect 654046 91432 654102 91488
rect 652758 90616 652814 90672
rect 656898 90344 656954 90400
rect 662234 95512 662290 95568
rect 657358 94696 657414 94752
rect 663246 93744 663302 93800
rect 663338 93064 663394 93120
rect 663430 92248 663486 92304
rect 663522 89528 663578 89584
rect 663706 90344 663762 90400
rect 662142 88712 662198 88768
rect 663890 91024 663946 91080
rect 646134 84632 646190 84688
rect 645858 82184 645914 82240
rect 643098 64368 643154 64424
rect 666742 168544 666798 168600
rect 666742 165144 666798 165200
rect 666742 163512 666798 163568
rect 666742 160112 666798 160168
rect 666742 158344 666798 158400
rect 666742 154944 666798 155000
rect 666742 153312 666798 153368
rect 666742 149912 666798 149968
rect 666742 148144 666798 148200
rect 666742 144880 666798 144936
rect 666742 143112 666798 143168
rect 666742 139712 666798 139768
rect 666742 132912 666798 132968
rect 670698 193976 670754 194032
rect 670698 190576 670754 190632
rect 670340 168282 670400 168342
rect 666742 129512 666798 129568
rect 666650 127880 666706 127936
rect 666650 124480 666706 124536
rect 666650 122848 666706 122904
rect 666650 119448 666706 119504
rect 670506 167872 670566 167932
rect 670346 117728 670402 117784
rect 670698 138080 670754 138136
rect 670698 134680 670754 134736
rect 670502 116098 670558 116154
rect 676126 896008 676182 896064
rect 676034 893036 676090 893072
rect 676034 893016 676036 893036
rect 676036 893016 676088 893036
rect 676088 893016 676090 893036
rect 679162 892608 679218 892664
rect 676034 892200 676090 892256
rect 676034 890976 676090 891032
rect 676034 890568 676090 890624
rect 676034 888936 676090 888992
rect 676034 888528 676090 888584
rect 679070 888120 679126 888176
rect 676034 887712 676090 887768
rect 676034 887304 676090 887360
rect 678978 885012 679034 885048
rect 678978 884992 678980 885012
rect 678980 884992 679032 885012
rect 679032 884992 679034 885012
rect 679438 891792 679494 891848
rect 679254 891384 679310 891440
rect 680266 890160 680322 890216
rect 679714 889752 679770 889808
rect 679530 889344 679586 889400
rect 675114 788296 675170 788352
rect 675206 787072 675262 787128
rect 675298 786800 675354 786856
rect 671986 178744 672042 178800
rect 673734 742736 673790 742792
rect 673734 728456 673790 728512
rect 672078 173576 672134 173632
rect 674286 742600 674342 742656
rect 673458 640192 673514 640248
rect 672170 168544 672226 168600
rect 673550 637608 673606 637664
rect 673550 629312 673606 629368
rect 674470 724648 674526 724704
rect 674470 721520 674526 721576
rect 674470 681128 674526 681184
rect 674470 674056 674526 674112
rect 673734 609184 673790 609240
rect 673734 593544 673790 593600
rect 672262 163512 672318 163568
rect 674838 728728 674894 728784
rect 675390 742872 675446 742928
rect 675666 742464 675722 742520
rect 675114 740288 675170 740344
rect 675114 740152 675170 740208
rect 675114 739608 675170 739664
rect 675390 738656 675446 738712
rect 675758 737976 675814 738032
rect 675298 729000 675354 729056
rect 674930 728592 674986 728648
rect 675022 728320 675078 728376
rect 675298 728184 675354 728240
rect 674286 553832 674342 553888
rect 672354 158344 672410 158400
rect 675942 716488 675998 716544
rect 675850 716080 675906 716136
rect 676034 715672 676090 715728
rect 676034 714892 676036 714912
rect 676036 714892 676088 714912
rect 676088 714892 676090 714912
rect 676034 714856 676090 714892
rect 675666 710776 675722 710832
rect 675942 714060 675998 714096
rect 675942 714040 675944 714060
rect 675944 714040 675996 714060
rect 675996 714040 675998 714060
rect 675942 713244 675998 713280
rect 675942 713224 675944 713244
rect 675944 713224 675996 713244
rect 675996 713224 675998 713244
rect 675942 712428 675998 712464
rect 675942 712408 675944 712428
rect 675944 712408 675996 712428
rect 675996 712408 675998 712428
rect 675758 710368 675814 710424
rect 675758 709180 675760 709200
rect 675760 709180 675812 709200
rect 675812 709180 675814 709200
rect 675758 709144 675814 709180
rect 675850 708328 675906 708384
rect 676034 711592 676090 711648
rect 676034 709960 676090 710016
rect 678978 714448 679034 714504
rect 679070 712816 679126 712872
rect 676034 708736 676090 708792
rect 675942 707920 675998 707976
rect 676034 707512 676090 707568
rect 676034 706288 676090 706344
rect 676034 705100 676036 705120
rect 676036 705100 676088 705120
rect 676088 705100 676090 705120
rect 676034 705064 676090 705100
rect 675574 699624 675630 699680
rect 675390 698128 675446 698184
rect 675758 697176 675814 697232
rect 675758 696632 675814 696688
rect 675758 694728 675814 694784
rect 675482 694320 675538 694376
rect 675758 693504 675814 693560
rect 675758 692960 675814 693016
rect 675390 690512 675446 690568
rect 675390 690104 675446 690160
rect 675942 678408 675998 678464
rect 675942 674736 675998 674792
rect 676218 671064 676274 671120
rect 676034 670928 676090 670984
rect 678978 670248 679034 670304
rect 676034 669704 676090 669760
rect 676034 668888 676090 668944
rect 675482 668072 675538 668128
rect 675390 667256 675446 667312
rect 675298 666440 675354 666496
rect 676218 668652 676220 668672
rect 676220 668652 676272 668672
rect 676272 668652 676274 668672
rect 676218 668616 676274 668652
rect 679162 670248 679218 670304
rect 679070 669432 679126 669488
rect 679254 667800 679310 667856
rect 676034 665216 676090 665272
rect 676034 664808 676090 664864
rect 676034 663176 676090 663232
rect 676034 662768 676090 662824
rect 676034 661544 676090 661600
rect 678978 660864 679034 660920
rect 678978 660048 679034 660104
rect 675666 652568 675722 652624
rect 675482 652160 675538 652216
rect 675390 651616 675446 651672
rect 675390 648896 675446 648952
rect 675390 648624 675446 648680
rect 675298 624688 675354 624744
rect 675206 617072 675262 617128
rect 675758 638152 675814 638208
rect 678978 626048 679034 626104
rect 676218 625640 676274 625696
rect 676126 625232 676182 625288
rect 676034 623908 676036 623928
rect 676036 623908 676088 623928
rect 676088 623908 676090 623928
rect 676034 623872 676090 623908
rect 679070 625232 679126 625288
rect 679162 624416 679218 624472
rect 679254 623600 679310 623656
rect 679346 622784 679402 622840
rect 676218 621988 676274 622024
rect 676218 621968 676220 621988
rect 676220 621968 676272 621988
rect 676272 621968 676274 621988
rect 676034 621424 676090 621480
rect 676034 621016 676090 621072
rect 676034 619792 676090 619848
rect 676034 618196 676036 618216
rect 676036 618196 676088 618216
rect 676088 618196 676090 618216
rect 676034 618160 676090 618196
rect 676126 617888 676182 617944
rect 676034 616528 676090 616584
rect 678978 615848 679034 615904
rect 678978 615032 679034 615088
rect 675390 607824 675446 607880
rect 675758 607280 675814 607336
rect 675206 604968 675262 605024
rect 675114 604424 675170 604480
rect 675298 604424 675354 604480
rect 675114 603744 675170 603800
rect 675114 601840 675170 601896
rect 675574 593136 675630 593192
rect 676034 587696 676090 587752
rect 676034 586200 676090 586256
rect 676126 580896 676182 580952
rect 676310 580488 676366 580544
rect 676218 580100 676274 580136
rect 676218 580080 676220 580100
rect 676220 580080 676272 580100
rect 676272 580080 676274 580100
rect 676034 579808 676090 579864
rect 678978 579264 679034 579320
rect 676034 578584 676090 578640
rect 679070 577632 679126 577688
rect 675942 576136 675998 576192
rect 676034 575728 676090 575784
rect 675574 575320 675630 575376
rect 676034 574912 676090 574968
rect 676034 574504 676090 574560
rect 676034 572872 676090 572928
rect 676034 572464 676090 572520
rect 675482 572056 675538 572112
rect 678978 570696 679034 570752
rect 678978 569880 679034 569936
rect 675482 562400 675538 562456
rect 675298 562264 675354 562320
rect 675482 561176 675538 561232
rect 675298 557504 675354 557560
rect 675482 547984 675538 548040
rect 679254 544040 679310 544096
rect 679070 543904 679126 543960
rect 678978 543768 679034 543824
rect 676126 542680 676182 542736
rect 676126 541184 676182 541240
rect 675482 531256 675538 531312
rect 675390 488824 675446 488880
rect 672446 153312 672502 153368
rect 675482 487192 675538 487248
rect 676218 535880 676274 535936
rect 676034 535712 676036 535732
rect 676036 535712 676088 535732
rect 676088 535712 676090 535732
rect 676034 535676 676090 535712
rect 678978 535064 679034 535120
rect 679162 535064 679218 535120
rect 679346 534248 679402 534304
rect 679530 534248 679586 534304
rect 679254 533432 679310 533488
rect 679070 532616 679126 532672
rect 678978 531800 679034 531856
rect 676034 529964 676090 530020
rect 676034 529556 676090 529612
rect 676034 527924 676090 527980
rect 676034 527516 676090 527572
rect 675942 526700 675998 526756
rect 676034 526292 676090 526348
rect 679070 525680 679126 525736
rect 679070 524864 679126 524920
rect 676034 492088 676090 492144
rect 675942 491680 675998 491736
rect 676034 491272 676090 491328
rect 679254 532616 679310 532672
rect 679438 533432 679494 533488
rect 675758 490456 675814 490512
rect 676034 490864 676090 490920
rect 676034 490048 676090 490104
rect 676034 489640 676090 489696
rect 676034 489232 676090 489288
rect 675942 488416 675998 488472
rect 675942 488008 675998 488064
rect 675850 486376 675906 486432
rect 675850 484336 675906 484392
rect 675574 482704 675630 482760
rect 675850 402600 675906 402656
rect 675298 402192 675354 402248
rect 672538 148144 672594 148200
rect 675758 401376 675814 401432
rect 675666 395664 675722 395720
rect 675666 395256 675722 395312
rect 675850 400968 675906 401024
rect 676034 485968 676090 486024
rect 676034 485560 676090 485616
rect 676034 483928 676090 483984
rect 676034 483520 676090 483576
rect 676034 483112 676090 483168
rect 676034 482296 676090 482352
rect 676034 481888 676090 481944
rect 676034 480700 676036 480720
rect 676036 480700 676088 480720
rect 676088 480700 676090 480720
rect 676034 480664 676090 480700
rect 676126 403688 676182 403744
rect 676218 403280 676274 403336
rect 676126 402872 676182 402928
rect 676034 401784 676090 401840
rect 675942 400152 675998 400208
rect 676034 399744 676090 399800
rect 676034 399336 676090 399392
rect 675850 398520 675906 398576
rect 676126 398792 676182 398848
rect 676034 398112 676090 398168
rect 675942 397704 675998 397760
rect 676034 397296 676090 397352
rect 676034 396888 676090 396944
rect 675942 396072 675998 396128
rect 675942 394848 675998 394904
rect 676126 396344 676182 396400
rect 676034 394440 676090 394496
rect 676034 394032 676090 394088
rect 678978 393488 679034 393544
rect 678978 392672 679034 392728
rect 675298 357448 675354 357504
rect 675206 357040 675262 357096
rect 672630 143112 672686 143168
rect 672722 138352 672778 138408
rect 675850 358672 675906 358728
rect 675758 356632 675814 356688
rect 676034 358264 676090 358320
rect 675942 357856 675998 357912
rect 676034 356224 676090 356280
rect 675758 355408 675814 355464
rect 675666 355000 675722 355056
rect 675298 354592 675354 354648
rect 675390 353776 675446 353832
rect 675666 350512 675722 350568
rect 676034 354184 676090 354240
rect 676034 353368 676090 353424
rect 676034 352960 676090 353016
rect 675942 352552 675998 352608
rect 675942 352144 675998 352200
rect 676034 351736 676090 351792
rect 675942 351328 675998 351384
rect 675850 350920 675906 350976
rect 676034 350104 676090 350160
rect 676034 349696 676090 349752
rect 675942 349288 675998 349344
rect 675850 348880 675906 348936
rect 676034 347268 676090 347304
rect 676034 347248 676036 347268
rect 676036 347248 676088 347268
rect 676088 347248 676090 347268
rect 676310 313520 676366 313576
rect 676126 313112 676182 313168
rect 676034 312432 676090 312488
rect 676218 312704 676274 312760
rect 676218 311908 676274 311944
rect 676218 311888 676220 311908
rect 676220 311888 676272 311908
rect 676272 311888 676274 311908
rect 676034 311652 676036 311672
rect 676036 311652 676088 311672
rect 676088 311652 676090 311672
rect 676034 311616 676090 311652
rect 675298 310800 675354 310856
rect 676218 311092 676274 311128
rect 676218 311072 676220 311092
rect 676220 311072 676272 311092
rect 676272 311072 676274 311092
rect 676218 310276 676274 310312
rect 676218 310256 676220 310276
rect 676220 310256 676272 310276
rect 676272 310256 676274 310276
rect 676034 309984 676090 310040
rect 676218 309460 676274 309496
rect 676218 309440 676220 309460
rect 676220 309440 676272 309460
rect 676272 309440 676274 309460
rect 676034 309188 676090 309224
rect 676034 309168 676036 309188
rect 676036 309168 676088 309188
rect 676088 309168 676090 309188
rect 676034 308760 676090 308816
rect 675758 308352 675814 308408
rect 675298 306312 675354 306368
rect 676034 307944 676090 308000
rect 676126 307400 676182 307456
rect 676034 307128 676090 307184
rect 676034 306720 676090 306776
rect 676034 305904 676090 305960
rect 676126 305360 676182 305416
rect 676126 304952 676182 305008
rect 676034 304680 676090 304736
rect 676126 304136 676182 304192
rect 676034 303864 676090 303920
rect 678978 303320 679034 303376
rect 678978 302504 679034 302560
rect 676126 268504 676182 268560
rect 676034 268232 676090 268288
rect 676218 268116 676274 268152
rect 676218 268096 676220 268116
rect 676220 268096 676272 268116
rect 676272 268096 676274 268116
rect 676034 267452 676036 267472
rect 676036 267452 676088 267472
rect 676088 267452 676090 267472
rect 676034 267416 676090 267452
rect 675666 267008 675722 267064
rect 676034 266636 676036 266656
rect 676036 266636 676088 266656
rect 676088 266636 676090 266656
rect 676034 266600 676090 266636
rect 675758 266192 675814 266248
rect 672814 132912 672870 132968
rect 671986 114280 672042 114336
rect 670882 107480 670938 107536
rect 672262 105848 672318 105904
rect 672170 104080 672226 104136
rect 675206 250144 675262 250200
rect 675206 246200 675262 246256
rect 675482 263336 675538 263392
rect 676034 265820 676036 265840
rect 676036 265820 676088 265840
rect 676088 265820 676090 265840
rect 676034 265784 676090 265820
rect 676218 264832 676274 264888
rect 676034 264560 676090 264616
rect 676034 264152 676090 264208
rect 676126 263608 676182 263664
rect 676034 262928 676090 262984
rect 675942 262520 675998 262576
rect 676034 262112 676090 262168
rect 675850 261704 675906 261760
rect 676034 261296 676090 261352
rect 675942 260480 675998 260536
rect 675942 260072 675998 260128
rect 676126 260752 676182 260808
rect 676034 259664 676090 259720
rect 676034 259256 676090 259312
rect 676126 258712 676182 258768
rect 678978 258304 679034 258360
rect 678978 257488 679034 257544
rect 675666 222264 675722 222320
rect 675298 221856 675354 221912
rect 675942 223488 675998 223544
rect 675850 223080 675906 223136
rect 675758 221448 675814 221504
rect 675758 221040 675814 221096
rect 675666 220224 675722 220280
rect 672906 127880 672962 127936
rect 675022 203768 675078 203824
rect 675022 203496 675078 203552
rect 675298 219408 675354 219464
rect 675390 218592 675446 218648
rect 675482 217368 675538 217424
rect 675574 215328 675630 215384
rect 676034 222672 676090 222728
rect 676034 219816 676090 219872
rect 676034 219000 676090 219056
rect 676034 218184 676090 218240
rect 676034 217776 676090 217832
rect 675942 216960 675998 217016
rect 676034 216552 676090 216608
rect 675942 216144 675998 216200
rect 675850 215736 675906 215792
rect 676034 214920 676090 214976
rect 676034 214512 676090 214568
rect 675942 214104 675998 214160
rect 675942 213696 675998 213752
rect 676034 212084 676090 212120
rect 676034 212064 676036 212084
rect 676036 212064 676088 212084
rect 676088 212064 676090 212084
rect 676218 178780 676220 178800
rect 676220 178780 676272 178800
rect 676272 178780 676274 178800
rect 676218 178744 676274 178780
rect 675942 178100 675944 178120
rect 675944 178100 675996 178120
rect 675996 178100 675998 178120
rect 675942 178064 675998 178100
rect 675942 177692 675944 177712
rect 675944 177692 675996 177712
rect 675996 177692 675998 177712
rect 675942 177656 675998 177692
rect 676034 177248 676090 177304
rect 676034 176860 676090 176896
rect 676034 176840 676036 176860
rect 676036 176840 676088 176860
rect 676088 176840 676090 176860
rect 676034 176432 676090 176488
rect 675942 176044 675998 176080
rect 675942 176024 675944 176044
rect 675944 176024 675996 176044
rect 675996 176024 675998 176044
rect 675298 175616 675354 175672
rect 675942 175228 675998 175264
rect 675942 175208 675944 175228
rect 675944 175208 675996 175228
rect 675996 175208 675998 175228
rect 676034 174800 676090 174856
rect 676034 174412 676090 174448
rect 676034 174392 676036 174412
rect 676036 174392 676088 174412
rect 676088 174392 676090 174412
rect 676034 173984 676090 174040
rect 676034 173576 676090 173632
rect 675298 173168 675354 173224
rect 676034 172760 676090 172816
rect 675942 172352 675998 172408
rect 675942 171944 675998 172000
rect 675942 171536 675998 171592
rect 676034 170720 676090 170776
rect 675942 170312 675998 170368
rect 675850 169904 675906 169960
rect 675942 169496 675998 169552
rect 675850 169088 675906 169144
rect 675758 168680 675814 168736
rect 676034 167068 676090 167104
rect 676034 167048 676036 167068
rect 676036 167048 676088 167068
rect 676088 167048 676090 167068
rect 675758 156984 675814 157040
rect 676126 133048 676182 133104
rect 676034 132932 676090 132968
rect 676034 132912 676036 132932
rect 676036 132912 676088 132932
rect 676088 132912 676090 132932
rect 676218 132640 676274 132696
rect 676218 132268 676220 132288
rect 676220 132268 676272 132288
rect 676272 132268 676274 132288
rect 676218 132232 676274 132268
rect 676034 131708 676090 131744
rect 676034 131688 676036 131708
rect 676036 131688 676088 131708
rect 676088 131688 676090 131708
rect 676218 131452 676220 131472
rect 676220 131452 676272 131472
rect 676272 131452 676274 131472
rect 676218 131416 676274 131452
rect 676034 130892 676090 130928
rect 676034 130872 676036 130892
rect 676036 130872 676088 130892
rect 676088 130872 676090 130892
rect 676218 130636 676220 130656
rect 676220 130636 676272 130656
rect 676272 130636 676274 130656
rect 676218 130600 676274 130636
rect 676034 130076 676090 130112
rect 676034 130056 676036 130076
rect 676036 130056 676088 130076
rect 676088 130056 676090 130076
rect 676034 129684 676036 129704
rect 676036 129684 676088 129704
rect 676088 129684 676090 129704
rect 676034 129648 676090 129684
rect 676218 129412 676220 129432
rect 676220 129412 676272 129432
rect 676272 129412 676274 129432
rect 676218 129376 676274 129412
rect 676034 128832 676090 128888
rect 675942 128424 675998 128480
rect 675574 128016 675630 128072
rect 673278 123072 673338 123132
rect 672998 122848 673054 122904
rect 673426 122670 673486 122730
rect 673284 112690 673340 112746
rect 673418 110926 673474 110982
rect 672446 109248 672502 109304
rect 675298 126384 675354 126440
rect 672354 102448 672410 102504
rect 676034 127608 676090 127664
rect 675942 127200 675998 127256
rect 676034 126792 676090 126848
rect 676034 125976 676090 126032
rect 675942 125568 675998 125624
rect 676126 124888 676182 124944
rect 676126 124480 676182 124536
rect 676034 124344 676090 124400
rect 676034 123936 676090 123992
rect 676034 123528 676090 123584
rect 676218 121644 676274 121680
rect 676218 121624 676220 121644
rect 676220 121624 676272 121644
rect 676272 121624 676274 121644
rect 672078 100816 672134 100872
rect 666558 49000 666614 49056
rect 543646 41248 543702 41304
<< metal3 >>
rect 676029 897154 676095 897157
rect 676029 897152 676292 897154
rect 676029 897096 676034 897152
rect 676090 897096 676292 897152
rect 676029 897094 676292 897096
rect 676029 897091 676095 897094
rect 676029 896746 676095 896749
rect 676029 896744 676292 896746
rect 676029 896688 676034 896744
rect 676090 896688 676292 896744
rect 676029 896686 676292 896688
rect 676029 896683 676095 896686
rect 676121 896066 676187 896069
rect 676262 896066 676322 896308
rect 676121 896064 676322 896066
rect 676121 896008 676126 896064
rect 676182 896008 676322 896064
rect 676121 896006 676322 896008
rect 676121 896003 676187 896006
rect 674414 895460 674420 895524
rect 674484 895522 674490 895524
rect 674484 895462 676292 895522
rect 674484 895460 674490 895462
rect 675937 894706 676003 894709
rect 675937 894704 676292 894706
rect 675937 894648 675942 894704
rect 675998 894648 676292 894704
rect 675937 894646 676292 894648
rect 675937 894643 676003 894646
rect 673862 893828 673868 893892
rect 673932 893890 673938 893892
rect 673932 893830 676292 893890
rect 673932 893828 673938 893830
rect 676029 893074 676095 893077
rect 676029 893072 676292 893074
rect 676029 893016 676034 893072
rect 676090 893016 676292 893072
rect 676029 893014 676292 893016
rect 676029 893011 676095 893014
rect 679157 892666 679223 892669
rect 679157 892664 679236 892666
rect 679157 892608 679162 892664
rect 679218 892608 679236 892664
rect 679157 892606 679236 892608
rect 679157 892603 679223 892606
rect 676029 892258 676095 892261
rect 676029 892256 676292 892258
rect 676029 892200 676034 892256
rect 676090 892200 676292 892256
rect 676029 892198 676292 892200
rect 676029 892195 676095 892198
rect 679433 891850 679499 891853
rect 679420 891848 679499 891850
rect 679420 891792 679438 891848
rect 679494 891792 679499 891848
rect 679420 891790 679499 891792
rect 679433 891787 679499 891790
rect 679249 891442 679315 891445
rect 679236 891440 679315 891442
rect 679236 891384 679254 891440
rect 679310 891384 679315 891440
rect 679236 891382 679315 891384
rect 679249 891379 679315 891382
rect 676029 891034 676095 891037
rect 676029 891032 676292 891034
rect 676029 890976 676034 891032
rect 676090 890976 676292 891032
rect 676029 890974 676292 890976
rect 676029 890971 676095 890974
rect 676029 890626 676095 890629
rect 676029 890624 676292 890626
rect 676029 890568 676034 890624
rect 676090 890568 676292 890624
rect 676029 890566 676292 890568
rect 676029 890563 676095 890566
rect 680261 890218 680327 890221
rect 680261 890216 680340 890218
rect 680261 890160 680266 890216
rect 680322 890160 680340 890216
rect 680261 890158 680340 890160
rect 680261 890155 680327 890158
rect 679709 889810 679775 889813
rect 679709 889808 679788 889810
rect 679709 889752 679714 889808
rect 679770 889752 679788 889808
rect 679709 889750 679788 889752
rect 679709 889747 679775 889750
rect 679525 889402 679591 889405
rect 679525 889400 679604 889402
rect 679525 889344 679530 889400
rect 679586 889344 679604 889400
rect 679525 889342 679604 889344
rect 679525 889339 679591 889342
rect 676029 888994 676095 888997
rect 676029 888992 676292 888994
rect 676029 888936 676034 888992
rect 676090 888936 676292 888992
rect 676029 888934 676292 888936
rect 676029 888931 676095 888934
rect 676029 888586 676095 888589
rect 676029 888584 676292 888586
rect 676029 888528 676034 888584
rect 676090 888528 676292 888584
rect 676029 888526 676292 888528
rect 676029 888523 676095 888526
rect 679065 888178 679131 888181
rect 679052 888176 679131 888178
rect 679052 888120 679070 888176
rect 679126 888120 679131 888176
rect 679052 888118 679131 888120
rect 679065 888115 679131 888118
rect 676029 887770 676095 887773
rect 676029 887768 676292 887770
rect 676029 887712 676034 887768
rect 676090 887712 676292 887768
rect 676029 887710 676292 887712
rect 676029 887707 676095 887710
rect 676029 887362 676095 887365
rect 676029 887360 676292 887362
rect 676029 887304 676034 887360
rect 676090 887304 676292 887360
rect 676029 887302 676292 887304
rect 676029 887299 676095 887302
rect 679206 886684 679266 886924
rect 679198 886620 679204 886684
rect 679268 886620 679274 886684
rect 684542 886108 684602 886516
rect 679198 885804 679204 885868
rect 679268 885804 679274 885868
rect 679206 885700 679266 885804
rect 678973 885050 679039 885053
rect 679198 885050 679204 885052
rect 678973 885048 679204 885050
rect 678973 884992 678978 885048
rect 679034 884992 679204 885048
rect 678973 884990 679204 884992
rect 678973 884987 679039 884990
rect 679198 884988 679204 884990
rect 679268 884988 679274 885052
rect 655605 868866 655671 868869
rect 649950 868864 655671 868866
rect 649950 868808 655610 868864
rect 655666 868808 655671 868864
rect 649950 868806 655671 868808
rect 649950 868246 650010 868806
rect 655605 868803 655671 868806
rect 655421 867642 655487 867645
rect 649950 867640 655487 867642
rect 649950 867584 655426 867640
rect 655482 867584 655487 867640
rect 649950 867582 655487 867584
rect 649950 867064 650010 867582
rect 655421 867579 655487 867582
rect 655513 866554 655579 866557
rect 649950 866552 655579 866554
rect 649950 866496 655518 866552
rect 655574 866496 655579 866552
rect 649950 866494 655579 866496
rect 649950 865882 650010 866494
rect 655513 866491 655579 866494
rect 655697 865330 655763 865333
rect 649950 865328 655763 865330
rect 649950 865272 655702 865328
rect 655758 865272 655763 865328
rect 649950 865270 655763 865272
rect 649950 864700 650010 865270
rect 655697 865267 655763 865270
rect 655789 863834 655855 863837
rect 649950 863832 655855 863834
rect 649950 863776 655794 863832
rect 655850 863776 655855 863832
rect 649950 863774 655855 863776
rect 649950 863518 650010 863774
rect 655789 863771 655855 863774
rect 656801 862610 656867 862613
rect 649950 862608 656867 862610
rect 649950 862552 656806 862608
rect 656862 862552 656867 862608
rect 649950 862550 656867 862552
rect 649950 862336 650010 862550
rect 656801 862547 656867 862550
rect 41781 817730 41847 817733
rect 41492 817728 41847 817730
rect 41492 817672 41786 817728
rect 41842 817672 41847 817728
rect 41492 817670 41847 817672
rect 41781 817667 41847 817670
rect 41781 817322 41847 817325
rect 41492 817320 41847 817322
rect 41492 817264 41786 817320
rect 41842 817264 41847 817320
rect 41492 817262 41847 817264
rect 41781 817259 41847 817262
rect 41781 816914 41847 816917
rect 41492 816912 41847 816914
rect 41492 816856 41786 816912
rect 41842 816856 41847 816912
rect 41492 816854 41847 816856
rect 41781 816851 41847 816854
rect 41781 816098 41847 816101
rect 41492 816096 41847 816098
rect 41492 816040 41786 816096
rect 41842 816040 41847 816096
rect 41492 816038 41847 816040
rect 41781 816035 41847 816038
rect 41781 815282 41847 815285
rect 41492 815280 41847 815282
rect 41492 815224 41786 815280
rect 41842 815224 41847 815280
rect 41492 815222 41847 815224
rect 41781 815219 41847 815222
rect 41781 814466 41847 814469
rect 41492 814464 41847 814466
rect 41492 814408 41786 814464
rect 41842 814408 41847 814464
rect 41492 814406 41847 814408
rect 41781 814403 41847 814406
rect 41781 813650 41847 813653
rect 41492 813648 41847 813650
rect 41492 813592 41786 813648
rect 41842 813592 41847 813648
rect 41492 813590 41847 813592
rect 41781 813587 41847 813590
rect 41781 813242 41847 813245
rect 41492 813240 41847 813242
rect 41492 813184 41786 813240
rect 41842 813184 41847 813240
rect 41492 813182 41847 813184
rect 41781 813179 41847 813182
rect 41781 812834 41847 812837
rect 41492 812832 41847 812834
rect 41492 812776 41786 812832
rect 41842 812776 41847 812832
rect 41492 812774 41847 812776
rect 41781 812771 41847 812774
rect 41781 812426 41847 812429
rect 41492 812424 41847 812426
rect 41492 812368 41786 812424
rect 41842 812368 41847 812424
rect 41492 812366 41847 812368
rect 41781 812363 41847 812366
rect 41278 811848 41338 811988
rect 43713 811882 43779 811885
rect 41692 811880 43779 811882
rect 41692 811848 43718 811880
rect 41278 811824 43718 811848
rect 43774 811824 43779 811880
rect 41278 811822 43779 811824
rect 41278 811788 41752 811822
rect 43713 811819 43779 811822
rect 41965 811610 42031 811613
rect 41492 811608 42031 811610
rect 41492 811552 41970 811608
rect 42026 811552 42031 811608
rect 41492 811550 42031 811552
rect 41965 811547 42031 811550
rect 42241 811202 42307 811205
rect 41492 811200 42307 811202
rect 41492 811144 42246 811200
rect 42302 811144 42307 811200
rect 41492 811142 42307 811144
rect 42241 811139 42307 811142
rect 41781 810794 41847 810797
rect 41492 810792 41847 810794
rect 41492 810736 41786 810792
rect 41842 810736 41847 810792
rect 41492 810734 41847 810736
rect 41781 810731 41847 810734
rect 41873 810386 41939 810389
rect 41492 810384 41939 810386
rect 41492 810328 41878 810384
rect 41934 810328 41939 810384
rect 41492 810326 41939 810328
rect 41873 810323 41939 810326
rect 42609 809978 42675 809981
rect 41492 809976 42675 809978
rect 41492 809920 42614 809976
rect 42670 809920 42675 809976
rect 41492 809918 42675 809920
rect 42609 809915 42675 809918
rect 41781 809570 41847 809573
rect 41492 809568 41847 809570
rect 41492 809512 41786 809568
rect 41842 809512 41847 809568
rect 41492 809510 41847 809512
rect 41781 809507 41847 809510
rect 41822 809162 41828 809164
rect 41492 809102 41828 809162
rect 41822 809100 41828 809102
rect 41892 809100 41898 809164
rect 41873 808754 41939 808757
rect 41492 808752 41939 808754
rect 41492 808696 41878 808752
rect 41934 808696 41939 808752
rect 41492 808694 41939 808696
rect 41873 808691 41939 808694
rect 41781 808346 41847 808349
rect 41492 808344 41847 808346
rect 41492 808288 41786 808344
rect 41842 808288 41847 808344
rect 41492 808286 41847 808288
rect 41781 808283 41847 808286
rect 41781 807938 41847 807941
rect 41492 807936 41847 807938
rect 41492 807880 41786 807936
rect 41842 807880 41847 807936
rect 41492 807878 41847 807880
rect 41781 807875 41847 807878
rect 42057 807530 42123 807533
rect 41492 807528 42123 807530
rect 41492 807472 42062 807528
rect 42118 807472 42123 807528
rect 41492 807470 42123 807472
rect 42057 807467 42123 807470
rect 30422 806684 30482 807092
rect 42057 806306 42123 806309
rect 41492 806304 42123 806306
rect 41492 806248 42062 806304
rect 42118 806248 42123 806304
rect 41492 806246 42123 806248
rect 42057 806243 42123 806246
rect 41873 794476 41939 794477
rect 41822 794474 41828 794476
rect 41782 794414 41828 794474
rect 41892 794472 41939 794476
rect 41934 794416 41939 794472
rect 41822 794412 41828 794414
rect 41892 794412 41939 794416
rect 41873 794411 41939 794412
rect 58249 790938 58315 790941
rect 58249 790936 64706 790938
rect 58249 790880 58254 790936
rect 58310 790880 64706 790936
rect 58249 790878 64706 790880
rect 58249 790875 58315 790878
rect 64646 790304 64706 790878
rect 58525 789306 58591 789309
rect 58525 789304 64706 789306
rect 58525 789248 58530 789304
rect 58586 789248 64706 789304
rect 58525 789246 64706 789248
rect 58525 789243 58591 789246
rect 64646 789122 64706 789246
rect 58157 788490 58223 788493
rect 58157 788488 64706 788490
rect 58157 788432 58162 788488
rect 58218 788432 64706 788488
rect 58157 788430 64706 788432
rect 58157 788427 58223 788430
rect 64646 787940 64706 788430
rect 674966 788292 674972 788356
rect 675036 788354 675042 788356
rect 675109 788354 675175 788357
rect 675036 788352 675175 788354
rect 675036 788296 675114 788352
rect 675170 788296 675175 788352
rect 675036 788294 675175 788296
rect 675036 788292 675042 788294
rect 675109 788291 675175 788294
rect 58433 787402 58499 787405
rect 58433 787400 64706 787402
rect 58433 787344 58438 787400
rect 58494 787344 64706 787400
rect 58433 787342 64706 787344
rect 58433 787339 58499 787342
rect 64646 786758 64706 787342
rect 675201 787132 675267 787133
rect 675150 787130 675156 787132
rect 675110 787070 675156 787130
rect 675220 787128 675267 787132
rect 675262 787072 675267 787128
rect 675150 787068 675156 787070
rect 675220 787068 675267 787072
rect 675201 787067 675267 787068
rect 674046 786796 674052 786860
rect 674116 786858 674122 786860
rect 675293 786858 675359 786861
rect 674116 786856 675359 786858
rect 674116 786800 675298 786856
rect 675354 786800 675359 786856
rect 674116 786798 675359 786800
rect 674116 786796 674122 786798
rect 675293 786795 675359 786798
rect 58525 786178 58591 786181
rect 58525 786176 64706 786178
rect 58525 786120 58530 786176
rect 58586 786120 64706 786176
rect 58525 786118 64706 786120
rect 58525 786115 58591 786118
rect 64646 785576 64706 786118
rect 58433 784954 58499 784957
rect 58433 784952 64706 784954
rect 58433 784896 58438 784952
rect 58494 784896 64706 784952
rect 58433 784894 64706 784896
rect 58433 784891 58499 784894
rect 64646 784394 64706 784894
rect 649950 778426 650010 778824
rect 655421 778426 655487 778429
rect 649950 778424 655487 778426
rect 649950 778368 655426 778424
rect 655482 778368 655487 778424
rect 649950 778366 655487 778368
rect 655421 778363 655487 778366
rect 649950 777066 650010 777642
rect 655789 777066 655855 777069
rect 649950 777064 655855 777066
rect 649950 777008 655794 777064
rect 655850 777008 655855 777064
rect 649950 777006 655855 777008
rect 655789 777003 655855 777006
rect 649950 775978 650010 776460
rect 655605 775978 655671 775981
rect 649950 775976 655671 775978
rect 649950 775920 655610 775976
rect 655666 775920 655671 775976
rect 649950 775918 655671 775920
rect 655605 775915 655671 775918
rect 655513 775570 655579 775573
rect 649950 775568 655579 775570
rect 649950 775512 655518 775568
rect 655574 775512 655579 775568
rect 649950 775510 655579 775512
rect 649950 775278 650010 775510
rect 655513 775507 655579 775510
rect 656525 774754 656591 774757
rect 649950 774752 656591 774754
rect 649950 774696 656530 774752
rect 656586 774696 656591 774752
rect 649950 774694 656591 774696
rect 41781 774482 41847 774485
rect 41492 774480 41847 774482
rect 41492 774424 41786 774480
rect 41842 774424 41847 774480
rect 41492 774422 41847 774424
rect 41781 774419 41847 774422
rect 649950 774096 650010 774694
rect 656525 774691 656591 774694
rect 41462 773941 41522 774044
rect 41413 773936 41522 773941
rect 41413 773880 41418 773936
rect 41474 773880 41522 773936
rect 41413 773878 41522 773880
rect 41413 773875 41479 773878
rect 41781 773666 41847 773669
rect 41492 773664 41847 773666
rect 41492 773608 41786 773664
rect 41842 773608 41847 773664
rect 41492 773606 41847 773608
rect 41781 773603 41847 773606
rect 41505 773530 41571 773533
rect 654961 773530 655027 773533
rect 41462 773528 41571 773530
rect 41462 773472 41510 773528
rect 41566 773472 41571 773528
rect 41462 773467 41571 773472
rect 649950 773528 655027 773530
rect 649950 773472 654966 773528
rect 655022 773472 655027 773528
rect 649950 773470 655027 773472
rect 41462 773228 41522 773467
rect 649950 772914 650010 773470
rect 654961 773467 655027 773470
rect 41873 772850 41939 772853
rect 41492 772848 41939 772850
rect 41492 772792 41878 772848
rect 41934 772792 41939 772848
rect 41492 772790 41939 772792
rect 41873 772787 41939 772790
rect 41505 772714 41571 772717
rect 41462 772712 41571 772714
rect 41462 772656 41510 772712
rect 41566 772656 41571 772712
rect 41462 772651 41571 772656
rect 41462 772412 41522 772651
rect 41462 771901 41522 772004
rect 41462 771896 41571 771901
rect 41462 771840 41510 771896
rect 41566 771840 41571 771896
rect 41462 771838 41571 771840
rect 41505 771835 41571 771838
rect 41781 771626 41847 771629
rect 41492 771624 41847 771626
rect 41492 771568 41786 771624
rect 41842 771568 41847 771624
rect 41492 771566 41847 771568
rect 41781 771563 41847 771566
rect 41462 771085 41522 771188
rect 41413 771080 41522 771085
rect 41413 771024 41418 771080
rect 41474 771024 41522 771080
rect 41413 771022 41522 771024
rect 41413 771019 41479 771022
rect 41781 770810 41847 770813
rect 41492 770808 41847 770810
rect 41492 770752 41786 770808
rect 41842 770752 41847 770808
rect 41492 770750 41847 770752
rect 41781 770747 41847 770750
rect 42149 770402 42215 770405
rect 41492 770400 42215 770402
rect 41492 770344 42154 770400
rect 42210 770344 42215 770400
rect 41492 770342 42215 770344
rect 42149 770339 42215 770342
rect 41462 769861 41522 769964
rect 41462 769856 41571 769861
rect 41462 769800 41510 769856
rect 41566 769800 41571 769856
rect 41462 769798 41571 769800
rect 41505 769795 41571 769798
rect 41462 769453 41522 769556
rect 41462 769448 41571 769453
rect 41462 769392 41510 769448
rect 41566 769392 41571 769448
rect 41462 769390 41571 769392
rect 41505 769387 41571 769390
rect 41462 769045 41522 769148
rect 41462 769040 41571 769045
rect 41462 768984 41510 769040
rect 41566 768984 41571 769040
rect 41462 768982 41571 768984
rect 41505 768979 41571 768982
rect 41462 768637 41522 768740
rect 41462 768632 41571 768637
rect 41462 768576 41510 768632
rect 41566 768576 41571 768632
rect 41462 768574 41571 768576
rect 41505 768571 41571 768574
rect 41462 768229 41522 768332
rect 41462 768224 41571 768229
rect 41462 768168 41510 768224
rect 41566 768168 41571 768224
rect 41462 768166 41571 768168
rect 41505 768163 41571 768166
rect 41781 767954 41847 767957
rect 41492 767952 41847 767954
rect 41492 767896 41786 767952
rect 41842 767896 41847 767952
rect 41492 767894 41847 767896
rect 41781 767891 41847 767894
rect 41462 767413 41522 767516
rect 41462 767408 41571 767413
rect 41462 767352 41510 767408
rect 41566 767352 41571 767408
rect 41462 767350 41571 767352
rect 41505 767347 41571 767350
rect 41462 767002 41522 767108
rect 41689 767002 41755 767005
rect 41462 767000 41755 767002
rect 41462 766944 41694 767000
rect 41750 766944 41755 767000
rect 41462 766942 41755 766944
rect 41689 766939 41755 766942
rect 41462 766597 41522 766700
rect 41413 766592 41522 766597
rect 41413 766536 41418 766592
rect 41474 766536 41522 766592
rect 41413 766534 41522 766536
rect 41413 766531 41479 766534
rect 41462 766189 41522 766292
rect 41462 766184 41571 766189
rect 41462 766128 41510 766184
rect 41566 766128 41571 766184
rect 41462 766126 41571 766128
rect 41505 766123 41571 766126
rect 41462 765781 41522 765884
rect 41462 765776 41571 765781
rect 41462 765720 41510 765776
rect 41566 765720 41571 765776
rect 41462 765718 41571 765720
rect 41505 765715 41571 765718
rect 41462 765370 41522 765476
rect 41597 765370 41663 765373
rect 41462 765368 41663 765370
rect 41462 765312 41602 765368
rect 41658 765312 41663 765368
rect 41462 765310 41663 765312
rect 41597 765307 41663 765310
rect 41462 764965 41522 765068
rect 41462 764960 41571 764965
rect 41462 764904 41510 764960
rect 41566 764904 41571 764960
rect 41462 764902 41571 764904
rect 41505 764899 41571 764902
rect 41462 764557 41522 764660
rect 41462 764552 41571 764557
rect 41462 764496 41510 764552
rect 41566 764496 41571 764552
rect 41462 764494 41571 764496
rect 41505 764491 41571 764494
rect 41462 764149 41522 764252
rect 41462 764144 41571 764149
rect 41462 764088 41510 764144
rect 41566 764088 41571 764144
rect 41462 764086 41571 764088
rect 41505 764083 41571 764086
rect 30422 763436 30482 763844
rect 41462 762925 41522 763028
rect 41462 762920 41571 762925
rect 41462 762864 41510 762920
rect 41566 762864 41571 762920
rect 41462 762862 41571 762864
rect 41505 762859 41571 762862
rect 41781 757074 41847 757077
rect 42006 757074 42012 757076
rect 41781 757072 42012 757074
rect 41781 757016 41786 757072
rect 41842 757016 42012 757072
rect 41781 757014 42012 757016
rect 41781 757011 41847 757014
rect 42006 757012 42012 757014
rect 42076 757012 42082 757076
rect 42149 757074 42215 757077
rect 42742 757074 42748 757076
rect 42149 757072 42748 757074
rect 42149 757016 42154 757072
rect 42210 757016 42748 757072
rect 42149 757014 42748 757016
rect 42149 757011 42215 757014
rect 42742 757012 42748 757014
rect 42812 757012 42818 757076
rect 42742 752932 42748 752996
rect 42812 752994 42818 752996
rect 43069 752994 43135 752997
rect 42812 752992 43135 752994
rect 42812 752936 43074 752992
rect 43130 752936 43135 752992
rect 42812 752934 43135 752936
rect 42812 752932 42818 752934
rect 43069 752931 43135 752934
rect 42006 748716 42012 748780
rect 42076 748778 42082 748780
rect 42425 748778 42491 748781
rect 42076 748776 42491 748778
rect 42076 748720 42430 748776
rect 42486 748720 42491 748776
rect 42076 748718 42491 748720
rect 42076 748716 42082 748718
rect 42425 748715 42491 748718
rect 58433 747690 58499 747693
rect 58433 747688 64706 747690
rect 58433 747632 58438 747688
rect 58494 747632 64706 747688
rect 58433 747630 64706 747632
rect 58433 747627 58499 747630
rect 64646 747082 64706 747630
rect 59261 746466 59327 746469
rect 59261 746464 64706 746466
rect 59261 746408 59266 746464
rect 59322 746408 64706 746464
rect 59261 746406 64706 746408
rect 59261 746403 59327 746406
rect 64646 745900 64706 746406
rect 58433 744970 58499 744973
rect 58433 744968 64706 744970
rect 58433 744912 58438 744968
rect 58494 744912 64706 744968
rect 58433 744910 64706 744912
rect 58433 744907 58499 744910
rect 64646 744718 64706 744910
rect 58525 744154 58591 744157
rect 58525 744152 64706 744154
rect 58525 744096 58530 744152
rect 58586 744096 64706 744152
rect 58525 744094 64706 744096
rect 58525 744091 58591 744094
rect 64646 743536 64706 744094
rect 675385 742932 675451 742933
rect 675334 742930 675340 742932
rect 675294 742870 675340 742930
rect 675404 742928 675451 742932
rect 675446 742872 675451 742928
rect 675334 742868 675340 742870
rect 675404 742868 675451 742872
rect 675385 742867 675451 742868
rect 673729 742794 673795 742797
rect 676642 742794 676648 742796
rect 673729 742792 676648 742794
rect 673729 742736 673734 742792
rect 673790 742736 676648 742792
rect 673729 742734 676648 742736
rect 673729 742731 673795 742734
rect 676642 742732 676648 742734
rect 676712 742732 676718 742796
rect 674281 742658 674347 742661
rect 676806 742658 676812 742660
rect 674281 742656 676812 742658
rect 674281 742600 674286 742656
rect 674342 742600 676812 742656
rect 674281 742598 676812 742600
rect 674281 742595 674347 742598
rect 676806 742596 676812 742598
rect 676876 742596 676882 742660
rect 675661 742524 675727 742525
rect 675661 742520 675708 742524
rect 675772 742522 675778 742524
rect 675661 742464 675666 742520
rect 675661 742460 675708 742464
rect 675772 742462 675818 742522
rect 675772 742460 675778 742462
rect 675661 742459 675727 742460
rect 57973 742386 58039 742389
rect 57973 742384 64706 742386
rect 57973 742328 57978 742384
rect 58034 742328 64706 742384
rect 57973 742326 64706 742328
rect 57973 742323 58039 742326
rect 58433 741842 58499 741845
rect 58433 741840 64706 741842
rect 58433 741784 58438 741840
rect 58494 741784 64706 741840
rect 58433 741782 64706 741784
rect 58433 741779 58499 741782
rect 64646 741172 64706 741782
rect 674230 740284 674236 740348
rect 674300 740346 674306 740348
rect 675109 740346 675175 740349
rect 674300 740344 675175 740346
rect 674300 740288 675114 740344
rect 675170 740288 675175 740344
rect 674300 740286 675175 740288
rect 674300 740284 674306 740286
rect 675109 740283 675175 740286
rect 674598 740148 674604 740212
rect 674668 740210 674674 740212
rect 675109 740210 675175 740213
rect 674668 740208 675175 740210
rect 674668 740152 675114 740208
rect 675170 740152 675175 740208
rect 674668 740150 675175 740152
rect 674668 740148 674674 740150
rect 675109 740147 675175 740150
rect 673494 739604 673500 739668
rect 673564 739666 673570 739668
rect 675109 739666 675175 739669
rect 673564 739664 675175 739666
rect 673564 739608 675114 739664
rect 675170 739608 675175 739664
rect 673564 739606 675175 739608
rect 673564 739604 673570 739606
rect 675109 739603 675175 739606
rect 674782 738652 674788 738716
rect 674852 738714 674858 738716
rect 675385 738714 675451 738717
rect 674852 738712 675451 738714
rect 674852 738656 675390 738712
rect 675446 738656 675451 738712
rect 674852 738654 675451 738656
rect 674852 738652 674858 738654
rect 675385 738651 675451 738654
rect 675753 738034 675819 738037
rect 677174 738034 677180 738036
rect 675753 738032 677180 738034
rect 675753 737976 675758 738032
rect 675814 737976 677180 738032
rect 675753 737974 677180 737976
rect 675753 737971 675819 737974
rect 677174 737972 677180 737974
rect 677244 737972 677250 738036
rect 649950 734362 650010 734402
rect 655513 734362 655579 734365
rect 649950 734360 655579 734362
rect 649950 734304 655518 734360
rect 655574 734304 655579 734360
rect 649950 734302 655579 734304
rect 655513 734299 655579 734302
rect 649950 732730 650010 733220
rect 655881 732730 655947 732733
rect 649950 732728 655947 732730
rect 649950 732672 655886 732728
rect 655942 732672 655947 732728
rect 649950 732670 655947 732672
rect 655881 732667 655947 732670
rect 649950 731506 650010 732038
rect 655697 731506 655763 731509
rect 649950 731504 655763 731506
rect 649950 731448 655702 731504
rect 655758 731448 655763 731504
rect 649950 731446 655763 731448
rect 655697 731443 655763 731446
rect 655973 731370 656039 731373
rect 649950 731368 656039 731370
rect 41462 731101 41522 731340
rect 649950 731312 655978 731368
rect 656034 731312 656039 731368
rect 649950 731310 656039 731312
rect 41462 731096 41571 731101
rect 41462 731040 41510 731096
rect 41566 731040 41571 731096
rect 41462 731038 41571 731040
rect 41505 731035 41571 731038
rect 41462 730693 41522 730932
rect 649950 730856 650010 731310
rect 655973 731307 656039 731310
rect 41462 730688 41571 730693
rect 41462 730632 41510 730688
rect 41566 730632 41571 730688
rect 41462 730630 41571 730632
rect 41505 730627 41571 730630
rect 41462 730285 41522 730524
rect 41462 730280 41571 730285
rect 654317 730282 654383 730285
rect 41462 730224 41510 730280
rect 41566 730224 41571 730280
rect 41462 730222 41571 730224
rect 41505 730219 41571 730222
rect 649950 730280 654383 730282
rect 649950 730224 654322 730280
rect 654378 730224 654383 730280
rect 649950 730222 654383 730224
rect 41873 730146 41939 730149
rect 41492 730144 41939 730146
rect 41492 730088 41878 730144
rect 41934 730088 41939 730144
rect 41492 730086 41939 730088
rect 41873 730083 41939 730086
rect 41462 729469 41522 729708
rect 649950 729674 650010 730222
rect 654317 730219 654383 730222
rect 41462 729464 41571 729469
rect 41462 729408 41510 729464
rect 41566 729408 41571 729464
rect 41462 729406 41571 729408
rect 41505 729403 41571 729406
rect 41781 729330 41847 729333
rect 41492 729328 41847 729330
rect 41492 729272 41786 729328
rect 41842 729272 41847 729328
rect 41492 729270 41847 729272
rect 41781 729267 41847 729270
rect 675293 729058 675359 729061
rect 675518 729058 675524 729060
rect 675293 729056 675524 729058
rect 675293 729000 675298 729056
rect 675354 729000 675524 729056
rect 675293 728998 675524 729000
rect 675293 728995 675359 728998
rect 675518 728996 675524 728998
rect 675588 728996 675594 729060
rect 42425 728922 42491 728925
rect 41492 728920 42491 728922
rect 41492 728864 42430 728920
rect 42486 728864 42491 728920
rect 41492 728862 42491 728864
rect 42425 728859 42491 728862
rect 674833 728786 674899 728789
rect 673502 728784 674899 728786
rect 673502 728728 674838 728784
rect 674894 728728 674899 728784
rect 673502 728726 674899 728728
rect 41505 728650 41571 728653
rect 656065 728650 656131 728653
rect 41462 728648 41571 728650
rect 41462 728592 41510 728648
rect 41566 728592 41571 728648
rect 41462 728587 41571 728592
rect 651330 728648 656131 728650
rect 651330 728592 656070 728648
rect 656126 728592 656131 728648
rect 651330 728590 656131 728592
rect 41462 728484 41522 728587
rect 651330 728514 651390 728590
rect 656065 728587 656131 728590
rect 649950 728454 651390 728514
rect 673502 728514 673562 728726
rect 674833 728723 674899 728726
rect 674925 728650 674991 728653
rect 674925 728648 675034 728650
rect 674925 728592 674930 728648
rect 674986 728592 675034 728648
rect 674925 728587 675034 728592
rect 673729 728514 673795 728517
rect 673502 728512 673795 728514
rect 673502 728456 673734 728512
rect 673790 728456 673795 728512
rect 673502 728454 673795 728456
rect 673729 728451 673795 728454
rect 674974 728381 675034 728587
rect 674974 728376 675083 728381
rect 674974 728320 675022 728376
rect 675078 728320 675083 728376
rect 674974 728318 675083 728320
rect 675017 728315 675083 728318
rect 675293 728242 675359 728245
rect 675518 728242 675524 728244
rect 675293 728240 675524 728242
rect 675293 728184 675298 728240
rect 675354 728184 675524 728240
rect 675293 728182 675524 728184
rect 675293 728179 675359 728182
rect 675518 728180 675524 728182
rect 675588 728180 675594 728244
rect 41781 728106 41847 728109
rect 41492 728104 41847 728106
rect 41492 728048 41786 728104
rect 41842 728048 41847 728104
rect 41492 728046 41847 728048
rect 41781 728043 41847 728046
rect 41505 727834 41571 727837
rect 41462 727832 41571 727834
rect 41462 727776 41510 727832
rect 41566 727776 41571 727832
rect 41462 727771 41571 727776
rect 41462 727668 41522 727771
rect 41965 727290 42031 727293
rect 41492 727288 42031 727290
rect 41492 727232 41970 727288
rect 42026 727232 42031 727288
rect 41492 727230 42031 727232
rect 41965 727227 42031 727230
rect 41462 726613 41522 726852
rect 41462 726608 41571 726613
rect 41462 726552 41510 726608
rect 41566 726552 41571 726608
rect 41462 726550 41571 726552
rect 41505 726547 41571 726550
rect 41462 726205 41522 726444
rect 41462 726200 41571 726205
rect 41462 726144 41510 726200
rect 41566 726144 41571 726200
rect 41462 726142 41571 726144
rect 41505 726139 41571 726142
rect 41781 726066 41847 726069
rect 41492 726064 41847 726066
rect 41492 726008 41786 726064
rect 41842 726008 41847 726064
rect 41492 726006 41847 726008
rect 41781 726003 41847 726006
rect 41462 725389 41522 725628
rect 41462 725384 41571 725389
rect 41462 725328 41510 725384
rect 41566 725328 41571 725384
rect 41462 725326 41571 725328
rect 41505 725323 41571 725326
rect 41781 725250 41847 725253
rect 41492 725248 41847 725250
rect 41492 725192 41786 725248
rect 41842 725192 41847 725248
rect 41492 725190 41847 725192
rect 41781 725187 41847 725190
rect 42241 724842 42307 724845
rect 41492 724840 42307 724842
rect 41492 724784 42246 724840
rect 42302 724784 42307 724840
rect 41492 724782 42307 724784
rect 42241 724779 42307 724782
rect 674046 724644 674052 724708
rect 674116 724706 674122 724708
rect 674465 724706 674531 724709
rect 674116 724704 674531 724706
rect 674116 724648 674470 724704
rect 674526 724648 674531 724704
rect 674116 724646 674531 724648
rect 674116 724644 674122 724646
rect 674465 724643 674531 724646
rect 41462 724165 41522 724404
rect 674046 724236 674052 724300
rect 674116 724298 674122 724300
rect 674414 724298 674420 724300
rect 674116 724238 674420 724298
rect 674116 724236 674122 724238
rect 674414 724236 674420 724238
rect 674484 724236 674490 724300
rect 41462 724160 41571 724165
rect 41462 724104 41510 724160
rect 41566 724104 41571 724160
rect 41462 724102 41571 724104
rect 41505 724099 41571 724102
rect 673862 724100 673868 724164
rect 673932 724162 673938 724164
rect 675150 724162 675156 724164
rect 673932 724102 675156 724162
rect 673932 724100 673938 724102
rect 675150 724100 675156 724102
rect 675220 724100 675226 724164
rect 30238 723757 30298 723996
rect 674414 723964 674420 724028
rect 674484 724026 674490 724028
rect 674966 724026 674972 724028
rect 674484 723966 674972 724026
rect 674484 723964 674490 723966
rect 674966 723964 674972 723966
rect 675036 723964 675042 724028
rect 30238 723752 30347 723757
rect 30238 723696 30286 723752
rect 30342 723696 30347 723752
rect 30238 723694 30347 723696
rect 30281 723691 30347 723694
rect 41462 723346 41522 723588
rect 41689 723346 41755 723349
rect 41462 723344 41755 723346
rect 41462 723288 41694 723344
rect 41750 723288 41755 723344
rect 41462 723286 41755 723288
rect 41689 723283 41755 723286
rect 41781 723210 41847 723213
rect 41492 723208 41847 723210
rect 41492 723152 41786 723208
rect 41842 723152 41847 723208
rect 41492 723150 41847 723152
rect 41781 723147 41847 723150
rect 41873 722802 41939 722805
rect 41492 722800 41939 722802
rect 41492 722744 41878 722800
rect 41934 722744 41939 722800
rect 41492 722742 41939 722744
rect 41873 722739 41939 722742
rect 41462 722125 41522 722364
rect 41462 722120 41571 722125
rect 41462 722064 41510 722120
rect 41566 722064 41571 722120
rect 41462 722062 41571 722064
rect 41505 722059 41571 722062
rect 41462 721717 41522 721956
rect 41462 721712 41571 721717
rect 41462 721656 41510 721712
rect 41566 721656 41571 721712
rect 41462 721654 41571 721656
rect 41505 721651 41571 721654
rect 674465 721578 674531 721581
rect 675886 721578 675892 721580
rect 674465 721576 675892 721578
rect 41462 721306 41522 721548
rect 674465 721520 674470 721576
rect 674526 721520 675892 721576
rect 674465 721518 675892 721520
rect 674465 721515 674531 721518
rect 675886 721516 675892 721518
rect 675956 721516 675962 721580
rect 41597 721306 41663 721309
rect 41462 721304 41663 721306
rect 41462 721248 41602 721304
rect 41658 721248 41663 721304
rect 41462 721246 41663 721248
rect 41597 721243 41663 721246
rect 41462 720901 41522 721140
rect 41413 720896 41522 720901
rect 41413 720840 41418 720896
rect 41474 720840 41522 720896
rect 41413 720838 41522 720840
rect 41413 720835 41479 720838
rect 24902 720324 24962 720732
rect 41462 719677 41522 719916
rect 41462 719672 41571 719677
rect 41462 719616 41510 719672
rect 41566 719616 41571 719672
rect 41462 719614 41571 719616
rect 41505 719611 41571 719614
rect 675937 716546 676003 716549
rect 675937 716544 676292 716546
rect 675937 716488 675942 716544
rect 675998 716488 676292 716544
rect 675937 716486 676292 716488
rect 675937 716483 676003 716486
rect 675845 716138 675911 716141
rect 675845 716136 676292 716138
rect 675845 716080 675850 716136
rect 675906 716080 676292 716136
rect 675845 716078 676292 716080
rect 675845 716075 675911 716078
rect 676029 715730 676095 715733
rect 676029 715728 676292 715730
rect 676029 715672 676034 715728
rect 676090 715672 676292 715728
rect 676029 715670 676292 715672
rect 676029 715667 676095 715670
rect 674046 715260 674052 715324
rect 674116 715322 674122 715324
rect 674116 715262 676292 715322
rect 674116 715260 674122 715262
rect 676029 714914 676095 714917
rect 676029 714912 676292 714914
rect 676029 714856 676034 714912
rect 676090 714856 676292 714912
rect 676029 714854 676292 714856
rect 676029 714851 676095 714854
rect 678973 714506 679039 714509
rect 678973 714504 679052 714506
rect 678973 714448 678978 714504
rect 679034 714448 679052 714504
rect 678973 714446 679052 714448
rect 678973 714443 679039 714446
rect 43069 714372 43135 714373
rect 43069 714370 43116 714372
rect 43024 714368 43116 714370
rect 43024 714312 43074 714368
rect 43024 714310 43116 714312
rect 43069 714308 43116 714310
rect 43180 714308 43186 714372
rect 43069 714307 43135 714308
rect 43161 714234 43227 714237
rect 43662 714234 43668 714236
rect 43161 714232 43668 714234
rect 43161 714176 43166 714232
rect 43222 714176 43668 714232
rect 43161 714174 43668 714176
rect 43161 714171 43227 714174
rect 43662 714172 43668 714174
rect 43732 714172 43738 714236
rect 675937 714098 676003 714101
rect 675937 714096 676292 714098
rect 675937 714040 675942 714096
rect 675998 714040 676292 714096
rect 675937 714038 676292 714040
rect 675937 714035 676003 714038
rect 673678 713628 673684 713692
rect 673748 713690 673754 713692
rect 673748 713630 676292 713690
rect 673748 713628 673754 713630
rect 675937 713282 676003 713285
rect 675937 713280 676292 713282
rect 675937 713224 675942 713280
rect 675998 713224 676292 713280
rect 675937 713222 676292 713224
rect 675937 713219 676003 713222
rect 679065 712874 679131 712877
rect 679052 712872 679131 712874
rect 679052 712816 679070 712872
rect 679126 712816 679131 712872
rect 679052 712814 679131 712816
rect 679065 712811 679131 712814
rect 675937 712466 676003 712469
rect 675937 712464 676292 712466
rect 675937 712408 675942 712464
rect 675998 712408 676292 712464
rect 675937 712406 676292 712408
rect 675937 712403 676003 712406
rect 675886 711996 675892 712060
rect 675956 712058 675962 712060
rect 675956 711998 676292 712058
rect 675956 711996 675962 711998
rect 676029 711650 676095 711653
rect 676029 711648 676292 711650
rect 676029 711592 676034 711648
rect 676090 711592 676292 711648
rect 676029 711590 676292 711592
rect 676029 711587 676095 711590
rect 43110 711452 43116 711516
rect 43180 711514 43186 711516
rect 43437 711514 43503 711517
rect 43180 711512 43503 711514
rect 43180 711456 43442 711512
rect 43498 711456 43503 711512
rect 43180 711454 43503 711456
rect 43180 711452 43186 711454
rect 43437 711451 43503 711454
rect 674414 711180 674420 711244
rect 674484 711242 674490 711244
rect 674484 711182 676292 711242
rect 674484 711180 674490 711182
rect 675661 710834 675727 710837
rect 675661 710832 676292 710834
rect 675661 710776 675666 710832
rect 675722 710776 676292 710832
rect 675661 710774 676292 710776
rect 675661 710771 675727 710774
rect 675753 710426 675819 710429
rect 675753 710424 676292 710426
rect 675753 710368 675758 710424
rect 675814 710368 676292 710424
rect 675753 710366 676292 710368
rect 675753 710363 675819 710366
rect 676029 710018 676095 710021
rect 676029 710016 676292 710018
rect 676029 709960 676034 710016
rect 676090 709960 676292 710016
rect 676029 709958 676292 709960
rect 676029 709955 676095 709958
rect 673862 709548 673868 709612
rect 673932 709610 673938 709612
rect 673932 709550 676292 709610
rect 673932 709548 673938 709550
rect 42742 709412 42748 709476
rect 42812 709474 42818 709476
rect 43713 709474 43779 709477
rect 42812 709472 43779 709474
rect 42812 709416 43718 709472
rect 43774 709416 43779 709472
rect 42812 709414 43779 709416
rect 42812 709412 42818 709414
rect 43713 709411 43779 709414
rect 675753 709202 675819 709205
rect 675753 709200 676292 709202
rect 675753 709144 675758 709200
rect 675814 709144 676292 709200
rect 675753 709142 676292 709144
rect 675753 709139 675819 709142
rect 42241 708930 42307 708933
rect 42742 708930 42748 708932
rect 42241 708928 42748 708930
rect 42241 708872 42246 708928
rect 42302 708872 42748 708928
rect 42241 708870 42748 708872
rect 42241 708867 42307 708870
rect 42742 708868 42748 708870
rect 42812 708868 42818 708932
rect 676029 708794 676095 708797
rect 676029 708792 676292 708794
rect 676029 708736 676034 708792
rect 676090 708736 676292 708792
rect 676029 708734 676292 708736
rect 676029 708731 676095 708734
rect 43662 708460 43668 708524
rect 43732 708522 43738 708524
rect 43805 708522 43871 708525
rect 43732 708520 43871 708522
rect 43732 708464 43810 708520
rect 43866 708464 43871 708520
rect 43732 708462 43871 708464
rect 43732 708460 43738 708462
rect 43805 708459 43871 708462
rect 675845 708386 675911 708389
rect 675845 708384 676292 708386
rect 675845 708328 675850 708384
rect 675906 708328 676292 708384
rect 675845 708326 676292 708328
rect 675845 708323 675911 708326
rect 675937 707978 676003 707981
rect 675937 707976 676292 707978
rect 675937 707920 675942 707976
rect 675998 707920 676292 707976
rect 675937 707918 676292 707920
rect 675937 707915 676003 707918
rect 676029 707570 676095 707573
rect 676029 707568 676292 707570
rect 676029 707512 676034 707568
rect 676090 707512 676292 707568
rect 676029 707510 676292 707512
rect 676029 707507 676095 707510
rect 676070 707236 676076 707300
rect 676140 707236 676146 707300
rect 676078 707162 676138 707236
rect 676078 707102 676292 707162
rect 675886 706692 675892 706756
rect 675956 706754 675962 706756
rect 675956 706694 676292 706754
rect 675956 706692 675962 706694
rect 676029 706346 676095 706349
rect 676029 706344 676292 706346
rect 676029 706288 676034 706344
rect 676090 706288 676292 706344
rect 676029 706286 676292 706288
rect 676029 706283 676095 706286
rect 684542 705500 684602 705908
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 59353 704442 59419 704445
rect 59353 704440 64706 704442
rect 59353 704384 59358 704440
rect 59414 704384 64706 704440
rect 59353 704382 64706 704384
rect 59353 704379 59419 704382
rect 64646 703860 64706 704382
rect 59261 703354 59327 703357
rect 59261 703352 64706 703354
rect 59261 703296 59266 703352
rect 59322 703296 64706 703352
rect 59261 703294 64706 703296
rect 59261 703291 59327 703294
rect 64646 702678 64706 703294
rect 58525 702130 58591 702133
rect 58525 702128 64706 702130
rect 58525 702072 58530 702128
rect 58586 702072 64706 702128
rect 58525 702070 64706 702072
rect 58525 702067 58591 702070
rect 64646 701496 64706 702070
rect 58249 700770 58315 700773
rect 58249 700768 64706 700770
rect 58249 700712 58254 700768
rect 58310 700712 64706 700768
rect 58249 700710 64706 700712
rect 58249 700707 58315 700710
rect 64646 700314 64706 700710
rect 58525 699682 58591 699685
rect 675569 699682 675635 699685
rect 676990 699682 676996 699684
rect 58525 699680 64706 699682
rect 58525 699624 58530 699680
rect 58586 699624 64706 699680
rect 58525 699622 64706 699624
rect 58525 699619 58591 699622
rect 64646 699132 64706 699622
rect 675569 699680 676996 699682
rect 675569 699624 675574 699680
rect 675630 699624 676996 699680
rect 675569 699622 676996 699624
rect 675569 699619 675635 699622
rect 676990 699620 676996 699622
rect 677060 699620 677066 699684
rect 58525 698186 58591 698189
rect 58525 698184 64706 698186
rect 58525 698128 58530 698184
rect 58586 698128 64706 698184
rect 58525 698126 64706 698128
rect 58525 698123 58591 698126
rect 64646 697950 64706 698126
rect 673862 698124 673868 698188
rect 673932 698186 673938 698188
rect 675385 698186 675451 698189
rect 673932 698184 675451 698186
rect 673932 698128 675390 698184
rect 675446 698128 675451 698184
rect 673932 698126 675451 698128
rect 673932 698124 673938 698126
rect 675385 698123 675451 698126
rect 675753 697234 675819 697237
rect 676070 697234 676076 697236
rect 675753 697232 676076 697234
rect 675753 697176 675758 697232
rect 675814 697176 676076 697232
rect 675753 697174 676076 697176
rect 675753 697171 675819 697174
rect 676070 697172 676076 697174
rect 676140 697172 676146 697236
rect 675753 696690 675819 696693
rect 676806 696690 676812 696692
rect 675753 696688 676812 696690
rect 675753 696632 675758 696688
rect 675814 696632 676812 696688
rect 675753 696630 676812 696632
rect 675753 696627 675819 696630
rect 676806 696628 676812 696630
rect 676876 696628 676882 696692
rect 675753 694786 675819 694789
rect 675886 694786 675892 694788
rect 675753 694784 675892 694786
rect 675753 694728 675758 694784
rect 675814 694728 675892 694784
rect 675753 694726 675892 694728
rect 675753 694723 675819 694726
rect 675886 694724 675892 694726
rect 675956 694724 675962 694788
rect 674046 694316 674052 694380
rect 674116 694378 674122 694380
rect 675477 694378 675543 694381
rect 674116 694376 675543 694378
rect 674116 694320 675482 694376
rect 675538 694320 675543 694376
rect 674116 694318 675543 694320
rect 674116 694316 674122 694318
rect 675477 694315 675543 694318
rect 675753 693562 675819 693565
rect 676642 693562 676648 693564
rect 675753 693560 676648 693562
rect 675753 693504 675758 693560
rect 675814 693504 676648 693560
rect 675753 693502 676648 693504
rect 675753 693499 675819 693502
rect 676642 693500 676648 693502
rect 676712 693500 676718 693564
rect 675753 693018 675819 693021
rect 677174 693018 677180 693020
rect 675753 693016 677180 693018
rect 675753 692960 675758 693016
rect 675814 692960 677180 693016
rect 675753 692958 677180 692960
rect 675753 692955 675819 692958
rect 677174 692956 677180 692958
rect 677244 692956 677250 693020
rect 673678 690508 673684 690572
rect 673748 690570 673754 690572
rect 675385 690570 675451 690573
rect 673748 690568 675451 690570
rect 673748 690512 675390 690568
rect 675446 690512 675451 690568
rect 673748 690510 675451 690512
rect 673748 690508 673754 690510
rect 675385 690507 675451 690510
rect 674414 690100 674420 690164
rect 674484 690162 674490 690164
rect 675385 690162 675451 690165
rect 674484 690160 675451 690162
rect 674484 690104 675390 690160
rect 675446 690104 675451 690160
rect 674484 690102 675451 690104
rect 674484 690100 674490 690102
rect 675385 690099 675451 690102
rect 649950 689482 650010 689980
rect 655789 689482 655855 689485
rect 649950 689480 655855 689482
rect 649950 689424 655794 689480
rect 655850 689424 655855 689480
rect 649950 689422 655855 689424
rect 655789 689419 655855 689422
rect 649950 688258 650010 688798
rect 655605 688258 655671 688261
rect 649950 688256 655671 688258
rect 649950 688200 655610 688256
rect 655666 688200 655671 688256
rect 649950 688198 655671 688200
rect 655605 688195 655671 688198
rect 41781 688122 41847 688125
rect 41492 688120 41847 688122
rect 41492 688064 41786 688120
rect 41842 688064 41847 688120
rect 41492 688062 41847 688064
rect 41781 688059 41847 688062
rect 41781 687714 41847 687717
rect 41492 687712 41847 687714
rect 41492 687656 41786 687712
rect 41842 687656 41847 687712
rect 41492 687654 41847 687656
rect 41781 687651 41847 687654
rect 41781 687306 41847 687309
rect 41492 687304 41847 687306
rect 41492 687248 41786 687304
rect 41842 687248 41847 687304
rect 41492 687246 41847 687248
rect 649950 687306 650010 687616
rect 655421 687306 655487 687309
rect 649950 687304 655487 687306
rect 649950 687248 655426 687304
rect 655482 687248 655487 687304
rect 649950 687246 655487 687248
rect 41781 687243 41847 687246
rect 655421 687243 655487 687246
rect 655973 687034 656039 687037
rect 649950 687032 656039 687034
rect 649950 686976 655978 687032
rect 656034 686976 656039 687032
rect 649950 686974 656039 686976
rect 41781 686898 41847 686901
rect 41492 686896 41847 686898
rect 41492 686840 41786 686896
rect 41842 686840 41847 686896
rect 41492 686838 41847 686840
rect 41781 686835 41847 686838
rect 41781 686490 41847 686493
rect 41492 686488 41847 686490
rect 41492 686432 41786 686488
rect 41842 686432 41847 686488
rect 649950 686434 650010 686974
rect 655973 686971 656039 686974
rect 41492 686430 41847 686432
rect 41781 686427 41847 686430
rect 42425 686082 42491 686085
rect 41492 686080 42491 686082
rect 41492 686024 42430 686080
rect 42486 686024 42491 686080
rect 41492 686022 42491 686024
rect 42425 686019 42491 686022
rect 654225 685810 654291 685813
rect 649950 685808 654291 685810
rect 649950 685752 654230 685808
rect 654286 685752 654291 685808
rect 649950 685750 654291 685752
rect 42057 685674 42123 685677
rect 41492 685672 42123 685674
rect 41492 685616 42062 685672
rect 42118 685616 42123 685672
rect 41492 685614 42123 685616
rect 42057 685611 42123 685614
rect 41781 685266 41847 685269
rect 41492 685264 41847 685266
rect 41492 685208 41786 685264
rect 41842 685208 41847 685264
rect 649950 685252 650010 685750
rect 654225 685747 654291 685750
rect 41492 685206 41847 685208
rect 41781 685203 41847 685206
rect 42425 684858 42491 684861
rect 41492 684856 42491 684858
rect 41492 684800 42430 684856
rect 42486 684800 42491 684856
rect 41492 684798 42491 684800
rect 42425 684795 42491 684798
rect 41781 684450 41847 684453
rect 654133 684450 654199 684453
rect 41492 684448 41847 684450
rect 41492 684392 41786 684448
rect 41842 684392 41847 684448
rect 41492 684390 41847 684392
rect 41781 684387 41847 684390
rect 649950 684448 654199 684450
rect 649950 684392 654138 684448
rect 654194 684392 654199 684448
rect 649950 684390 654199 684392
rect 649950 684070 650010 684390
rect 654133 684387 654199 684390
rect 41781 684042 41847 684045
rect 41492 684040 41847 684042
rect 41492 683984 41786 684040
rect 41842 683984 41847 684040
rect 41492 683982 41847 683984
rect 41781 683979 41847 683982
rect 41781 683634 41847 683637
rect 41492 683632 41847 683634
rect 41492 683576 41786 683632
rect 41842 683576 41847 683632
rect 41492 683574 41847 683576
rect 41781 683571 41847 683574
rect 42241 683226 42307 683229
rect 41492 683224 42307 683226
rect 41492 683168 42246 683224
rect 42302 683168 42307 683224
rect 41492 683166 42307 683168
rect 42241 683163 42307 683166
rect 41462 682682 41522 682788
rect 41689 682682 41755 682685
rect 41462 682680 41755 682682
rect 41462 682624 41694 682680
rect 41750 682624 41755 682680
rect 41462 682622 41755 682624
rect 41689 682619 41755 682622
rect 41462 682274 41522 682380
rect 41689 682274 41755 682277
rect 41462 682272 41755 682274
rect 41462 682216 41694 682272
rect 41750 682216 41755 682272
rect 41462 682214 41755 682216
rect 41689 682211 41755 682214
rect 30281 682002 30347 682005
rect 30268 682000 30347 682002
rect 30268 681944 30286 682000
rect 30342 681944 30347 682000
rect 30268 681942 30347 681944
rect 30281 681939 30347 681942
rect 42333 681594 42399 681597
rect 41492 681592 42399 681594
rect 41492 681536 42338 681592
rect 42394 681536 42399 681592
rect 41492 681534 42399 681536
rect 42333 681531 42399 681534
rect 41781 681186 41847 681189
rect 41492 681184 41847 681186
rect 41492 681128 41786 681184
rect 41842 681128 41847 681184
rect 41492 681126 41847 681128
rect 41781 681123 41847 681126
rect 674230 681124 674236 681188
rect 674300 681186 674306 681188
rect 674465 681186 674531 681189
rect 674300 681184 674531 681186
rect 674300 681128 674470 681184
rect 674526 681128 674531 681184
rect 674300 681126 674531 681128
rect 674300 681124 674306 681126
rect 674465 681123 674531 681126
rect 41965 680778 42031 680781
rect 41492 680776 42031 680778
rect 41492 680720 41970 680776
rect 42026 680720 42031 680776
rect 41492 680718 42031 680720
rect 41965 680715 42031 680718
rect 27429 680370 27495 680373
rect 27429 680368 27508 680370
rect 27429 680312 27434 680368
rect 27490 680312 27508 680368
rect 27429 680310 27508 680312
rect 27429 680307 27495 680310
rect 674230 680308 674236 680372
rect 674300 680370 674306 680372
rect 674598 680370 674604 680372
rect 674300 680310 674604 680370
rect 674300 680308 674306 680310
rect 674598 680308 674604 680310
rect 674668 680308 674674 680372
rect 674598 680172 674604 680236
rect 674668 680234 674674 680236
rect 675334 680234 675340 680236
rect 674668 680174 675340 680234
rect 674668 680172 674674 680174
rect 675334 680172 675340 680174
rect 675404 680172 675410 680236
rect 41781 679962 41847 679965
rect 41492 679960 41847 679962
rect 41492 679904 41786 679960
rect 41842 679904 41847 679960
rect 41492 679902 41847 679904
rect 41781 679899 41847 679902
rect 41462 679418 41522 679524
rect 41689 679418 41755 679421
rect 41462 679416 41755 679418
rect 41462 679360 41694 679416
rect 41750 679360 41755 679416
rect 41462 679358 41755 679360
rect 41689 679355 41755 679358
rect 27521 679146 27587 679149
rect 27508 679144 27587 679146
rect 27508 679088 27526 679144
rect 27582 679088 27587 679144
rect 27508 679086 27587 679088
rect 27521 679083 27587 679086
rect 41781 678738 41847 678741
rect 41492 678736 41847 678738
rect 41492 678680 41786 678736
rect 41842 678680 41847 678736
rect 41492 678678 41847 678680
rect 41781 678675 41847 678678
rect 675937 678468 676003 678469
rect 675886 678404 675892 678468
rect 675956 678466 676003 678468
rect 675956 678464 676048 678466
rect 675998 678408 676048 678464
rect 675956 678406 676048 678408
rect 675956 678404 676003 678406
rect 675937 678403 676003 678404
rect 41462 678194 41522 678300
rect 41689 678194 41755 678197
rect 41462 678192 41755 678194
rect 41462 678136 41694 678192
rect 41750 678136 41755 678192
rect 41462 678134 41755 678136
rect 41689 678131 41755 678134
rect 41462 677788 41522 677892
rect 41454 677724 41460 677788
rect 41524 677724 41530 677788
rect 30422 677076 30482 677484
rect 41454 676908 41460 676972
rect 41524 676908 41530 676972
rect 41462 676562 41522 676908
rect 41689 676562 41755 676565
rect 41462 676560 41755 676562
rect 41462 676504 41694 676560
rect 41750 676504 41755 676560
rect 41462 676502 41755 676504
rect 41689 676499 41755 676502
rect 675937 674796 676003 674797
rect 674598 674732 674604 674796
rect 674668 674794 674674 674796
rect 675334 674794 675340 674796
rect 674668 674734 675340 674794
rect 674668 674732 674674 674734
rect 675334 674732 675340 674734
rect 675404 674732 675410 674796
rect 675886 674794 675892 674796
rect 675846 674734 675892 674794
rect 675956 674792 676003 674796
rect 675998 674736 676003 674792
rect 675886 674732 675892 674734
rect 675956 674732 676003 674736
rect 675937 674731 676003 674732
rect 674230 674596 674236 674660
rect 674300 674658 674306 674660
rect 674598 674658 674604 674660
rect 674300 674598 674604 674658
rect 674300 674596 674306 674598
rect 674598 674596 674604 674598
rect 674668 674596 674674 674660
rect 674230 674052 674236 674116
rect 674300 674114 674306 674116
rect 674465 674114 674531 674117
rect 674300 674112 674531 674114
rect 674300 674056 674470 674112
rect 674526 674056 674531 674112
rect 674300 674054 674531 674056
rect 674300 674052 674306 674054
rect 674465 674051 674531 674054
rect 676262 671125 676322 671364
rect 43294 671060 43300 671124
rect 43364 671122 43370 671124
rect 43437 671122 43503 671125
rect 43364 671120 43503 671122
rect 43364 671064 43442 671120
rect 43498 671064 43503 671120
rect 43364 671062 43503 671064
rect 43364 671060 43370 671062
rect 43437 671059 43503 671062
rect 676213 671120 676322 671125
rect 676213 671064 676218 671120
rect 676274 671064 676322 671120
rect 676213 671062 676322 671064
rect 676213 671059 676279 671062
rect 42425 670986 42491 670989
rect 676029 670986 676095 670989
rect 42425 670984 44098 670986
rect 42425 670928 42430 670984
rect 42486 670928 44098 670984
rect 42425 670926 44098 670928
rect 42425 670923 42491 670926
rect 43621 670850 43687 670853
rect 43621 670848 43914 670850
rect 43621 670792 43626 670848
rect 43682 670792 43914 670848
rect 43621 670790 43914 670792
rect 43621 670787 43687 670790
rect 41965 670714 42031 670717
rect 42926 670714 42932 670716
rect 41965 670712 42932 670714
rect 41965 670656 41970 670712
rect 42026 670656 42932 670712
rect 41965 670654 42932 670656
rect 41965 670651 42031 670654
rect 42926 670652 42932 670654
rect 42996 670652 43002 670716
rect 43253 670714 43319 670717
rect 43253 670712 43546 670714
rect 43253 670656 43258 670712
rect 43314 670656 43546 670712
rect 43253 670654 43546 670656
rect 43253 670651 43319 670654
rect 42926 670516 42932 670580
rect 42996 670578 43002 670580
rect 43253 670578 43319 670581
rect 42996 670576 43319 670578
rect 42996 670520 43258 670576
rect 43314 670520 43319 670576
rect 42996 670518 43319 670520
rect 43486 670578 43546 670654
rect 43713 670578 43779 670581
rect 43854 670580 43914 670790
rect 44038 670717 44098 670926
rect 676029 670984 676292 670986
rect 676029 670928 676034 670984
rect 676090 670928 676292 670984
rect 676029 670926 676292 670928
rect 676029 670923 676095 670926
rect 44038 670712 44147 670717
rect 44038 670656 44086 670712
rect 44142 670656 44147 670712
rect 44038 670654 44147 670656
rect 44081 670651 44147 670654
rect 43486 670576 43779 670578
rect 43486 670520 43718 670576
rect 43774 670520 43779 670576
rect 43486 670518 43779 670520
rect 42996 670516 43002 670518
rect 43253 670515 43319 670518
rect 43713 670515 43779 670518
rect 43846 670516 43852 670580
rect 43916 670516 43922 670580
rect 43294 670380 43300 670444
rect 43364 670442 43370 670444
rect 43897 670442 43963 670445
rect 43364 670440 43963 670442
rect 43364 670384 43902 670440
rect 43958 670384 43963 670440
rect 43364 670382 43963 670384
rect 43364 670380 43370 670382
rect 43897 670379 43963 670382
rect 679022 670309 679082 670548
rect 678973 670304 679082 670309
rect 678973 670248 678978 670304
rect 679034 670248 679082 670304
rect 678973 670246 679082 670248
rect 679157 670306 679223 670309
rect 679157 670304 679266 670306
rect 679157 670248 679162 670304
rect 679218 670248 679266 670304
rect 678973 670243 679039 670246
rect 679157 670243 679266 670248
rect 679206 670140 679266 670243
rect 676029 669762 676095 669765
rect 676029 669760 676292 669762
rect 676029 669704 676034 669760
rect 676090 669704 676292 669760
rect 676029 669702 676292 669704
rect 676029 669699 676095 669702
rect 679065 669490 679131 669493
rect 679022 669488 679131 669490
rect 679022 669432 679070 669488
rect 679126 669432 679131 669488
rect 679022 669427 679131 669432
rect 679022 669324 679082 669427
rect 676029 668946 676095 668949
rect 676029 668944 676292 668946
rect 676029 668888 676034 668944
rect 676090 668888 676292 668944
rect 676029 668886 676292 668888
rect 676029 668883 676095 668886
rect 676213 668674 676279 668677
rect 676213 668672 676322 668674
rect 676213 668616 676218 668672
rect 676274 668616 676322 668672
rect 676213 668611 676322 668616
rect 676262 668508 676322 668611
rect 675477 668130 675543 668133
rect 675477 668128 676292 668130
rect 675477 668072 675482 668128
rect 675538 668072 676292 668128
rect 675477 668070 676292 668072
rect 675477 668067 675543 668070
rect 679249 667858 679315 667861
rect 679206 667856 679315 667858
rect 679206 667800 679254 667856
rect 679310 667800 679315 667856
rect 679206 667795 679315 667800
rect 679206 667692 679266 667795
rect 675385 667314 675451 667317
rect 675385 667312 676292 667314
rect 675385 667256 675390 667312
rect 675446 667256 676292 667312
rect 675385 667254 676292 667256
rect 675385 667251 675451 667254
rect 674230 666844 674236 666908
rect 674300 666906 674306 666908
rect 674300 666846 676292 666906
rect 674300 666844 674306 666846
rect 675293 666498 675359 666501
rect 675293 666496 676292 666498
rect 675293 666440 675298 666496
rect 675354 666440 676292 666496
rect 675293 666438 676292 666440
rect 675293 666435 675359 666438
rect 675334 666028 675340 666092
rect 675404 666090 675410 666092
rect 675404 666030 676292 666090
rect 675404 666028 675410 666030
rect 674598 665620 674604 665684
rect 674668 665682 674674 665684
rect 674668 665622 676292 665682
rect 674668 665620 674674 665622
rect 43069 665274 43135 665277
rect 43846 665274 43852 665276
rect 43069 665272 43852 665274
rect 43069 665216 43074 665272
rect 43130 665216 43852 665272
rect 43069 665214 43852 665216
rect 43069 665211 43135 665214
rect 43846 665212 43852 665214
rect 43916 665212 43922 665276
rect 676029 665274 676095 665277
rect 676029 665272 676292 665274
rect 676029 665216 676034 665272
rect 676090 665216 676292 665272
rect 676029 665214 676292 665216
rect 676029 665211 676095 665214
rect 676029 664866 676095 664869
rect 676029 664864 676292 664866
rect 676029 664808 676034 664864
rect 676090 664808 676292 664864
rect 676029 664806 676292 664808
rect 676029 664803 676095 664806
rect 675702 664396 675708 664460
rect 675772 664458 675778 664460
rect 675772 664398 676292 664458
rect 675772 664396 675778 664398
rect 673494 663988 673500 664052
rect 673564 664050 673570 664052
rect 673564 663990 676292 664050
rect 673564 663988 673570 663990
rect 674782 663580 674788 663644
rect 674852 663642 674858 663644
rect 674852 663582 676292 663642
rect 674852 663580 674858 663582
rect 676029 663234 676095 663237
rect 676029 663232 676292 663234
rect 676029 663176 676034 663232
rect 676090 663176 676292 663232
rect 676029 663174 676292 663176
rect 676029 663171 676095 663174
rect 676029 662826 676095 662829
rect 676029 662824 676292 662826
rect 676029 662768 676034 662824
rect 676090 662768 676292 662824
rect 676029 662766 676292 662768
rect 676029 662763 676095 662766
rect 677358 662492 677364 662556
rect 677428 662492 677434 662556
rect 677366 662388 677426 662492
rect 676990 662084 676996 662148
rect 677060 662084 677066 662148
rect 676998 661980 677058 662084
rect 676029 661602 676095 661605
rect 676029 661600 676292 661602
rect 676029 661544 676034 661600
rect 676090 661544 676292 661600
rect 676029 661542 676292 661544
rect 676029 661539 676095 661542
rect 60641 661194 60707 661197
rect 60641 661192 64706 661194
rect 60641 661136 60646 661192
rect 60702 661136 64706 661192
rect 60641 661134 64706 661136
rect 60641 661131 60707 661134
rect 64646 660638 64706 661134
rect 679022 660925 679082 661164
rect 678973 660920 679082 660925
rect 678973 660864 678978 660920
rect 679034 660864 679082 660920
rect 678973 660862 679082 660864
rect 678973 660859 679039 660862
rect 684542 660348 684602 660756
rect 678973 660106 679039 660109
rect 678973 660104 679082 660106
rect 678973 660048 678978 660104
rect 679034 660048 679082 660104
rect 678973 660043 679082 660048
rect 679022 659940 679082 660043
rect 58525 659562 58591 659565
rect 58525 659560 64706 659562
rect 58525 659504 58530 659560
rect 58586 659504 64706 659560
rect 58525 659502 64706 659504
rect 58525 659499 58591 659502
rect 64646 659456 64706 659502
rect 58433 658882 58499 658885
rect 58433 658880 64706 658882
rect 58433 658824 58438 658880
rect 58494 658824 64706 658880
rect 58433 658822 64706 658824
rect 58433 658819 58499 658822
rect 64646 658274 64706 658822
rect 58617 657658 58683 657661
rect 58617 657656 64706 657658
rect 58617 657600 58622 657656
rect 58678 657600 64706 657656
rect 58617 657598 64706 657600
rect 58617 657595 58683 657598
rect 64646 657092 64706 657598
rect 58433 656570 58499 656573
rect 58433 656568 64706 656570
rect 58433 656512 58438 656568
rect 58494 656512 64706 656568
rect 58433 656510 64706 656512
rect 58433 656507 58499 656510
rect 64646 655910 64706 656510
rect 58065 655346 58131 655349
rect 58065 655344 64706 655346
rect 58065 655288 58070 655344
rect 58126 655288 64706 655344
rect 58065 655286 64706 655288
rect 58065 655283 58131 655286
rect 64646 654728 64706 655286
rect 675661 652628 675727 652629
rect 675661 652624 675708 652628
rect 675772 652626 675778 652628
rect 675661 652568 675666 652624
rect 675661 652564 675708 652568
rect 675772 652566 675818 652626
rect 675772 652564 675778 652566
rect 675661 652563 675727 652564
rect 675150 652156 675156 652220
rect 675220 652218 675226 652220
rect 675477 652218 675543 652221
rect 675220 652216 675543 652218
rect 675220 652160 675482 652216
rect 675538 652160 675543 652216
rect 675220 652158 675543 652160
rect 675220 652156 675226 652158
rect 675477 652155 675543 652158
rect 675385 651676 675451 651677
rect 675334 651674 675340 651676
rect 675294 651614 675340 651674
rect 675404 651672 675451 651676
rect 675446 651616 675451 651672
rect 675334 651612 675340 651614
rect 675404 651612 675451 651616
rect 675385 651611 675451 651612
rect 674966 648892 674972 648956
rect 675036 648954 675042 648956
rect 675385 648954 675451 648957
rect 675036 648952 675451 648954
rect 675036 648896 675390 648952
rect 675446 648896 675451 648952
rect 675036 648894 675451 648896
rect 675036 648892 675042 648894
rect 675385 648891 675451 648894
rect 673494 648620 673500 648684
rect 673564 648682 673570 648684
rect 675385 648682 675451 648685
rect 673564 648680 675451 648682
rect 673564 648624 675390 648680
rect 675446 648624 675451 648680
rect 673564 648622 675451 648624
rect 673564 648620 673570 648622
rect 675385 648619 675451 648622
rect 41462 644741 41522 644912
rect 41462 644736 41571 644741
rect 41462 644680 41510 644736
rect 41566 644680 41571 644736
rect 41462 644678 41571 644680
rect 41505 644675 41571 644678
rect 41462 644333 41522 644504
rect 41462 644328 41571 644333
rect 41462 644272 41510 644328
rect 41566 644272 41571 644328
rect 41462 644270 41571 644272
rect 41505 644267 41571 644270
rect 41781 644126 41847 644129
rect 41492 644124 41847 644126
rect 41492 644068 41786 644124
rect 41842 644068 41847 644124
rect 41492 644066 41847 644068
rect 41781 644063 41847 644066
rect 41505 643922 41571 643925
rect 41462 643920 41571 643922
rect 41462 643864 41510 643920
rect 41566 643864 41571 643920
rect 41462 643859 41571 643864
rect 41462 643688 41522 643859
rect 41781 643310 41847 643313
rect 41492 643308 41847 643310
rect 41492 643252 41786 643308
rect 41842 643252 41847 643308
rect 41492 643250 41847 643252
rect 41781 643247 41847 643250
rect 649950 643242 650010 643558
rect 655513 643242 655579 643245
rect 649950 643240 655579 643242
rect 649950 643184 655518 643240
rect 655574 643184 655579 643240
rect 649950 643182 655579 643184
rect 655513 643179 655579 643182
rect 41505 643106 41571 643109
rect 41462 643104 41571 643106
rect 41462 643048 41510 643104
rect 41566 643048 41571 643104
rect 41462 643043 41571 643048
rect 41462 642872 41522 643043
rect 41462 642290 41522 642464
rect 41597 642290 41663 642293
rect 41462 642288 41663 642290
rect 41462 642232 41602 642288
rect 41658 642232 41663 642288
rect 41462 642230 41663 642232
rect 41597 642227 41663 642230
rect 41781 642086 41847 642089
rect 41492 642084 41847 642086
rect 41492 642028 41786 642084
rect 41842 642028 41847 642084
rect 41492 642026 41847 642028
rect 41781 642023 41847 642026
rect 649950 641882 650010 642376
rect 655881 641882 655947 641885
rect 649950 641880 655947 641882
rect 649950 641824 655886 641880
rect 655942 641824 655947 641880
rect 649950 641822 655947 641824
rect 655881 641819 655947 641822
rect 674782 641684 674788 641748
rect 674852 641746 674858 641748
rect 676070 641746 676076 641748
rect 674852 641686 676076 641746
rect 674852 641684 674858 641686
rect 676070 641684 676076 641686
rect 676140 641684 676146 641748
rect 41781 641678 41847 641681
rect 41492 641676 41847 641678
rect 41492 641620 41786 641676
rect 41842 641620 41847 641676
rect 41492 641618 41847 641620
rect 41781 641615 41847 641618
rect 674598 641548 674604 641612
rect 674668 641610 674674 641612
rect 675886 641610 675892 641612
rect 674668 641550 675892 641610
rect 674668 641548 674674 641550
rect 675886 641548 675892 641550
rect 675956 641548 675962 641612
rect 41505 641474 41571 641477
rect 41462 641472 41571 641474
rect 41462 641416 41510 641472
rect 41566 641416 41571 641472
rect 41462 641411 41571 641416
rect 41462 641240 41522 641411
rect 41462 640661 41522 640832
rect 41462 640656 41571 640661
rect 41462 640600 41510 640656
rect 41566 640600 41571 640656
rect 41462 640598 41571 640600
rect 649950 640658 650010 641194
rect 656065 640658 656131 640661
rect 649950 640656 656131 640658
rect 649950 640600 656070 640656
rect 656126 640600 656131 640656
rect 649950 640598 656131 640600
rect 41505 640595 41571 640598
rect 656065 640595 656131 640598
rect 41781 640454 41847 640457
rect 41492 640452 41847 640454
rect 41492 640396 41786 640452
rect 41842 640396 41847 640452
rect 41492 640394 41847 640396
rect 41781 640391 41847 640394
rect 655697 640250 655763 640253
rect 649950 640248 655763 640250
rect 649950 640192 655702 640248
rect 655758 640192 655763 640248
rect 649950 640190 655763 640192
rect 41462 639978 41522 640016
rect 649950 640012 650010 640190
rect 655697 640187 655763 640190
rect 673453 640250 673519 640253
rect 673862 640250 673868 640252
rect 673453 640248 673868 640250
rect 673453 640192 673458 640248
rect 673514 640192 673868 640248
rect 673453 640190 673868 640192
rect 673453 640187 673519 640190
rect 673862 640188 673868 640190
rect 673932 640188 673938 640252
rect 42333 639978 42399 639981
rect 41462 639976 42399 639978
rect 41462 639920 42338 639976
rect 42394 639920 42399 639976
rect 41462 639918 42399 639920
rect 42333 639915 42399 639918
rect 41462 639437 41522 639608
rect 41462 639432 41571 639437
rect 654409 639434 654475 639437
rect 41462 639376 41510 639432
rect 41566 639376 41571 639432
rect 41462 639374 41571 639376
rect 41505 639371 41571 639374
rect 649950 639432 654475 639434
rect 649950 639376 654414 639432
rect 654470 639376 654475 639432
rect 649950 639374 654475 639376
rect 41462 639029 41522 639200
rect 41462 639024 41571 639029
rect 41462 638968 41510 639024
rect 41566 638968 41571 639024
rect 41462 638966 41571 638968
rect 41505 638963 41571 638966
rect 649950 638830 650010 639374
rect 654409 639371 654475 639374
rect 41781 638822 41847 638825
rect 41492 638820 41847 638822
rect 41492 638764 41786 638820
rect 41842 638764 41847 638820
rect 41492 638762 41847 638764
rect 41781 638759 41847 638762
rect 41781 638414 41847 638417
rect 41492 638412 41847 638414
rect 41492 638356 41786 638412
rect 41842 638356 41847 638412
rect 41492 638354 41847 638356
rect 41781 638351 41847 638354
rect 656433 638210 656499 638213
rect 675753 638212 675819 638213
rect 675702 638210 675708 638212
rect 649950 638208 656499 638210
rect 649950 638152 656438 638208
rect 656494 638152 656499 638208
rect 649950 638150 656499 638152
rect 675662 638150 675708 638210
rect 675772 638208 675819 638212
rect 675814 638152 675819 638208
rect 41462 637805 41522 637976
rect 41462 637800 41571 637805
rect 41462 637744 41510 637800
rect 41566 637744 41571 637800
rect 41462 637742 41571 637744
rect 41505 637739 41571 637742
rect 649950 637648 650010 638150
rect 656433 638147 656499 638150
rect 675702 638148 675708 638150
rect 675772 638148 675819 638152
rect 675753 638147 675819 638148
rect 673545 637666 673611 637669
rect 675334 637666 675340 637668
rect 673545 637664 675340 637666
rect 673545 637608 673550 637664
rect 673606 637608 675340 637664
rect 673545 637606 675340 637608
rect 673545 637603 673611 637606
rect 675334 637604 675340 637606
rect 675404 637604 675410 637668
rect 41873 637598 41939 637601
rect 41492 637596 41939 637598
rect 41492 637540 41878 637596
rect 41934 637540 41939 637596
rect 41492 637538 41939 637540
rect 41873 637535 41939 637538
rect 38150 636989 38210 637160
rect 38101 636984 38210 636989
rect 38101 636928 38106 636984
rect 38162 636928 38210 636984
rect 38101 636926 38210 636928
rect 38101 636923 38167 636926
rect 41462 636581 41522 636752
rect 41462 636576 41571 636581
rect 41462 636520 41510 636576
rect 41566 636520 41571 636576
rect 41462 636518 41571 636520
rect 41505 636515 41571 636518
rect 41462 636170 41522 636344
rect 41597 636170 41663 636173
rect 41462 636168 41663 636170
rect 41462 636112 41602 636168
rect 41658 636112 41663 636168
rect 41462 636110 41663 636112
rect 41597 636107 41663 636110
rect 38150 635765 38210 635936
rect 38150 635760 38259 635765
rect 38150 635704 38198 635760
rect 38254 635704 38259 635760
rect 38150 635702 38259 635704
rect 38193 635699 38259 635702
rect 41462 635354 41522 635528
rect 41597 635354 41663 635357
rect 41462 635352 41663 635354
rect 41462 635296 41602 635352
rect 41658 635296 41663 635352
rect 41462 635294 41663 635296
rect 41597 635291 41663 635294
rect 41462 634946 41522 635120
rect 41597 634946 41663 634949
rect 41462 634944 41663 634946
rect 41462 634888 41602 634944
rect 41658 634888 41663 634944
rect 41462 634886 41663 634888
rect 41597 634883 41663 634886
rect 41462 634541 41522 634712
rect 41462 634536 41571 634541
rect 41462 634480 41510 634536
rect 41566 634480 41571 634536
rect 41462 634478 41571 634480
rect 41505 634475 41571 634478
rect 30422 633896 30482 634304
rect 41462 633317 41522 633488
rect 41462 633312 41571 633317
rect 41462 633256 41510 633312
rect 41566 633256 41571 633312
rect 41462 633254 41571 633256
rect 41505 633251 41571 633254
rect 43897 632090 43963 632093
rect 43854 632088 43963 632090
rect 43854 632032 43902 632088
rect 43958 632032 43963 632088
rect 43854 632027 43963 632032
rect 41689 631954 41755 631957
rect 43854 631954 43914 632027
rect 41689 631952 43914 631954
rect 41689 631896 41694 631952
rect 41750 631896 43914 631952
rect 41689 631894 43914 631896
rect 41689 631891 41755 631894
rect 673545 629370 673611 629373
rect 674782 629370 674788 629372
rect 673545 629368 674788 629370
rect 673545 629312 673550 629368
rect 673606 629312 674788 629368
rect 673545 629310 674788 629312
rect 673545 629307 673611 629310
rect 674782 629308 674788 629310
rect 674852 629308 674858 629372
rect 41781 627468 41847 627469
rect 42425 627468 42491 627469
rect 41781 627464 41828 627468
rect 41892 627466 41898 627468
rect 42374 627466 42380 627468
rect 41781 627408 41786 627464
rect 41781 627404 41828 627408
rect 41892 627406 41938 627466
rect 42334 627406 42380 627466
rect 42444 627464 42491 627468
rect 42486 627408 42491 627464
rect 41892 627404 41898 627406
rect 42374 627404 42380 627406
rect 42444 627404 42491 627408
rect 41781 627403 41847 627404
rect 42425 627403 42491 627404
rect 679022 626109 679082 626348
rect 678973 626104 679082 626109
rect 678973 626048 678978 626104
rect 679034 626048 679082 626104
rect 678973 626046 679082 626048
rect 678973 626043 679039 626046
rect 676262 625701 676322 625940
rect 676213 625696 676322 625701
rect 676213 625640 676218 625696
rect 676274 625640 676322 625696
rect 676213 625638 676322 625640
rect 676213 625635 676279 625638
rect 676121 625290 676187 625293
rect 676262 625290 676322 625532
rect 679065 625290 679131 625293
rect 676121 625288 676322 625290
rect 676121 625232 676126 625288
rect 676182 625232 676322 625288
rect 676121 625230 676322 625232
rect 679022 625288 679131 625290
rect 679022 625232 679070 625288
rect 679126 625232 679131 625288
rect 676121 625227 676187 625230
rect 679022 625227 679131 625232
rect 679022 625124 679082 625227
rect 675293 624746 675359 624749
rect 675293 624744 676292 624746
rect 675293 624688 675298 624744
rect 675354 624688 676292 624744
rect 675293 624686 676292 624688
rect 675293 624683 675359 624686
rect 679157 624474 679223 624477
rect 679157 624472 679266 624474
rect 679157 624416 679162 624472
rect 679218 624416 679266 624472
rect 679157 624411 679266 624416
rect 679206 624308 679266 624411
rect 676029 623930 676095 623933
rect 676029 623928 676292 623930
rect 676029 623872 676034 623928
rect 676090 623872 676292 623928
rect 676029 623870 676292 623872
rect 676029 623867 676095 623870
rect 679249 623658 679315 623661
rect 679206 623656 679315 623658
rect 679206 623600 679254 623656
rect 679310 623600 679315 623656
rect 679206 623595 679315 623600
rect 679206 623492 679266 623595
rect 677550 622844 677610 623084
rect 677542 622780 677548 622844
rect 677612 622780 677618 622844
rect 679341 622842 679407 622845
rect 679341 622840 679450 622842
rect 679341 622784 679346 622840
rect 679402 622784 679450 622840
rect 679341 622779 679450 622784
rect 679390 622676 679450 622779
rect 676262 622029 676322 622268
rect 42057 622026 42123 622029
rect 42374 622026 42380 622028
rect 42057 622024 42380 622026
rect 42057 621968 42062 622024
rect 42118 621968 42380 622024
rect 42057 621966 42380 621968
rect 42057 621963 42123 621966
rect 42374 621964 42380 621966
rect 42444 621964 42450 622028
rect 676213 622024 676322 622029
rect 676213 621968 676218 622024
rect 676274 621968 676322 622024
rect 676213 621966 676322 621968
rect 676213 621963 676279 621966
rect 676806 621964 676812 622028
rect 676876 621964 676882 622028
rect 676814 621860 676874 621964
rect 41873 621484 41939 621485
rect 41822 621420 41828 621484
rect 41892 621482 41939 621484
rect 676029 621482 676095 621485
rect 41892 621480 41984 621482
rect 41934 621424 41984 621480
rect 41892 621422 41984 621424
rect 676029 621480 676292 621482
rect 676029 621424 676034 621480
rect 676090 621424 676292 621480
rect 676029 621422 676292 621424
rect 41892 621420 41939 621422
rect 41873 621419 41939 621420
rect 676029 621419 676095 621422
rect 676029 621074 676095 621077
rect 676029 621072 676292 621074
rect 676029 621016 676034 621072
rect 676090 621016 676292 621072
rect 676029 621014 676292 621016
rect 676029 621011 676095 621014
rect 674414 620604 674420 620668
rect 674484 620666 674490 620668
rect 674484 620606 676292 620666
rect 674484 620604 674490 620606
rect 673678 620196 673684 620260
rect 673748 620258 673754 620260
rect 673748 620198 676292 620258
rect 673748 620196 673754 620198
rect 676029 619850 676095 619853
rect 676029 619848 676292 619850
rect 676029 619792 676034 619848
rect 676090 619792 676292 619848
rect 676029 619790 676292 619792
rect 676029 619787 676095 619790
rect 674598 619380 674604 619444
rect 674668 619442 674674 619444
rect 674668 619382 676292 619442
rect 674668 619380 674674 619382
rect 674046 618972 674052 619036
rect 674116 619034 674122 619036
rect 674116 618974 676292 619034
rect 674116 618972 674122 618974
rect 676642 618700 676648 618764
rect 676712 618700 676718 618764
rect 676650 618596 676710 618700
rect 676029 618218 676095 618221
rect 676029 618216 676292 618218
rect 676029 618160 676034 618216
rect 676090 618160 676292 618216
rect 676029 618158 676292 618160
rect 676029 618155 676095 618158
rect 676121 617946 676187 617949
rect 676121 617944 676322 617946
rect 676121 617888 676126 617944
rect 676182 617888 676322 617944
rect 676121 617886 676322 617888
rect 676121 617883 676187 617886
rect 58157 617810 58223 617813
rect 58157 617808 64706 617810
rect 58157 617752 58162 617808
rect 58218 617752 64706 617808
rect 676262 617780 676322 617886
rect 58157 617750 64706 617752
rect 58157 617747 58223 617750
rect 64646 617416 64706 617750
rect 677174 617476 677180 617540
rect 677244 617476 677250 617540
rect 677182 617372 677242 617476
rect 675201 617130 675267 617133
rect 677358 617130 677364 617132
rect 675201 617128 677364 617130
rect 675201 617072 675206 617128
rect 675262 617072 677364 617128
rect 675201 617070 677364 617072
rect 675201 617067 675267 617070
rect 677358 617068 677364 617070
rect 677428 617068 677434 617132
rect 674230 616932 674236 616996
rect 674300 616994 674306 616996
rect 674300 616934 676292 616994
rect 674300 616932 674306 616934
rect 58525 616858 58591 616861
rect 58525 616856 64706 616858
rect 58525 616800 58530 616856
rect 58586 616800 64706 616856
rect 58525 616798 64706 616800
rect 58525 616795 58591 616798
rect 64646 616234 64706 616798
rect 676029 616586 676095 616589
rect 676029 616584 676292 616586
rect 676029 616528 676034 616584
rect 676090 616528 676292 616584
rect 676029 616526 676292 616528
rect 676029 616523 676095 616526
rect 679022 615909 679082 616148
rect 678973 615904 679082 615909
rect 678973 615848 678978 615904
rect 679034 615848 679082 615904
rect 678973 615846 679082 615848
rect 678973 615843 679039 615846
rect 58525 615498 58591 615501
rect 58525 615496 64706 615498
rect 58525 615440 58530 615496
rect 58586 615440 64706 615496
rect 58525 615438 64706 615440
rect 58525 615435 58591 615438
rect 64646 615052 64706 615438
rect 679022 615332 679082 615740
rect 678973 615090 679039 615093
rect 678973 615088 679082 615090
rect 678973 615032 678978 615088
rect 679034 615032 679082 615088
rect 678973 615027 679082 615032
rect 679022 614924 679082 615027
rect 58157 614546 58223 614549
rect 58157 614544 64706 614546
rect 58157 614488 58162 614544
rect 58218 614488 64706 614544
rect 58157 614486 64706 614488
rect 58157 614483 58223 614486
rect 64646 613870 64706 614486
rect 58525 612642 58591 612645
rect 64646 612642 64706 612688
rect 58525 612640 64706 612642
rect 58525 612584 58530 612640
rect 58586 612584 64706 612640
rect 58525 612582 64706 612584
rect 58525 612579 58591 612582
rect 58341 612098 58407 612101
rect 58341 612096 64706 612098
rect 58341 612040 58346 612096
rect 58402 612040 64706 612096
rect 58341 612038 64706 612040
rect 58341 612035 58407 612038
rect 64646 611506 64706 612038
rect 673729 609242 673795 609245
rect 676662 609242 676668 609244
rect 673729 609240 676668 609242
rect 673729 609184 673734 609240
rect 673790 609184 676668 609240
rect 673729 609182 676668 609184
rect 673729 609179 673795 609182
rect 676662 609180 676668 609182
rect 676732 609180 676738 609244
rect 673678 607820 673684 607884
rect 673748 607882 673754 607884
rect 675385 607882 675451 607885
rect 673748 607880 675451 607882
rect 673748 607824 675390 607880
rect 675446 607824 675451 607880
rect 673748 607822 675451 607824
rect 673748 607820 673754 607822
rect 675385 607819 675451 607822
rect 675753 607338 675819 607341
rect 676070 607338 676076 607340
rect 675753 607336 676076 607338
rect 675753 607280 675758 607336
rect 675814 607280 676076 607336
rect 675753 607278 676076 607280
rect 675753 607275 675819 607278
rect 676070 607276 676076 607278
rect 676140 607276 676146 607340
rect 674230 604964 674236 605028
rect 674300 605026 674306 605028
rect 675201 605026 675267 605029
rect 674300 605024 675267 605026
rect 674300 604968 675206 605024
rect 675262 604968 675267 605024
rect 674300 604966 675267 604968
rect 674300 604964 674306 604966
rect 675201 604963 675267 604966
rect 674598 604420 674604 604484
rect 674668 604482 674674 604484
rect 675109 604482 675175 604485
rect 674668 604480 675175 604482
rect 674668 604424 675114 604480
rect 675170 604424 675175 604480
rect 674668 604422 675175 604424
rect 674668 604420 674674 604422
rect 675109 604419 675175 604422
rect 675293 604484 675359 604485
rect 675293 604480 675340 604484
rect 675404 604482 675410 604484
rect 675293 604424 675298 604480
rect 675293 604420 675340 604424
rect 675404 604422 675450 604482
rect 675404 604420 675410 604422
rect 675293 604419 675359 604420
rect 674414 603740 674420 603804
rect 674484 603802 674490 603804
rect 675109 603802 675175 603805
rect 674484 603800 675175 603802
rect 674484 603744 675114 603800
rect 675170 603744 675175 603800
rect 674484 603742 675175 603744
rect 674484 603740 674490 603742
rect 675109 603739 675175 603742
rect 673862 601836 673868 601900
rect 673932 601898 673938 601900
rect 675109 601898 675175 601901
rect 673932 601896 675175 601898
rect 673932 601840 675114 601896
rect 675170 601840 675175 601896
rect 673932 601838 675175 601840
rect 673932 601836 673938 601838
rect 675109 601835 675175 601838
rect 41781 601762 41847 601765
rect 41492 601760 41847 601762
rect 41492 601704 41786 601760
rect 41842 601704 41847 601760
rect 41492 601702 41847 601704
rect 41781 601699 41847 601702
rect 41781 601354 41847 601357
rect 41492 601352 41847 601354
rect 41492 601296 41786 601352
rect 41842 601296 41847 601352
rect 41492 601294 41847 601296
rect 41781 601291 41847 601294
rect 41781 600946 41847 600949
rect 41492 600944 41847 600946
rect 41492 600888 41786 600944
rect 41842 600888 41847 600944
rect 41492 600886 41847 600888
rect 41781 600883 41847 600886
rect 41505 600674 41571 600677
rect 41462 600672 41571 600674
rect 41462 600616 41510 600672
rect 41566 600616 41571 600672
rect 41462 600611 41571 600616
rect 41462 600508 41522 600611
rect 41781 600130 41847 600133
rect 41492 600128 41847 600130
rect 41492 600072 41786 600128
rect 41842 600072 41847 600128
rect 41492 600070 41847 600072
rect 41781 600067 41847 600070
rect 41505 599858 41571 599861
rect 41462 599856 41571 599858
rect 41462 599800 41510 599856
rect 41566 599800 41571 599856
rect 41462 599795 41571 599800
rect 41462 599692 41522 599795
rect 41462 599045 41522 599284
rect 41462 599040 41571 599045
rect 41462 598984 41510 599040
rect 41566 598984 41571 599040
rect 41462 598982 41571 598984
rect 41505 598979 41571 598982
rect 41781 598906 41847 598909
rect 41492 598904 41847 598906
rect 41492 598848 41786 598904
rect 41842 598848 41847 598904
rect 41492 598846 41847 598848
rect 41781 598843 41847 598846
rect 42425 598498 42491 598501
rect 41492 598496 42491 598498
rect 41492 598440 42430 598496
rect 42486 598440 42491 598496
rect 41492 598438 42491 598440
rect 42425 598435 42491 598438
rect 41505 598226 41571 598229
rect 41462 598224 41571 598226
rect 41462 598168 41510 598224
rect 41566 598168 41571 598224
rect 41462 598163 41571 598168
rect 41462 598060 41522 598163
rect 649950 597818 650010 598336
rect 655973 597818 656039 597821
rect 649950 597816 656039 597818
rect 649950 597760 655978 597816
rect 656034 597760 656039 597816
rect 649950 597758 656039 597760
rect 655973 597755 656039 597758
rect 41462 597413 41522 597652
rect 41462 597408 41571 597413
rect 41462 597352 41510 597408
rect 41566 597352 41571 597408
rect 41462 597350 41571 597352
rect 41505 597347 41571 597350
rect 41462 597005 41522 597244
rect 41462 597000 41571 597005
rect 41462 596944 41510 597000
rect 41566 596944 41571 597000
rect 41462 596942 41571 596944
rect 41505 596939 41571 596942
rect 41462 596597 41522 596836
rect 41462 596592 41571 596597
rect 41462 596536 41510 596592
rect 41566 596536 41571 596592
rect 41462 596534 41571 596536
rect 649950 596594 650010 597154
rect 655697 596594 655763 596597
rect 649950 596592 655763 596594
rect 649950 596536 655702 596592
rect 655758 596536 655763 596592
rect 649950 596534 655763 596536
rect 41505 596531 41571 596534
rect 655697 596531 655763 596534
rect 42149 596458 42215 596461
rect 41492 596456 42215 596458
rect 41492 596400 42154 596456
rect 42210 596400 42215 596456
rect 41492 596398 42215 596400
rect 42149 596395 42215 596398
rect 41462 595781 41522 596020
rect 41462 595776 41571 595781
rect 41462 595720 41510 595776
rect 41566 595720 41571 595776
rect 41462 595718 41571 595720
rect 41505 595715 41571 595718
rect 41462 595373 41522 595612
rect 649950 595506 650010 595972
rect 655789 595506 655855 595509
rect 649950 595504 655855 595506
rect 649950 595448 655794 595504
rect 655850 595448 655855 595504
rect 649950 595446 655855 595448
rect 655789 595443 655855 595446
rect 41462 595368 41571 595373
rect 655421 595370 655487 595373
rect 41462 595312 41510 595368
rect 41566 595312 41571 595368
rect 41462 595310 41571 595312
rect 41505 595307 41571 595310
rect 649950 595368 655487 595370
rect 649950 595312 655426 595368
rect 655482 595312 655487 595368
rect 649950 595310 655487 595312
rect 41873 595234 41939 595237
rect 41492 595232 41939 595234
rect 41492 595176 41878 595232
rect 41934 595176 41939 595232
rect 41492 595174 41939 595176
rect 41873 595171 41939 595174
rect 41462 594557 41522 594796
rect 649950 594790 650010 595310
rect 655421 595307 655487 595310
rect 41462 594552 41571 594557
rect 41462 594496 41510 594552
rect 41566 594496 41571 594552
rect 41462 594494 41571 594496
rect 41505 594491 41571 594494
rect 37966 594149 38026 594388
rect 655237 594282 655303 594285
rect 649950 594280 655303 594282
rect 649950 594224 655242 594280
rect 655298 594224 655303 594280
rect 649950 594222 655303 594224
rect 37966 594144 38075 594149
rect 37966 594088 38014 594144
rect 38070 594088 38075 594144
rect 37966 594086 38075 594088
rect 38009 594083 38075 594086
rect 38150 593741 38210 593980
rect 38101 593736 38210 593741
rect 38101 593680 38106 593736
rect 38162 593680 38210 593736
rect 38101 593678 38210 593680
rect 38101 593675 38167 593678
rect 649950 593608 650010 594222
rect 655237 594219 655303 594222
rect 41781 593602 41847 593605
rect 41492 593600 41847 593602
rect 41492 593544 41786 593600
rect 41842 593544 41847 593600
rect 41492 593542 41847 593544
rect 41781 593539 41847 593542
rect 673729 593602 673795 593605
rect 673729 593600 675218 593602
rect 673729 593544 673734 593600
rect 673790 593544 675218 593600
rect 673729 593542 675218 593544
rect 673729 593539 673795 593542
rect 675158 593194 675218 593542
rect 675569 593194 675635 593197
rect 675158 593192 675635 593194
rect 41462 592925 41522 593164
rect 675158 593136 675574 593192
rect 675630 593136 675635 593192
rect 675158 593134 675635 593136
rect 675569 593131 675635 593134
rect 655605 593058 655671 593061
rect 649950 593056 655671 593058
rect 649950 593000 655610 593056
rect 655666 593000 655671 593056
rect 649950 592998 655671 593000
rect 41462 592920 41571 592925
rect 41462 592864 41510 592920
rect 41566 592864 41571 592920
rect 41462 592862 41571 592864
rect 41505 592859 41571 592862
rect 41462 592514 41522 592756
rect 41689 592514 41755 592517
rect 41462 592512 41755 592514
rect 41462 592456 41694 592512
rect 41750 592456 41755 592512
rect 41462 592454 41755 592456
rect 41689 592451 41755 592454
rect 649950 592426 650010 592998
rect 655605 592995 655671 592998
rect 41462 592109 41522 592348
rect 41462 592104 41571 592109
rect 41462 592048 41510 592104
rect 41566 592048 41571 592104
rect 41462 592046 41571 592048
rect 41505 592043 41571 592046
rect 41462 591701 41522 591940
rect 41462 591696 41571 591701
rect 41462 591640 41510 591696
rect 41566 591640 41571 591696
rect 41462 591638 41571 591640
rect 41505 591635 41571 591638
rect 41462 591293 41522 591532
rect 41413 591288 41522 591293
rect 41413 591232 41418 591288
rect 41474 591232 41522 591288
rect 41413 591230 41522 591232
rect 41413 591227 41479 591230
rect 30422 590716 30482 591124
rect 41462 590069 41522 590308
rect 41462 590064 41571 590069
rect 41462 590008 41510 590064
rect 41566 590008 41571 590064
rect 41462 590006 41571 590008
rect 41505 590003 41571 590006
rect 674046 587964 674052 588028
rect 674116 588026 674122 588028
rect 675150 588026 675156 588028
rect 674116 587966 675156 588026
rect 674116 587964 674122 587966
rect 675150 587964 675156 587966
rect 675220 587964 675226 588028
rect 676029 587756 676095 587757
rect 676029 587754 676076 587756
rect 675984 587752 676076 587754
rect 675984 587696 676034 587752
rect 675984 587694 676076 587696
rect 676029 587692 676076 587694
rect 676140 587692 676146 587756
rect 676029 587691 676095 587692
rect 676029 586260 676095 586261
rect 676029 586256 676076 586260
rect 676140 586258 676146 586260
rect 676029 586200 676034 586256
rect 676029 586196 676076 586200
rect 676140 586198 676186 586258
rect 676140 586196 676146 586198
rect 676029 586195 676095 586196
rect 42190 585244 42196 585308
rect 42260 585306 42266 585308
rect 42333 585306 42399 585309
rect 42260 585304 42399 585306
rect 42260 585248 42338 585304
rect 42394 585248 42399 585304
rect 42260 585246 42399 585248
rect 42260 585244 42266 585246
rect 42333 585243 42399 585246
rect 41781 584220 41847 584221
rect 41781 584218 41828 584220
rect 41736 584216 41828 584218
rect 41736 584160 41786 584216
rect 41736 584158 41828 584160
rect 41781 584156 41828 584158
rect 41892 584156 41898 584220
rect 41781 584155 41847 584156
rect 42701 583946 42767 583949
rect 42926 583946 42932 583948
rect 42701 583944 42932 583946
rect 42701 583888 42706 583944
rect 42762 583888 42932 583944
rect 42701 583886 42932 583888
rect 42701 583883 42767 583886
rect 42926 583884 42932 583886
rect 42996 583884 43002 583948
rect 43897 583810 43963 583813
rect 44081 583810 44147 583813
rect 43897 583808 44147 583810
rect 43897 583752 43902 583808
rect 43958 583752 44086 583808
rect 44142 583752 44147 583808
rect 43897 583750 44147 583752
rect 43897 583747 43963 583750
rect 44081 583747 44147 583750
rect 42926 581844 42932 581908
rect 42996 581906 43002 581908
rect 43161 581906 43227 581909
rect 42996 581904 43227 581906
rect 42996 581848 43166 581904
rect 43222 581848 43227 581904
rect 42996 581846 43227 581848
rect 42996 581844 43002 581846
rect 43161 581843 43227 581846
rect 676121 580954 676187 580957
rect 676262 580954 676322 581060
rect 676121 580952 676322 580954
rect 676121 580896 676126 580952
rect 676182 580896 676322 580952
rect 676121 580894 676322 580896
rect 676121 580891 676187 580894
rect 41822 580620 41828 580684
rect 41892 580682 41898 580684
rect 42241 580682 42307 580685
rect 41892 580680 42307 580682
rect 41892 580624 42246 580680
rect 42302 580624 42307 580680
rect 41892 580622 42307 580624
rect 41892 580620 41898 580622
rect 42241 580619 42307 580622
rect 676262 580549 676322 580652
rect 676262 580544 676371 580549
rect 676262 580488 676310 580544
rect 676366 580488 676371 580544
rect 676262 580486 676371 580488
rect 676305 580483 676371 580486
rect 676262 580141 676322 580244
rect 676213 580136 676322 580141
rect 676213 580080 676218 580136
rect 676274 580080 676322 580136
rect 676213 580078 676322 580080
rect 676213 580075 676279 580078
rect 676029 579866 676095 579869
rect 676029 579864 676292 579866
rect 676029 579808 676034 579864
rect 676090 579808 676292 579864
rect 676029 579806 676292 579808
rect 676029 579803 676095 579806
rect 676998 579324 677058 579428
rect 676990 579260 676996 579324
rect 677060 579260 677066 579324
rect 678973 579322 679039 579325
rect 678973 579320 679082 579322
rect 678973 579264 678978 579320
rect 679034 579264 679082 579320
rect 678973 579259 679082 579264
rect 679022 579020 679082 579259
rect 676029 578642 676095 578645
rect 676029 578640 676292 578642
rect 676029 578584 676034 578640
rect 676090 578584 676292 578640
rect 676029 578582 676292 578584
rect 676029 578579 676095 578582
rect 677542 578444 677548 578508
rect 677612 578444 677618 578508
rect 677550 578204 677610 578444
rect 677182 577692 677242 577796
rect 677174 577628 677180 577692
rect 677244 577628 677250 577692
rect 679065 577690 679131 577693
rect 679022 577688 679131 577690
rect 679022 577632 679070 577688
rect 679126 577632 679131 577688
rect 679022 577627 679131 577632
rect 679022 577388 679082 577627
rect 42149 577012 42215 577013
rect 42149 577010 42196 577012
rect 42104 577008 42196 577010
rect 42104 576952 42154 577008
rect 42104 576950 42196 576952
rect 42149 576948 42196 576950
rect 42260 576948 42266 577012
rect 42149 576947 42215 576948
rect 676814 576876 676874 576980
rect 676806 576812 676812 576876
rect 676876 576812 676882 576876
rect 674782 576540 674788 576604
rect 674852 576602 674858 576604
rect 674852 576542 676292 576602
rect 674852 576540 674858 576542
rect 675937 576194 676003 576197
rect 675937 576192 676292 576194
rect 675937 576136 675942 576192
rect 675998 576136 676292 576192
rect 675937 576134 676292 576136
rect 675937 576131 676003 576134
rect 676029 575786 676095 575789
rect 676029 575784 676292 575786
rect 676029 575728 676034 575784
rect 676090 575728 676292 575784
rect 676029 575726 676292 575728
rect 676029 575723 676095 575726
rect 675569 575378 675635 575381
rect 675569 575376 676292 575378
rect 675569 575320 675574 575376
rect 675630 575320 676292 575376
rect 675569 575318 676292 575320
rect 675569 575315 675635 575318
rect 676029 574970 676095 574973
rect 676029 574968 676292 574970
rect 676029 574912 676034 574968
rect 676090 574912 676292 574968
rect 676029 574910 676292 574912
rect 676029 574907 676095 574910
rect 58525 574834 58591 574837
rect 58525 574832 64706 574834
rect 58525 574776 58530 574832
rect 58586 574776 64706 574832
rect 58525 574774 64706 574776
rect 58525 574771 58591 574774
rect 64646 574194 64706 574774
rect 676029 574562 676095 574565
rect 676029 574560 676292 574562
rect 676029 574504 676034 574560
rect 676090 574504 676292 574560
rect 676029 574502 676292 574504
rect 676029 574499 676095 574502
rect 674046 574092 674052 574156
rect 674116 574154 674122 574156
rect 674116 574094 676292 574154
rect 674116 574092 674122 574094
rect 674966 573684 674972 573748
rect 675036 573746 675042 573748
rect 675036 573686 676292 573746
rect 675036 573684 675042 573686
rect 59261 573610 59327 573613
rect 59261 573608 64706 573610
rect 59261 573552 59266 573608
rect 59322 573552 64706 573608
rect 59261 573550 64706 573552
rect 59261 573547 59327 573550
rect 64646 573012 64706 573550
rect 673494 573276 673500 573340
rect 673564 573338 673570 573340
rect 673564 573278 676292 573338
rect 673564 573276 673570 573278
rect 676029 572930 676095 572933
rect 676029 572928 676292 572930
rect 676029 572872 676034 572928
rect 676090 572872 676292 572928
rect 676029 572870 676292 572872
rect 676029 572867 676095 572870
rect 676029 572522 676095 572525
rect 676029 572520 676292 572522
rect 676029 572464 676034 572520
rect 676090 572464 676292 572520
rect 676029 572462 676292 572464
rect 676029 572459 676095 572462
rect 60641 572386 60707 572389
rect 60641 572384 64706 572386
rect 60641 572328 60646 572384
rect 60702 572328 64706 572384
rect 60641 572326 64706 572328
rect 60641 572323 60707 572326
rect 64646 571830 64706 572326
rect 675477 572114 675543 572117
rect 675477 572112 676292 572114
rect 675477 572056 675482 572112
rect 675538 572056 676292 572112
rect 675477 572054 676292 572056
rect 675477 572051 675543 572054
rect 676662 571916 676668 571980
rect 676732 571916 676738 571980
rect 676670 571676 676730 571916
rect 677358 571508 677364 571572
rect 677428 571508 677434 571572
rect 677366 571268 677426 571508
rect 58065 571026 58131 571029
rect 58065 571024 64706 571026
rect 58065 570968 58070 571024
rect 58126 570968 64706 571024
rect 58065 570966 64706 570968
rect 58065 570963 58131 570966
rect 64646 570648 64706 570966
rect 679022 570757 679082 570860
rect 678973 570752 679082 570757
rect 678973 570696 678978 570752
rect 679034 570696 679082 570752
rect 678973 570694 679082 570696
rect 678973 570691 679039 570694
rect 58341 570074 58407 570077
rect 58341 570072 64706 570074
rect 58341 570016 58346 570072
rect 58402 570016 64706 570072
rect 684542 570044 684602 570452
rect 58341 570014 64706 570016
rect 58341 570011 58407 570014
rect 64646 569466 64706 570014
rect 678973 569938 679039 569941
rect 678973 569936 679082 569938
rect 678973 569880 678978 569936
rect 679034 569880 679082 569936
rect 678973 569875 679082 569880
rect 679022 569636 679082 569875
rect 58249 568306 58315 568309
rect 58249 568304 64706 568306
rect 58249 568248 58254 568304
rect 58310 568248 64706 568304
rect 58249 568246 64706 568248
rect 58249 568243 58315 568246
rect 675150 562396 675156 562460
rect 675220 562458 675226 562460
rect 675477 562458 675543 562461
rect 675220 562456 675543 562458
rect 675220 562400 675482 562456
rect 675538 562400 675543 562456
rect 675220 562398 675543 562400
rect 675220 562396 675226 562398
rect 675477 562395 675543 562398
rect 674046 562260 674052 562324
rect 674116 562322 674122 562324
rect 675293 562322 675359 562325
rect 674116 562320 675359 562322
rect 674116 562264 675298 562320
rect 675354 562264 675359 562320
rect 674116 562262 675359 562264
rect 674116 562260 674122 562262
rect 675293 562259 675359 562262
rect 674966 561172 674972 561236
rect 675036 561234 675042 561236
rect 675477 561234 675543 561237
rect 675036 561232 675543 561234
rect 675036 561176 675482 561232
rect 675538 561176 675543 561232
rect 675036 561174 675543 561176
rect 675036 561172 675042 561174
rect 675477 561171 675543 561174
rect 41462 558381 41522 558484
rect 41462 558376 41571 558381
rect 41462 558320 41510 558376
rect 41566 558320 41571 558376
rect 41462 558318 41571 558320
rect 41505 558315 41571 558318
rect 41462 557973 41522 558076
rect 41462 557968 41571 557973
rect 41462 557912 41510 557968
rect 41566 557912 41571 557968
rect 41462 557910 41571 557912
rect 41505 557907 41571 557910
rect 41462 557565 41522 557668
rect 41462 557560 41571 557565
rect 41462 557504 41510 557560
rect 41566 557504 41571 557560
rect 41462 557502 41571 557504
rect 41505 557499 41571 557502
rect 674782 557500 674788 557564
rect 674852 557562 674858 557564
rect 675293 557562 675359 557565
rect 674852 557560 675359 557562
rect 674852 557504 675298 557560
rect 675354 557504 675359 557560
rect 674852 557502 675359 557504
rect 674852 557500 674858 557502
rect 675293 557499 675359 557502
rect 41781 557290 41847 557293
rect 41492 557288 41847 557290
rect 41492 557232 41786 557288
rect 41842 557232 41847 557288
rect 41492 557230 41847 557232
rect 41781 557227 41847 557230
rect 41462 556746 41522 556852
rect 41638 556746 41644 556748
rect 41462 556686 41644 556746
rect 41638 556684 41644 556686
rect 41708 556684 41714 556748
rect 41781 556474 41847 556477
rect 41492 556472 41847 556474
rect 41492 556416 41786 556472
rect 41842 556416 41847 556472
rect 41492 556414 41847 556416
rect 41781 556411 41847 556414
rect 42374 556066 42380 556068
rect 41492 556006 42380 556066
rect 42374 556004 42380 556006
rect 42444 556004 42450 556068
rect 41505 555930 41571 555933
rect 41462 555928 41571 555930
rect 41462 555872 41510 555928
rect 41566 555872 41571 555928
rect 41462 555867 41571 555872
rect 41462 555628 41522 555867
rect 44030 555250 44036 555252
rect 41492 555190 44036 555250
rect 44030 555188 44036 555190
rect 44100 555188 44106 555252
rect 38518 554709 38578 554812
rect 38518 554704 38627 554709
rect 38518 554648 38566 554704
rect 38622 554648 38627 554704
rect 38518 554646 38627 554648
rect 38561 554643 38627 554646
rect 39990 554300 40050 554404
rect 39982 554236 39988 554300
rect 40052 554236 40058 554300
rect 42558 554026 42564 554028
rect 41492 553966 42564 554026
rect 42558 553964 42564 553966
rect 42628 553964 42634 554028
rect 41462 553485 41522 553588
rect 41462 553480 41571 553485
rect 41462 553424 41510 553480
rect 41566 553424 41571 553480
rect 41462 553422 41571 553424
rect 41505 553419 41571 553422
rect 649950 553346 650010 553914
rect 674281 553890 674347 553893
rect 675518 553890 675524 553892
rect 674281 553888 675524 553890
rect 674281 553832 674286 553888
rect 674342 553832 675524 553888
rect 674281 553830 675524 553832
rect 674281 553827 674347 553830
rect 675518 553828 675524 553830
rect 675588 553828 675594 553892
rect 655421 553346 655487 553349
rect 649950 553344 655487 553346
rect 649950 553288 655426 553344
rect 655482 553288 655487 553344
rect 649950 553286 655487 553288
rect 655421 553283 655487 553286
rect 42742 553210 42748 553212
rect 41492 553150 42748 553210
rect 42742 553148 42748 553150
rect 42812 553148 42818 553212
rect 42190 552802 42196 552804
rect 41492 552742 42196 552802
rect 42190 552740 42196 552742
rect 42260 552740 42266 552804
rect 42926 552394 42932 552396
rect 41492 552334 42932 552394
rect 42926 552332 42932 552334
rect 42996 552332 43002 552396
rect 649950 552122 650010 552732
rect 655605 552122 655671 552125
rect 649950 552120 655671 552122
rect 649950 552064 655610 552120
rect 655666 552064 655671 552120
rect 649950 552062 655671 552064
rect 655605 552059 655671 552062
rect 41781 551986 41847 551989
rect 41492 551984 41847 551986
rect 41492 551928 41786 551984
rect 41842 551928 41847 551984
rect 41492 551926 41847 551928
rect 41781 551923 41847 551926
rect 41822 551578 41828 551580
rect 41492 551518 41828 551578
rect 41822 551516 41828 551518
rect 41892 551516 41898 551580
rect 41462 551036 41522 551140
rect 41454 550972 41460 551036
rect 41524 550972 41530 551036
rect 649950 551034 650010 551550
rect 655513 551034 655579 551037
rect 649950 551032 655579 551034
rect 649950 550976 655518 551032
rect 655574 550976 655579 551032
rect 649950 550974 655579 550976
rect 655513 550971 655579 550974
rect 655881 550898 655947 550901
rect 649950 550896 655947 550898
rect 649950 550840 655886 550896
rect 655942 550840 655947 550896
rect 649950 550838 655947 550840
rect 42006 550762 42012 550764
rect 41492 550702 42012 550762
rect 42006 550700 42012 550702
rect 42076 550700 42082 550764
rect 649950 550368 650010 550838
rect 655881 550835 655947 550838
rect 41462 550221 41522 550324
rect 41462 550216 41571 550221
rect 41462 550160 41510 550216
rect 41566 550160 41571 550216
rect 41462 550158 41571 550160
rect 41505 550155 41571 550158
rect 41462 549813 41522 549916
rect 41413 549808 41522 549813
rect 41413 549752 41418 549808
rect 41474 549752 41522 549808
rect 41413 549750 41522 549752
rect 41413 549747 41479 549750
rect 41462 549405 41522 549508
rect 41462 549400 41571 549405
rect 41462 549344 41510 549400
rect 41566 549344 41571 549400
rect 41462 549342 41571 549344
rect 41505 549339 41571 549342
rect 654225 549266 654291 549269
rect 649950 549264 654291 549266
rect 649950 549208 654230 549264
rect 654286 549208 654291 549264
rect 649950 549206 654291 549208
rect 649950 549186 650010 549206
rect 654225 549203 654291 549206
rect 41462 548997 41522 549100
rect 41462 548992 41571 548997
rect 41462 548936 41510 548992
rect 41566 548936 41571 548992
rect 41462 548934 41571 548936
rect 41505 548931 41571 548934
rect 41462 548589 41522 548692
rect 41462 548584 41571 548589
rect 654133 548586 654199 548589
rect 41462 548528 41510 548584
rect 41566 548528 41571 548584
rect 41462 548526 41571 548528
rect 41505 548523 41571 548526
rect 649950 548584 654199 548586
rect 649950 548528 654138 548584
rect 654194 548528 654199 548584
rect 649950 548526 654199 548528
rect 41462 548181 41522 548284
rect 41413 548176 41522 548181
rect 41413 548120 41418 548176
rect 41474 548120 41522 548176
rect 41413 548118 41522 548120
rect 41413 548115 41479 548118
rect 649950 548004 650010 548526
rect 654133 548523 654199 548526
rect 675477 548044 675543 548045
rect 675477 548040 675524 548044
rect 675588 548042 675594 548044
rect 675477 547984 675482 548040
rect 675477 547980 675524 547984
rect 675588 547982 675634 548042
rect 675588 547980 675594 547982
rect 675477 547979 675543 547980
rect 30422 547468 30482 547876
rect 41462 546957 41522 547060
rect 41462 546952 41571 546957
rect 41462 546896 41510 546952
rect 41566 546896 41571 546952
rect 41462 546894 41571 546896
rect 41505 546891 41571 546894
rect 677174 544036 677180 544100
rect 677244 544098 677250 544100
rect 679249 544098 679315 544101
rect 677244 544096 679315 544098
rect 677244 544040 679254 544096
rect 679310 544040 679315 544096
rect 677244 544038 679315 544040
rect 677244 544036 677250 544038
rect 679249 544035 679315 544038
rect 676806 543900 676812 543964
rect 676876 543962 676882 543964
rect 679065 543962 679131 543965
rect 676876 543960 679131 543962
rect 676876 543904 679070 543960
rect 679126 543904 679131 543960
rect 676876 543902 679131 543904
rect 676876 543900 676882 543902
rect 679065 543899 679131 543902
rect 676990 543764 676996 543828
rect 677060 543826 677066 543828
rect 678973 543826 679039 543829
rect 677060 543824 679039 543826
rect 677060 543768 678978 543824
rect 679034 543768 679039 543824
rect 677060 543766 679039 543768
rect 677060 543764 677066 543766
rect 678973 543763 679039 543766
rect 673678 543084 673684 543148
rect 673748 543146 673754 543148
rect 674414 543146 674420 543148
rect 673748 543086 674420 543146
rect 673748 543084 673754 543086
rect 674414 543084 674420 543086
rect 674484 543084 674490 543148
rect 676121 542740 676187 542741
rect 674598 542676 674604 542740
rect 674668 542738 674674 542740
rect 675334 542738 675340 542740
rect 674668 542678 675340 542738
rect 674668 542676 674674 542678
rect 675334 542676 675340 542678
rect 675404 542676 675410 542740
rect 676070 542738 676076 542740
rect 676030 542678 676076 542738
rect 676140 542736 676187 542740
rect 676182 542680 676187 542736
rect 676070 542676 676076 542678
rect 676140 542676 676187 542680
rect 676121 542675 676187 542676
rect 676121 541244 676187 541245
rect 676070 541180 676076 541244
rect 676140 541242 676187 541244
rect 676140 541240 676232 541242
rect 676182 541184 676232 541240
rect 676140 541182 676232 541184
rect 676140 541180 676187 541182
rect 676121 541179 676187 541180
rect 41638 538460 41644 538524
rect 41708 538522 41714 538524
rect 43621 538522 43687 538525
rect 41708 538520 43687 538522
rect 41708 538464 43626 538520
rect 43682 538464 43687 538520
rect 41708 538462 43687 538464
rect 41708 538460 41714 538462
rect 43621 538459 43687 538462
rect 42926 538324 42932 538388
rect 42996 538386 43002 538388
rect 43069 538386 43135 538389
rect 42996 538384 43135 538386
rect 42996 538328 43074 538384
rect 43130 538328 43135 538384
rect 42996 538326 43135 538328
rect 42996 538324 43002 538326
rect 43069 538323 43135 538326
rect 42374 538188 42380 538252
rect 42444 538250 42450 538252
rect 43713 538250 43779 538253
rect 42444 538248 43779 538250
rect 42444 538192 43718 538248
rect 43774 538192 43779 538248
rect 42444 538190 43779 538192
rect 42444 538188 42450 538190
rect 43713 538187 43779 538190
rect 42006 538052 42012 538116
rect 42076 538114 42082 538116
rect 42701 538114 42767 538117
rect 42076 538112 42767 538114
rect 42076 538056 42706 538112
rect 42762 538056 42767 538112
rect 42076 538054 42767 538056
rect 42076 538052 42082 538054
rect 42701 538051 42767 538054
rect 676262 535941 676322 536112
rect 676213 535936 676322 535941
rect 676213 535880 676218 535936
rect 676274 535880 676322 535936
rect 676213 535878 676322 535880
rect 676213 535875 676279 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 41454 535332 41460 535396
rect 41524 535394 41530 535396
rect 42241 535394 42307 535397
rect 41524 535392 42307 535394
rect 41524 535336 42246 535392
rect 42302 535336 42307 535392
rect 41524 535334 42307 535336
rect 41524 535332 41530 535334
rect 42241 535331 42307 535334
rect 42558 535332 42564 535396
rect 42628 535394 42634 535396
rect 43161 535394 43227 535397
rect 42628 535392 43227 535394
rect 42628 535336 43166 535392
rect 43222 535336 43227 535392
rect 42628 535334 43227 535336
rect 42628 535332 42634 535334
rect 43161 535331 43227 535334
rect 679206 535125 679266 535296
rect 678973 535122 679039 535125
rect 678973 535120 679082 535122
rect 678973 535064 678978 535120
rect 679034 535064 679082 535120
rect 678973 535059 679082 535064
rect 679157 535120 679266 535125
rect 679157 535064 679162 535120
rect 679218 535064 679266 535120
rect 679157 535062 679266 535064
rect 679157 535059 679223 535062
rect 679022 534888 679082 535059
rect 679574 534309 679634 534480
rect 679341 534306 679407 534309
rect 679341 534304 679450 534306
rect 679341 534248 679346 534304
rect 679402 534248 679450 534304
rect 679341 534243 679450 534248
rect 679525 534304 679634 534309
rect 679525 534248 679530 534304
rect 679586 534248 679634 534304
rect 679525 534246 679634 534248
rect 679525 534243 679591 534246
rect 679390 534072 679450 534243
rect 679390 533493 679450 533664
rect 679249 533490 679315 533493
rect 679206 533488 679315 533490
rect 679206 533432 679254 533488
rect 679310 533432 679315 533488
rect 679206 533427 679315 533432
rect 679390 533488 679499 533493
rect 679390 533432 679438 533488
rect 679494 533432 679499 533488
rect 679390 533430 679499 533432
rect 679433 533427 679499 533430
rect 679206 533256 679266 533427
rect 42190 532748 42196 532812
rect 42260 532810 42266 532812
rect 42425 532810 42491 532813
rect 42260 532808 42491 532810
rect 42260 532752 42430 532808
rect 42486 532752 42491 532808
rect 42260 532750 42491 532752
rect 42260 532748 42266 532750
rect 42425 532747 42491 532750
rect 679206 532677 679266 532848
rect 41822 532612 41828 532676
rect 41892 532674 41898 532676
rect 42333 532674 42399 532677
rect 41892 532672 42399 532674
rect 41892 532616 42338 532672
rect 42394 532616 42399 532672
rect 41892 532614 42399 532616
rect 41892 532612 41898 532614
rect 42333 532611 42399 532614
rect 42742 532612 42748 532676
rect 42812 532674 42818 532676
rect 43069 532674 43135 532677
rect 679065 532674 679131 532677
rect 42812 532672 43135 532674
rect 42812 532616 43074 532672
rect 43130 532616 43135 532672
rect 42812 532614 43135 532616
rect 42812 532612 42818 532614
rect 43069 532611 43135 532614
rect 679022 532672 679131 532674
rect 679022 532616 679070 532672
rect 679126 532616 679131 532672
rect 679022 532611 679131 532616
rect 679206 532672 679315 532677
rect 679206 532616 679254 532672
rect 679310 532616 679315 532672
rect 679206 532614 679315 532616
rect 679249 532611 679315 532614
rect 679022 532440 679082 532611
rect 679022 531861 679082 532032
rect 674414 531796 674420 531860
rect 674484 531858 674490 531860
rect 674484 531798 676322 531858
rect 674484 531796 674490 531798
rect 59445 531722 59511 531725
rect 59445 531720 64706 531722
rect 59445 531664 59450 531720
rect 59506 531664 64706 531720
rect 59445 531662 64706 531664
rect 59445 531659 59511 531662
rect 64646 531172 64706 531662
rect 676262 531624 676322 531798
rect 678973 531856 679082 531861
rect 678973 531800 678978 531856
rect 679034 531800 679082 531856
rect 678973 531798 679082 531800
rect 678973 531795 679039 531798
rect 675477 531314 675543 531317
rect 675477 531312 676322 531314
rect 675477 531256 675482 531312
rect 675538 531256 676322 531312
rect 675477 531254 676322 531256
rect 675477 531251 675543 531254
rect 676262 531216 676322 531254
rect 673494 530980 673500 531044
rect 673564 531042 673570 531044
rect 673564 530982 676322 531042
rect 673564 530980 673570 530982
rect 676262 530808 676322 530982
rect 59261 530634 59327 530637
rect 59261 530632 64706 530634
rect 59261 530576 59266 530632
rect 59322 530576 64706 530632
rect 59261 530574 64706 530576
rect 59261 530571 59327 530574
rect 64646 529990 64706 530574
rect 674230 530572 674236 530636
rect 674300 530634 674306 530636
rect 674300 530574 676322 530634
rect 674300 530572 674306 530574
rect 676262 530400 676322 530574
rect 676029 530022 676095 530025
rect 676029 530020 676292 530022
rect 676029 529964 676034 530020
rect 676090 529964 676292 530020
rect 676029 529962 676292 529964
rect 676029 529959 676095 529962
rect 676029 529614 676095 529617
rect 676029 529612 676292 529614
rect 676029 529556 676034 529612
rect 676090 529556 676292 529612
rect 676029 529554 676292 529556
rect 676029 529551 676095 529554
rect 58525 529410 58591 529413
rect 58525 529408 64706 529410
rect 58525 529352 58530 529408
rect 58586 529352 64706 529408
rect 58525 529350 64706 529352
rect 58525 529347 58591 529350
rect 64646 528808 64706 529350
rect 676070 529348 676076 529412
rect 676140 529410 676146 529412
rect 676140 529350 676322 529410
rect 676140 529348 676146 529350
rect 676262 529176 676322 529350
rect 674598 528940 674604 529004
rect 674668 529002 674674 529004
rect 674668 528942 676322 529002
rect 674668 528940 674674 528942
rect 676262 528768 676322 528942
rect 673678 528532 673684 528596
rect 673748 528594 673754 528596
rect 673748 528534 676322 528594
rect 673748 528532 673754 528534
rect 676262 528360 676322 528534
rect 58341 528186 58407 528189
rect 58341 528184 64706 528186
rect 58341 528128 58346 528184
rect 58402 528128 64706 528184
rect 58341 528126 64706 528128
rect 58341 528123 58407 528126
rect 64646 527626 64706 528126
rect 676029 527982 676095 527985
rect 676029 527980 676292 527982
rect 676029 527924 676034 527980
rect 676090 527924 676292 527980
rect 676029 527922 676292 527924
rect 676029 527919 676095 527922
rect 676029 527574 676095 527577
rect 676029 527572 676292 527574
rect 676029 527516 676034 527572
rect 676090 527516 676292 527572
rect 676029 527514 676292 527516
rect 676029 527511 676095 527514
rect 673862 527036 673868 527100
rect 673932 527098 673938 527100
rect 676262 527098 676322 527136
rect 673932 527038 676322 527098
rect 673932 527036 673938 527038
rect 57973 526962 58039 526965
rect 57973 526960 64706 526962
rect 57973 526904 57978 526960
rect 58034 526904 64706 526960
rect 57973 526902 64706 526904
rect 57973 526899 58039 526902
rect 64646 526444 64706 526902
rect 675937 526758 676003 526761
rect 675937 526756 676292 526758
rect 675937 526700 675942 526756
rect 675998 526700 676292 526756
rect 675937 526698 676292 526700
rect 675937 526695 676003 526698
rect 676029 526350 676095 526353
rect 676029 526348 676292 526350
rect 676029 526292 676034 526348
rect 676090 526292 676292 526348
rect 676029 526290 676292 526292
rect 676029 526287 676095 526290
rect 58065 525874 58131 525877
rect 58065 525872 64706 525874
rect 58065 525816 58070 525872
rect 58126 525816 64706 525872
rect 58065 525814 64706 525816
rect 58065 525811 58131 525814
rect 64646 525262 64706 525814
rect 679022 525741 679082 525912
rect 679022 525736 679131 525741
rect 679022 525680 679070 525736
rect 679126 525680 679131 525736
rect 679022 525678 679131 525680
rect 679065 525675 679131 525678
rect 684542 525096 684602 525504
rect 679065 524922 679131 524925
rect 679022 524920 679131 524922
rect 679022 524864 679070 524920
rect 679126 524864 679131 524920
rect 679022 524859 679131 524864
rect 679022 524688 679082 524859
rect 676029 492146 676095 492149
rect 676029 492144 676292 492146
rect 676029 492088 676034 492144
rect 676090 492088 676292 492144
rect 676029 492086 676292 492088
rect 676029 492083 676095 492086
rect 675937 491738 676003 491741
rect 675937 491736 676292 491738
rect 675937 491680 675942 491736
rect 675998 491680 676292 491736
rect 675937 491678 676292 491680
rect 675937 491675 676003 491678
rect 676029 491330 676095 491333
rect 676029 491328 676292 491330
rect 676029 491272 676034 491328
rect 676090 491272 676292 491328
rect 676029 491270 676292 491272
rect 676029 491267 676095 491270
rect 676029 490922 676095 490925
rect 676029 490920 676292 490922
rect 676029 490864 676034 490920
rect 676090 490864 676292 490920
rect 676029 490862 676292 490864
rect 676029 490859 676095 490862
rect 675753 490514 675819 490517
rect 675753 490512 676292 490514
rect 675753 490456 675758 490512
rect 675814 490456 676292 490512
rect 675753 490454 676292 490456
rect 675753 490451 675819 490454
rect 676029 490106 676095 490109
rect 676029 490104 676292 490106
rect 676029 490048 676034 490104
rect 676090 490048 676292 490104
rect 676029 490046 676292 490048
rect 676029 490043 676095 490046
rect 676029 489698 676095 489701
rect 676029 489696 676292 489698
rect 676029 489640 676034 489696
rect 676090 489640 676292 489696
rect 676029 489638 676292 489640
rect 676029 489635 676095 489638
rect 676029 489290 676095 489293
rect 676029 489288 676292 489290
rect 676029 489232 676034 489288
rect 676090 489232 676292 489288
rect 676029 489230 676292 489232
rect 676029 489227 676095 489230
rect 675385 488882 675451 488885
rect 675385 488880 676292 488882
rect 675385 488824 675390 488880
rect 675446 488824 676292 488880
rect 675385 488822 676292 488824
rect 675385 488819 675451 488822
rect 675937 488474 676003 488477
rect 675937 488472 676292 488474
rect 675937 488416 675942 488472
rect 675998 488416 676292 488472
rect 675937 488414 676292 488416
rect 675937 488411 676003 488414
rect 675937 488066 676003 488069
rect 675937 488064 676292 488066
rect 675937 488008 675942 488064
rect 675998 488008 676292 488064
rect 675937 488006 676292 488008
rect 675937 488003 676003 488006
rect 674966 487596 674972 487660
rect 675036 487658 675042 487660
rect 675036 487598 676292 487658
rect 675036 487596 675042 487598
rect 675477 487250 675543 487253
rect 675477 487248 676292 487250
rect 675477 487192 675482 487248
rect 675538 487192 676292 487248
rect 675477 487190 676292 487192
rect 675477 487187 675543 487190
rect 675150 486780 675156 486844
rect 675220 486842 675226 486844
rect 675220 486782 676292 486842
rect 675220 486780 675226 486782
rect 675845 486434 675911 486437
rect 675845 486432 676292 486434
rect 675845 486376 675850 486432
rect 675906 486376 676292 486432
rect 675845 486374 676292 486376
rect 675845 486371 675911 486374
rect 676029 486026 676095 486029
rect 676029 486024 676292 486026
rect 676029 485968 676034 486024
rect 676090 485968 676292 486024
rect 676029 485966 676292 485968
rect 676029 485963 676095 485966
rect 676029 485618 676095 485621
rect 676029 485616 676292 485618
rect 676029 485560 676034 485616
rect 676090 485560 676292 485616
rect 676029 485558 676292 485560
rect 676029 485555 676095 485558
rect 674046 485148 674052 485212
rect 674116 485210 674122 485212
rect 674116 485150 676292 485210
rect 674116 485148 674122 485150
rect 674782 484740 674788 484804
rect 674852 484802 674858 484804
rect 674852 484742 676292 484802
rect 674852 484740 674858 484742
rect 675845 484394 675911 484397
rect 675845 484392 676292 484394
rect 675845 484336 675850 484392
rect 675906 484336 676292 484392
rect 675845 484334 676292 484336
rect 675845 484331 675911 484334
rect 676029 483986 676095 483989
rect 676029 483984 676292 483986
rect 676029 483928 676034 483984
rect 676090 483928 676292 483984
rect 676029 483926 676292 483928
rect 676029 483923 676095 483926
rect 676029 483578 676095 483581
rect 676029 483576 676292 483578
rect 676029 483520 676034 483576
rect 676090 483520 676292 483576
rect 676029 483518 676292 483520
rect 676029 483515 676095 483518
rect 676029 483170 676095 483173
rect 676029 483168 676292 483170
rect 676029 483112 676034 483168
rect 676090 483112 676292 483168
rect 676029 483110 676292 483112
rect 676029 483107 676095 483110
rect 675569 482762 675635 482765
rect 675569 482760 676292 482762
rect 675569 482704 675574 482760
rect 675630 482704 676292 482760
rect 675569 482702 676292 482704
rect 675569 482699 675635 482702
rect 676029 482354 676095 482357
rect 676029 482352 676292 482354
rect 676029 482296 676034 482352
rect 676090 482296 676292 482352
rect 676029 482294 676292 482296
rect 676029 482291 676095 482294
rect 676029 481946 676095 481949
rect 676029 481944 676292 481946
rect 676029 481888 676034 481944
rect 676090 481888 676292 481944
rect 676029 481886 676292 481888
rect 676029 481883 676095 481886
rect 684542 481100 684602 481508
rect 676029 480722 676095 480725
rect 676029 480720 676292 480722
rect 676029 480664 676034 480720
rect 676090 480664 676292 480720
rect 676029 480662 676292 480664
rect 676029 480659 676095 480662
rect 39982 435916 39988 435980
rect 40052 435978 40058 435980
rect 41873 435978 41939 435981
rect 40052 435976 41939 435978
rect 40052 435920 41878 435976
rect 41934 435920 41939 435976
rect 40052 435918 41939 435920
rect 40052 435916 40058 435918
rect 41873 435915 41939 435918
rect 41781 430946 41847 430949
rect 41492 430944 41847 430946
rect 41492 430888 41786 430944
rect 41842 430888 41847 430944
rect 41492 430886 41847 430888
rect 41781 430883 41847 430886
rect 41781 430538 41847 430541
rect 41492 430536 41847 430538
rect 41492 430480 41786 430536
rect 41842 430480 41847 430536
rect 41492 430478 41847 430480
rect 41781 430475 41847 430478
rect 41781 430130 41847 430133
rect 41492 430128 41847 430130
rect 41492 430072 41786 430128
rect 41842 430072 41847 430128
rect 41492 430070 41847 430072
rect 41781 430067 41847 430070
rect 41781 429722 41847 429725
rect 41492 429720 41847 429722
rect 41492 429664 41786 429720
rect 41842 429664 41847 429720
rect 41492 429662 41847 429664
rect 41781 429659 41847 429662
rect 41781 429314 41847 429317
rect 41492 429312 41847 429314
rect 41492 429256 41786 429312
rect 41842 429256 41847 429312
rect 41492 429254 41847 429256
rect 41781 429251 41847 429254
rect 41781 428906 41847 428909
rect 41492 428904 41847 428906
rect 41492 428848 41786 428904
rect 41842 428848 41847 428904
rect 41492 428846 41847 428848
rect 41781 428843 41847 428846
rect 42425 428498 42491 428501
rect 41492 428496 42491 428498
rect 41492 428440 42430 428496
rect 42486 428440 42491 428496
rect 41492 428438 42491 428440
rect 42425 428435 42491 428438
rect 44030 428090 44036 428092
rect 41492 428030 44036 428090
rect 44030 428028 44036 428030
rect 44100 428028 44106 428092
rect 42057 427682 42123 427685
rect 41492 427680 42123 427682
rect 41492 427624 42062 427680
rect 42118 427624 42123 427680
rect 41492 427622 42123 427624
rect 42057 427619 42123 427622
rect 41873 427274 41939 427277
rect 41492 427272 41939 427274
rect 41492 427216 41878 427272
rect 41934 427216 41939 427272
rect 41492 427214 41939 427216
rect 41873 427211 41939 427214
rect 41781 426866 41847 426869
rect 41492 426864 41847 426866
rect 41492 426808 41786 426864
rect 41842 426808 41847 426864
rect 41492 426806 41847 426808
rect 41781 426803 41847 426806
rect 41781 426458 41847 426461
rect 41492 426456 41847 426458
rect 41492 426400 41786 426456
rect 41842 426400 41847 426456
rect 41492 426398 41847 426400
rect 41781 426395 41847 426398
rect 41965 426050 42031 426053
rect 41492 426048 42031 426050
rect 41492 425992 41970 426048
rect 42026 425992 42031 426048
rect 41492 425990 42031 425992
rect 41965 425987 42031 425990
rect 41781 425642 41847 425645
rect 41492 425640 41847 425642
rect 41492 425584 41786 425640
rect 41842 425584 41847 425640
rect 41492 425582 41847 425584
rect 41781 425579 41847 425582
rect 41781 425234 41847 425237
rect 41492 425232 41847 425234
rect 41492 425176 41786 425232
rect 41842 425176 41847 425232
rect 41492 425174 41847 425176
rect 41781 425171 41847 425174
rect 41781 424826 41847 424829
rect 41492 424824 41847 424826
rect 41492 424768 41786 424824
rect 41842 424768 41847 424824
rect 41492 424766 41847 424768
rect 41781 424763 41847 424766
rect 42241 424418 42307 424421
rect 41492 424416 42307 424418
rect 41492 424360 42246 424416
rect 42302 424360 42307 424416
rect 41492 424358 42307 424360
rect 42241 424355 42307 424358
rect 41873 424010 41939 424013
rect 41492 424008 41939 424010
rect 41492 423952 41878 424008
rect 41934 423952 41939 424008
rect 41492 423950 41939 423952
rect 41873 423947 41939 423950
rect 41873 423602 41939 423605
rect 41492 423600 41939 423602
rect 41492 423544 41878 423600
rect 41934 423544 41939 423600
rect 41492 423542 41939 423544
rect 41873 423539 41939 423542
rect 41873 423194 41939 423197
rect 41492 423192 41939 423194
rect 41492 423136 41878 423192
rect 41934 423136 41939 423192
rect 41492 423134 41939 423136
rect 41873 423131 41939 423134
rect 41873 422786 41939 422789
rect 41492 422784 41939 422786
rect 41492 422728 41878 422784
rect 41934 422728 41939 422784
rect 41492 422726 41939 422728
rect 41873 422723 41939 422726
rect 41781 422378 41847 422381
rect 41492 422376 41847 422378
rect 41492 422320 41786 422376
rect 41842 422320 41847 422376
rect 41492 422318 41847 422320
rect 41781 422315 41847 422318
rect 41781 421970 41847 421973
rect 41492 421968 41847 421970
rect 41492 421912 41786 421968
rect 41842 421912 41847 421968
rect 41492 421910 41847 421912
rect 41781 421907 41847 421910
rect 41873 421562 41939 421565
rect 41492 421560 41939 421562
rect 41492 421504 41878 421560
rect 41934 421504 41939 421560
rect 41492 421502 41939 421504
rect 41873 421499 41939 421502
rect 42333 421154 42399 421157
rect 41492 421152 42399 421154
rect 41492 421096 42338 421152
rect 42394 421096 42399 421152
rect 41492 421094 42399 421096
rect 42333 421091 42399 421094
rect 41781 420746 41847 420749
rect 41492 420744 41847 420746
rect 41492 420688 41786 420744
rect 41842 420688 41847 420744
rect 41492 420686 41847 420688
rect 41781 420683 41847 420686
rect 30422 419900 30482 420308
rect 41781 419522 41847 419525
rect 41492 419520 41847 419522
rect 41492 419464 41786 419520
rect 41842 419464 41847 419520
rect 41492 419462 41847 419464
rect 41781 419459 41847 419462
rect 43110 411436 43116 411500
rect 43180 411498 43186 411500
rect 43253 411498 43319 411501
rect 43180 411496 43319 411498
rect 43180 411440 43258 411496
rect 43314 411440 43319 411496
rect 43180 411438 43319 411440
rect 43180 411436 43186 411438
rect 43253 411435 43319 411438
rect 43161 406876 43227 406877
rect 43110 406812 43116 406876
rect 43180 406874 43227 406876
rect 43180 406872 43272 406874
rect 43222 406816 43272 406872
rect 43180 406814 43272 406816
rect 43180 406812 43227 406814
rect 43161 406811 43227 406812
rect 58433 404154 58499 404157
rect 58433 404152 64706 404154
rect 58433 404096 58438 404152
rect 58494 404096 64706 404152
rect 58433 404094 64706 404096
rect 58433 404091 58499 404094
rect 64646 403550 64706 404094
rect 676121 403746 676187 403749
rect 676262 403746 676322 403852
rect 676121 403744 676322 403746
rect 676121 403688 676126 403744
rect 676182 403688 676322 403744
rect 676121 403686 676322 403688
rect 676121 403683 676187 403686
rect 676262 403341 676322 403444
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 676213 403275 676279 403278
rect 58525 402930 58591 402933
rect 676121 402930 676187 402933
rect 676262 402930 676322 403036
rect 58525 402928 64706 402930
rect 58525 402872 58530 402928
rect 58586 402872 64706 402928
rect 58525 402870 64706 402872
rect 58525 402867 58591 402870
rect 64646 402368 64706 402870
rect 676121 402928 676322 402930
rect 676121 402872 676126 402928
rect 676182 402872 676322 402928
rect 676121 402870 676322 402872
rect 676121 402867 676187 402870
rect 675845 402658 675911 402661
rect 675845 402656 676292 402658
rect 675845 402600 675850 402656
rect 675906 402600 676292 402656
rect 675845 402598 676292 402600
rect 675845 402595 675911 402598
rect 675293 402250 675359 402253
rect 675293 402248 676292 402250
rect 675293 402192 675298 402248
rect 675354 402192 676292 402248
rect 675293 402190 676292 402192
rect 675293 402187 675359 402190
rect 676029 401842 676095 401845
rect 676029 401840 676292 401842
rect 676029 401784 676034 401840
rect 676090 401784 676292 401840
rect 676029 401782 676292 401784
rect 676029 401779 676095 401782
rect 675753 401434 675819 401437
rect 675753 401432 676292 401434
rect 675753 401376 675758 401432
rect 675814 401376 676292 401432
rect 675753 401374 676292 401376
rect 675753 401371 675819 401374
rect 60365 400754 60431 400757
rect 64646 400754 64706 401186
rect 675845 401026 675911 401029
rect 675845 401024 676292 401026
rect 675845 400968 675850 401024
rect 675906 400968 676292 401024
rect 675845 400966 676292 400968
rect 675845 400963 675911 400966
rect 60365 400752 64706 400754
rect 60365 400696 60370 400752
rect 60426 400696 64706 400752
rect 60365 400694 64706 400696
rect 60365 400691 60431 400694
rect 675150 400556 675156 400620
rect 675220 400618 675226 400620
rect 675220 400558 676292 400618
rect 675220 400556 675226 400558
rect 675937 400210 676003 400213
rect 675937 400208 676292 400210
rect 675937 400152 675942 400208
rect 675998 400152 676292 400208
rect 675937 400150 676292 400152
rect 675937 400147 676003 400150
rect 58433 400074 58499 400077
rect 58433 400072 64706 400074
rect 58433 400016 58438 400072
rect 58494 400016 64706 400072
rect 58433 400014 64706 400016
rect 58433 400011 58499 400014
rect 64646 400004 64706 400014
rect 676029 399802 676095 399805
rect 676029 399800 676292 399802
rect 676029 399744 676034 399800
rect 676090 399744 676292 399800
rect 676029 399742 676292 399744
rect 676029 399739 676095 399742
rect 58525 399394 58591 399397
rect 676029 399394 676095 399397
rect 58525 399392 64706 399394
rect 58525 399336 58530 399392
rect 58586 399336 64706 399392
rect 58525 399334 64706 399336
rect 58525 399331 58591 399334
rect 64646 398822 64706 399334
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 676121 398850 676187 398853
rect 676262 398850 676322 398956
rect 676121 398848 676322 398850
rect 676121 398792 676126 398848
rect 676182 398792 676322 398848
rect 676121 398790 676322 398792
rect 676121 398787 676187 398790
rect 675845 398578 675911 398581
rect 675845 398576 676292 398578
rect 675845 398520 675850 398576
rect 675906 398520 676292 398576
rect 675845 398518 676292 398520
rect 675845 398515 675911 398518
rect 58341 398306 58407 398309
rect 58341 398304 64706 398306
rect 58341 398248 58346 398304
rect 58402 398248 64706 398304
rect 58341 398246 64706 398248
rect 58341 398243 58407 398246
rect 64646 397640 64706 398246
rect 676029 398170 676095 398173
rect 676029 398168 676292 398170
rect 676029 398112 676034 398168
rect 676090 398112 676292 398168
rect 676029 398110 676292 398112
rect 676029 398107 676095 398110
rect 675937 397762 676003 397765
rect 675937 397760 676292 397762
rect 675937 397704 675942 397760
rect 675998 397704 676292 397760
rect 675937 397702 676292 397704
rect 675937 397699 676003 397702
rect 676029 397354 676095 397357
rect 676029 397352 676292 397354
rect 676029 397296 676034 397352
rect 676090 397296 676292 397352
rect 676029 397294 676292 397296
rect 676029 397291 676095 397294
rect 676029 396946 676095 396949
rect 676029 396944 676292 396946
rect 676029 396888 676034 396944
rect 676090 396888 676292 396944
rect 676029 396886 676292 396888
rect 676029 396883 676095 396886
rect 676121 396402 676187 396405
rect 676262 396402 676322 396508
rect 676121 396400 676322 396402
rect 676121 396344 676126 396400
rect 676182 396344 676322 396400
rect 676121 396342 676322 396344
rect 676121 396339 676187 396342
rect 675937 396130 676003 396133
rect 675937 396128 676292 396130
rect 675937 396072 675942 396128
rect 675998 396072 676292 396128
rect 675937 396070 676292 396072
rect 675937 396067 676003 396070
rect 675661 395722 675727 395725
rect 675661 395720 676292 395722
rect 675661 395664 675666 395720
rect 675722 395664 676292 395720
rect 675661 395662 676292 395664
rect 675661 395659 675727 395662
rect 675661 395314 675727 395317
rect 675661 395312 676292 395314
rect 675661 395256 675666 395312
rect 675722 395256 676292 395312
rect 675661 395254 676292 395256
rect 675661 395251 675727 395254
rect 675937 394906 676003 394909
rect 675937 394904 676292 394906
rect 675937 394848 675942 394904
rect 675998 394848 676292 394904
rect 675937 394846 676292 394848
rect 675937 394843 676003 394846
rect 676029 394498 676095 394501
rect 676029 394496 676292 394498
rect 676029 394440 676034 394496
rect 676090 394440 676292 394496
rect 676029 394438 676292 394440
rect 676029 394435 676095 394438
rect 676029 394090 676095 394093
rect 676029 394088 676292 394090
rect 676029 394032 676034 394088
rect 676090 394032 676292 394088
rect 676029 394030 676292 394032
rect 676029 394027 676095 394030
rect 679022 393549 679082 393652
rect 678973 393544 679082 393549
rect 678973 393488 678978 393544
rect 679034 393488 679082 393544
rect 678973 393486 679082 393488
rect 678973 393483 679039 393486
rect 684542 392836 684602 393244
rect 678973 392730 679039 392733
rect 678973 392728 679082 392730
rect 678973 392672 678978 392728
rect 679034 392672 679082 392728
rect 678973 392667 679082 392672
rect 679022 392428 679082 392667
rect 41462 387565 41522 387668
rect 41413 387560 41522 387565
rect 41413 387504 41418 387560
rect 41474 387504 41522 387560
rect 41413 387502 41522 387504
rect 41413 387499 41479 387502
rect 41462 387157 41522 387260
rect 41413 387152 41522 387157
rect 41413 387096 41418 387152
rect 41474 387096 41522 387152
rect 41413 387094 41522 387096
rect 41413 387091 41479 387094
rect 41781 386882 41847 386885
rect 41492 386880 41847 386882
rect 41492 386824 41786 386880
rect 41842 386824 41847 386880
rect 41492 386822 41847 386824
rect 41781 386819 41847 386822
rect 41505 386746 41571 386749
rect 41462 386744 41571 386746
rect 41462 386688 41510 386744
rect 41566 386688 41571 386744
rect 41462 386683 41571 386688
rect 41462 386444 41522 386683
rect 42425 386066 42491 386069
rect 41492 386064 42491 386066
rect 41492 386008 42430 386064
rect 42486 386008 42491 386064
rect 41492 386006 42491 386008
rect 42425 386003 42491 386006
rect 41505 385930 41571 385933
rect 41462 385928 41571 385930
rect 41462 385872 41510 385928
rect 41566 385872 41571 385928
rect 41462 385867 41571 385872
rect 41462 385628 41522 385867
rect 41873 385250 41939 385253
rect 41492 385248 41939 385250
rect 41492 385192 41878 385248
rect 41934 385192 41939 385248
rect 41492 385190 41939 385192
rect 41873 385187 41939 385190
rect 41505 385114 41571 385117
rect 41462 385112 41571 385114
rect 41462 385056 41510 385112
rect 41566 385056 41571 385112
rect 41462 385051 41571 385056
rect 41462 384812 41522 385051
rect 41462 384301 41522 384404
rect 41462 384296 41571 384301
rect 41462 384240 41510 384296
rect 41566 384240 41571 384296
rect 41462 384238 41571 384240
rect 41505 384235 41571 384238
rect 41781 384026 41847 384029
rect 41492 384024 41847 384026
rect 41492 383968 41786 384024
rect 41842 383968 41847 384024
rect 41492 383966 41847 383968
rect 41781 383963 41847 383966
rect 41462 383485 41522 383588
rect 41462 383480 41571 383485
rect 41462 383424 41510 383480
rect 41566 383424 41571 383480
rect 41462 383422 41571 383424
rect 41505 383419 41571 383422
rect 41462 383074 41522 383180
rect 41638 383074 41644 383076
rect 41462 383014 41644 383074
rect 41638 383012 41644 383014
rect 41708 383012 41714 383076
rect 41462 382669 41522 382772
rect 41462 382664 41571 382669
rect 41462 382608 41510 382664
rect 41566 382608 41571 382664
rect 41462 382606 41571 382608
rect 41505 382603 41571 382606
rect 41462 382260 41522 382364
rect 41454 382196 41460 382260
rect 41524 382196 41530 382260
rect 41462 381853 41522 381956
rect 41462 381848 41571 381853
rect 41462 381792 41510 381848
rect 41566 381792 41571 381848
rect 41462 381790 41571 381792
rect 41505 381787 41571 381790
rect 41462 381445 41522 381548
rect 41462 381440 41571 381445
rect 41462 381384 41510 381440
rect 41566 381384 41571 381440
rect 41462 381382 41571 381384
rect 41505 381379 41571 381382
rect 42333 381170 42399 381173
rect 41492 381168 42399 381170
rect 41492 381112 42338 381168
rect 42394 381112 42399 381168
rect 41492 381110 42399 381112
rect 42333 381107 42399 381110
rect 41965 380762 42031 380765
rect 41492 380760 42031 380762
rect 41492 380704 41970 380760
rect 42026 380704 42031 380760
rect 41492 380702 42031 380704
rect 41965 380699 42031 380702
rect 41462 380221 41522 380324
rect 41462 380216 41571 380221
rect 41462 380160 41510 380216
rect 41566 380160 41571 380216
rect 41462 380158 41571 380160
rect 41505 380155 41571 380158
rect 41462 379813 41522 379916
rect 41462 379808 41571 379813
rect 41462 379752 41510 379808
rect 41566 379752 41571 379808
rect 41462 379750 41571 379752
rect 41505 379747 41571 379750
rect 41462 379405 41522 379508
rect 41462 379400 41571 379405
rect 41462 379344 41510 379400
rect 41566 379344 41571 379400
rect 41462 379342 41571 379344
rect 41505 379339 41571 379342
rect 41462 378997 41522 379100
rect 41413 378992 41522 378997
rect 41413 378936 41418 378992
rect 41474 378936 41522 378992
rect 41413 378934 41522 378936
rect 41413 378931 41479 378934
rect 41462 378586 41522 378692
rect 41597 378586 41663 378589
rect 41462 378584 41663 378586
rect 41462 378528 41602 378584
rect 41658 378528 41663 378584
rect 41462 378526 41663 378528
rect 41597 378523 41663 378526
rect 41462 378181 41522 378284
rect 41462 378176 41571 378181
rect 41462 378120 41510 378176
rect 41566 378120 41571 378176
rect 41462 378118 41571 378120
rect 41505 378115 41571 378118
rect 41278 377773 41338 377876
rect 41278 377768 41387 377773
rect 41278 377712 41326 377768
rect 41382 377712 41387 377768
rect 41278 377710 41387 377712
rect 41321 377707 41387 377710
rect 41462 377365 41522 377468
rect 41413 377360 41522 377365
rect 41413 377304 41418 377360
rect 41474 377304 41522 377360
rect 41413 377302 41522 377304
rect 41413 377299 41479 377302
rect 30422 376652 30482 377060
rect 41462 376141 41522 376244
rect 41413 376136 41522 376141
rect 41413 376080 41418 376136
rect 41474 376080 41522 376136
rect 41413 376078 41522 376080
rect 41413 376075 41479 376078
rect 655513 374506 655579 374509
rect 649950 374504 655579 374506
rect 649950 374448 655518 374504
rect 655574 374448 655579 374504
rect 649950 374446 655579 374448
rect 649950 373892 650010 374446
rect 655513 374443 655579 374446
rect 655697 373282 655763 373285
rect 649950 373280 655763 373282
rect 649950 373224 655702 373280
rect 655758 373224 655763 373280
rect 649950 373222 655763 373224
rect 649950 372710 650010 373222
rect 655697 373219 655763 373222
rect 655421 372194 655487 372197
rect 649950 372192 655487 372194
rect 649950 372136 655426 372192
rect 655482 372136 655487 372192
rect 649950 372134 655487 372136
rect 649950 371528 650010 372134
rect 655421 372131 655487 372134
rect 654501 370970 654567 370973
rect 649950 370968 654567 370970
rect 649950 370912 654506 370968
rect 654562 370912 654567 370968
rect 649950 370910 654567 370912
rect 649950 370346 650010 370910
rect 654501 370907 654567 370910
rect 58157 360906 58223 360909
rect 58157 360904 64706 360906
rect 58157 360848 58162 360904
rect 58218 360848 64706 360904
rect 58157 360846 64706 360848
rect 58157 360843 58223 360846
rect 64646 360328 64706 360846
rect 58525 359818 58591 359821
rect 58525 359816 64706 359818
rect 58525 359760 58530 359816
rect 58586 359760 64706 359816
rect 58525 359758 64706 359760
rect 58525 359755 58591 359758
rect 64646 359146 64706 359758
rect 675845 358730 675911 358733
rect 675845 358728 676292 358730
rect 675845 358672 675850 358728
rect 675906 358672 676292 358728
rect 675845 358670 676292 358672
rect 675845 358667 675911 358670
rect 676029 358322 676095 358325
rect 676029 358320 676292 358322
rect 676029 358264 676034 358320
rect 676090 358264 676292 358320
rect 676029 358262 676292 358264
rect 676029 358259 676095 358262
rect 57973 357506 58039 357509
rect 64646 357506 64706 357964
rect 675937 357914 676003 357917
rect 675937 357912 676292 357914
rect 675937 357856 675942 357912
rect 675998 357856 676292 357912
rect 675937 357854 676292 357856
rect 675937 357851 676003 357854
rect 57973 357504 64706 357506
rect 57973 357448 57978 357504
rect 58034 357448 64706 357504
rect 57973 357446 64706 357448
rect 675293 357506 675359 357509
rect 675293 357504 676292 357506
rect 675293 357448 675298 357504
rect 675354 357448 676292 357504
rect 675293 357446 676292 357448
rect 57973 357443 58039 357446
rect 675293 357443 675359 357446
rect 58525 357370 58591 357373
rect 58525 357368 64706 357370
rect 58525 357312 58530 357368
rect 58586 357312 64706 357368
rect 58525 357310 64706 357312
rect 58525 357307 58591 357310
rect 41638 356900 41644 356964
rect 41708 356962 41714 356964
rect 41781 356962 41847 356965
rect 41708 356960 41847 356962
rect 41708 356904 41786 356960
rect 41842 356904 41847 356960
rect 41708 356902 41847 356904
rect 41708 356900 41714 356902
rect 41781 356899 41847 356902
rect 64646 356782 64706 357310
rect 675201 357098 675267 357101
rect 675201 357096 676292 357098
rect 675201 357040 675206 357096
rect 675262 357040 676292 357096
rect 675201 357038 676292 357040
rect 675201 357035 675267 357038
rect 675753 356690 675819 356693
rect 675753 356688 676292 356690
rect 675753 356632 675758 356688
rect 675814 356632 676292 356688
rect 675753 356630 676292 356632
rect 675753 356627 675819 356630
rect 676029 356282 676095 356285
rect 676029 356280 676292 356282
rect 676029 356224 676034 356280
rect 676090 356224 676292 356280
rect 676029 356222 676292 356224
rect 676029 356219 676095 356222
rect 58525 355874 58591 355877
rect 58525 355872 64706 355874
rect 58525 355816 58530 355872
rect 58586 355816 64706 355872
rect 58525 355814 64706 355816
rect 58525 355811 58591 355814
rect 41454 355676 41460 355740
rect 41524 355738 41530 355740
rect 41781 355738 41847 355741
rect 41524 355736 41847 355738
rect 41524 355680 41786 355736
rect 41842 355680 41847 355736
rect 41524 355678 41847 355680
rect 41524 355676 41530 355678
rect 41781 355675 41847 355678
rect 64646 355600 64706 355814
rect 675150 355812 675156 355876
rect 675220 355874 675226 355876
rect 675220 355814 676292 355874
rect 675220 355812 675226 355814
rect 675753 355466 675819 355469
rect 675753 355464 676292 355466
rect 675753 355408 675758 355464
rect 675814 355408 676292 355464
rect 675753 355406 676292 355408
rect 675753 355403 675819 355406
rect 58433 355058 58499 355061
rect 675661 355058 675727 355061
rect 58433 355056 64706 355058
rect 58433 355000 58438 355056
rect 58494 355000 64706 355056
rect 58433 354998 64706 355000
rect 58433 354995 58499 354998
rect 64646 354418 64706 354998
rect 675661 355056 676292 355058
rect 675661 355000 675666 355056
rect 675722 355000 676292 355056
rect 675661 354998 676292 355000
rect 675661 354995 675727 354998
rect 675293 354650 675359 354653
rect 675293 354648 676292 354650
rect 675293 354592 675298 354648
rect 675354 354592 676292 354648
rect 675293 354590 676292 354592
rect 675293 354587 675359 354590
rect 676029 354242 676095 354245
rect 676029 354240 676292 354242
rect 676029 354184 676034 354240
rect 676090 354184 676292 354240
rect 676029 354182 676292 354184
rect 676029 354179 676095 354182
rect 675385 353834 675451 353837
rect 675385 353832 676292 353834
rect 675385 353776 675390 353832
rect 675446 353776 676292 353832
rect 675385 353774 676292 353776
rect 675385 353771 675451 353774
rect 676029 353426 676095 353429
rect 676029 353424 676292 353426
rect 676029 353368 676034 353424
rect 676090 353368 676292 353424
rect 676029 353366 676292 353368
rect 676029 353363 676095 353366
rect 676029 353018 676095 353021
rect 676029 353016 676292 353018
rect 676029 352960 676034 353016
rect 676090 352960 676292 353016
rect 676029 352958 676292 352960
rect 676029 352955 676095 352958
rect 675937 352610 676003 352613
rect 675937 352608 676292 352610
rect 675937 352552 675942 352608
rect 675998 352552 676292 352608
rect 675937 352550 676292 352552
rect 675937 352547 676003 352550
rect 675937 352202 676003 352205
rect 675937 352200 676292 352202
rect 675937 352144 675942 352200
rect 675998 352144 676292 352200
rect 675937 352142 676292 352144
rect 675937 352139 676003 352142
rect 676029 351794 676095 351797
rect 676029 351792 676292 351794
rect 676029 351736 676034 351792
rect 676090 351736 676292 351792
rect 676029 351734 676292 351736
rect 676029 351731 676095 351734
rect 675937 351386 676003 351389
rect 675937 351384 676292 351386
rect 675937 351328 675942 351384
rect 675998 351328 676292 351384
rect 675937 351326 676292 351328
rect 675937 351323 676003 351326
rect 675845 350978 675911 350981
rect 675845 350976 676292 350978
rect 675845 350920 675850 350976
rect 675906 350920 676292 350976
rect 675845 350918 676292 350920
rect 675845 350915 675911 350918
rect 675661 350570 675727 350573
rect 675661 350568 676292 350570
rect 675661 350512 675666 350568
rect 675722 350512 676292 350568
rect 675661 350510 676292 350512
rect 675661 350507 675727 350510
rect 676029 350162 676095 350165
rect 676029 350160 676292 350162
rect 676029 350104 676034 350160
rect 676090 350104 676292 350160
rect 676029 350102 676292 350104
rect 676029 350099 676095 350102
rect 676029 349754 676095 349757
rect 676029 349752 676292 349754
rect 676029 349696 676034 349752
rect 676090 349696 676292 349752
rect 676029 349694 676292 349696
rect 676029 349691 676095 349694
rect 675937 349346 676003 349349
rect 675937 349344 676292 349346
rect 675937 349288 675942 349344
rect 675998 349288 676292 349344
rect 675937 349286 676292 349288
rect 675937 349283 676003 349286
rect 675845 348938 675911 348941
rect 675845 348936 676292 348938
rect 675845 348880 675850 348936
rect 675906 348880 676292 348936
rect 675845 348878 676292 348880
rect 675845 348875 675911 348878
rect 676078 348470 676292 348530
rect 676078 347309 676138 348470
rect 679022 347684 679082 348092
rect 676029 347306 676138 347309
rect 675948 347304 676292 347306
rect 675948 347248 676034 347304
rect 676090 347248 676292 347304
rect 675948 347246 676292 347248
rect 676029 347243 676095 347246
rect 41462 344317 41522 344556
rect 41462 344312 41571 344317
rect 41462 344256 41510 344312
rect 41566 344256 41571 344312
rect 41462 344254 41571 344256
rect 41505 344251 41571 344254
rect 41462 343909 41522 344148
rect 41462 343904 41571 343909
rect 41462 343848 41510 343904
rect 41566 343848 41571 343904
rect 41462 343846 41571 343848
rect 41505 343843 41571 343846
rect 41462 343501 41522 343740
rect 41462 343496 41571 343501
rect 41462 343440 41510 343496
rect 41566 343440 41571 343496
rect 41462 343438 41571 343440
rect 41505 343435 41571 343438
rect 41873 343362 41939 343365
rect 41492 343360 41939 343362
rect 41492 343304 41878 343360
rect 41934 343304 41939 343360
rect 41492 343302 41939 343304
rect 41873 343299 41939 343302
rect 41462 342685 41522 342924
rect 41462 342680 41571 342685
rect 41462 342624 41510 342680
rect 41566 342624 41571 342680
rect 41462 342622 41571 342624
rect 41505 342619 41571 342622
rect 41781 342546 41847 342549
rect 41492 342544 41847 342546
rect 41492 342488 41786 342544
rect 41842 342488 41847 342544
rect 41492 342486 41847 342488
rect 41781 342483 41847 342486
rect 41781 342138 41847 342141
rect 41492 342136 41847 342138
rect 41492 342080 41786 342136
rect 41842 342080 41847 342136
rect 41492 342078 41847 342080
rect 41781 342075 41847 342078
rect 41505 341866 41571 341869
rect 41462 341864 41571 341866
rect 41462 341808 41510 341864
rect 41566 341808 41571 341864
rect 41462 341803 41571 341808
rect 41462 341700 41522 341803
rect 41781 341322 41847 341325
rect 41492 341320 41847 341322
rect 41492 341264 41786 341320
rect 41842 341264 41847 341320
rect 41492 341262 41847 341264
rect 41781 341259 41847 341262
rect 41505 341050 41571 341053
rect 41462 341048 41571 341050
rect 41462 340992 41510 341048
rect 41566 340992 41571 341048
rect 41462 340987 41571 340992
rect 41462 340884 41522 340987
rect 41462 340236 41522 340476
rect 41454 340172 41460 340236
rect 41524 340172 41530 340236
rect 29870 339829 29930 340068
rect 29870 339824 29979 339829
rect 33041 339826 33107 339829
rect 29870 339768 29918 339824
rect 29974 339768 29979 339824
rect 29870 339766 29979 339768
rect 29913 339763 29979 339766
rect 32998 339824 33107 339826
rect 32998 339768 33046 339824
rect 33102 339768 33107 339824
rect 32998 339763 33107 339768
rect 32998 339660 33058 339763
rect 30054 339013 30114 339252
rect 30054 339008 30163 339013
rect 30054 338952 30102 339008
rect 30158 338952 30163 339008
rect 30054 338950 30163 338952
rect 30097 338947 30163 338950
rect 30054 338605 30114 338844
rect 30005 338600 30114 338605
rect 30005 338544 30010 338600
rect 30066 338544 30114 338600
rect 30005 338542 30114 338544
rect 30005 338539 30071 338542
rect 30238 338197 30298 338436
rect 30189 338192 30298 338197
rect 30189 338136 30194 338192
rect 30250 338136 30298 338192
rect 30189 338134 30298 338136
rect 30189 338131 30255 338134
rect 30238 337789 30298 338028
rect 30238 337784 30347 337789
rect 30238 337728 30286 337784
rect 30342 337728 30347 337784
rect 30238 337726 30347 337728
rect 30281 337723 30347 337726
rect 41462 337378 41522 337620
rect 41638 337378 41644 337380
rect 41462 337318 41644 337378
rect 41638 337316 41644 337318
rect 41708 337316 41714 337380
rect 41822 337242 41828 337244
rect 41492 337182 41828 337242
rect 41822 337180 41828 337182
rect 41892 337180 41898 337244
rect 42558 336834 42564 336836
rect 41492 336774 42564 336834
rect 42558 336772 42564 336774
rect 42628 336772 42634 336836
rect 41462 336157 41522 336396
rect 41462 336152 41571 336157
rect 41462 336096 41510 336152
rect 41566 336096 41571 336152
rect 41462 336094 41571 336096
rect 41505 336091 41571 336094
rect 41781 336018 41847 336021
rect 41492 336016 41847 336018
rect 41492 335960 41786 336016
rect 41842 335960 41847 336016
rect 41492 335958 41847 335960
rect 41781 335955 41847 335958
rect 41462 335338 41522 335580
rect 41597 335338 41663 335341
rect 41462 335336 41663 335338
rect 41462 335280 41602 335336
rect 41658 335280 41663 335336
rect 41462 335278 41663 335280
rect 41597 335275 41663 335278
rect 41462 334933 41522 335172
rect 41413 334928 41522 334933
rect 41413 334872 41418 334928
rect 41474 334872 41522 334928
rect 41413 334870 41522 334872
rect 41413 334867 41479 334870
rect 41462 334522 41522 334764
rect 41689 334522 41755 334525
rect 41462 334520 41755 334522
rect 41462 334464 41694 334520
rect 41750 334464 41755 334520
rect 41462 334462 41755 334464
rect 41689 334459 41755 334462
rect 41873 334386 41939 334389
rect 41492 334384 41939 334386
rect 41492 334328 41878 334384
rect 41934 334328 41939 334384
rect 41492 334326 41939 334328
rect 41873 334323 41939 334326
rect 30422 333540 30482 333948
rect 41873 333162 41939 333165
rect 41492 333160 41939 333162
rect 41492 333104 41878 333160
rect 41934 333104 41939 333160
rect 41492 333102 41939 333104
rect 41873 333099 41939 333102
rect 30097 330170 30163 330173
rect 42190 330170 42196 330172
rect 30097 330168 42196 330170
rect 30097 330112 30102 330168
rect 30158 330112 42196 330168
rect 30097 330110 42196 330112
rect 30097 330107 30163 330110
rect 42190 330108 42196 330110
rect 42260 330108 42266 330172
rect 29913 330034 29979 330037
rect 42006 330034 42012 330036
rect 29913 330032 42012 330034
rect 29913 329976 29918 330032
rect 29974 329976 42012 330032
rect 29913 329974 42012 329976
rect 29913 329971 29979 329974
rect 42006 329972 42012 329974
rect 42076 329972 42082 330036
rect 30005 329898 30071 329901
rect 42374 329898 42380 329900
rect 30005 329896 42380 329898
rect 30005 329840 30010 329896
rect 30066 329840 42380 329896
rect 30005 329838 42380 329840
rect 30005 329835 30071 329838
rect 42374 329836 42380 329838
rect 42444 329836 42450 329900
rect 655513 329898 655579 329901
rect 649950 329896 655579 329898
rect 649950 329840 655518 329896
rect 655574 329840 655579 329896
rect 649950 329838 655579 329840
rect 649950 329234 650010 329838
rect 655513 329835 655579 329838
rect 655421 328266 655487 328269
rect 649950 328264 655487 328266
rect 649950 328208 655426 328264
rect 655482 328208 655487 328264
rect 649950 328206 655487 328208
rect 649950 328052 650010 328206
rect 655421 328203 655487 328206
rect 655605 327450 655671 327453
rect 649950 327448 655671 327450
rect 649950 327392 655610 327448
rect 655666 327392 655671 327448
rect 649950 327390 655671 327392
rect 649950 326870 650010 327390
rect 655605 327387 655671 327390
rect 649950 325682 650010 325688
rect 655973 325682 656039 325685
rect 649950 325680 656039 325682
rect 649950 325624 655978 325680
rect 656034 325624 656039 325680
rect 649950 325622 656039 325624
rect 655973 325619 656039 325622
rect 58525 317386 58591 317389
rect 58525 317384 64706 317386
rect 58525 317328 58530 317384
rect 58586 317328 64706 317384
rect 58525 317326 64706 317328
rect 58525 317323 58591 317326
rect 64646 317106 64706 317326
rect 58065 316570 58131 316573
rect 58065 316568 64706 316570
rect 58065 316512 58070 316568
rect 58126 316512 64706 316568
rect 58065 316510 64706 316512
rect 58065 316507 58131 316510
rect 42425 316434 42491 316437
rect 42558 316434 42564 316436
rect 42425 316432 42564 316434
rect 42425 316376 42430 316432
rect 42486 316376 42564 316432
rect 42425 316374 42564 316376
rect 42425 316371 42491 316374
rect 42558 316372 42564 316374
rect 42628 316372 42634 316436
rect 41781 316300 41847 316301
rect 41781 316296 41828 316300
rect 41892 316298 41898 316300
rect 41781 316240 41786 316296
rect 41781 316236 41828 316240
rect 41892 316238 41938 316298
rect 41892 316236 41898 316238
rect 41781 316235 41847 316236
rect 64646 315924 64706 316510
rect 42149 315482 42215 315485
rect 42374 315482 42380 315484
rect 42149 315480 42380 315482
rect 42149 315424 42154 315480
rect 42210 315424 42380 315480
rect 42149 315422 42380 315424
rect 42149 315419 42215 315422
rect 42374 315420 42380 315422
rect 42444 315420 42450 315484
rect 58341 314802 58407 314805
rect 58341 314800 64706 314802
rect 58341 314744 58346 314800
rect 58402 314744 64706 314800
rect 58341 314742 64706 314744
rect 58341 314739 58407 314742
rect 58525 314122 58591 314125
rect 58525 314120 64706 314122
rect 58525 314064 58530 314120
rect 58586 314064 64706 314120
rect 58525 314062 64706 314064
rect 58525 314059 58591 314062
rect 41965 313852 42031 313853
rect 41965 313848 42012 313852
rect 42076 313850 42082 313852
rect 41965 313792 41970 313848
rect 41965 313788 42012 313792
rect 42076 313790 42122 313850
rect 42076 313788 42082 313790
rect 41965 313787 42031 313788
rect 64646 313560 64706 314062
rect 676262 313581 676322 313684
rect 676262 313576 676371 313581
rect 676262 313520 676310 313576
rect 676366 313520 676371 313576
rect 676262 313518 676371 313520
rect 676305 313515 676371 313518
rect 676121 313170 676187 313173
rect 676262 313170 676322 313276
rect 676121 313168 676322 313170
rect 676121 313112 676126 313168
rect 676182 313112 676322 313168
rect 676121 313110 676322 313112
rect 676121 313107 676187 313110
rect 41638 312972 41644 313036
rect 41708 313034 41714 313036
rect 41781 313034 41847 313037
rect 41708 313032 41847 313034
rect 41708 312976 41786 313032
rect 41842 312976 41847 313032
rect 41708 312974 41847 312976
rect 41708 312972 41714 312974
rect 41781 312971 41847 312974
rect 58157 313034 58223 313037
rect 58157 313032 64706 313034
rect 58157 312976 58162 313032
rect 58218 312976 64706 313032
rect 58157 312974 64706 312976
rect 58157 312971 58223 312974
rect 64646 312378 64706 312974
rect 676262 312765 676322 312868
rect 676213 312760 676322 312765
rect 676213 312704 676218 312760
rect 676274 312704 676322 312760
rect 676213 312702 676322 312704
rect 676213 312699 676279 312702
rect 676029 312490 676095 312493
rect 676029 312488 676292 312490
rect 676029 312432 676034 312488
rect 676090 312432 676292 312488
rect 676029 312430 676292 312432
rect 676029 312427 676095 312430
rect 42149 312356 42215 312357
rect 42149 312354 42196 312356
rect 42104 312352 42196 312354
rect 42104 312296 42154 312352
rect 42104 312294 42196 312296
rect 42149 312292 42196 312294
rect 42260 312292 42266 312356
rect 42149 312291 42215 312292
rect 676262 311949 676322 312052
rect 676213 311944 676322 311949
rect 676213 311888 676218 311944
rect 676274 311888 676322 311944
rect 676213 311886 676322 311888
rect 676213 311883 676279 311886
rect 58525 311810 58591 311813
rect 58525 311808 64706 311810
rect 58525 311752 58530 311808
rect 58586 311752 64706 311808
rect 58525 311750 64706 311752
rect 58525 311747 58591 311750
rect 64646 311196 64706 311750
rect 676029 311674 676095 311677
rect 676029 311672 676292 311674
rect 676029 311616 676034 311672
rect 676090 311616 676292 311672
rect 676029 311614 676292 311616
rect 676029 311611 676095 311614
rect 676262 311133 676322 311236
rect 676213 311128 676322 311133
rect 676213 311072 676218 311128
rect 676274 311072 676322 311128
rect 676213 311070 676322 311072
rect 676213 311067 676279 311070
rect 675293 310858 675359 310861
rect 675293 310856 676292 310858
rect 675293 310800 675298 310856
rect 675354 310800 676292 310856
rect 675293 310798 676292 310800
rect 675293 310795 675359 310798
rect 676262 310317 676322 310420
rect 676213 310312 676322 310317
rect 676213 310256 676218 310312
rect 676274 310256 676322 310312
rect 676213 310254 676322 310256
rect 676213 310251 676279 310254
rect 676029 310042 676095 310045
rect 676029 310040 676292 310042
rect 676029 309984 676034 310040
rect 676090 309984 676292 310040
rect 676029 309982 676292 309984
rect 676029 309979 676095 309982
rect 676262 309501 676322 309604
rect 676213 309496 676322 309501
rect 676213 309440 676218 309496
rect 676274 309440 676322 309496
rect 676213 309438 676322 309440
rect 676213 309435 676279 309438
rect 676029 309226 676095 309229
rect 676029 309224 676292 309226
rect 676029 309168 676034 309224
rect 676090 309168 676292 309224
rect 676029 309166 676292 309168
rect 676029 309163 676095 309166
rect 676029 308818 676095 308821
rect 676029 308816 676292 308818
rect 676029 308760 676034 308816
rect 676090 308760 676292 308816
rect 676029 308758 676292 308760
rect 676029 308755 676095 308758
rect 675753 308410 675819 308413
rect 675753 308408 676292 308410
rect 675753 308352 675758 308408
rect 675814 308352 676292 308408
rect 675753 308350 676292 308352
rect 675753 308347 675819 308350
rect 676029 308002 676095 308005
rect 676029 308000 676292 308002
rect 676029 307944 676034 308000
rect 676090 307944 676292 308000
rect 676029 307942 676292 307944
rect 676029 307939 676095 307942
rect 676121 307458 676187 307461
rect 676262 307458 676322 307564
rect 676121 307456 676322 307458
rect 676121 307400 676126 307456
rect 676182 307400 676322 307456
rect 676121 307398 676322 307400
rect 676121 307395 676187 307398
rect 676029 307186 676095 307189
rect 676029 307184 676292 307186
rect 676029 307128 676034 307184
rect 676090 307128 676292 307184
rect 676029 307126 676292 307128
rect 676029 307123 676095 307126
rect 676029 306778 676095 306781
rect 676029 306776 676292 306778
rect 676029 306720 676034 306776
rect 676090 306720 676292 306776
rect 676029 306718 676292 306720
rect 676029 306715 676095 306718
rect 675293 306370 675359 306373
rect 675293 306368 676292 306370
rect 675293 306312 675298 306368
rect 675354 306312 676292 306368
rect 675293 306310 676292 306312
rect 675293 306307 675359 306310
rect 676029 305962 676095 305965
rect 676029 305960 676292 305962
rect 676029 305904 676034 305960
rect 676090 305904 676292 305960
rect 676029 305902 676292 305904
rect 676029 305899 676095 305902
rect 676121 305418 676187 305421
rect 676262 305418 676322 305524
rect 676121 305416 676322 305418
rect 676121 305360 676126 305416
rect 676182 305360 676322 305416
rect 676121 305358 676322 305360
rect 676121 305355 676187 305358
rect 676121 305010 676187 305013
rect 676262 305010 676322 305116
rect 676121 305008 676322 305010
rect 676121 304952 676126 305008
rect 676182 304952 676322 305008
rect 676121 304950 676322 304952
rect 676121 304947 676187 304950
rect 676029 304738 676095 304741
rect 676029 304736 676292 304738
rect 676029 304680 676034 304736
rect 676090 304680 676292 304736
rect 676029 304678 676292 304680
rect 676029 304675 676095 304678
rect 676121 304194 676187 304197
rect 676262 304194 676322 304300
rect 676121 304192 676322 304194
rect 676121 304136 676126 304192
rect 676182 304136 676322 304192
rect 676121 304134 676322 304136
rect 676121 304131 676187 304134
rect 676029 303922 676095 303925
rect 676029 303920 676292 303922
rect 676029 303864 676034 303920
rect 676090 303864 676292 303920
rect 676029 303862 676292 303864
rect 676029 303859 676095 303862
rect 679022 303381 679082 303484
rect 655513 303378 655579 303381
rect 649950 303376 655579 303378
rect 649950 303320 655518 303376
rect 655574 303320 655579 303376
rect 649950 303318 655579 303320
rect 649950 302776 650010 303318
rect 655513 303315 655579 303318
rect 678973 303376 679082 303381
rect 678973 303320 678978 303376
rect 679034 303320 679082 303376
rect 678973 303318 679082 303320
rect 678973 303315 679039 303318
rect 684542 302668 684602 303076
rect 678973 302562 679039 302565
rect 678973 302560 679082 302562
rect 678973 302504 678978 302560
rect 679034 302504 679082 302560
rect 678973 302499 679082 302504
rect 679022 302260 679082 302499
rect 655697 302154 655763 302157
rect 649950 302152 655763 302154
rect 649950 302096 655702 302152
rect 655758 302096 655763 302152
rect 649950 302094 655763 302096
rect 649950 301594 650010 302094
rect 655697 302091 655763 302094
rect 41965 301338 42031 301341
rect 41492 301336 42031 301338
rect 41492 301280 41970 301336
rect 42026 301280 42031 301336
rect 41492 301278 42031 301280
rect 41965 301275 42031 301278
rect 27521 300930 27587 300933
rect 27508 300928 27587 300930
rect 27508 300872 27526 300928
rect 27582 300872 27587 300928
rect 27508 300870 27587 300872
rect 27521 300867 27587 300870
rect 655421 300794 655487 300797
rect 649950 300792 655487 300794
rect 649950 300736 655426 300792
rect 655482 300736 655487 300792
rect 649950 300734 655487 300736
rect 41873 300522 41939 300525
rect 41492 300520 41939 300522
rect 41492 300464 41878 300520
rect 41934 300464 41939 300520
rect 41492 300462 41939 300464
rect 41873 300459 41939 300462
rect 649950 300412 650010 300734
rect 655421 300731 655487 300734
rect 41781 300114 41847 300117
rect 41492 300112 41847 300114
rect 41492 300056 41786 300112
rect 41842 300056 41847 300112
rect 41492 300054 41847 300056
rect 41781 300051 41847 300054
rect 42057 299706 42123 299709
rect 41492 299704 42123 299706
rect 41492 299648 42062 299704
rect 42118 299648 42123 299704
rect 41492 299646 42123 299648
rect 42057 299643 42123 299646
rect 41781 299298 41847 299301
rect 41492 299296 41847 299298
rect 41492 299240 41786 299296
rect 41842 299240 41847 299296
rect 41492 299238 41847 299240
rect 41781 299235 41847 299238
rect 42425 298890 42491 298893
rect 41492 298888 42491 298890
rect 41492 298832 42430 298888
rect 42486 298832 42491 298888
rect 41492 298830 42491 298832
rect 42425 298827 42491 298830
rect 649950 298754 650010 299230
rect 655053 298754 655119 298757
rect 649950 298752 655119 298754
rect 649950 298696 655058 298752
rect 655114 298696 655119 298752
rect 649950 298694 655119 298696
rect 655053 298691 655119 298694
rect 41781 298482 41847 298485
rect 41492 298480 41847 298482
rect 41492 298424 41786 298480
rect 41842 298424 41847 298480
rect 41492 298422 41847 298424
rect 41781 298419 41847 298422
rect 41781 298074 41847 298077
rect 41492 298072 41847 298074
rect 41492 298016 41786 298072
rect 41842 298016 41847 298072
rect 41492 298014 41847 298016
rect 41781 298011 41847 298014
rect 41822 297666 41828 297668
rect 41492 297606 41828 297666
rect 41822 297604 41828 297606
rect 41892 297604 41898 297668
rect 649950 297530 650010 298048
rect 656065 297530 656131 297533
rect 649950 297528 656131 297530
rect 649950 297472 656070 297528
rect 656126 297472 656131 297528
rect 649950 297470 656131 297472
rect 656065 297467 656131 297470
rect 41781 297258 41847 297261
rect 41492 297256 41847 297258
rect 41492 297200 41786 297256
rect 41842 297200 41847 297256
rect 41492 297198 41847 297200
rect 41781 297195 41847 297198
rect 41822 296850 41828 296852
rect 41492 296790 41828 296850
rect 41822 296788 41828 296790
rect 41892 296788 41898 296852
rect 35801 296442 35867 296445
rect 35788 296440 35867 296442
rect 35788 296384 35806 296440
rect 35862 296384 35867 296440
rect 35788 296382 35867 296384
rect 35801 296379 35867 296382
rect 649950 296306 650010 296866
rect 655881 296306 655947 296309
rect 649950 296304 655947 296306
rect 649950 296248 655886 296304
rect 655942 296248 655947 296304
rect 649950 296246 655947 296248
rect 655881 296243 655947 296246
rect 41822 296034 41828 296036
rect 41492 295974 41828 296034
rect 41822 295972 41828 295974
rect 41892 295972 41898 296036
rect 41822 295626 41828 295628
rect 41492 295566 41828 295626
rect 41822 295564 41828 295566
rect 41892 295564 41898 295628
rect 58525 295490 58591 295493
rect 64646 295490 64706 295684
rect 58525 295488 64706 295490
rect 58525 295432 58530 295488
rect 58586 295432 64706 295488
rect 58525 295430 64706 295432
rect 58525 295427 58591 295430
rect 649950 295354 650010 295684
rect 656249 295354 656315 295357
rect 649950 295352 656315 295354
rect 649950 295296 656254 295352
rect 656310 295296 656315 295352
rect 649950 295294 656315 295296
rect 656249 295291 656315 295294
rect 41492 295158 41752 295218
rect 41692 295085 41752 295158
rect 41689 295080 41755 295085
rect 41689 295024 41694 295080
rect 41750 295024 41755 295080
rect 41689 295019 41755 295024
rect 41781 294810 41847 294813
rect 41492 294808 41847 294810
rect 41492 294752 41786 294808
rect 41842 294752 41847 294808
rect 41492 294750 41847 294752
rect 41781 294747 41847 294750
rect 42006 294402 42012 294404
rect 41492 294342 42012 294402
rect 42006 294340 42012 294342
rect 42076 294340 42082 294404
rect 42057 293994 42123 293997
rect 41492 293992 42123 293994
rect 41492 293936 42062 293992
rect 42118 293936 42123 293992
rect 41492 293934 42123 293936
rect 42057 293931 42123 293934
rect 58433 293994 58499 293997
rect 64646 293994 64706 294502
rect 58433 293992 64706 293994
rect 58433 293936 58438 293992
rect 58494 293936 64706 293992
rect 58433 293934 64706 293936
rect 649950 293994 650010 294502
rect 655697 293994 655763 293997
rect 649950 293992 655763 293994
rect 649950 293936 655702 293992
rect 655758 293936 655763 293992
rect 649950 293934 655763 293936
rect 58433 293931 58499 293934
rect 655697 293931 655763 293934
rect 42057 293586 42123 293589
rect 41492 293584 42123 293586
rect 41492 293528 42062 293584
rect 42118 293528 42123 293584
rect 41492 293526 42123 293528
rect 42057 293523 42123 293526
rect 42057 293178 42123 293181
rect 41492 293176 42123 293178
rect 41492 293120 42062 293176
rect 42118 293120 42123 293176
rect 41492 293118 42123 293120
rect 42057 293115 42123 293118
rect 42149 292770 42215 292773
rect 41492 292768 42215 292770
rect 41492 292712 42154 292768
rect 42210 292712 42215 292768
rect 41492 292710 42215 292712
rect 42149 292707 42215 292710
rect 59261 292770 59327 292773
rect 64646 292770 64706 293320
rect 59261 292768 64706 292770
rect 59261 292712 59266 292768
rect 59322 292712 64706 292768
rect 59261 292710 64706 292712
rect 649950 292770 650010 293320
rect 655513 292770 655579 292773
rect 649950 292768 655579 292770
rect 649950 292712 655518 292768
rect 655574 292712 655579 292768
rect 649950 292710 655579 292712
rect 59261 292707 59327 292710
rect 655513 292707 655579 292710
rect 41873 292362 41939 292365
rect 41492 292360 41939 292362
rect 41492 292304 41878 292360
rect 41934 292304 41939 292360
rect 41492 292302 41939 292304
rect 41873 292299 41939 292302
rect 58525 292362 58591 292365
rect 58525 292360 64706 292362
rect 58525 292304 58530 292360
rect 58586 292304 64706 292360
rect 58525 292302 64706 292304
rect 58525 292299 58591 292302
rect 64646 292138 64706 292302
rect 41965 291954 42031 291957
rect 41492 291952 42031 291954
rect 41492 291896 41970 291952
rect 42026 291896 42031 291952
rect 41492 291894 42031 291896
rect 41965 291891 42031 291894
rect 42701 291546 42767 291549
rect 41492 291544 42767 291546
rect 41492 291488 42706 291544
rect 42762 291488 42767 291544
rect 41492 291486 42767 291488
rect 42701 291483 42767 291486
rect 57973 291546 58039 291549
rect 649950 291546 650010 292138
rect 655789 291546 655855 291549
rect 57973 291544 64706 291546
rect 57973 291488 57978 291544
rect 58034 291488 64706 291544
rect 57973 291486 64706 291488
rect 649950 291544 655855 291546
rect 649950 291488 655794 291544
rect 655850 291488 655855 291544
rect 649950 291486 655855 291488
rect 57973 291483 58039 291486
rect 41781 291138 41847 291141
rect 41492 291136 41847 291138
rect 41492 291080 41786 291136
rect 41842 291080 41847 291136
rect 41492 291078 41847 291080
rect 41781 291075 41847 291078
rect 64646 290956 64706 291486
rect 655789 291483 655855 291486
rect 41781 290730 41847 290733
rect 41492 290728 41847 290730
rect 41492 290672 41786 290728
rect 41842 290672 41847 290728
rect 41492 290670 41847 290672
rect 41781 290667 41847 290670
rect 649950 290458 650010 290956
rect 655605 290458 655671 290461
rect 649950 290456 655671 290458
rect 649950 290400 655610 290456
rect 655666 290400 655671 290456
rect 649950 290398 655671 290400
rect 655605 290395 655671 290398
rect 41781 289914 41847 289917
rect 41492 289912 41847 289914
rect 41492 289856 41786 289912
rect 41842 289856 41847 289912
rect 41492 289854 41847 289856
rect 41781 289851 41847 289854
rect 57973 289778 58039 289781
rect 57973 289776 64706 289778
rect 57973 289720 57978 289776
rect 58034 289720 64706 289776
rect 57973 289718 64706 289720
rect 57973 289715 58039 289718
rect 649950 289234 650010 289774
rect 654501 289234 654567 289237
rect 649950 289232 654567 289234
rect 649950 289176 654506 289232
rect 654562 289176 654567 289232
rect 649950 289174 654567 289176
rect 654501 289171 654567 289174
rect 58157 288010 58223 288013
rect 64646 288010 64706 288592
rect 58157 288008 64706 288010
rect 58157 287952 58162 288008
rect 58218 287952 64706 288008
rect 58157 287950 64706 287952
rect 649950 288010 650010 288592
rect 654869 288010 654935 288013
rect 649950 288008 654935 288010
rect 649950 287952 654874 288008
rect 654930 287952 654935 288008
rect 649950 287950 654935 287952
rect 58157 287947 58223 287950
rect 654869 287947 654935 287950
rect 58525 287194 58591 287197
rect 64646 287194 64706 287410
rect 649766 287406 651390 287466
rect 651330 287330 651390 287406
rect 656801 287330 656867 287333
rect 651330 287328 656867 287330
rect 651330 287272 656806 287328
rect 656862 287272 656867 287328
rect 651330 287270 656867 287272
rect 656801 287267 656867 287270
rect 58525 287192 64706 287194
rect 58525 287136 58530 287192
rect 58586 287136 64706 287192
rect 58525 287134 64706 287136
rect 58525 287131 58591 287134
rect 57973 285698 58039 285701
rect 64646 285698 64706 286228
rect 57973 285696 64706 285698
rect 57973 285640 57978 285696
rect 58034 285640 64706 285696
rect 57973 285638 64706 285640
rect 649950 285698 650010 286228
rect 655421 285698 655487 285701
rect 649950 285696 655487 285698
rect 649950 285640 655426 285696
rect 655482 285640 655487 285696
rect 649950 285638 655487 285640
rect 57973 285635 58039 285638
rect 655421 285635 655487 285638
rect 58525 284474 58591 284477
rect 64646 284474 64706 285046
rect 649950 284746 650010 285046
rect 654869 284746 654935 284749
rect 649950 284744 654935 284746
rect 649950 284688 654874 284744
rect 654930 284688 654935 284744
rect 649950 284686 654935 284688
rect 654869 284683 654935 284686
rect 58525 284472 64706 284474
rect 58525 284416 58530 284472
rect 58586 284416 64706 284472
rect 58525 284414 64706 284416
rect 58525 284411 58591 284414
rect 58525 283250 58591 283253
rect 64646 283250 64706 283864
rect 58525 283248 64706 283250
rect 58525 283192 58530 283248
rect 58586 283192 64706 283248
rect 58525 283190 64706 283192
rect 649950 283250 650010 283864
rect 655421 283250 655487 283253
rect 649950 283248 655487 283250
rect 649950 283192 655426 283248
rect 655482 283192 655487 283248
rect 649950 283190 655487 283192
rect 58525 283187 58591 283190
rect 655421 283187 655487 283190
rect 58249 282162 58315 282165
rect 64646 282162 64706 282682
rect 58249 282160 64706 282162
rect 58249 282104 58254 282160
rect 58310 282104 64706 282160
rect 58249 282102 64706 282104
rect 649950 282162 650010 282682
rect 656801 282162 656867 282165
rect 649950 282160 656867 282162
rect 649950 282104 656806 282160
rect 656862 282104 656867 282160
rect 649950 282102 656867 282104
rect 58249 282099 58315 282102
rect 656801 282099 656867 282102
rect 58157 280938 58223 280941
rect 64646 280938 64706 281500
rect 58157 280936 64706 280938
rect 58157 280880 58162 280936
rect 58218 280880 64706 280936
rect 58157 280878 64706 280880
rect 649950 280938 650010 281500
rect 654685 280938 654751 280941
rect 649950 280936 654751 280938
rect 649950 280880 654690 280936
rect 654746 280880 654751 280936
rect 649950 280878 654751 280880
rect 58157 280875 58223 280878
rect 654685 280875 654751 280878
rect 58249 279714 58315 279717
rect 64646 279714 64706 280318
rect 649950 279986 650010 280318
rect 654869 279986 654935 279989
rect 649950 279984 654935 279986
rect 649950 279928 654874 279984
rect 654930 279928 654935 279984
rect 649950 279926 654935 279928
rect 654869 279923 654935 279926
rect 58249 279712 64706 279714
rect 58249 279656 58254 279712
rect 58310 279656 64706 279712
rect 58249 279654 64706 279656
rect 58249 279651 58315 279654
rect 394969 275906 395035 275909
rect 603625 275906 603691 275909
rect 394969 275904 603691 275906
rect 394969 275848 394974 275904
rect 395030 275848 603630 275904
rect 603686 275848 603691 275904
rect 394969 275846 603691 275848
rect 394969 275843 395035 275846
rect 603625 275843 603691 275846
rect 397361 275770 397427 275773
rect 609605 275770 609671 275773
rect 397361 275768 609671 275770
rect 397361 275712 397366 275768
rect 397422 275712 609610 275768
rect 609666 275712 609671 275768
rect 397361 275710 609671 275712
rect 397361 275707 397427 275710
rect 609605 275707 609671 275710
rect 398465 275634 398531 275637
rect 613101 275634 613167 275637
rect 398465 275632 613167 275634
rect 398465 275576 398470 275632
rect 398526 275576 613106 275632
rect 613162 275576 613167 275632
rect 398465 275574 613167 275576
rect 398465 275571 398531 275574
rect 613101 275571 613167 275574
rect 400397 275498 400463 275501
rect 617793 275498 617859 275501
rect 400397 275496 617859 275498
rect 400397 275440 400402 275496
rect 400458 275440 617798 275496
rect 617854 275440 617859 275496
rect 400397 275438 617859 275440
rect 400397 275435 400463 275438
rect 617793 275435 617859 275438
rect 401133 275362 401199 275365
rect 620185 275362 620251 275365
rect 401133 275360 620251 275362
rect 401133 275304 401138 275360
rect 401194 275304 620190 275360
rect 620246 275304 620251 275360
rect 401133 275302 620251 275304
rect 401133 275299 401199 275302
rect 620185 275299 620251 275302
rect 399845 275226 399911 275229
rect 616689 275226 616755 275229
rect 399845 275224 616755 275226
rect 399845 275168 399850 275224
rect 399906 275168 616694 275224
rect 616750 275168 616755 275224
rect 399845 275166 616755 275168
rect 399845 275163 399911 275166
rect 616689 275163 616755 275166
rect 402605 275090 402671 275093
rect 623773 275090 623839 275093
rect 402605 275088 623839 275090
rect 402605 275032 402610 275088
rect 402666 275032 623778 275088
rect 623834 275032 623839 275088
rect 402605 275030 623839 275032
rect 402605 275027 402671 275030
rect 623773 275027 623839 275030
rect 403985 274954 404051 274957
rect 627269 274954 627335 274957
rect 403985 274952 627335 274954
rect 403985 274896 403990 274952
rect 404046 274896 627274 274952
rect 627330 274896 627335 274952
rect 403985 274894 627335 274896
rect 403985 274891 404051 274894
rect 627269 274891 627335 274894
rect 405181 274818 405247 274821
rect 630857 274818 630923 274821
rect 405181 274816 630923 274818
rect 405181 274760 405186 274816
rect 405242 274760 630862 274816
rect 630918 274760 630923 274816
rect 405181 274758 630923 274760
rect 405181 274755 405247 274758
rect 630857 274755 630923 274758
rect 406929 274682 406995 274685
rect 635549 274682 635615 274685
rect 406929 274680 635615 274682
rect 406929 274624 406934 274680
rect 406990 274624 635554 274680
rect 635610 274624 635615 274680
rect 406929 274622 635615 274624
rect 406929 274619 406995 274622
rect 635549 274619 635615 274622
rect 408125 274546 408191 274549
rect 637941 274546 638007 274549
rect 408125 274544 638007 274546
rect 408125 274488 408130 274544
rect 408186 274488 637946 274544
rect 638002 274488 638007 274544
rect 408125 274486 638007 274488
rect 408125 274483 408191 274486
rect 637941 274483 638007 274486
rect 391013 274410 391079 274413
rect 593045 274410 593111 274413
rect 391013 274408 593111 274410
rect 391013 274352 391018 274408
rect 391074 274352 593050 274408
rect 593106 274352 593111 274408
rect 391013 274350 593111 274352
rect 391013 274347 391079 274350
rect 593045 274347 593111 274350
rect 388253 274274 388319 274277
rect 585961 274274 586027 274277
rect 388253 274272 586027 274274
rect 388253 274216 388258 274272
rect 388314 274216 585966 274272
rect 586022 274216 586027 274272
rect 388253 274214 586027 274216
rect 388253 274211 388319 274214
rect 585961 274211 586027 274214
rect 385585 274138 385651 274141
rect 578877 274138 578943 274141
rect 385585 274136 578943 274138
rect 385585 274080 385590 274136
rect 385646 274080 578882 274136
rect 578938 274080 578943 274136
rect 385585 274078 578943 274080
rect 385585 274075 385651 274078
rect 578877 274075 578943 274078
rect 110781 273186 110847 273189
rect 209405 273186 209471 273189
rect 110781 273184 209471 273186
rect 110781 273128 110786 273184
rect 110842 273128 209410 273184
rect 209466 273128 209471 273184
rect 110781 273126 209471 273128
rect 110781 273123 110847 273126
rect 209405 273123 209471 273126
rect 365989 273186 366055 273189
rect 526805 273186 526871 273189
rect 365989 273184 526871 273186
rect 365989 273128 365994 273184
rect 366050 273128 526810 273184
rect 526866 273128 526871 273184
rect 365989 273126 526871 273128
rect 365989 273123 366055 273126
rect 526805 273123 526871 273126
rect 109585 273050 109651 273053
rect 206737 273050 206803 273053
rect 109585 273048 206803 273050
rect 109585 272992 109590 273048
rect 109646 272992 206742 273048
rect 206798 272992 206803 273048
rect 109585 272990 206803 272992
rect 109585 272987 109651 272990
rect 206737 272987 206803 272990
rect 365529 273050 365595 273053
rect 525609 273050 525675 273053
rect 365529 273048 525675 273050
rect 365529 272992 365534 273048
rect 365590 272992 525614 273048
rect 525670 272992 525675 273048
rect 365529 272990 525675 272992
rect 365529 272987 365595 272990
rect 525609 272987 525675 272990
rect 104893 272914 104959 272917
rect 206461 272914 206527 272917
rect 104893 272912 206527 272914
rect 104893 272856 104898 272912
rect 104954 272856 206466 272912
rect 206522 272856 206527 272912
rect 104893 272854 206527 272856
rect 104893 272851 104959 272854
rect 206461 272851 206527 272854
rect 368657 272914 368723 272917
rect 533889 272914 533955 272917
rect 368657 272912 533955 272914
rect 368657 272856 368662 272912
rect 368718 272856 533894 272912
rect 533950 272856 533955 272912
rect 368657 272854 533955 272856
rect 368657 272851 368723 272854
rect 533889 272851 533955 272854
rect 103697 272778 103763 272781
rect 207381 272778 207447 272781
rect 103697 272776 207447 272778
rect 103697 272720 103702 272776
rect 103758 272720 207386 272776
rect 207442 272720 207447 272776
rect 103697 272718 207447 272720
rect 103697 272715 103763 272718
rect 207381 272715 207447 272718
rect 370865 272778 370931 272781
rect 539869 272778 539935 272781
rect 370865 272776 539935 272778
rect 370865 272720 370870 272776
rect 370926 272720 539874 272776
rect 539930 272720 539935 272776
rect 370865 272718 539935 272720
rect 370865 272715 370931 272718
rect 539869 272715 539935 272718
rect 95417 272642 95483 272645
rect 203517 272642 203583 272645
rect 95417 272640 203583 272642
rect 95417 272584 95422 272640
rect 95478 272584 203522 272640
rect 203578 272584 203583 272640
rect 95417 272582 203583 272584
rect 95417 272579 95483 272582
rect 203517 272579 203583 272582
rect 371325 272642 371391 272645
rect 540973 272642 541039 272645
rect 371325 272640 541039 272642
rect 371325 272584 371330 272640
rect 371386 272584 540978 272640
rect 541034 272584 541039 272640
rect 371325 272582 541039 272584
rect 371325 272579 371391 272582
rect 540973 272579 541039 272582
rect 90725 272506 90791 272509
rect 201953 272506 202019 272509
rect 90725 272504 202019 272506
rect 90725 272448 90730 272504
rect 90786 272448 201958 272504
rect 202014 272448 202019 272504
rect 90725 272446 202019 272448
rect 90725 272443 90791 272446
rect 201953 272443 202019 272446
rect 373993 272506 374059 272509
rect 548057 272506 548123 272509
rect 373993 272504 548123 272506
rect 373993 272448 373998 272504
rect 374054 272448 548062 272504
rect 548118 272448 548123 272504
rect 373993 272446 548123 272448
rect 373993 272443 374059 272446
rect 548057 272443 548123 272446
rect 41781 272372 41847 272373
rect 41781 272368 41828 272372
rect 41892 272370 41898 272372
rect 84745 272370 84811 272373
rect 199101 272370 199167 272373
rect 41781 272312 41786 272368
rect 41781 272308 41828 272312
rect 41892 272310 41938 272370
rect 84745 272368 199167 272370
rect 84745 272312 84750 272368
rect 84806 272312 199106 272368
rect 199162 272312 199167 272368
rect 84745 272310 199167 272312
rect 41892 272308 41898 272310
rect 41781 272307 41847 272308
rect 84745 272307 84811 272310
rect 199101 272307 199167 272310
rect 387425 272370 387491 272373
rect 583569 272370 583635 272373
rect 387425 272368 583635 272370
rect 387425 272312 387430 272368
rect 387486 272312 583574 272368
rect 583630 272312 583635 272368
rect 387425 272310 583635 272312
rect 387425 272307 387491 272310
rect 583569 272307 583635 272310
rect 81249 272234 81315 272237
rect 198089 272234 198155 272237
rect 81249 272232 198155 272234
rect 81249 272176 81254 272232
rect 81310 272176 198094 272232
rect 198150 272176 198155 272232
rect 81249 272174 198155 272176
rect 81249 272171 81315 272174
rect 198089 272171 198155 272174
rect 395429 272234 395495 272237
rect 604821 272234 604887 272237
rect 395429 272232 604887 272234
rect 395429 272176 395434 272232
rect 395490 272176 604826 272232
rect 604882 272176 604887 272232
rect 395429 272174 604887 272176
rect 395429 272171 395495 272174
rect 604821 272171 604887 272174
rect 80053 272098 80119 272101
rect 196893 272098 196959 272101
rect 80053 272096 196959 272098
rect 80053 272040 80058 272096
rect 80114 272040 196898 272096
rect 196954 272040 196959 272096
rect 80053 272038 196959 272040
rect 80053 272035 80119 272038
rect 196893 272035 196959 272038
rect 403433 272098 403499 272101
rect 626073 272098 626139 272101
rect 403433 272096 626139 272098
rect 403433 272040 403438 272096
rect 403494 272040 626078 272096
rect 626134 272040 626139 272096
rect 403433 272038 626139 272040
rect 403433 272035 403499 272038
rect 626073 272035 626139 272038
rect 83641 271962 83707 271965
rect 199377 271962 199443 271965
rect 83641 271960 199443 271962
rect 83641 271904 83646 271960
rect 83702 271904 199382 271960
rect 199438 271904 199443 271960
rect 83641 271902 199443 271904
rect 83641 271899 83707 271902
rect 199377 271899 199443 271902
rect 408769 271962 408835 271965
rect 640333 271962 640399 271965
rect 408769 271960 640399 271962
rect 408769 271904 408774 271960
rect 408830 271904 640338 271960
rect 640394 271904 640399 271960
rect 408769 271902 640399 271904
rect 408769 271899 408835 271902
rect 640333 271899 640399 271902
rect 69381 271826 69447 271829
rect 193673 271826 193739 271829
rect 69381 271824 193739 271826
rect 69381 271768 69386 271824
rect 69442 271768 193678 271824
rect 193734 271768 193739 271824
rect 69381 271766 193739 271768
rect 69381 271763 69447 271766
rect 193673 271763 193739 271766
rect 410517 271826 410583 271829
rect 645025 271826 645091 271829
rect 410517 271824 645091 271826
rect 410517 271768 410522 271824
rect 410578 271768 645030 271824
rect 645086 271768 645091 271824
rect 410517 271766 645091 271768
rect 410517 271763 410583 271766
rect 645025 271763 645091 271766
rect 120257 271690 120323 271693
rect 212349 271690 212415 271693
rect 120257 271688 212415 271690
rect 120257 271632 120262 271688
rect 120318 271632 212354 271688
rect 212410 271632 212415 271688
rect 120257 271630 212415 271632
rect 120257 271627 120323 271630
rect 212349 271627 212415 271630
rect 363321 271690 363387 271693
rect 519721 271690 519787 271693
rect 363321 271688 519787 271690
rect 363321 271632 363326 271688
rect 363382 271632 519726 271688
rect 519782 271632 519787 271688
rect 363321 271630 519787 271632
rect 363321 271627 363387 271630
rect 519721 271627 519787 271630
rect 124949 271554 125015 271557
rect 215017 271554 215083 271557
rect 124949 271552 215083 271554
rect 124949 271496 124954 271552
rect 125010 271496 215022 271552
rect 215078 271496 215083 271552
rect 124949 271494 215083 271496
rect 124949 271491 125015 271494
rect 215017 271491 215083 271494
rect 360653 271554 360719 271557
rect 512637 271554 512703 271557
rect 360653 271552 512703 271554
rect 360653 271496 360658 271552
rect 360714 271496 512642 271552
rect 512698 271496 512703 271552
rect 360653 271494 512703 271496
rect 360653 271491 360719 271494
rect 512637 271491 512703 271494
rect 134425 271418 134491 271421
rect 218145 271418 218211 271421
rect 134425 271416 218211 271418
rect 134425 271360 134430 271416
rect 134486 271360 218150 271416
rect 218206 271360 218211 271416
rect 134425 271358 218211 271360
rect 134425 271355 134491 271358
rect 218145 271355 218211 271358
rect 357985 271418 358051 271421
rect 505553 271418 505619 271421
rect 357985 271416 505619 271418
rect 357985 271360 357990 271416
rect 358046 271360 505558 271416
rect 505614 271360 505619 271416
rect 357985 271358 505619 271360
rect 357985 271355 358051 271358
rect 505553 271355 505619 271358
rect 132033 271282 132099 271285
rect 217685 271282 217751 271285
rect 132033 271280 217751 271282
rect 132033 271224 132038 271280
rect 132094 271224 217690 271280
rect 217746 271224 217751 271280
rect 132033 271222 217751 271224
rect 132033 271219 132099 271222
rect 217685 271219 217751 271222
rect 357525 271282 357591 271285
rect 504357 271282 504423 271285
rect 357525 271280 504423 271282
rect 357525 271224 357530 271280
rect 357586 271224 504362 271280
rect 504418 271224 504423 271280
rect 357525 271222 504423 271224
rect 357525 271219 357591 271222
rect 504357 271219 504423 271222
rect 133229 271146 133295 271149
rect 217317 271146 217383 271149
rect 133229 271144 217383 271146
rect 133229 271088 133234 271144
rect 133290 271088 217322 271144
rect 217378 271088 217383 271144
rect 133229 271086 217383 271088
rect 133229 271083 133295 271086
rect 217317 271083 217383 271086
rect 355317 271146 355383 271149
rect 498469 271146 498535 271149
rect 355317 271144 498535 271146
rect 355317 271088 355322 271144
rect 355378 271088 498474 271144
rect 498530 271088 498535 271144
rect 355317 271086 498535 271088
rect 355317 271083 355383 271086
rect 498469 271083 498535 271086
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 114369 270466 114435 270469
rect 210693 270466 210759 270469
rect 114369 270464 210759 270466
rect 114369 270408 114374 270464
rect 114430 270408 210698 270464
rect 210754 270408 210759 270464
rect 114369 270406 210759 270408
rect 114369 270403 114435 270406
rect 210693 270403 210759 270406
rect 364241 270466 364307 270469
rect 522113 270466 522179 270469
rect 364241 270464 522179 270466
rect 364241 270408 364246 270464
rect 364302 270408 522118 270464
rect 522174 270408 522179 270464
rect 364241 270406 522179 270408
rect 364241 270403 364307 270406
rect 522113 270403 522179 270406
rect 108389 270330 108455 270333
rect 207933 270330 207999 270333
rect 108389 270328 207999 270330
rect 108389 270272 108394 270328
rect 108450 270272 207938 270328
rect 207994 270272 207999 270328
rect 108389 270270 207999 270272
rect 108389 270267 108455 270270
rect 207933 270267 207999 270270
rect 366909 270330 366975 270333
rect 529197 270330 529263 270333
rect 366909 270328 529263 270330
rect 366909 270272 366914 270328
rect 366970 270272 529202 270328
rect 529258 270272 529263 270328
rect 366909 270270 529263 270272
rect 366909 270267 366975 270270
rect 529197 270267 529263 270270
rect 107193 270194 107259 270197
rect 208393 270194 208459 270197
rect 107193 270192 208459 270194
rect 107193 270136 107198 270192
rect 107254 270136 208398 270192
rect 208454 270136 208459 270192
rect 107193 270134 208459 270136
rect 107193 270131 107259 270134
rect 208393 270131 208459 270134
rect 369577 270194 369643 270197
rect 536281 270194 536347 270197
rect 369577 270192 536347 270194
rect 369577 270136 369582 270192
rect 369638 270136 536286 270192
rect 536342 270136 536347 270192
rect 369577 270134 536347 270136
rect 369577 270131 369643 270134
rect 536281 270131 536347 270134
rect 106089 270058 106155 270061
rect 207473 270058 207539 270061
rect 106089 270056 207539 270058
rect 106089 270000 106094 270056
rect 106150 270000 207478 270056
rect 207534 270000 207539 270056
rect 106089 269998 207539 270000
rect 106089 269995 106155 269998
rect 207473 269995 207539 269998
rect 372245 270058 372311 270061
rect 543365 270058 543431 270061
rect 372245 270056 543431 270058
rect 372245 270000 372250 270056
rect 372306 270000 543370 270056
rect 543426 270000 543431 270056
rect 372245 269998 543431 270000
rect 372245 269995 372311 269998
rect 543365 269995 543431 269998
rect 99005 269922 99071 269925
rect 204805 269922 204871 269925
rect 99005 269920 204871 269922
rect 99005 269864 99010 269920
rect 99066 269864 204810 269920
rect 204866 269864 204871 269920
rect 99005 269862 204871 269864
rect 99005 269859 99071 269862
rect 204805 269859 204871 269862
rect 380709 269922 380775 269925
rect 565813 269922 565879 269925
rect 380709 269920 565879 269922
rect 380709 269864 380714 269920
rect 380770 269864 565818 269920
rect 565874 269864 565879 269920
rect 380709 269862 565879 269864
rect 380709 269859 380775 269862
rect 565813 269859 565879 269862
rect 41965 269788 42031 269789
rect 41965 269784 42012 269788
rect 42076 269786 42082 269788
rect 93025 269786 93091 269789
rect 203057 269786 203123 269789
rect 41965 269728 41970 269784
rect 41965 269724 42012 269728
rect 42076 269726 42122 269786
rect 93025 269784 203123 269786
rect 93025 269728 93030 269784
rect 93086 269728 203062 269784
rect 203118 269728 203123 269784
rect 93025 269726 203123 269728
rect 42076 269724 42082 269726
rect 41965 269723 42031 269724
rect 93025 269723 93091 269726
rect 203057 269723 203123 269726
rect 383377 269786 383443 269789
rect 572897 269786 572963 269789
rect 383377 269784 572963 269786
rect 383377 269728 383382 269784
rect 383438 269728 572902 269784
rect 572958 269728 572963 269784
rect 383377 269726 572963 269728
rect 383377 269723 383443 269726
rect 572897 269723 572963 269726
rect 85941 269650 86007 269653
rect 199929 269650 199995 269653
rect 85941 269648 199995 269650
rect 85941 269592 85946 269648
rect 86002 269592 199934 269648
rect 199990 269592 199995 269648
rect 85941 269590 199995 269592
rect 85941 269587 86007 269590
rect 199929 269587 199995 269590
rect 399385 269650 399451 269653
rect 615493 269650 615559 269653
rect 399385 269648 615559 269650
rect 399385 269592 399390 269648
rect 399446 269592 615498 269648
rect 615554 269592 615559 269648
rect 399385 269590 615559 269592
rect 399385 269587 399451 269590
rect 615493 269587 615559 269590
rect 87137 269514 87203 269517
rect 200389 269514 200455 269517
rect 87137 269512 200455 269514
rect 87137 269456 87142 269512
rect 87198 269456 200394 269512
rect 200450 269456 200455 269512
rect 87137 269454 200455 269456
rect 87137 269451 87203 269454
rect 200389 269451 200455 269454
rect 404721 269514 404787 269517
rect 629661 269514 629727 269517
rect 404721 269512 629727 269514
rect 404721 269456 404726 269512
rect 404782 269456 629666 269512
rect 629722 269456 629727 269512
rect 404721 269454 629727 269456
rect 404721 269451 404787 269454
rect 629661 269451 629727 269454
rect 41638 269316 41644 269380
rect 41708 269378 41714 269380
rect 41781 269378 41847 269381
rect 41708 269376 41847 269378
rect 41708 269320 41786 269376
rect 41842 269320 41847 269376
rect 41708 269318 41847 269320
rect 41708 269316 41714 269318
rect 41781 269315 41847 269318
rect 78857 269378 78923 269381
rect 197721 269378 197787 269381
rect 78857 269376 197787 269378
rect 78857 269320 78862 269376
rect 78918 269320 197726 269376
rect 197782 269320 197787 269376
rect 78857 269318 197787 269320
rect 78857 269315 78923 269318
rect 197721 269315 197787 269318
rect 198733 269378 198799 269381
rect 204345 269378 204411 269381
rect 198733 269376 204411 269378
rect 198733 269320 198738 269376
rect 198794 269320 204350 269376
rect 204406 269320 204411 269376
rect 198733 269318 204411 269320
rect 198733 269315 198799 269318
rect 204345 269315 204411 269318
rect 407389 269378 407455 269381
rect 636745 269378 636811 269381
rect 407389 269376 636811 269378
rect 407389 269320 407394 269376
rect 407450 269320 636750 269376
rect 636806 269320 636811 269376
rect 407389 269318 636811 269320
rect 407389 269315 407455 269318
rect 636745 269315 636811 269318
rect 76465 269242 76531 269245
rect 195973 269242 196039 269245
rect 76465 269240 196039 269242
rect 76465 269184 76470 269240
rect 76526 269184 195978 269240
rect 196034 269184 196039 269240
rect 76465 269182 196039 269184
rect 76465 269179 76531 269182
rect 195973 269179 196039 269182
rect 410793 269242 410859 269245
rect 646221 269242 646287 269245
rect 410793 269240 646287 269242
rect 410793 269184 410798 269240
rect 410854 269184 646226 269240
rect 646282 269184 646287 269240
rect 410793 269182 646287 269184
rect 410793 269179 410859 269182
rect 646221 269179 646287 269182
rect 70577 269106 70643 269109
rect 194133 269106 194199 269109
rect 70577 269104 194199 269106
rect 70577 269048 70582 269104
rect 70638 269048 194138 269104
rect 194194 269048 194199 269104
rect 70577 269046 194199 269048
rect 70577 269043 70643 269046
rect 194133 269043 194199 269046
rect 411897 269106 411963 269109
rect 648613 269106 648679 269109
rect 411897 269104 648679 269106
rect 411897 269048 411902 269104
rect 411958 269048 648618 269104
rect 648674 269048 648679 269104
rect 411897 269046 648679 269048
rect 411897 269043 411963 269046
rect 648613 269043 648679 269046
rect 121453 268970 121519 268973
rect 213729 268970 213795 268973
rect 121453 268968 213795 268970
rect 121453 268912 121458 268968
rect 121514 268912 213734 268968
rect 213790 268912 213795 268968
rect 121453 268910 213795 268912
rect 121453 268907 121519 268910
rect 213729 268907 213795 268910
rect 362033 268970 362099 268973
rect 516225 268970 516291 268973
rect 362033 268968 516291 268970
rect 362033 268912 362038 268968
rect 362094 268912 516230 268968
rect 516286 268912 516291 268968
rect 362033 268910 516291 268912
rect 362033 268907 362099 268910
rect 516225 268907 516291 268910
rect 184933 268834 184999 268837
rect 201217 268834 201283 268837
rect 184933 268832 201283 268834
rect 184933 268776 184938 268832
rect 184994 268776 201222 268832
rect 201278 268776 201283 268832
rect 184933 268774 201283 268776
rect 184933 268771 184999 268774
rect 201217 268771 201283 268774
rect 359365 268834 359431 268837
rect 509049 268834 509115 268837
rect 359365 268832 509115 268834
rect 359365 268776 359370 268832
rect 359426 268776 509054 268832
rect 509110 268776 509115 268832
rect 359365 268774 509115 268776
rect 359365 268771 359431 268774
rect 509049 268771 509115 268774
rect 356605 268698 356671 268701
rect 501965 268698 502031 268701
rect 356605 268696 502031 268698
rect 356605 268640 356610 268696
rect 356666 268640 501970 268696
rect 502026 268640 502031 268696
rect 356605 268638 502031 268640
rect 356605 268635 356671 268638
rect 501965 268635 502031 268638
rect 676121 268562 676187 268565
rect 676262 268562 676322 268668
rect 676121 268560 676322 268562
rect 676121 268504 676126 268560
rect 676182 268504 676322 268560
rect 676121 268502 676322 268504
rect 676121 268499 676187 268502
rect 676029 268290 676095 268293
rect 676029 268288 676292 268290
rect 676029 268232 676034 268288
rect 676090 268232 676292 268288
rect 676029 268230 676292 268232
rect 676029 268227 676095 268230
rect 676213 268154 676279 268157
rect 676213 268152 676322 268154
rect 676213 268096 676218 268152
rect 676274 268096 676322 268152
rect 676213 268091 676322 268096
rect 676262 267852 676322 268091
rect 405457 267746 405523 267749
rect 477309 267746 477375 267749
rect 405457 267744 477375 267746
rect 405457 267688 405462 267744
rect 405518 267688 477314 267744
rect 477370 267688 477375 267744
rect 405457 267686 477375 267688
rect 405457 267683 405523 267686
rect 477309 267683 477375 267686
rect 398925 267610 398991 267613
rect 471973 267610 472039 267613
rect 398925 267608 472039 267610
rect 398925 267552 398930 267608
rect 398986 267552 471978 267608
rect 472034 267552 472039 267608
rect 398925 267550 472039 267552
rect 398925 267547 398991 267550
rect 471973 267547 472039 267550
rect 396257 267474 396323 267477
rect 485681 267474 485747 267477
rect 396257 267472 485747 267474
rect 396257 267416 396262 267472
rect 396318 267416 485686 267472
rect 485742 267416 485747 267472
rect 396257 267414 485747 267416
rect 396257 267411 396323 267414
rect 485681 267411 485747 267414
rect 676029 267474 676095 267477
rect 676029 267472 676292 267474
rect 676029 267416 676034 267472
rect 676090 267416 676292 267472
rect 676029 267414 676292 267416
rect 676029 267411 676095 267414
rect 393589 267338 393655 267341
rect 497917 267338 497983 267341
rect 393589 267336 497983 267338
rect 393589 267280 393594 267336
rect 393650 267280 497922 267336
rect 497978 267280 497983 267336
rect 393589 267278 497983 267280
rect 393589 267275 393655 267278
rect 497917 267275 497983 267278
rect 387793 267202 387859 267205
rect 584765 267202 584831 267205
rect 387793 267200 584831 267202
rect 387793 267144 387798 267200
rect 387854 267144 584770 267200
rect 584826 267144 584831 267200
rect 387793 267142 584831 267144
rect 387793 267139 387859 267142
rect 584765 267139 584831 267142
rect 386965 267066 387031 267069
rect 582373 267066 582439 267069
rect 386965 267064 582439 267066
rect 386965 267008 386970 267064
rect 387026 267008 582378 267064
rect 582434 267008 582439 267064
rect 386965 267006 582439 267008
rect 386965 267003 387031 267006
rect 582373 267003 582439 267006
rect 675661 267066 675727 267069
rect 675661 267064 676292 267066
rect 675661 267008 675666 267064
rect 675722 267008 676292 267064
rect 675661 267006 676292 267008
rect 675661 267003 675727 267006
rect 389633 266930 389699 266933
rect 589457 266930 589523 266933
rect 389633 266928 589523 266930
rect 389633 266872 389638 266928
rect 389694 266872 589462 266928
rect 589518 266872 589523 266928
rect 389633 266870 589523 266872
rect 389633 266867 389699 266870
rect 589457 266867 589523 266870
rect 390461 266794 390527 266797
rect 591849 266794 591915 266797
rect 390461 266792 591915 266794
rect 390461 266736 390466 266792
rect 390522 266736 591854 266792
rect 591910 266736 591915 266792
rect 390461 266734 591915 266736
rect 390461 266731 390527 266734
rect 591849 266731 591915 266734
rect 391841 266658 391907 266661
rect 595345 266658 595411 266661
rect 391841 266656 595411 266658
rect 391841 266600 391846 266656
rect 391902 266600 595350 266656
rect 595406 266600 595411 266656
rect 391841 266598 595411 266600
rect 391841 266595 391907 266598
rect 595345 266595 595411 266598
rect 676029 266658 676095 266661
rect 676029 266656 676292 266658
rect 676029 266600 676034 266656
rect 676090 266600 676292 266656
rect 676029 266598 676292 266600
rect 676029 266595 676095 266598
rect 393129 266522 393195 266525
rect 598933 266522 598999 266525
rect 393129 266520 598999 266522
rect 393129 266464 393134 266520
rect 393190 266464 598938 266520
rect 598994 266464 598999 266520
rect 393129 266462 598999 266464
rect 393129 266459 393195 266462
rect 598933 266459 598999 266462
rect 394509 266386 394575 266389
rect 602429 266386 602495 266389
rect 394509 266384 602495 266386
rect 394509 266328 394514 266384
rect 394570 266328 602434 266384
rect 602490 266328 602495 266384
rect 394509 266326 602495 266328
rect 394509 266323 394575 266326
rect 602429 266323 602495 266326
rect 408309 266250 408375 266253
rect 436093 266250 436159 266253
rect 408309 266248 436159 266250
rect 408309 266192 408314 266248
rect 408370 266192 436098 266248
rect 436154 266192 436159 266248
rect 408309 266190 436159 266192
rect 408309 266187 408375 266190
rect 436093 266187 436159 266190
rect 675753 266250 675819 266253
rect 675753 266248 676292 266250
rect 675753 266192 675758 266248
rect 675814 266192 676292 266248
rect 675753 266190 676292 266192
rect 675753 266187 675819 266190
rect 676029 265842 676095 265845
rect 676029 265840 676292 265842
rect 676029 265784 676034 265840
rect 676090 265784 676292 265840
rect 676029 265782 676292 265784
rect 676029 265779 676095 265782
rect 676070 265236 676076 265300
rect 676140 265298 676146 265300
rect 676262 265298 676322 265404
rect 676140 265238 676322 265298
rect 676140 265236 676146 265238
rect 676262 264893 676322 264996
rect 676213 264888 676322 264893
rect 676213 264832 676218 264888
rect 676274 264832 676322 264888
rect 676213 264830 676322 264832
rect 676213 264827 676279 264830
rect 676029 264618 676095 264621
rect 676029 264616 676292 264618
rect 676029 264560 676034 264616
rect 676090 264560 676292 264616
rect 676029 264558 676292 264560
rect 676029 264555 676095 264558
rect 676029 264210 676095 264213
rect 676029 264208 676292 264210
rect 676029 264152 676034 264208
rect 676090 264152 676292 264208
rect 676029 264150 676292 264152
rect 676029 264147 676095 264150
rect 676121 263666 676187 263669
rect 676262 263666 676322 263772
rect 676121 263664 676322 263666
rect 676121 263608 676126 263664
rect 676182 263608 676322 263664
rect 676121 263606 676322 263608
rect 676121 263603 676187 263606
rect 675477 263394 675543 263397
rect 675477 263392 676292 263394
rect 675477 263336 675482 263392
rect 675538 263336 676292 263392
rect 675477 263334 676292 263336
rect 675477 263331 675543 263334
rect 676029 262986 676095 262989
rect 676029 262984 676292 262986
rect 676029 262928 676034 262984
rect 676090 262928 676292 262984
rect 676029 262926 676292 262928
rect 676029 262923 676095 262926
rect 675937 262578 676003 262581
rect 675937 262576 676292 262578
rect 675937 262520 675942 262576
rect 675998 262520 676292 262576
rect 675937 262518 676292 262520
rect 675937 262515 676003 262518
rect 412380 262320 573116 262334
rect 412380 262274 573044 262320
rect 573039 262260 573044 262274
rect 573104 262274 573116 262320
rect 573104 262260 573109 262274
rect 573039 262255 573109 262260
rect 676029 262170 676095 262173
rect 676029 262168 676292 262170
rect 676029 262112 676034 262168
rect 676090 262112 676292 262168
rect 676029 262110 676292 262112
rect 676029 262107 676095 262110
rect 675845 261762 675911 261765
rect 675845 261760 676292 261762
rect 675845 261704 675850 261760
rect 675906 261704 676292 261760
rect 675845 261702 676292 261704
rect 675845 261699 675911 261702
rect 676029 261354 676095 261357
rect 676029 261352 676292 261354
rect 676029 261296 676034 261352
rect 676090 261296 676292 261352
rect 676029 261294 676292 261296
rect 676029 261291 676095 261294
rect 676121 260810 676187 260813
rect 676262 260810 676322 260916
rect 676121 260808 676322 260810
rect 676121 260752 676126 260808
rect 676182 260752 676322 260808
rect 676121 260750 676322 260752
rect 676121 260747 676187 260750
rect 675937 260538 676003 260541
rect 675937 260536 676292 260538
rect 675937 260480 675942 260536
rect 675998 260480 676292 260536
rect 675937 260478 676292 260480
rect 675937 260475 676003 260478
rect 675937 260130 676003 260133
rect 675937 260128 676292 260130
rect 675937 260072 675942 260128
rect 675998 260072 676292 260128
rect 675937 260070 676292 260072
rect 675937 260067 676003 260070
rect 676029 259722 676095 259725
rect 676029 259720 676292 259722
rect 676029 259664 676034 259720
rect 676090 259664 676292 259720
rect 676029 259662 676292 259664
rect 676029 259659 676095 259662
rect 676029 259314 676095 259317
rect 676029 259312 676292 259314
rect 676029 259256 676034 259312
rect 676090 259256 676292 259312
rect 676029 259254 676292 259256
rect 676029 259251 676095 259254
rect 572213 259186 572283 259189
rect 412380 259184 572292 259186
rect 412380 259126 572218 259184
rect 572213 259124 572218 259126
rect 572278 259126 572292 259184
rect 572278 259124 572283 259126
rect 572213 259119 572283 259124
rect 676121 258770 676187 258773
rect 676262 258770 676322 258876
rect 676121 258768 676322 258770
rect 676121 258712 676126 258768
rect 676182 258712 676322 258768
rect 676121 258710 676322 258712
rect 676121 258707 676187 258710
rect 184933 258634 184999 258637
rect 184933 258632 191820 258634
rect 184933 258576 184938 258632
rect 184994 258576 191820 258632
rect 184933 258574 191820 258576
rect 184933 258571 184999 258574
rect 679022 258365 679082 258468
rect 678973 258360 679082 258365
rect 678973 258304 678978 258360
rect 679034 258304 679082 258360
rect 678973 258302 679082 258304
rect 678973 258299 679039 258302
rect 41462 257957 41522 258060
rect 41462 257952 41571 257957
rect 41462 257896 41510 257952
rect 41566 257896 41571 257952
rect 41462 257894 41571 257896
rect 41505 257891 41571 257894
rect 41873 257682 41939 257685
rect 41492 257680 41939 257682
rect 41492 257624 41878 257680
rect 41934 257624 41939 257680
rect 684542 257652 684602 258060
rect 41492 257622 41939 257624
rect 41873 257619 41939 257622
rect 41597 257546 41663 257549
rect 41462 257544 41663 257546
rect 41462 257488 41602 257544
rect 41658 257488 41663 257544
rect 41462 257486 41663 257488
rect 41462 257244 41522 257486
rect 41597 257483 41663 257486
rect 678973 257546 679039 257549
rect 678973 257544 679082 257546
rect 678973 257488 678978 257544
rect 679034 257488 679082 257544
rect 678973 257483 679082 257488
rect 679022 257244 679082 257483
rect 41781 256866 41847 256869
rect 41492 256864 41847 256866
rect 41492 256808 41786 256864
rect 41842 256808 41847 256864
rect 41492 256806 41847 256808
rect 41781 256803 41847 256806
rect 41873 256458 41939 256461
rect 41492 256456 41939 256458
rect 41492 256400 41878 256456
rect 41934 256400 41939 256456
rect 41492 256398 41939 256400
rect 41873 256395 41939 256398
rect 41505 256322 41571 256325
rect 41462 256320 41571 256322
rect 41462 256264 41510 256320
rect 41566 256264 41571 256320
rect 41462 256259 41571 256264
rect 41462 256020 41522 256259
rect 412336 255912 571470 255924
rect 412336 255864 571394 255912
rect 571389 255852 571394 255864
rect 571454 255864 571470 255912
rect 571454 255852 571459 255864
rect 571389 255847 571459 255852
rect 39990 255508 40050 255612
rect 39982 255444 39988 255508
rect 40052 255444 40058 255508
rect 41505 255506 41571 255509
rect 41462 255504 41571 255506
rect 41462 255448 41510 255504
rect 41566 255448 41571 255504
rect 41462 255443 41571 255448
rect 41462 255204 41522 255443
rect 41781 254826 41847 254829
rect 41492 254824 41847 254826
rect 41492 254768 41786 254824
rect 41842 254768 41847 254824
rect 41492 254766 41847 254768
rect 41781 254763 41847 254766
rect 41505 254690 41571 254693
rect 41462 254688 41571 254690
rect 41462 254632 41510 254688
rect 41566 254632 41571 254688
rect 41462 254627 41571 254632
rect 41462 254388 41522 254627
rect 41873 254010 41939 254013
rect 41492 254008 41939 254010
rect 41492 253952 41878 254008
rect 41934 253952 41939 254008
rect 41492 253950 41939 253952
rect 41873 253947 41939 253950
rect 42057 253602 42123 253605
rect 41492 253600 42123 253602
rect 41492 253544 42062 253600
rect 42118 253544 42123 253600
rect 41492 253542 42123 253544
rect 42057 253539 42123 253542
rect 41462 253058 41522 253164
rect 41689 253058 41755 253061
rect 41462 253056 41755 253058
rect 41462 253000 41694 253056
rect 41750 253000 41755 253056
rect 41462 252998 41755 253000
rect 41689 252995 41755 252998
rect 41873 252786 41939 252789
rect 416773 252786 416839 252789
rect 41492 252784 41939 252786
rect 41492 252728 41878 252784
rect 41934 252728 41939 252784
rect 41492 252726 41939 252728
rect 412436 252784 416839 252786
rect 412436 252728 416778 252784
rect 416834 252728 416839 252784
rect 412436 252726 416839 252728
rect 41873 252723 41939 252726
rect 416773 252723 416839 252726
rect 41965 252378 42031 252381
rect 41492 252376 42031 252378
rect 41492 252320 41970 252376
rect 42026 252320 42031 252376
rect 41492 252318 42031 252320
rect 41965 252315 42031 252318
rect 41781 251970 41847 251973
rect 41492 251968 41847 251970
rect 41492 251912 41786 251968
rect 41842 251912 41847 251968
rect 41492 251910 41847 251912
rect 41781 251907 41847 251910
rect 41094 251429 41154 251532
rect 41094 251424 41203 251429
rect 41094 251368 41142 251424
rect 41198 251368 41203 251424
rect 41094 251366 41203 251368
rect 41137 251363 41203 251366
rect 35758 251021 35818 251124
rect 35758 251016 35867 251021
rect 35758 250960 35806 251016
rect 35862 250960 35867 251016
rect 35758 250958 35867 250960
rect 35801 250955 35867 250958
rect 38518 250613 38578 250716
rect 38469 250608 38578 250613
rect 38469 250552 38474 250608
rect 38530 250552 38578 250608
rect 38469 250550 38578 250552
rect 38469 250547 38535 250550
rect 38518 250205 38578 250308
rect 38518 250200 38627 250205
rect 38518 250144 38566 250200
rect 38622 250144 38627 250200
rect 38518 250142 38627 250144
rect 38561 250139 38627 250142
rect 675201 250202 675267 250205
rect 676070 250202 676076 250204
rect 675201 250200 676076 250202
rect 675201 250144 675206 250200
rect 675262 250144 676076 250200
rect 675201 250142 676076 250144
rect 675201 250139 675267 250142
rect 676070 250140 676076 250142
rect 676140 250140 676146 250204
rect 41278 249797 41338 249900
rect 41229 249792 41338 249797
rect 41229 249736 41234 249792
rect 41290 249736 41338 249792
rect 41229 249734 41338 249736
rect 41229 249731 41295 249734
rect 42333 249522 42399 249525
rect 416773 249522 416839 249525
rect 41492 249520 42399 249522
rect 41492 249464 42338 249520
rect 42394 249464 42399 249520
rect 41492 249462 42399 249464
rect 412436 249520 416839 249522
rect 412436 249464 416778 249520
rect 416834 249464 416839 249520
rect 412436 249462 416839 249464
rect 42333 249459 42399 249462
rect 416773 249459 416839 249462
rect 41462 248978 41522 249084
rect 41597 248978 41663 248981
rect 41462 248976 41663 248978
rect 41462 248920 41602 248976
rect 41658 248920 41663 248976
rect 41462 248918 41663 248920
rect 41597 248915 41663 248918
rect 41462 248573 41522 248676
rect 41413 248568 41522 248573
rect 41413 248512 41418 248568
rect 41474 248512 41522 248568
rect 41413 248510 41522 248512
rect 41413 248507 41479 248510
rect 41278 248165 41338 248268
rect 41278 248160 41387 248165
rect 41278 248104 41326 248160
rect 41382 248104 41387 248160
rect 41278 248102 41387 248104
rect 41321 248099 41387 248102
rect 187601 248026 187667 248029
rect 187601 248024 191820 248026
rect 187601 247968 187606 248024
rect 187662 247968 191820 248024
rect 187601 247966 191820 247968
rect 187601 247963 187667 247966
rect 41462 247757 41522 247860
rect 41462 247752 41571 247757
rect 41462 247696 41510 247752
rect 41566 247696 41571 247752
rect 41462 247694 41571 247696
rect 41505 247691 41571 247694
rect 41462 247349 41522 247452
rect 41462 247344 41571 247349
rect 41462 247288 41510 247344
rect 41566 247288 41571 247344
rect 41462 247286 41571 247288
rect 41505 247283 41571 247286
rect 41462 246533 41522 246636
rect 41462 246528 41571 246533
rect 41462 246472 41510 246528
rect 41566 246472 41571 246528
rect 41462 246470 41571 246472
rect 41505 246467 41571 246470
rect 416773 246394 416839 246397
rect 412436 246392 416839 246394
rect 412436 246336 416778 246392
rect 416834 246336 416839 246392
rect 412436 246334 416839 246336
rect 416773 246331 416839 246334
rect 675201 246260 675267 246261
rect 675150 246258 675156 246260
rect 675110 246198 675156 246258
rect 675220 246256 675267 246260
rect 675262 246200 675267 246256
rect 675150 246196 675156 246198
rect 675220 246196 675267 246200
rect 675201 246195 675267 246196
rect 418061 243130 418127 243133
rect 412436 243128 418127 243130
rect 412436 243072 418066 243128
rect 418122 243072 418127 243128
rect 412436 243070 418127 243072
rect 418061 243067 418127 243070
rect 41965 242314 42031 242317
rect 43846 242314 43852 242316
rect 41965 242312 43852 242314
rect 41965 242256 41970 242312
rect 42026 242256 43852 242312
rect 41965 242254 43852 242256
rect 41965 242251 42031 242254
rect 43846 242252 43852 242254
rect 43916 242252 43922 242316
rect 42057 242178 42123 242181
rect 44030 242178 44036 242180
rect 42057 242176 44036 242178
rect 42057 242120 42062 242176
rect 42118 242120 44036 242176
rect 42057 242118 44036 242120
rect 42057 242115 42123 242118
rect 44030 242116 44036 242118
rect 44100 242116 44106 242180
rect 418153 240002 418219 240005
rect 412436 240000 418219 240002
rect 412436 239944 418158 240000
rect 418214 239944 418219 240000
rect 412436 239942 418219 239944
rect 418153 239939 418219 239942
rect 43529 238098 43595 238101
rect 43662 238098 43668 238100
rect 43529 238096 43668 238098
rect 43529 238040 43534 238096
rect 43590 238040 43668 238096
rect 43529 238038 43668 238040
rect 43529 238035 43595 238038
rect 43662 238036 43668 238038
rect 43732 238036 43738 238100
rect 184933 237418 184999 237421
rect 184933 237416 191820 237418
rect 184933 237360 184938 237416
rect 184994 237360 191820 237416
rect 184933 237358 191820 237360
rect 184933 237355 184999 237358
rect 418429 236738 418495 236741
rect 412436 236736 418495 236738
rect 412436 236680 418434 236736
rect 418490 236680 418495 236736
rect 412436 236678 418495 236680
rect 418429 236675 418495 236678
rect 418521 233610 418587 233613
rect 412436 233608 418587 233610
rect 412436 233552 418526 233608
rect 418582 233552 418587 233608
rect 412436 233550 418587 233552
rect 418521 233547 418587 233550
rect 93025 228986 93091 228989
rect 210049 228986 210115 228989
rect 93025 228984 210115 228986
rect 93025 228928 93030 228984
rect 93086 228928 210054 228984
rect 210110 228928 210115 228984
rect 93025 228926 210115 228928
rect 93025 228923 93091 228926
rect 210049 228923 210115 228926
rect 256693 228986 256759 228989
rect 261753 228986 261819 228989
rect 256693 228984 261819 228986
rect 256693 228928 256698 228984
rect 256754 228928 261758 228984
rect 261814 228928 261819 228984
rect 256693 228926 261819 228928
rect 256693 228923 256759 228926
rect 261753 228923 261819 228926
rect 384757 228986 384823 228989
rect 507393 228986 507459 228989
rect 384757 228984 507459 228986
rect 384757 228928 384762 228984
rect 384818 228928 507398 228984
rect 507454 228928 507459 228984
rect 384757 228926 507459 228928
rect 384757 228923 384823 228926
rect 507393 228923 507459 228926
rect 42425 228850 42491 228853
rect 43846 228850 43852 228852
rect 42425 228848 43852 228850
rect 42425 228792 42430 228848
rect 42486 228792 43852 228848
rect 42425 228790 43852 228792
rect 42425 228787 42491 228790
rect 43846 228788 43852 228790
rect 43916 228788 43922 228852
rect 84653 228850 84719 228853
rect 206185 228850 206251 228853
rect 84653 228848 206251 228850
rect 84653 228792 84658 228848
rect 84714 228792 206190 228848
rect 206246 228792 206251 228848
rect 84653 228790 206251 228792
rect 84653 228787 84719 228790
rect 206185 228787 206251 228790
rect 245837 228850 245903 228853
rect 261385 228850 261451 228853
rect 245837 228848 261451 228850
rect 245837 228792 245842 228848
rect 245898 228792 261390 228848
rect 261446 228792 261451 228848
rect 245837 228790 261451 228792
rect 245837 228787 245903 228790
rect 261385 228787 261451 228790
rect 386873 228850 386939 228853
rect 512177 228850 512243 228853
rect 386873 228848 512243 228850
rect 386873 228792 386878 228848
rect 386934 228792 512182 228848
rect 512238 228792 512243 228848
rect 386873 228790 512243 228792
rect 386873 228787 386939 228790
rect 512177 228787 512243 228790
rect 42425 228714 42491 228717
rect 44030 228714 44036 228716
rect 42425 228712 44036 228714
rect 42425 228656 42430 228712
rect 42486 228656 44036 228712
rect 42425 228654 44036 228656
rect 42425 228651 42491 228654
rect 44030 228652 44036 228654
rect 44100 228652 44106 228716
rect 88057 228714 88123 228717
rect 207565 228714 207631 228717
rect 88057 228712 207631 228714
rect 88057 228656 88062 228712
rect 88118 228656 207570 228712
rect 207626 228656 207631 228712
rect 88057 228654 207631 228656
rect 88057 228651 88123 228654
rect 207565 228651 207631 228654
rect 390093 228714 390159 228717
rect 518985 228714 519051 228717
rect 390093 228712 519051 228714
rect 390093 228656 390098 228712
rect 390154 228656 518990 228712
rect 519046 228656 519051 228712
rect 390093 228654 519051 228656
rect 390093 228651 390159 228654
rect 518985 228651 519051 228654
rect 86309 228578 86375 228581
rect 207197 228578 207263 228581
rect 86309 228576 207263 228578
rect 86309 228520 86314 228576
rect 86370 228520 207202 228576
rect 207258 228520 207263 228576
rect 86309 228518 207263 228520
rect 86309 228515 86375 228518
rect 207197 228515 207263 228518
rect 234797 228578 234863 228581
rect 259637 228578 259703 228581
rect 234797 228576 259703 228578
rect 234797 228520 234802 228576
rect 234858 228520 259642 228576
rect 259698 228520 259703 228576
rect 234797 228518 259703 228520
rect 234797 228515 234863 228518
rect 259637 228515 259703 228518
rect 392209 228578 392275 228581
rect 525057 228578 525123 228581
rect 392209 228576 525123 228578
rect 392209 228520 392214 228576
rect 392270 228520 525062 228576
rect 525118 228520 525123 228576
rect 392209 228518 525123 228520
rect 392209 228515 392275 228518
rect 525057 228515 525123 228518
rect 82721 228442 82787 228445
rect 205817 228442 205883 228445
rect 82721 228440 205883 228442
rect 82721 228384 82726 228440
rect 82782 228384 205822 228440
rect 205878 228384 205883 228440
rect 82721 228382 205883 228384
rect 82721 228379 82787 228382
rect 205817 228379 205883 228382
rect 234613 228442 234679 228445
rect 262489 228442 262555 228445
rect 234613 228440 262555 228442
rect 234613 228384 234618 228440
rect 234674 228384 262494 228440
rect 262550 228384 262555 228440
rect 234613 228382 262555 228384
rect 234613 228379 234679 228382
rect 262489 228379 262555 228382
rect 394417 228442 394483 228445
rect 530117 228442 530183 228445
rect 394417 228440 530183 228442
rect 394417 228384 394422 228440
rect 394478 228384 530122 228440
rect 530178 228384 530183 228440
rect 394417 228382 530183 228384
rect 394417 228379 394483 228382
rect 530117 228379 530183 228382
rect 76281 228306 76347 228309
rect 202965 228306 203031 228309
rect 76281 228304 203031 228306
rect 76281 228248 76286 228304
rect 76342 228248 202970 228304
rect 203026 228248 203031 228304
rect 76281 228246 203031 228248
rect 76281 228243 76347 228246
rect 202965 228243 203031 228246
rect 225965 228306 226031 228309
rect 266077 228306 266143 228309
rect 225965 228304 266143 228306
rect 225965 228248 225970 228304
rect 226026 228248 266082 228304
rect 266138 228248 266143 228304
rect 225965 228246 266143 228248
rect 225965 228243 226031 228246
rect 266077 228243 266143 228246
rect 396533 228306 396599 228309
rect 534901 228306 534967 228309
rect 396533 228304 534967 228306
rect 396533 228248 396538 228304
rect 396594 228248 534906 228304
rect 534962 228248 534967 228304
rect 396533 228246 534967 228248
rect 396533 228243 396599 228246
rect 534901 228243 534967 228246
rect 69473 228170 69539 228173
rect 200113 228170 200179 228173
rect 69473 228168 200179 228170
rect 69473 228112 69478 228168
rect 69534 228112 200118 228168
rect 200174 228112 200179 228168
rect 69473 228110 200179 228112
rect 69473 228107 69539 228110
rect 200113 228107 200179 228110
rect 219249 228170 219315 228173
rect 263225 228170 263291 228173
rect 219249 228168 263291 228170
rect 219249 228112 219254 228168
rect 219310 228112 263230 228168
rect 263286 228112 263291 228168
rect 219249 228110 263291 228112
rect 219249 228107 219315 228110
rect 263225 228107 263291 228110
rect 398649 228170 398715 228173
rect 538305 228170 538371 228173
rect 398649 228168 538371 228170
rect 398649 228112 398654 228168
rect 398710 228112 538310 228168
rect 538366 228112 538371 228168
rect 398649 228110 538371 228112
rect 398649 228107 398715 228110
rect 538305 228107 538371 228110
rect 71221 228034 71287 228037
rect 200481 228034 200547 228037
rect 71221 228032 200547 228034
rect 71221 227976 71226 228032
rect 71282 227976 200486 228032
rect 200542 227976 200547 228032
rect 71221 227974 200547 227976
rect 71221 227971 71287 227974
rect 200481 227971 200547 227974
rect 220721 228034 220787 228037
rect 264237 228034 264303 228037
rect 220721 228032 264303 228034
rect 220721 227976 220726 228032
rect 220782 227976 264242 228032
rect 264298 227976 264303 228032
rect 220721 227974 264303 227976
rect 220721 227971 220787 227974
rect 264237 227971 264303 227974
rect 399753 228034 399819 228037
rect 542721 228034 542787 228037
rect 399753 228032 542787 228034
rect 399753 227976 399758 228032
rect 399814 227976 542726 228032
rect 542782 227976 542787 228032
rect 399753 227974 542787 227976
rect 399753 227971 399819 227974
rect 542721 227971 542787 227974
rect 62757 227898 62823 227901
rect 197261 227898 197327 227901
rect 62757 227896 197327 227898
rect 62757 227840 62762 227896
rect 62818 227840 197266 227896
rect 197322 227840 197327 227896
rect 62757 227838 197327 227840
rect 62757 227835 62823 227838
rect 197261 227835 197327 227838
rect 217593 227898 217659 227901
rect 262857 227898 262923 227901
rect 217593 227896 262923 227898
rect 217593 227840 217598 227896
rect 217654 227840 262862 227896
rect 262918 227840 262923 227896
rect 217593 227838 262923 227840
rect 217593 227835 217659 227838
rect 262857 227835 262923 227838
rect 403985 227898 404051 227901
rect 552565 227898 552631 227901
rect 403985 227896 552631 227898
rect 403985 227840 403990 227896
rect 404046 227840 552570 227896
rect 552626 227840 552631 227896
rect 403985 227838 552631 227840
rect 403985 227835 404051 227838
rect 552565 227835 552631 227838
rect 57605 227762 57671 227765
rect 194777 227762 194843 227765
rect 57605 227760 194843 227762
rect 57605 227704 57610 227760
rect 57666 227704 194782 227760
rect 194838 227704 194843 227760
rect 57605 227702 194843 227704
rect 57605 227699 57671 227702
rect 194777 227699 194843 227702
rect 212349 227762 212415 227765
rect 260373 227762 260439 227765
rect 212349 227760 260439 227762
rect 212349 227704 212354 227760
rect 212410 227704 260378 227760
rect 260434 227704 260439 227760
rect 212349 227702 260439 227704
rect 212349 227699 212415 227702
rect 260373 227699 260439 227702
rect 410057 227762 410123 227765
rect 566825 227762 566891 227765
rect 410057 227760 566891 227762
rect 410057 227704 410062 227760
rect 410118 227704 566830 227760
rect 566886 227704 566891 227760
rect 410057 227702 566891 227704
rect 410057 227699 410123 227702
rect 566825 227699 566891 227702
rect 56041 227626 56107 227629
rect 194409 227626 194475 227629
rect 56041 227624 194475 227626
rect 56041 227568 56046 227624
rect 56102 227568 194414 227624
rect 194470 227568 194475 227624
rect 56041 227566 194475 227568
rect 56041 227563 56107 227566
rect 194409 227563 194475 227566
rect 210693 227626 210759 227629
rect 260005 227626 260071 227629
rect 210693 227624 260071 227626
rect 210693 227568 210698 227624
rect 210754 227568 260010 227624
rect 260066 227568 260071 227624
rect 210693 227566 260071 227568
rect 210693 227563 210759 227566
rect 260005 227563 260071 227566
rect 411161 227626 411227 227629
rect 569309 227626 569375 227629
rect 411161 227624 569375 227626
rect 411161 227568 411166 227624
rect 411222 227568 569314 227624
rect 569370 227568 569375 227624
rect 411161 227566 569375 227568
rect 411161 227563 411227 227566
rect 569309 227563 569375 227566
rect 94773 227490 94839 227493
rect 210417 227490 210483 227493
rect 94773 227488 210483 227490
rect 94773 227432 94778 227488
rect 94834 227432 210422 227488
rect 210478 227432 210483 227488
rect 94773 227430 210483 227432
rect 94773 227427 94839 227430
rect 210417 227427 210483 227430
rect 380157 227490 380223 227493
rect 496169 227490 496235 227493
rect 380157 227488 496235 227490
rect 380157 227432 380162 227488
rect 380218 227432 496174 227488
rect 496230 227432 496235 227488
rect 380157 227430 496235 227432
rect 380157 227427 380223 227430
rect 496169 227427 496235 227430
rect 99833 227354 99899 227357
rect 212901 227354 212967 227357
rect 99833 227352 212967 227354
rect 99833 227296 99838 227352
rect 99894 227296 212906 227352
rect 212962 227296 212967 227352
rect 99833 227294 212967 227296
rect 99833 227291 99899 227294
rect 212901 227291 212967 227294
rect 376937 227354 377003 227357
rect 488901 227354 488967 227357
rect 376937 227352 488967 227354
rect 376937 227296 376942 227352
rect 376998 227296 488906 227352
rect 488962 227296 488967 227352
rect 376937 227294 488967 227296
rect 376937 227291 377003 227294
rect 488901 227291 488967 227294
rect 101489 227218 101555 227221
rect 213269 227218 213335 227221
rect 101489 227216 213335 227218
rect 101489 227160 101494 227216
rect 101550 227160 213274 227216
rect 213330 227160 213335 227216
rect 101489 227158 213335 227160
rect 101489 227155 101555 227158
rect 213269 227155 213335 227158
rect 377305 227218 377371 227221
rect 488441 227218 488507 227221
rect 377305 227216 488507 227218
rect 377305 227160 377310 227216
rect 377366 227160 488446 227216
rect 488502 227160 488507 227216
rect 377305 227158 488507 227160
rect 377305 227155 377371 227158
rect 488441 227155 488507 227158
rect 106549 227082 106615 227085
rect 215753 227082 215819 227085
rect 106549 227080 215819 227082
rect 106549 227024 106554 227080
rect 106610 227024 215758 227080
rect 215814 227024 215819 227080
rect 106549 227022 215819 227024
rect 106549 227019 106615 227022
rect 215753 227019 215819 227022
rect 382641 227082 382707 227085
rect 480253 227082 480319 227085
rect 382641 227080 480319 227082
rect 382641 227024 382646 227080
rect 382702 227024 480258 227080
rect 480314 227024 480319 227080
rect 382641 227022 480319 227024
rect 382641 227019 382707 227022
rect 480253 227019 480319 227022
rect 113081 226946 113147 226949
rect 218605 226946 218671 226949
rect 113081 226944 218671 226946
rect 113081 226888 113086 226944
rect 113142 226888 218610 226944
rect 218666 226888 218671 226944
rect 113081 226886 218671 226888
rect 113081 226883 113147 226886
rect 218605 226883 218671 226886
rect 114921 226810 114987 226813
rect 218973 226810 219039 226813
rect 114921 226808 219039 226810
rect 114921 226752 114926 226808
rect 114982 226752 218978 226808
rect 219034 226752 219039 226808
rect 114921 226750 219039 226752
rect 114921 226747 114987 226750
rect 218973 226747 219039 226750
rect 98913 226266 98979 226269
rect 211153 226266 211219 226269
rect 98913 226264 211219 226266
rect 98913 226208 98918 226264
rect 98974 226208 211158 226264
rect 211214 226208 211219 226264
rect 98913 226206 211219 226208
rect 98913 226203 98979 226206
rect 211153 226203 211219 226206
rect 373717 226266 373783 226269
rect 481909 226266 481975 226269
rect 373717 226264 481975 226266
rect 373717 226208 373722 226264
rect 373778 226208 481914 226264
rect 481970 226208 481975 226264
rect 373717 226206 481975 226208
rect 373717 226203 373783 226206
rect 481909 226203 481975 226206
rect 97257 226130 97323 226133
rect 210785 226130 210851 226133
rect 97257 226128 210851 226130
rect 97257 226072 97262 226128
rect 97318 226072 210790 226128
rect 210846 226072 210851 226128
rect 97257 226070 210851 226072
rect 97257 226067 97323 226070
rect 210785 226067 210851 226070
rect 411161 226130 411227 226133
rect 518617 226130 518683 226133
rect 411161 226128 518683 226130
rect 411161 226072 411166 226128
rect 411222 226072 518622 226128
rect 518678 226072 518683 226128
rect 411161 226070 518683 226072
rect 411161 226067 411227 226070
rect 518617 226067 518683 226070
rect 92197 225994 92263 225997
rect 208301 225994 208367 225997
rect 92197 225992 208367 225994
rect 92197 225936 92202 225992
rect 92258 225936 208306 225992
rect 208362 225936 208367 225992
rect 92197 225934 208367 225936
rect 92197 225931 92263 225934
rect 208301 225931 208367 225934
rect 390461 225994 390527 225997
rect 520825 225994 520891 225997
rect 390461 225992 520891 225994
rect 390461 225936 390466 225992
rect 390522 225936 520830 225992
rect 520886 225936 520891 225992
rect 390461 225934 520891 225936
rect 390461 225931 390527 225934
rect 520825 225931 520891 225934
rect 83825 225858 83891 225861
rect 205081 225858 205147 225861
rect 83825 225856 205147 225858
rect 83825 225800 83830 225856
rect 83886 225800 205086 225856
rect 205142 225800 205147 225856
rect 83825 225798 205147 225800
rect 83825 225795 83891 225798
rect 205081 225795 205147 225798
rect 392577 225858 392643 225861
rect 525793 225858 525859 225861
rect 392577 225856 525859 225858
rect 392577 225800 392582 225856
rect 392638 225800 525798 225856
rect 525854 225800 525859 225856
rect 392577 225798 525859 225800
rect 392577 225795 392643 225798
rect 525793 225795 525859 225798
rect 42425 225722 42491 225725
rect 43662 225722 43668 225724
rect 42425 225720 43668 225722
rect 42425 225664 42430 225720
rect 42486 225664 43668 225720
rect 42425 225662 43668 225664
rect 42425 225659 42491 225662
rect 43662 225660 43668 225662
rect 43732 225660 43738 225724
rect 80421 225722 80487 225725
rect 203701 225722 203767 225725
rect 80421 225720 203767 225722
rect 80421 225664 80426 225720
rect 80482 225664 203706 225720
rect 203762 225664 203767 225720
rect 80421 225662 203767 225664
rect 80421 225659 80487 225662
rect 203701 225659 203767 225662
rect 391565 225722 391631 225725
rect 523401 225722 523467 225725
rect 391565 225720 523467 225722
rect 391565 225664 391570 225720
rect 391626 225664 523406 225720
rect 523462 225664 523467 225720
rect 391565 225662 523467 225664
rect 391565 225659 391631 225662
rect 523401 225659 523467 225662
rect 77109 225586 77175 225589
rect 202229 225586 202295 225589
rect 77109 225584 202295 225586
rect 77109 225528 77114 225584
rect 77170 225528 202234 225584
rect 202290 225528 202295 225584
rect 77109 225526 202295 225528
rect 77109 225523 77175 225526
rect 202229 225523 202295 225526
rect 393681 225586 393747 225589
rect 528093 225586 528159 225589
rect 393681 225584 528159 225586
rect 393681 225528 393686 225584
rect 393742 225528 528098 225584
rect 528154 225528 528159 225584
rect 393681 225526 528159 225528
rect 393681 225523 393747 225526
rect 528093 225523 528159 225526
rect 70393 225450 70459 225453
rect 199377 225450 199443 225453
rect 70393 225448 199443 225450
rect 70393 225392 70398 225448
rect 70454 225392 199382 225448
rect 199438 225392 199443 225448
rect 70393 225390 199443 225392
rect 70393 225387 70459 225390
rect 199377 225387 199443 225390
rect 394785 225450 394851 225453
rect 530669 225450 530735 225453
rect 394785 225448 530735 225450
rect 394785 225392 394790 225448
rect 394846 225392 530674 225448
rect 530730 225392 530735 225448
rect 394785 225390 530735 225392
rect 394785 225387 394851 225390
rect 530669 225387 530735 225390
rect 66989 225314 67055 225317
rect 197997 225314 198063 225317
rect 66989 225312 198063 225314
rect 66989 225256 66994 225312
rect 67050 225256 198002 225312
rect 198058 225256 198063 225312
rect 66989 225254 198063 225256
rect 66989 225251 67055 225254
rect 197997 225251 198063 225254
rect 397913 225314 397979 225317
rect 539317 225314 539383 225317
rect 397913 225312 539383 225314
rect 397913 225256 397918 225312
rect 397974 225256 539322 225312
rect 539378 225256 539383 225312
rect 397913 225254 539383 225256
rect 397913 225251 397979 225254
rect 539317 225251 539383 225254
rect 63401 225178 63467 225181
rect 196525 225178 196591 225181
rect 63401 225176 196591 225178
rect 63401 225120 63406 225176
rect 63462 225120 196530 225176
rect 196586 225120 196591 225176
rect 63401 225118 196591 225120
rect 63401 225115 63467 225118
rect 196525 225115 196591 225118
rect 401133 225178 401199 225181
rect 545757 225178 545823 225181
rect 401133 225176 545823 225178
rect 401133 225120 401138 225176
rect 401194 225120 545762 225176
rect 545818 225120 545823 225176
rect 401133 225118 545823 225120
rect 401133 225115 401199 225118
rect 545757 225115 545823 225118
rect 56869 225042 56935 225045
rect 193673 225042 193739 225045
rect 56869 225040 193739 225042
rect 56869 224984 56874 225040
rect 56930 224984 193678 225040
rect 193734 224984 193739 225040
rect 56869 224982 193739 224984
rect 56869 224979 56935 224982
rect 193673 224979 193739 224982
rect 407573 225042 407639 225045
rect 561213 225042 561279 225045
rect 407573 225040 561279 225042
rect 407573 224984 407578 225040
rect 407634 224984 561218 225040
rect 561274 224984 561279 225040
rect 407573 224982 561279 224984
rect 407573 224979 407639 224982
rect 561213 224979 561279 224982
rect 55121 224906 55187 224909
rect 192569 224906 192635 224909
rect 55121 224904 192635 224906
rect 55121 224848 55126 224904
rect 55182 224848 192574 224904
rect 192630 224848 192635 224904
rect 55121 224846 192635 224848
rect 55121 224843 55187 224846
rect 192569 224843 192635 224846
rect 410793 224906 410859 224909
rect 568573 224906 568639 224909
rect 410793 224904 568639 224906
rect 410793 224848 410798 224904
rect 410854 224848 568578 224904
rect 568634 224848 568639 224904
rect 410793 224846 568639 224848
rect 410793 224843 410859 224846
rect 568573 224843 568639 224846
rect 102041 224770 102107 224773
rect 212533 224770 212599 224773
rect 102041 224768 212599 224770
rect 102041 224712 102046 224768
rect 102102 224712 212538 224768
rect 212594 224712 212599 224768
rect 102041 224710 212599 224712
rect 102041 224707 102107 224710
rect 212533 224707 212599 224710
rect 372245 224770 372311 224773
rect 478505 224770 478571 224773
rect 372245 224768 478571 224770
rect 372245 224712 372250 224768
rect 372306 224712 478510 224768
rect 478566 224712 478571 224768
rect 372245 224710 478571 224712
rect 372245 224707 372311 224710
rect 478505 224707 478571 224710
rect 109033 224634 109099 224637
rect 215385 224634 215451 224637
rect 109033 224632 215451 224634
rect 109033 224576 109038 224632
rect 109094 224576 215390 224632
rect 215446 224576 215451 224632
rect 109033 224574 215451 224576
rect 109033 224571 109099 224574
rect 215385 224571 215451 224574
rect 369393 224634 369459 224637
rect 471973 224634 472039 224637
rect 369393 224632 472039 224634
rect 369393 224576 369398 224632
rect 369454 224576 471978 224632
rect 472034 224576 472039 224632
rect 369393 224574 472039 224576
rect 369393 224571 369459 224574
rect 471973 224571 472039 224574
rect 110689 224498 110755 224501
rect 216489 224498 216555 224501
rect 110689 224496 216555 224498
rect 110689 224440 110694 224496
rect 110750 224440 216494 224496
rect 216550 224440 216555 224496
rect 110689 224438 216555 224440
rect 110689 224435 110755 224438
rect 216489 224435 216555 224438
rect 370865 224498 370931 224501
rect 475101 224498 475167 224501
rect 370865 224496 475167 224498
rect 370865 224440 370870 224496
rect 370926 224440 475106 224496
rect 475162 224440 475167 224496
rect 370865 224438 475167 224440
rect 370865 224435 370931 224438
rect 475101 224435 475167 224438
rect 115749 224362 115815 224365
rect 218237 224362 218303 224365
rect 115749 224360 218303 224362
rect 115749 224304 115754 224360
rect 115810 224304 218242 224360
rect 218298 224304 218303 224360
rect 115749 224302 218303 224304
rect 115749 224299 115815 224302
rect 218237 224299 218303 224302
rect 372613 224362 372679 224365
rect 476021 224362 476087 224365
rect 372613 224360 476087 224362
rect 372613 224304 372618 224360
rect 372674 224304 476026 224360
rect 476082 224304 476087 224360
rect 372613 224302 476087 224304
rect 372613 224299 372679 224302
rect 476021 224299 476087 224302
rect 112437 224226 112503 224229
rect 216857 224226 216923 224229
rect 112437 224224 216923 224226
rect 112437 224168 112442 224224
rect 112498 224168 216862 224224
rect 216918 224168 216923 224224
rect 112437 224166 216923 224168
rect 112437 224163 112503 224166
rect 216857 224163 216923 224166
rect 120809 224090 120875 224093
rect 220813 224090 220879 224093
rect 120809 224088 220879 224090
rect 120809 224032 120814 224088
rect 120870 224032 220818 224088
rect 220874 224032 220879 224088
rect 120809 224030 220879 224032
rect 120809 224027 120875 224030
rect 220813 224027 220879 224030
rect 104801 223546 104867 223549
rect 214741 223546 214807 223549
rect 104801 223544 214807 223546
rect 104801 223488 104806 223544
rect 104862 223488 214746 223544
rect 214802 223488 214807 223544
rect 104801 223486 214807 223488
rect 104801 223483 104867 223486
rect 214741 223483 214807 223486
rect 222101 223546 222167 223549
rect 227805 223546 227871 223549
rect 222101 223544 227871 223546
rect 222101 223488 222106 223544
rect 222162 223488 227810 223544
rect 227866 223488 227871 223544
rect 222101 223486 227871 223488
rect 222101 223483 222167 223486
rect 227805 223483 227871 223486
rect 378317 223546 378383 223549
rect 491937 223546 492003 223549
rect 378317 223544 492003 223546
rect 378317 223488 378322 223544
rect 378378 223488 491942 223544
rect 491998 223488 492003 223544
rect 378317 223486 492003 223488
rect 378317 223483 378383 223486
rect 491937 223483 492003 223486
rect 675937 223546 676003 223549
rect 675937 223544 676292 223546
rect 675937 223488 675942 223544
rect 675998 223488 676292 223544
rect 675937 223486 676292 223488
rect 675937 223483 676003 223486
rect 98085 223410 98151 223413
rect 211889 223410 211955 223413
rect 98085 223408 211955 223410
rect 98085 223352 98090 223408
rect 98146 223352 211894 223408
rect 211950 223352 211955 223408
rect 98085 223350 211955 223352
rect 98085 223347 98151 223350
rect 211889 223347 211955 223350
rect 378685 223410 378751 223413
rect 492765 223410 492831 223413
rect 378685 223408 492831 223410
rect 378685 223352 378690 223408
rect 378746 223352 492770 223408
rect 492826 223352 492831 223408
rect 378685 223350 492831 223352
rect 378685 223347 378751 223350
rect 492765 223347 492831 223350
rect 96429 223274 96495 223277
rect 211521 223274 211587 223277
rect 96429 223272 211587 223274
rect 96429 223216 96434 223272
rect 96490 223216 211526 223272
rect 211582 223216 211587 223272
rect 96429 223214 211587 223216
rect 96429 223211 96495 223214
rect 211521 223211 211587 223214
rect 381169 223274 381235 223277
rect 499297 223274 499363 223277
rect 381169 223272 499363 223274
rect 381169 223216 381174 223272
rect 381230 223216 499302 223272
rect 499358 223216 499363 223272
rect 381169 223214 499363 223216
rect 381169 223211 381235 223214
rect 499297 223211 499363 223214
rect 89713 223138 89779 223141
rect 208669 223138 208735 223141
rect 89713 223136 208735 223138
rect 89713 223080 89718 223136
rect 89774 223080 208674 223136
rect 208730 223080 208735 223136
rect 89713 223078 208735 223080
rect 89713 223075 89779 223078
rect 208669 223075 208735 223078
rect 381537 223138 381603 223141
rect 500217 223138 500283 223141
rect 381537 223136 500283 223138
rect 381537 223080 381542 223136
rect 381598 223080 500222 223136
rect 500278 223080 500283 223136
rect 381537 223078 500283 223080
rect 381537 223075 381603 223078
rect 500217 223075 500283 223078
rect 675845 223138 675911 223141
rect 675845 223136 676292 223138
rect 675845 223080 675850 223136
rect 675906 223080 676292 223136
rect 675845 223078 676292 223080
rect 675845 223075 675911 223078
rect 81249 223002 81315 223005
rect 204713 223002 204779 223005
rect 81249 223000 204779 223002
rect 81249 222944 81254 223000
rect 81310 222944 204718 223000
rect 204774 222944 204779 223000
rect 81249 222942 204779 222944
rect 81249 222939 81315 222942
rect 204713 222939 204779 222942
rect 330937 223002 331003 223005
rect 381077 223002 381143 223005
rect 330937 223000 381143 223002
rect 330937 222944 330942 223000
rect 330998 222944 381082 223000
rect 381138 222944 381143 223000
rect 330937 222942 381143 222944
rect 330937 222939 331003 222942
rect 381077 222939 381143 222942
rect 383929 223002 383995 223005
rect 504817 223002 504883 223005
rect 383929 223000 504883 223002
rect 383929 222944 383934 223000
rect 383990 222944 504822 223000
rect 504878 222944 504883 223000
rect 383929 222942 504883 222944
rect 383929 222939 383995 222942
rect 504817 222939 504883 222942
rect 79593 222866 79659 222869
rect 204437 222866 204503 222869
rect 79593 222864 204503 222866
rect 79593 222808 79598 222864
rect 79654 222808 204442 222864
rect 204498 222808 204503 222864
rect 79593 222806 204503 222808
rect 79593 222803 79659 222806
rect 204437 222803 204503 222806
rect 333053 222866 333119 222869
rect 383653 222866 383719 222869
rect 333053 222864 383719 222866
rect 333053 222808 333058 222864
rect 333114 222808 383658 222864
rect 383714 222808 383719 222864
rect 333053 222806 383719 222808
rect 333053 222803 333119 222806
rect 383653 222803 383719 222806
rect 385861 222866 385927 222869
rect 509601 222866 509667 222869
rect 385861 222864 509667 222866
rect 385861 222808 385866 222864
rect 385922 222808 509606 222864
rect 509662 222808 509667 222864
rect 385861 222806 509667 222808
rect 385861 222803 385927 222806
rect 509601 222803 509667 222806
rect 74441 222730 74507 222733
rect 201861 222730 201927 222733
rect 74441 222728 201927 222730
rect 74441 222672 74446 222728
rect 74502 222672 201866 222728
rect 201922 222672 201927 222728
rect 74441 222670 201927 222672
rect 74441 222667 74507 222670
rect 201861 222667 201927 222670
rect 334525 222730 334591 222733
rect 386781 222730 386847 222733
rect 334525 222728 386847 222730
rect 334525 222672 334530 222728
rect 334586 222672 386786 222728
rect 386842 222672 386847 222728
rect 334525 222670 386847 222672
rect 334525 222667 334591 222670
rect 386781 222667 386847 222670
rect 387977 222730 388043 222733
rect 513373 222730 513439 222733
rect 387977 222728 513439 222730
rect 387977 222672 387982 222728
rect 388038 222672 513378 222728
rect 513434 222672 513439 222728
rect 387977 222670 513439 222672
rect 387977 222667 388043 222670
rect 513373 222667 513439 222670
rect 676029 222730 676095 222733
rect 676029 222728 676292 222730
rect 676029 222672 676034 222728
rect 676090 222672 676292 222728
rect 676029 222670 676292 222672
rect 676029 222667 676095 222670
rect 67817 222594 67883 222597
rect 198733 222594 198799 222597
rect 67817 222592 198799 222594
rect 67817 222536 67822 222592
rect 67878 222536 198738 222592
rect 198794 222536 198799 222592
rect 67817 222534 198799 222536
rect 67817 222531 67883 222534
rect 198733 222531 198799 222534
rect 332317 222594 332383 222597
rect 384297 222594 384363 222597
rect 332317 222592 384363 222594
rect 332317 222536 332322 222592
rect 332378 222536 384302 222592
rect 384358 222536 384363 222592
rect 332317 222534 384363 222536
rect 332317 222531 332383 222534
rect 384297 222531 384363 222534
rect 388989 222594 389055 222597
rect 517237 222594 517303 222597
rect 388989 222592 517303 222594
rect 388989 222536 388994 222592
rect 389050 222536 517242 222592
rect 517298 222536 517303 222592
rect 388989 222534 517303 222536
rect 388989 222531 389055 222534
rect 517237 222531 517303 222534
rect 66161 222458 66227 222461
rect 198641 222458 198707 222461
rect 66161 222456 198707 222458
rect 66161 222400 66166 222456
rect 66222 222400 198646 222456
rect 198702 222400 198707 222456
rect 66161 222398 198707 222400
rect 66161 222395 66227 222398
rect 198641 222395 198707 222398
rect 333789 222458 333855 222461
rect 387701 222458 387767 222461
rect 333789 222456 387767 222458
rect 333789 222400 333794 222456
rect 333850 222400 387706 222456
rect 387762 222400 387767 222456
rect 333789 222398 387767 222400
rect 333789 222395 333855 222398
rect 387701 222395 387767 222398
rect 391197 222458 391263 222461
rect 522205 222458 522271 222461
rect 391197 222456 522271 222458
rect 391197 222400 391202 222456
rect 391258 222400 522210 222456
rect 522266 222400 522271 222456
rect 391197 222398 522271 222400
rect 391197 222395 391263 222398
rect 522205 222395 522271 222398
rect 61101 222322 61167 222325
rect 196157 222322 196223 222325
rect 61101 222320 196223 222322
rect 61101 222264 61106 222320
rect 61162 222264 196162 222320
rect 196218 222264 196223 222320
rect 61101 222262 196223 222264
rect 61101 222259 61167 222262
rect 196157 222259 196223 222262
rect 335905 222322 335971 222325
rect 390185 222322 390251 222325
rect 335905 222320 390251 222322
rect 335905 222264 335910 222320
rect 335966 222264 390190 222320
rect 390246 222264 390251 222320
rect 335905 222262 390251 222264
rect 335905 222259 335971 222262
rect 390185 222259 390251 222262
rect 393313 222322 393379 222325
rect 527265 222322 527331 222325
rect 393313 222320 527331 222322
rect 393313 222264 393318 222320
rect 393374 222264 527270 222320
rect 527326 222264 527331 222320
rect 393313 222262 527331 222264
rect 393313 222259 393379 222262
rect 527265 222259 527331 222262
rect 675661 222322 675727 222325
rect 675661 222320 676292 222322
rect 675661 222264 675666 222320
rect 675722 222264 676292 222320
rect 675661 222262 676292 222264
rect 675661 222259 675727 222262
rect 54385 222186 54451 222189
rect 193305 222186 193371 222189
rect 54385 222184 193371 222186
rect 54385 222128 54390 222184
rect 54446 222128 193310 222184
rect 193366 222128 193371 222184
rect 54385 222126 193371 222128
rect 54385 222123 54451 222126
rect 193305 222123 193371 222126
rect 338757 222186 338823 222189
rect 396901 222186 396967 222189
rect 338757 222184 396967 222186
rect 338757 222128 338762 222184
rect 338818 222128 396906 222184
rect 396962 222128 396967 222184
rect 338757 222126 396967 222128
rect 338757 222123 338823 222126
rect 396901 222123 396967 222126
rect 397637 222186 397703 222189
rect 537385 222186 537451 222189
rect 397637 222184 537451 222186
rect 397637 222128 397642 222184
rect 397698 222128 537390 222184
rect 537446 222128 537451 222184
rect 397637 222126 537451 222128
rect 397637 222123 397703 222126
rect 537385 222123 537451 222126
rect 567285 222186 567351 222189
rect 574369 222186 574435 222189
rect 567285 222184 574435 222186
rect 567285 222128 567290 222184
rect 567346 222128 574374 222184
rect 574430 222128 574435 222184
rect 567285 222126 574435 222128
rect 567285 222123 567351 222126
rect 574369 222123 574435 222126
rect 103145 222050 103211 222053
rect 214373 222050 214439 222053
rect 103145 222048 214439 222050
rect 103145 221992 103150 222048
rect 103206 221992 214378 222048
rect 214434 221992 214439 222048
rect 103145 221990 214439 221992
rect 103145 221987 103211 221990
rect 214373 221987 214439 221990
rect 375833 222050 375899 222053
rect 486325 222050 486391 222053
rect 375833 222048 486391 222050
rect 375833 221992 375838 222048
rect 375894 221992 486330 222048
rect 486386 221992 486391 222048
rect 375833 221990 486391 221992
rect 375833 221987 375899 221990
rect 486325 221987 486391 221990
rect 109861 221914 109927 221917
rect 217225 221914 217291 221917
rect 109861 221912 217291 221914
rect 109861 221856 109866 221912
rect 109922 221856 217230 221912
rect 217286 221856 217291 221912
rect 109861 221854 217291 221856
rect 109861 221851 109927 221854
rect 217225 221851 217291 221854
rect 335813 221914 335879 221917
rect 388529 221914 388595 221917
rect 335813 221912 388595 221914
rect 335813 221856 335818 221912
rect 335874 221856 388534 221912
rect 388590 221856 388595 221912
rect 335813 221854 388595 221856
rect 335813 221851 335879 221854
rect 388529 221851 388595 221854
rect 391749 221914 391815 221917
rect 495617 221914 495683 221917
rect 675293 221914 675359 221917
rect 391749 221912 496830 221914
rect 391749 221856 391754 221912
rect 391810 221856 495622 221912
rect 495678 221856 496830 221912
rect 391749 221854 496830 221856
rect 391749 221851 391815 221854
rect 495617 221851 495683 221854
rect 111609 221778 111675 221781
rect 217317 221778 217383 221781
rect 111609 221776 217383 221778
rect 111609 221720 111614 221776
rect 111670 221720 217322 221776
rect 217378 221720 217383 221776
rect 111609 221718 217383 221720
rect 111609 221715 111675 221718
rect 217317 221715 217383 221718
rect 118325 221642 118391 221645
rect 220445 221642 220511 221645
rect 118325 221640 220511 221642
rect 118325 221584 118330 221640
rect 118386 221584 220450 221640
rect 220506 221584 220511 221640
rect 118325 221582 220511 221584
rect 118325 221579 118391 221582
rect 220445 221579 220511 221582
rect 121361 221506 121427 221509
rect 221825 221506 221891 221509
rect 121361 221504 221891 221506
rect 121361 221448 121366 221504
rect 121422 221448 221830 221504
rect 221886 221448 221891 221504
rect 121361 221446 221891 221448
rect 121361 221443 121427 221446
rect 221825 221443 221891 221446
rect 496770 221370 496830 221854
rect 675293 221912 676292 221914
rect 675293 221856 675298 221912
rect 675354 221856 676292 221912
rect 675293 221854 676292 221856
rect 675293 221851 675359 221854
rect 567101 221778 567167 221781
rect 575197 221778 575263 221781
rect 567101 221776 575263 221778
rect 567101 221720 567106 221776
rect 567162 221720 575202 221776
rect 575258 221720 575263 221776
rect 567101 221718 575263 221720
rect 567101 221715 567167 221718
rect 575197 221715 575263 221718
rect 564341 221506 564407 221509
rect 573541 221506 573607 221509
rect 564341 221504 573607 221506
rect 564341 221448 564346 221504
rect 564402 221448 573546 221504
rect 573602 221448 573607 221504
rect 564341 221446 573607 221448
rect 564341 221443 564407 221446
rect 573541 221443 573607 221446
rect 675753 221506 675819 221509
rect 675753 221504 676292 221506
rect 675753 221448 675758 221504
rect 675814 221448 676292 221504
rect 675753 221446 676292 221448
rect 675753 221443 675819 221446
rect 622485 221370 622551 221373
rect 496770 221368 622551 221370
rect 496770 221312 622490 221368
rect 622546 221312 622551 221368
rect 496770 221310 622551 221312
rect 622485 221307 622551 221310
rect 488901 221234 488967 221237
rect 621473 221234 621539 221237
rect 488901 221232 621539 221234
rect 488901 221176 488906 221232
rect 488962 221176 621478 221232
rect 621534 221176 621539 221232
rect 488901 221174 621539 221176
rect 488901 221171 488967 221174
rect 621473 221171 621539 221174
rect 500217 221098 500283 221101
rect 637849 221098 637915 221101
rect 500217 221096 637915 221098
rect 500217 221040 500222 221096
rect 500278 221040 637854 221096
rect 637910 221040 637915 221096
rect 500217 221038 637915 221040
rect 500217 221035 500283 221038
rect 637849 221035 637915 221038
rect 675753 221098 675819 221101
rect 675753 221096 676292 221098
rect 675753 221040 675758 221096
rect 675814 221040 676292 221096
rect 675753 221038 676292 221040
rect 675753 221035 675819 221038
rect 496169 220962 496235 220965
rect 637389 220962 637455 220965
rect 496169 220960 637455 220962
rect 496169 220904 496174 220960
rect 496230 220904 637394 220960
rect 637450 220904 637455 220960
rect 496169 220902 637455 220904
rect 496169 220899 496235 220902
rect 637389 220899 637455 220902
rect 675150 220628 675156 220692
rect 675220 220690 675226 220692
rect 675220 220630 676292 220690
rect 675220 220628 675226 220630
rect 675661 220282 675727 220285
rect 675661 220280 676292 220282
rect 675661 220224 675666 220280
rect 675722 220224 676292 220280
rect 675661 220222 676292 220224
rect 675661 220219 675727 220222
rect 676029 219874 676095 219877
rect 676029 219872 676292 219874
rect 676029 219816 676034 219872
rect 676090 219816 676292 219872
rect 676029 219814 676292 219816
rect 676029 219811 676095 219814
rect 675293 219466 675359 219469
rect 675293 219464 676292 219466
rect 675293 219408 675298 219464
rect 675354 219408 676292 219464
rect 675293 219406 676292 219408
rect 675293 219403 675359 219406
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 675385 218650 675451 218653
rect 675385 218648 676292 218650
rect 675385 218592 675390 218648
rect 675446 218592 676292 218648
rect 675385 218590 676292 218592
rect 675385 218587 675451 218590
rect 676029 218242 676095 218245
rect 676029 218240 676292 218242
rect 676029 218184 676034 218240
rect 676090 218184 676292 218240
rect 676029 218182 676292 218184
rect 676029 218179 676095 218182
rect 676029 217834 676095 217837
rect 676029 217832 676292 217834
rect 676029 217776 676034 217832
rect 676090 217776 676292 217832
rect 676029 217774 676292 217776
rect 676029 217771 676095 217774
rect 675477 217426 675543 217429
rect 675477 217424 676292 217426
rect 675477 217368 675482 217424
rect 675538 217368 676292 217424
rect 675477 217366 676292 217368
rect 675477 217363 675543 217366
rect 675937 217018 676003 217021
rect 675937 217016 676292 217018
rect 675937 216960 675942 217016
rect 675998 216960 676292 217016
rect 675937 216958 676292 216960
rect 675937 216955 676003 216958
rect 676029 216610 676095 216613
rect 676029 216608 676292 216610
rect 676029 216552 676034 216608
rect 676090 216552 676292 216608
rect 676029 216550 676292 216552
rect 676029 216547 676095 216550
rect 582281 216202 582347 216205
rect 576380 216200 582347 216202
rect 576380 216144 582286 216200
rect 582342 216144 582347 216200
rect 576380 216142 582347 216144
rect 582281 216139 582347 216142
rect 675937 216202 676003 216205
rect 675937 216200 676292 216202
rect 675937 216144 675942 216200
rect 675998 216144 676292 216200
rect 675937 216142 676292 216144
rect 675937 216139 676003 216142
rect 675845 215794 675911 215797
rect 675845 215792 676292 215794
rect 675845 215736 675850 215792
rect 675906 215736 676292 215792
rect 675845 215734 676292 215736
rect 675845 215731 675911 215734
rect 675569 215386 675635 215389
rect 675569 215384 676292 215386
rect 675569 215328 675574 215384
rect 675630 215328 676292 215384
rect 675569 215326 676292 215328
rect 675569 215323 675635 215326
rect 41505 215114 41571 215117
rect 41462 215112 41571 215114
rect 41462 215056 41510 215112
rect 41566 215056 41571 215112
rect 41462 215051 41571 215056
rect 41462 214948 41522 215051
rect 676029 214978 676095 214981
rect 676029 214976 676292 214978
rect 676029 214920 676034 214976
rect 676090 214920 676292 214976
rect 676029 214918 676292 214920
rect 676029 214915 676095 214918
rect 41505 214706 41571 214709
rect 580441 214706 580507 214709
rect 41462 214704 41571 214706
rect 41462 214648 41510 214704
rect 41566 214648 41571 214704
rect 41462 214643 41571 214648
rect 576380 214704 580507 214706
rect 576380 214648 580446 214704
rect 580502 214648 580507 214704
rect 576380 214646 580507 214648
rect 580441 214643 580507 214646
rect 41462 214540 41522 214643
rect 676029 214570 676095 214573
rect 676029 214568 676292 214570
rect 676029 214512 676034 214568
rect 676090 214512 676292 214568
rect 676029 214510 676292 214512
rect 676029 214507 676095 214510
rect 41505 214298 41571 214301
rect 41462 214296 41571 214298
rect 41462 214240 41510 214296
rect 41566 214240 41571 214296
rect 41462 214235 41571 214240
rect 41462 214132 41522 214235
rect 675937 214162 676003 214165
rect 675937 214160 676292 214162
rect 675937 214104 675942 214160
rect 675998 214104 676292 214160
rect 675937 214102 676292 214104
rect 675937 214099 676003 214102
rect 41505 213890 41571 213893
rect 41462 213888 41571 213890
rect 41462 213832 41510 213888
rect 41566 213832 41571 213888
rect 41462 213827 41571 213832
rect 41462 213724 41522 213827
rect 675937 213754 676003 213757
rect 675937 213752 676292 213754
rect 675937 213696 675942 213752
rect 675998 213696 676292 213752
rect 675937 213694 676292 213696
rect 675937 213691 676003 213694
rect 41505 213482 41571 213485
rect 41462 213480 41571 213482
rect 41462 213424 41510 213480
rect 41566 213424 41571 213480
rect 41462 213419 41571 213424
rect 41462 213316 41522 213419
rect 676078 213286 676292 213346
rect 580165 213210 580231 213213
rect 576380 213208 580231 213210
rect 576380 213152 580170 213208
rect 580226 213152 580231 213208
rect 576380 213150 580231 213152
rect 580165 213147 580231 213150
rect 39982 213012 39988 213076
rect 40052 213012 40058 213076
rect 39990 212908 40050 213012
rect 33041 212666 33107 212669
rect 32998 212664 33107 212666
rect 32998 212608 33046 212664
rect 33102 212608 33107 212664
rect 32998 212603 33107 212608
rect 32998 212500 33058 212603
rect 41505 212258 41571 212261
rect 41462 212256 41571 212258
rect 41462 212200 41510 212256
rect 41566 212200 41571 212256
rect 41462 212195 41571 212200
rect 41462 212092 41522 212195
rect 676078 212125 676138 213286
rect 679022 212500 679082 212908
rect 676029 212122 676138 212125
rect 675948 212120 676292 212122
rect 675948 212064 676034 212120
rect 676090 212064 676292 212120
rect 675948 212062 676292 212064
rect 676029 212059 676095 212062
rect 32949 211850 33015 211853
rect 32949 211848 33058 211850
rect 32949 211792 32954 211848
rect 33010 211792 33058 211848
rect 32949 211787 33058 211792
rect 32998 211684 33058 211787
rect 580073 211714 580139 211717
rect 576380 211712 580139 211714
rect 576380 211656 580078 211712
rect 580134 211656 580139 211712
rect 576380 211654 580139 211656
rect 580073 211651 580139 211654
rect 41505 211442 41571 211445
rect 41462 211440 41571 211442
rect 41462 211384 41510 211440
rect 41566 211384 41571 211440
rect 41462 211379 41571 211384
rect 41462 211276 41522 211379
rect 32857 211034 32923 211037
rect 32814 211032 32923 211034
rect 32814 210976 32862 211032
rect 32918 210976 32923 211032
rect 32814 210971 32923 210976
rect 32814 210868 32874 210971
rect 30054 210221 30114 210460
rect 30005 210216 30114 210221
rect 582281 210218 582347 210221
rect 30005 210160 30010 210216
rect 30066 210160 30114 210216
rect 30005 210158 30114 210160
rect 576380 210216 582347 210218
rect 576380 210160 582286 210216
rect 582342 210160 582347 210216
rect 576380 210158 582347 210160
rect 30005 210155 30071 210158
rect 582281 210155 582347 210158
rect 30238 209813 30298 210052
rect 30189 209808 30298 209813
rect 30189 209752 30194 209808
rect 30250 209752 30298 209808
rect 30189 209750 30298 209752
rect 30189 209747 30255 209750
rect 30054 209405 30114 209644
rect 599853 209538 599919 209541
rect 599853 209536 606556 209538
rect 599853 209480 599858 209536
rect 599914 209480 606556 209536
rect 599853 209478 606556 209480
rect 599853 209475 599919 209478
rect 30054 209400 30163 209405
rect 30054 209344 30102 209400
rect 30158 209344 30163 209400
rect 30054 209342 30163 209344
rect 30097 209339 30163 209342
rect 666553 209266 666619 209269
rect 666356 209264 666619 209266
rect 41462 208997 41522 209236
rect 666356 209208 666558 209264
rect 666614 209208 666619 209264
rect 666356 209206 666619 209208
rect 666553 209203 666619 209206
rect 41462 208992 41571 208997
rect 41462 208936 41510 208992
rect 41566 208936 41571 208992
rect 41462 208934 41571 208936
rect 41505 208931 41571 208934
rect 37966 208589 38026 208828
rect 579797 208722 579863 208725
rect 576380 208720 579863 208722
rect 576380 208664 579802 208720
rect 579858 208664 579863 208720
rect 576380 208662 579863 208664
rect 579797 208659 579863 208662
rect 37966 208584 38075 208589
rect 37966 208528 38014 208584
rect 38070 208528 38075 208584
rect 37966 208526 38075 208528
rect 38009 208523 38075 208526
rect 599945 208586 600011 208589
rect 599945 208584 606556 208586
rect 599945 208528 599950 208584
rect 600006 208528 606556 208584
rect 599945 208526 606556 208528
rect 599945 208523 600011 208526
rect 30238 208181 30298 208420
rect 30238 208176 30347 208181
rect 30238 208120 30286 208176
rect 30342 208120 30347 208176
rect 30238 208118 30347 208120
rect 30281 208115 30347 208118
rect 38150 207773 38210 208012
rect 38101 207768 38210 207773
rect 38101 207712 38106 207768
rect 38162 207712 38210 207768
rect 38101 207710 38210 207712
rect 38101 207707 38167 207710
rect 41462 207365 41522 207604
rect 598933 207498 598999 207501
rect 598933 207496 606556 207498
rect 598933 207440 598938 207496
rect 598994 207440 606556 207496
rect 598933 207438 606556 207440
rect 598933 207435 598999 207438
rect 41462 207360 41571 207365
rect 41462 207304 41510 207360
rect 41566 207304 41571 207360
rect 41462 207302 41571 207304
rect 41505 207299 41571 207302
rect 41781 207226 41847 207229
rect 582281 207226 582347 207229
rect 41492 207224 41847 207226
rect 41492 207168 41786 207224
rect 41842 207168 41847 207224
rect 41492 207166 41847 207168
rect 576380 207224 582347 207226
rect 576380 207168 582286 207224
rect 582342 207168 582347 207224
rect 576380 207166 582347 207168
rect 41781 207163 41847 207166
rect 582281 207163 582347 207166
rect 41462 206549 41522 206788
rect 41413 206544 41522 206549
rect 41413 206488 41418 206544
rect 41474 206488 41522 206544
rect 41413 206486 41522 206488
rect 601141 206546 601207 206549
rect 601141 206544 606556 206546
rect 601141 206488 601146 206544
rect 601202 206488 606556 206544
rect 601141 206486 606556 206488
rect 41413 206483 41479 206486
rect 601141 206483 601207 206486
rect 41462 206138 41522 206380
rect 41689 206138 41755 206141
rect 41462 206136 41755 206138
rect 41462 206080 41694 206136
rect 41750 206080 41755 206136
rect 41462 206078 41755 206080
rect 41689 206075 41755 206078
rect 41781 206002 41847 206005
rect 41492 206000 41847 206002
rect 41492 205944 41786 206000
rect 41842 205944 41847 206000
rect 41492 205942 41847 205944
rect 41781 205939 41847 205942
rect 666553 205866 666619 205869
rect 666356 205864 666619 205866
rect 666356 205808 666558 205864
rect 666614 205808 666619 205864
rect 666356 205806 666619 205808
rect 666553 205803 666619 205806
rect 581453 205730 581519 205733
rect 576380 205728 581519 205730
rect 576380 205672 581458 205728
rect 581514 205672 581519 205728
rect 576380 205670 581519 205672
rect 581453 205667 581519 205670
rect 41462 205322 41522 205564
rect 599117 205458 599183 205461
rect 599117 205456 606556 205458
rect 599117 205400 599122 205456
rect 599178 205400 606556 205456
rect 599117 205398 606556 205400
rect 599117 205395 599183 205398
rect 41597 205322 41663 205325
rect 41462 205320 41663 205322
rect 41462 205264 41602 205320
rect 41658 205264 41663 205320
rect 41462 205262 41663 205264
rect 41597 205259 41663 205262
rect 41462 204917 41522 205156
rect 25129 204914 25195 204917
rect 25086 204912 25195 204914
rect 25086 204856 25134 204912
rect 25190 204856 25195 204912
rect 25086 204851 25195 204856
rect 41462 204912 41571 204917
rect 41462 204856 41510 204912
rect 41566 204856 41571 204912
rect 41462 204854 41571 204856
rect 41505 204851 41571 204854
rect 25086 204748 25146 204851
rect 24945 204506 25011 204509
rect 24902 204504 25011 204506
rect 24902 204448 24950 204504
rect 25006 204448 25011 204504
rect 24902 204443 25011 204448
rect 600957 204506 601023 204509
rect 600957 204504 606556 204506
rect 600957 204448 600962 204504
rect 601018 204448 606556 204504
rect 600957 204446 606556 204448
rect 600957 204443 601023 204446
rect 24902 204340 24962 204443
rect 580625 204234 580691 204237
rect 666553 204234 666619 204237
rect 576380 204232 580691 204234
rect 576380 204176 580630 204232
rect 580686 204176 580691 204232
rect 576380 204174 580691 204176
rect 666356 204232 666619 204234
rect 666356 204176 666558 204232
rect 666614 204176 666619 204232
rect 666356 204174 666619 204176
rect 580625 204171 580691 204174
rect 666553 204171 666619 204174
rect 675017 203826 675083 203829
rect 674974 203824 675083 203826
rect 674974 203768 675022 203824
rect 675078 203768 675083 203824
rect 674974 203763 675083 203768
rect 24853 203690 24919 203693
rect 24853 203688 24962 203690
rect 24853 203632 24858 203688
rect 24914 203632 24962 203688
rect 24853 203627 24962 203632
rect 24902 203524 24962 203627
rect 674974 203557 675034 203763
rect 674974 203552 675083 203557
rect 674974 203496 675022 203552
rect 675078 203496 675083 203552
rect 674974 203494 675083 203496
rect 675017 203491 675083 203494
rect 601509 203418 601575 203421
rect 601509 203416 606556 203418
rect 601509 203360 601514 203416
rect 601570 203360 606556 203416
rect 601509 203358 606556 203360
rect 601509 203355 601575 203358
rect 582281 202738 582347 202741
rect 576380 202736 582347 202738
rect 576380 202680 582286 202736
rect 582342 202680 582347 202736
rect 576380 202678 582347 202680
rect 582281 202675 582347 202678
rect 599945 202466 600011 202469
rect 599945 202464 606556 202466
rect 599945 202408 599950 202464
rect 600006 202408 606556 202464
rect 599945 202406 606556 202408
rect 599945 202403 600011 202406
rect 38101 201378 38167 201381
rect 41454 201378 41460 201380
rect 38101 201376 41460 201378
rect 38101 201320 38106 201376
rect 38162 201320 41460 201376
rect 38101 201318 41460 201320
rect 38101 201315 38167 201318
rect 41454 201316 41460 201318
rect 41524 201316 41530 201380
rect 598933 201378 598999 201381
rect 598933 201376 606556 201378
rect 598933 201320 598938 201376
rect 598994 201320 606556 201376
rect 598933 201318 606556 201320
rect 598933 201315 598999 201318
rect 582281 201242 582347 201245
rect 576380 201240 582347 201242
rect 576380 201184 582286 201240
rect 582342 201184 582347 201240
rect 576380 201182 582347 201184
rect 582281 201179 582347 201182
rect 666553 200834 666619 200837
rect 666356 200832 666619 200834
rect 666356 200776 666558 200832
rect 666614 200776 666619 200832
rect 666356 200774 666619 200776
rect 666553 200771 666619 200774
rect 599945 200426 600011 200429
rect 599945 200424 606556 200426
rect 599945 200368 599950 200424
rect 600006 200368 606556 200424
rect 599945 200366 606556 200368
rect 599945 200363 600011 200366
rect 30097 200290 30163 200293
rect 41638 200290 41644 200292
rect 30097 200288 41644 200290
rect 30097 200232 30102 200288
rect 30158 200232 41644 200288
rect 30097 200230 41644 200232
rect 30097 200227 30163 200230
rect 41638 200228 41644 200230
rect 41708 200228 41714 200292
rect 30005 200154 30071 200157
rect 41822 200154 41828 200156
rect 30005 200152 41828 200154
rect 30005 200096 30010 200152
rect 30066 200096 41828 200152
rect 30005 200094 41828 200096
rect 30005 200091 30071 200094
rect 41822 200092 41828 200094
rect 41892 200092 41898 200156
rect 581085 199746 581151 199749
rect 576380 199744 581151 199746
rect 576380 199688 581090 199744
rect 581146 199688 581151 199744
rect 576380 199686 581151 199688
rect 581085 199683 581151 199686
rect 599945 199338 600011 199341
rect 599945 199336 606556 199338
rect 599945 199280 599950 199336
rect 600006 199280 606556 199336
rect 599945 199278 606556 199280
rect 599945 199275 600011 199278
rect 666553 199066 666619 199069
rect 666356 199064 666619 199066
rect 666356 199008 666558 199064
rect 666614 199008 666619 199064
rect 666356 199006 666619 199008
rect 666553 199003 666619 199006
rect 599117 198386 599183 198389
rect 599117 198384 606556 198386
rect 599117 198328 599122 198384
rect 599178 198328 606556 198384
rect 599117 198326 606556 198328
rect 599117 198323 599183 198326
rect 580717 198250 580783 198253
rect 576380 198248 580783 198250
rect 576380 198192 580722 198248
rect 580778 198192 580783 198248
rect 576380 198190 580783 198192
rect 580717 198187 580783 198190
rect 599301 197298 599367 197301
rect 599301 197296 606556 197298
rect 599301 197240 599306 197296
rect 599362 197240 606556 197296
rect 599301 197238 606556 197240
rect 599301 197235 599367 197238
rect 582281 196754 582347 196757
rect 576380 196752 582347 196754
rect 576380 196696 582286 196752
rect 582342 196696 582347 196752
rect 576380 196694 582347 196696
rect 582281 196691 582347 196694
rect 599945 196346 600011 196349
rect 599945 196344 606556 196346
rect 599945 196288 599950 196344
rect 600006 196288 606556 196344
rect 599945 196286 606556 196288
rect 599945 196283 600011 196286
rect 666553 195666 666619 195669
rect 666356 195664 666619 195666
rect 666356 195608 666558 195664
rect 666614 195608 666619 195664
rect 666356 195606 666619 195608
rect 666553 195603 666619 195606
rect 582281 195258 582347 195261
rect 576380 195256 582347 195258
rect 576380 195200 582286 195256
rect 582342 195200 582347 195256
rect 576380 195198 582347 195200
rect 582281 195195 582347 195198
rect 599945 195258 600011 195261
rect 599945 195256 606556 195258
rect 599945 195200 599950 195256
rect 600006 195200 606556 195256
rect 599945 195198 606556 195200
rect 599945 195195 600011 195198
rect 599117 194306 599183 194309
rect 599117 194304 606556 194306
rect 599117 194248 599122 194304
rect 599178 194248 606556 194304
rect 599117 194246 606556 194248
rect 599117 194243 599183 194246
rect 670693 194034 670759 194037
rect 666356 194032 670759 194034
rect 666356 193976 670698 194032
rect 670754 193976 670759 194032
rect 666356 193974 670759 193976
rect 670693 193971 670759 193974
rect 582189 193626 582255 193629
rect 576380 193624 582255 193626
rect 576380 193568 582194 193624
rect 582250 193568 582255 193624
rect 576380 193566 582255 193568
rect 582189 193563 582255 193566
rect 599945 193218 600011 193221
rect 599945 193216 606556 193218
rect 599945 193160 599950 193216
rect 600006 193160 606556 193216
rect 599945 193158 606556 193160
rect 599945 193155 600011 193158
rect 599117 192266 599183 192269
rect 599117 192264 606556 192266
rect 599117 192208 599122 192264
rect 599178 192208 606556 192264
rect 599117 192206 606556 192208
rect 599117 192203 599183 192206
rect 582281 192130 582347 192133
rect 576380 192128 582347 192130
rect 576380 192072 582286 192128
rect 582342 192072 582347 192128
rect 576380 192070 582347 192072
rect 582281 192067 582347 192070
rect 599853 191178 599919 191181
rect 599853 191176 606556 191178
rect 599853 191120 599858 191176
rect 599914 191120 606556 191176
rect 599853 191118 606556 191120
rect 599853 191115 599919 191118
rect 582189 190634 582255 190637
rect 670693 190634 670759 190637
rect 576380 190632 582255 190634
rect 576380 190576 582194 190632
rect 582250 190576 582255 190632
rect 576380 190574 582255 190576
rect 666356 190632 670759 190634
rect 666356 190576 670698 190632
rect 670754 190576 670759 190632
rect 666356 190574 670759 190576
rect 582189 190571 582255 190574
rect 670693 190571 670759 190574
rect 600957 190226 601023 190229
rect 600957 190224 606556 190226
rect 600957 190168 600962 190224
rect 601018 190168 606556 190224
rect 600957 190166 606556 190168
rect 600957 190163 601023 190166
rect 581361 189138 581427 189141
rect 576380 189136 581427 189138
rect 576380 189080 581366 189136
rect 581422 189080 581427 189136
rect 576380 189078 581427 189080
rect 581361 189075 581427 189078
rect 601601 189138 601667 189141
rect 601601 189136 606556 189138
rect 601601 189080 601606 189136
rect 601662 189080 606556 189136
rect 601601 189078 606556 189080
rect 601601 189075 601667 189078
rect 666553 189002 666619 189005
rect 666356 189000 666619 189002
rect 666356 188944 666558 189000
rect 666614 188944 666619 189000
rect 666356 188942 666619 188944
rect 666553 188939 666619 188942
rect 601509 188186 601575 188189
rect 601509 188184 606556 188186
rect 601509 188128 601514 188184
rect 601570 188128 606556 188184
rect 601509 188126 606556 188128
rect 601509 188123 601575 188126
rect 582281 187642 582347 187645
rect 576380 187640 582347 187642
rect 576380 187584 582286 187640
rect 582342 187584 582347 187640
rect 576380 187582 582347 187584
rect 582281 187579 582347 187582
rect 599945 187098 600011 187101
rect 599945 187096 606556 187098
rect 599945 187040 599950 187096
rect 600006 187040 606556 187096
rect 599945 187038 606556 187040
rect 599945 187035 600011 187038
rect 582189 186146 582255 186149
rect 576380 186144 582255 186146
rect 576380 186088 582194 186144
rect 582250 186088 582255 186144
rect 576380 186086 582255 186088
rect 582189 186083 582255 186086
rect 600037 186146 600103 186149
rect 600037 186144 606556 186146
rect 600037 186088 600042 186144
rect 600098 186088 606556 186144
rect 600037 186086 606556 186088
rect 600037 186083 600103 186086
rect 666553 185602 666619 185605
rect 666356 185600 666619 185602
rect 666356 185544 666558 185600
rect 666614 185544 666619 185600
rect 666356 185542 666619 185544
rect 666553 185539 666619 185542
rect 599853 185058 599919 185061
rect 599853 185056 606556 185058
rect 599853 185000 599858 185056
rect 599914 185000 606556 185056
rect 599853 184998 606556 185000
rect 599853 184995 599919 184998
rect 582281 184650 582347 184653
rect 576380 184648 582347 184650
rect 576380 184592 582286 184648
rect 582342 184592 582347 184648
rect 576380 184590 582347 184592
rect 582281 184587 582347 184590
rect 41873 184244 41939 184245
rect 41822 184242 41828 184244
rect 41782 184182 41828 184242
rect 41892 184240 41939 184244
rect 41934 184184 41939 184240
rect 41822 184180 41828 184182
rect 41892 184180 41939 184184
rect 41873 184179 41939 184180
rect 599761 184106 599827 184109
rect 599761 184104 606556 184106
rect 599761 184048 599766 184104
rect 599822 184048 606556 184104
rect 599761 184046 606556 184048
rect 599761 184043 599827 184046
rect 666553 183834 666619 183837
rect 666356 183832 666619 183834
rect 666356 183776 666558 183832
rect 666614 183776 666619 183832
rect 666356 183774 666619 183776
rect 666553 183771 666619 183774
rect 41454 183364 41460 183428
rect 41524 183426 41530 183428
rect 41781 183426 41847 183429
rect 41524 183424 41847 183426
rect 41524 183368 41786 183424
rect 41842 183368 41847 183424
rect 41524 183366 41847 183368
rect 41524 183364 41530 183366
rect 41781 183363 41847 183366
rect 579797 183154 579863 183157
rect 576380 183152 579863 183154
rect 576380 183096 579802 183152
rect 579858 183096 579863 183152
rect 576380 183094 579863 183096
rect 579797 183091 579863 183094
rect 41638 182956 41644 183020
rect 41708 183018 41714 183020
rect 41781 183018 41847 183021
rect 41708 183016 41847 183018
rect 41708 182960 41786 183016
rect 41842 182960 41847 183016
rect 41708 182958 41847 182960
rect 41708 182956 41714 182958
rect 41781 182955 41847 182958
rect 599945 183018 600011 183021
rect 599945 183016 606556 183018
rect 599945 182960 599950 183016
rect 600006 182960 606556 183016
rect 599945 182958 606556 182960
rect 599945 182955 600011 182958
rect 600129 182066 600195 182069
rect 600129 182064 606556 182066
rect 600129 182008 600134 182064
rect 600190 182008 606556 182064
rect 600129 182006 606556 182008
rect 600129 182003 600195 182006
rect 582281 181658 582347 181661
rect 576380 181656 582347 181658
rect 576380 181600 582286 181656
rect 582342 181600 582347 181656
rect 576380 181598 582347 181600
rect 582281 181595 582347 181598
rect 599853 180978 599919 180981
rect 599853 180976 606556 180978
rect 599853 180920 599858 180976
rect 599914 180920 606556 180976
rect 599853 180918 606556 180920
rect 599853 180915 599919 180918
rect 666553 180434 666619 180437
rect 666356 180432 666619 180434
rect 666356 180376 666558 180432
rect 666614 180376 666619 180432
rect 666356 180374 666619 180376
rect 666553 180371 666619 180374
rect 580165 180162 580231 180165
rect 576380 180160 580231 180162
rect 576380 180104 580170 180160
rect 580226 180104 580231 180160
rect 576380 180102 580231 180104
rect 580165 180099 580231 180102
rect 599669 180026 599735 180029
rect 599669 180024 606556 180026
rect 599669 179968 599674 180024
rect 599730 179968 606556 180024
rect 599669 179966 606556 179968
rect 599669 179963 599735 179966
rect 600037 178938 600103 178941
rect 600037 178936 606556 178938
rect 600037 178880 600042 178936
rect 600098 178880 606556 178936
rect 600037 178878 606556 178880
rect 600037 178875 600103 178878
rect 666553 178802 666619 178805
rect 671981 178802 672047 178805
rect 666356 178800 672047 178802
rect 666356 178744 666558 178800
rect 666614 178744 671986 178800
rect 672042 178744 672047 178800
rect 666356 178742 672047 178744
rect 666553 178739 666619 178742
rect 671981 178739 672047 178742
rect 676213 178802 676279 178805
rect 676213 178800 676322 178802
rect 676213 178744 676218 178800
rect 676274 178744 676322 178800
rect 676213 178739 676322 178744
rect 580533 178666 580599 178669
rect 576380 178664 580599 178666
rect 576380 178608 580538 178664
rect 580594 178608 580599 178664
rect 576380 178606 580599 178608
rect 580533 178603 580599 178606
rect 676262 178500 676322 178739
rect 675937 178122 676003 178125
rect 675937 178120 676292 178122
rect 675937 178064 675942 178120
rect 675998 178064 676292 178120
rect 675937 178062 676292 178064
rect 675937 178059 676003 178062
rect 599761 177986 599827 177989
rect 599761 177984 606556 177986
rect 599761 177928 599766 177984
rect 599822 177928 606556 177984
rect 599761 177926 606556 177928
rect 599761 177923 599827 177926
rect 675937 177714 676003 177717
rect 675937 177712 676292 177714
rect 675937 177656 675942 177712
rect 675998 177656 676292 177712
rect 675937 177654 676292 177656
rect 675937 177651 676003 177654
rect 676029 177306 676095 177309
rect 676029 177304 676292 177306
rect 676029 177248 676034 177304
rect 676090 177248 676292 177304
rect 676029 177246 676292 177248
rect 676029 177243 676095 177246
rect 580257 177170 580323 177173
rect 576380 177168 580323 177170
rect 576380 177112 580262 177168
rect 580318 177112 580323 177168
rect 576380 177110 580323 177112
rect 580257 177107 580323 177110
rect 598933 176898 598999 176901
rect 676029 176898 676095 176901
rect 598933 176896 606556 176898
rect 598933 176840 598938 176896
rect 598994 176840 606556 176896
rect 598933 176838 606556 176840
rect 676029 176896 676292 176898
rect 676029 176840 676034 176896
rect 676090 176840 676292 176896
rect 676029 176838 676292 176840
rect 598933 176835 598999 176838
rect 676029 176835 676095 176838
rect 676029 176490 676095 176493
rect 676029 176488 676292 176490
rect 676029 176432 676034 176488
rect 676090 176432 676292 176488
rect 676029 176430 676292 176432
rect 676029 176427 676095 176430
rect 675937 176082 676003 176085
rect 675937 176080 676292 176082
rect 675937 176024 675942 176080
rect 675998 176024 676292 176080
rect 675937 176022 676292 176024
rect 675937 176019 676003 176022
rect 600313 175946 600379 175949
rect 600313 175944 606556 175946
rect 600313 175888 600318 175944
rect 600374 175888 606556 175944
rect 600313 175886 606556 175888
rect 600313 175883 600379 175886
rect 580809 175674 580875 175677
rect 576380 175672 580875 175674
rect 576380 175616 580814 175672
rect 580870 175616 580875 175672
rect 576380 175614 580875 175616
rect 580809 175611 580875 175614
rect 675293 175674 675359 175677
rect 675293 175672 676292 175674
rect 675293 175616 675298 175672
rect 675354 175616 676292 175672
rect 675293 175614 676292 175616
rect 675293 175611 675359 175614
rect 666553 175402 666619 175405
rect 666356 175400 666619 175402
rect 666356 175344 666558 175400
rect 666614 175344 666619 175400
rect 666356 175342 666619 175344
rect 666553 175339 666619 175342
rect 675937 175266 676003 175269
rect 675937 175264 676292 175266
rect 675937 175208 675942 175264
rect 675998 175208 676292 175264
rect 675937 175206 676292 175208
rect 675937 175203 676003 175206
rect 599945 174858 600011 174861
rect 676029 174858 676095 174861
rect 599945 174856 606556 174858
rect 599945 174800 599950 174856
rect 600006 174800 606556 174856
rect 599945 174798 606556 174800
rect 676029 174856 676292 174858
rect 676029 174800 676034 174856
rect 676090 174800 676292 174856
rect 676029 174798 676292 174800
rect 599945 174795 600011 174798
rect 676029 174795 676095 174798
rect 676029 174450 676095 174453
rect 676029 174448 676292 174450
rect 676029 174392 676034 174448
rect 676090 174392 676292 174448
rect 676029 174390 676292 174392
rect 676029 174387 676095 174390
rect 580533 174178 580599 174181
rect 576380 174176 580599 174178
rect 576380 174120 580538 174176
rect 580594 174120 580599 174176
rect 576380 174118 580599 174120
rect 580533 174115 580599 174118
rect 676029 174042 676095 174045
rect 676029 174040 676292 174042
rect 676029 173984 676034 174040
rect 676090 173984 676292 174040
rect 676029 173982 676292 173984
rect 676029 173979 676095 173982
rect 600129 173906 600195 173909
rect 600129 173904 606556 173906
rect 600129 173848 600134 173904
rect 600190 173848 606556 173904
rect 600129 173846 606556 173848
rect 600129 173843 600195 173846
rect 666553 173634 666619 173637
rect 672073 173634 672139 173637
rect 666356 173632 672139 173634
rect 666356 173576 666558 173632
rect 666614 173576 672078 173632
rect 672134 173576 672139 173632
rect 666356 173574 672139 173576
rect 666553 173571 666619 173574
rect 672073 173571 672139 173574
rect 676029 173634 676095 173637
rect 676029 173632 676292 173634
rect 676029 173576 676034 173632
rect 676090 173576 676292 173632
rect 676029 173574 676292 173576
rect 676029 173571 676095 173574
rect 675293 173226 675359 173229
rect 675293 173224 676292 173226
rect 675293 173168 675298 173224
rect 675354 173168 676292 173224
rect 675293 173166 676292 173168
rect 675293 173163 675359 173166
rect 599853 172818 599919 172821
rect 676029 172818 676095 172821
rect 599853 172816 606556 172818
rect 599853 172760 599858 172816
rect 599914 172760 606556 172816
rect 599853 172758 606556 172760
rect 676029 172816 676292 172818
rect 676029 172760 676034 172816
rect 676090 172760 676292 172816
rect 676029 172758 676292 172760
rect 599853 172755 599919 172758
rect 676029 172755 676095 172758
rect 582281 172682 582347 172685
rect 576380 172680 582347 172682
rect 576380 172624 582286 172680
rect 582342 172624 582347 172680
rect 576380 172622 582347 172624
rect 582281 172619 582347 172622
rect 675937 172410 676003 172413
rect 675937 172408 676292 172410
rect 675937 172352 675942 172408
rect 675998 172352 676292 172408
rect 675937 172350 676292 172352
rect 675937 172347 676003 172350
rect 675937 172002 676003 172005
rect 675937 172000 676292 172002
rect 675937 171944 675942 172000
rect 675998 171944 676292 172000
rect 675937 171942 676292 171944
rect 675937 171939 676003 171942
rect 599945 171866 600011 171869
rect 599945 171864 606556 171866
rect 599945 171808 599950 171864
rect 600006 171808 606556 171864
rect 599945 171806 606556 171808
rect 599945 171803 600011 171806
rect 675937 171594 676003 171597
rect 675937 171592 676292 171594
rect 675937 171536 675942 171592
rect 675998 171536 676292 171592
rect 675937 171534 676292 171536
rect 675937 171531 676003 171534
rect 582189 171186 582255 171189
rect 576380 171184 582255 171186
rect 576380 171128 582194 171184
rect 582250 171128 582255 171184
rect 576380 171126 582255 171128
rect 582189 171123 582255 171126
rect 675886 171124 675892 171188
rect 675956 171186 675962 171188
rect 675956 171126 676292 171186
rect 675956 171124 675962 171126
rect 599945 170778 600011 170781
rect 676029 170778 676095 170781
rect 599945 170776 606556 170778
rect 599945 170720 599950 170776
rect 600006 170720 606556 170776
rect 599945 170718 606556 170720
rect 676029 170776 676292 170778
rect 676029 170720 676034 170776
rect 676090 170720 676292 170776
rect 676029 170718 676292 170720
rect 599945 170715 600011 170718
rect 676029 170715 676095 170718
rect 675937 170370 676003 170373
rect 675937 170368 676292 170370
rect 675937 170312 675942 170368
rect 675998 170312 676292 170368
rect 675937 170310 676292 170312
rect 675937 170307 676003 170310
rect 666553 170234 666619 170237
rect 666356 170232 666619 170234
rect 666356 170176 666558 170232
rect 666614 170176 666619 170232
rect 666356 170174 666619 170176
rect 666553 170171 666619 170174
rect 675845 169962 675911 169965
rect 675845 169960 676292 169962
rect 675845 169904 675850 169960
rect 675906 169904 676292 169960
rect 675845 169902 676292 169904
rect 675845 169899 675911 169902
rect 599853 169826 599919 169829
rect 599853 169824 606556 169826
rect 599853 169768 599858 169824
rect 599914 169768 606556 169824
rect 599853 169766 606556 169768
rect 599853 169763 599919 169766
rect 582281 169554 582347 169557
rect 576380 169552 582347 169554
rect 576380 169496 582286 169552
rect 582342 169496 582347 169552
rect 576380 169494 582347 169496
rect 582281 169491 582347 169494
rect 675937 169554 676003 169557
rect 675937 169552 676292 169554
rect 675937 169496 675942 169552
rect 675998 169496 676292 169552
rect 675937 169494 676292 169496
rect 675937 169491 676003 169494
rect 675845 169146 675911 169149
rect 675845 169144 676292 169146
rect 675845 169088 675850 169144
rect 675906 169088 676292 169144
rect 675845 169086 676292 169088
rect 675845 169083 675911 169086
rect 599025 168738 599091 168741
rect 675753 168738 675819 168741
rect 599025 168736 606556 168738
rect 599025 168680 599030 168736
rect 599086 168680 606556 168736
rect 599025 168678 606556 168680
rect 675753 168736 676292 168738
rect 675753 168680 675758 168736
rect 675814 168680 676292 168736
rect 675753 168678 676292 168680
rect 599025 168675 599091 168678
rect 675753 168675 675819 168678
rect 666737 168602 666803 168605
rect 672165 168602 672231 168605
rect 666356 168600 672231 168602
rect 666356 168544 666742 168600
rect 666798 168544 672170 168600
rect 672226 168544 672231 168600
rect 666356 168542 672231 168544
rect 666737 168539 666803 168542
rect 672165 168539 672231 168542
rect 670335 168342 670405 168347
rect 670335 168282 670340 168342
rect 670400 168282 676576 168342
rect 670335 168277 670405 168282
rect 581269 168058 581335 168061
rect 576380 168056 581335 168058
rect 576380 168000 581274 168056
rect 581330 168000 581335 168056
rect 576380 167998 581335 168000
rect 581269 167995 581335 167998
rect 670501 167932 670571 167937
rect 670501 167872 670506 167932
rect 670566 167872 676414 167932
rect 670501 167867 670571 167872
rect 599853 167786 599919 167789
rect 599853 167784 606556 167786
rect 599853 167728 599858 167784
rect 599914 167728 606556 167784
rect 599853 167726 606556 167728
rect 599853 167723 599919 167726
rect 676029 167106 676095 167109
rect 676029 167104 676292 167106
rect 676029 167048 676034 167104
rect 676090 167048 676292 167104
rect 676029 167046 676292 167048
rect 676029 167043 676095 167046
rect 600037 166698 600103 166701
rect 600037 166696 606556 166698
rect 600037 166640 600042 166696
rect 600098 166640 606556 166696
rect 600037 166638 606556 166640
rect 600037 166635 600103 166638
rect 581453 166562 581519 166565
rect 576380 166560 581519 166562
rect 576380 166504 581458 166560
rect 581514 166504 581519 166560
rect 576380 166502 581519 166504
rect 581453 166499 581519 166502
rect 599945 165746 600011 165749
rect 599945 165744 606556 165746
rect 599945 165688 599950 165744
rect 600006 165688 606556 165744
rect 599945 165686 606556 165688
rect 599945 165683 600011 165686
rect 666737 165202 666803 165205
rect 666356 165200 666803 165202
rect 666356 165144 666742 165200
rect 666798 165144 666803 165200
rect 666356 165142 666803 165144
rect 666737 165139 666803 165142
rect 580993 165066 581059 165069
rect 576380 165064 581059 165066
rect 576380 165008 580998 165064
rect 581054 165008 581059 165064
rect 576380 165006 581059 165008
rect 580993 165003 581059 165006
rect 599853 164658 599919 164661
rect 599853 164656 606556 164658
rect 599853 164600 599858 164656
rect 599914 164600 606556 164656
rect 599853 164598 606556 164600
rect 599853 164595 599919 164598
rect 599945 163706 600011 163709
rect 599945 163704 606556 163706
rect 599945 163648 599950 163704
rect 600006 163648 606556 163704
rect 599945 163646 606556 163648
rect 599945 163643 600011 163646
rect 580257 163570 580323 163573
rect 666737 163570 666803 163573
rect 672257 163570 672323 163573
rect 576380 163568 580323 163570
rect 576380 163512 580262 163568
rect 580318 163512 580323 163568
rect 576380 163510 580323 163512
rect 666356 163568 672323 163570
rect 666356 163512 666742 163568
rect 666798 163512 672262 163568
rect 672318 163512 672323 163568
rect 666356 163510 672323 163512
rect 580257 163507 580323 163510
rect 666737 163507 666803 163510
rect 672257 163507 672323 163510
rect 599853 162618 599919 162621
rect 599853 162616 606556 162618
rect 599853 162560 599858 162616
rect 599914 162560 606556 162616
rect 599853 162558 606556 162560
rect 599853 162555 599919 162558
rect 579889 162074 579955 162077
rect 576380 162072 579955 162074
rect 576380 162016 579894 162072
rect 579950 162016 579955 162072
rect 576380 162014 579955 162016
rect 579889 162011 579955 162014
rect 599945 161666 600011 161669
rect 599945 161664 606556 161666
rect 599945 161608 599950 161664
rect 600006 161608 606556 161664
rect 599945 161606 606556 161608
rect 599945 161603 600011 161606
rect 582005 160578 582071 160581
rect 576380 160576 582071 160578
rect 576380 160520 582010 160576
rect 582066 160520 582071 160576
rect 576380 160518 582071 160520
rect 582005 160515 582071 160518
rect 599301 160578 599367 160581
rect 599301 160576 606556 160578
rect 599301 160520 599306 160576
rect 599362 160520 606556 160576
rect 599301 160518 606556 160520
rect 599301 160515 599367 160518
rect 666737 160170 666803 160173
rect 666356 160168 666803 160170
rect 666356 160112 666742 160168
rect 666798 160112 666803 160168
rect 666356 160110 666803 160112
rect 666737 160107 666803 160110
rect 600037 159626 600103 159629
rect 600037 159624 606556 159626
rect 600037 159568 600042 159624
rect 600098 159568 606556 159624
rect 600037 159566 606556 159568
rect 600037 159563 600103 159566
rect 579797 159082 579863 159085
rect 576380 159080 579863 159082
rect 576380 159024 579802 159080
rect 579858 159024 579863 159080
rect 576380 159022 579863 159024
rect 579797 159019 579863 159022
rect 599945 158538 600011 158541
rect 599945 158536 606556 158538
rect 599945 158480 599950 158536
rect 600006 158480 606556 158536
rect 599945 158478 606556 158480
rect 599945 158475 600011 158478
rect 666737 158402 666803 158405
rect 672349 158402 672415 158405
rect 666356 158400 672415 158402
rect 666356 158344 666742 158400
rect 666798 158344 672354 158400
rect 672410 158344 672415 158400
rect 666356 158342 672415 158344
rect 666737 158339 666803 158342
rect 672349 158339 672415 158342
rect 579705 157586 579771 157589
rect 576380 157584 579771 157586
rect 576380 157528 579710 157584
rect 579766 157528 579771 157584
rect 576380 157526 579771 157528
rect 579705 157523 579771 157526
rect 599853 157586 599919 157589
rect 599853 157584 606556 157586
rect 599853 157528 599858 157584
rect 599914 157528 606556 157584
rect 599853 157526 606556 157528
rect 599853 157523 599919 157526
rect 675753 157042 675819 157045
rect 675886 157042 675892 157044
rect 675753 157040 675892 157042
rect 675753 156984 675758 157040
rect 675814 156984 675892 157040
rect 675753 156982 675892 156984
rect 675753 156979 675819 156982
rect 675886 156980 675892 156982
rect 675956 156980 675962 157044
rect 599853 156498 599919 156501
rect 599853 156496 606556 156498
rect 599853 156440 599858 156496
rect 599914 156440 606556 156496
rect 599853 156438 606556 156440
rect 599853 156435 599919 156438
rect 581729 156090 581795 156093
rect 576380 156088 581795 156090
rect 576380 156032 581734 156088
rect 581790 156032 581795 156088
rect 576380 156030 581795 156032
rect 581729 156027 581795 156030
rect 599945 155546 600011 155549
rect 599945 155544 606556 155546
rect 599945 155488 599950 155544
rect 600006 155488 606556 155544
rect 599945 155486 606556 155488
rect 599945 155483 600011 155486
rect 666737 155002 666803 155005
rect 666356 155000 666803 155002
rect 666356 154944 666742 155000
rect 666798 154944 666803 155000
rect 666356 154942 666803 154944
rect 666737 154939 666803 154942
rect 582281 154594 582347 154597
rect 576380 154592 582347 154594
rect 576380 154536 582286 154592
rect 582342 154536 582347 154592
rect 576380 154534 582347 154536
rect 582281 154531 582347 154534
rect 599853 154458 599919 154461
rect 599853 154456 606556 154458
rect 599853 154400 599858 154456
rect 599914 154400 606556 154456
rect 599853 154398 606556 154400
rect 599853 154395 599919 154398
rect 599945 153506 600011 153509
rect 599945 153504 606556 153506
rect 599945 153448 599950 153504
rect 600006 153448 606556 153504
rect 599945 153446 606556 153448
rect 599945 153443 600011 153446
rect 666737 153370 666803 153373
rect 672441 153370 672507 153373
rect 666356 153368 672507 153370
rect 666356 153312 666742 153368
rect 666798 153312 672446 153368
rect 672502 153312 672507 153368
rect 666356 153310 672507 153312
rect 666737 153307 666803 153310
rect 672441 153307 672507 153310
rect 581913 153098 581979 153101
rect 576380 153096 581979 153098
rect 576380 153040 581918 153096
rect 581974 153040 581979 153096
rect 576380 153038 581979 153040
rect 581913 153035 581979 153038
rect 599301 152418 599367 152421
rect 599301 152416 606556 152418
rect 599301 152360 599306 152416
rect 599362 152360 606556 152416
rect 599301 152358 606556 152360
rect 599301 152355 599367 152358
rect 581821 151602 581887 151605
rect 576380 151600 581887 151602
rect 576380 151544 581826 151600
rect 581882 151544 581887 151600
rect 576380 151542 581887 151544
rect 581821 151539 581887 151542
rect 598933 151466 598999 151469
rect 598933 151464 606556 151466
rect 598933 151408 598938 151464
rect 598994 151408 606556 151464
rect 598933 151406 606556 151408
rect 598933 151403 598999 151406
rect 599761 150378 599827 150381
rect 599761 150376 606556 150378
rect 599761 150320 599766 150376
rect 599822 150320 606556 150376
rect 599761 150318 606556 150320
rect 599761 150315 599827 150318
rect 582097 150106 582163 150109
rect 576380 150104 582163 150106
rect 576380 150048 582102 150104
rect 582158 150048 582163 150104
rect 576380 150046 582163 150048
rect 582097 150043 582163 150046
rect 666737 149970 666803 149973
rect 666356 149968 666803 149970
rect 666356 149912 666742 149968
rect 666798 149912 666803 149968
rect 666356 149910 666803 149912
rect 666737 149907 666803 149910
rect 599945 149426 600011 149429
rect 599945 149424 606556 149426
rect 599945 149368 599950 149424
rect 600006 149368 606556 149424
rect 599945 149366 606556 149368
rect 599945 149363 600011 149366
rect 581453 148610 581519 148613
rect 576380 148608 581519 148610
rect 576380 148552 581458 148608
rect 581514 148552 581519 148608
rect 576380 148550 581519 148552
rect 581453 148547 581519 148550
rect 599853 148338 599919 148341
rect 599853 148336 606556 148338
rect 599853 148280 599858 148336
rect 599914 148280 606556 148336
rect 599853 148278 606556 148280
rect 599853 148275 599919 148278
rect 666737 148202 666803 148205
rect 672533 148202 672599 148205
rect 666356 148200 672599 148202
rect 666356 148144 666742 148200
rect 666798 148144 672538 148200
rect 672594 148144 672599 148200
rect 666356 148142 672599 148144
rect 666737 148139 666803 148142
rect 672533 148139 672599 148142
rect 599945 147386 600011 147389
rect 599945 147384 606556 147386
rect 599945 147328 599950 147384
rect 600006 147328 606556 147384
rect 599945 147326 606556 147328
rect 599945 147323 600011 147326
rect 580901 146978 580967 146981
rect 576380 146976 580967 146978
rect 576380 146920 580906 146976
rect 580962 146920 580967 146976
rect 576380 146918 580967 146920
rect 580901 146915 580967 146918
rect 600037 146298 600103 146301
rect 600037 146296 606556 146298
rect 600037 146240 600042 146296
rect 600098 146240 606556 146296
rect 600037 146238 606556 146240
rect 600037 146235 600103 146238
rect 581269 145482 581335 145485
rect 576380 145480 581335 145482
rect 576380 145424 581274 145480
rect 581330 145424 581335 145480
rect 576380 145422 581335 145424
rect 581269 145419 581335 145422
rect 599853 145346 599919 145349
rect 599853 145344 606556 145346
rect 599853 145288 599858 145344
rect 599914 145288 606556 145344
rect 599853 145286 606556 145288
rect 599853 145283 599919 145286
rect 666737 144938 666803 144941
rect 666356 144936 666803 144938
rect 666356 144880 666742 144936
rect 666798 144880 666803 144936
rect 666356 144878 666803 144880
rect 666737 144875 666803 144878
rect 599945 144258 600011 144261
rect 599945 144256 606556 144258
rect 599945 144200 599950 144256
rect 600006 144200 606556 144256
rect 599945 144198 606556 144200
rect 599945 144195 600011 144198
rect 580993 143986 581059 143989
rect 576380 143984 581059 143986
rect 576380 143928 580998 143984
rect 581054 143928 581059 143984
rect 576380 143926 581059 143928
rect 580993 143923 581059 143926
rect 599853 143306 599919 143309
rect 599853 143304 606556 143306
rect 599853 143248 599858 143304
rect 599914 143248 606556 143304
rect 599853 143246 606556 143248
rect 599853 143243 599919 143246
rect 666737 143170 666803 143173
rect 672625 143170 672691 143173
rect 666356 143168 672691 143170
rect 666356 143112 666742 143168
rect 666798 143112 672630 143168
rect 672686 143112 672691 143168
rect 666356 143110 672691 143112
rect 666737 143107 666803 143110
rect 672625 143107 672691 143110
rect 581545 142490 581611 142493
rect 576380 142488 581611 142490
rect 576380 142432 581550 142488
rect 581606 142432 581611 142488
rect 576380 142430 581611 142432
rect 581545 142427 581611 142430
rect 599945 142218 600011 142221
rect 599945 142216 606556 142218
rect 599945 142160 599950 142216
rect 600006 142160 606556 142216
rect 599945 142158 606556 142160
rect 599945 142155 600011 142158
rect 599301 141266 599367 141269
rect 599301 141264 606556 141266
rect 599301 141208 599306 141264
rect 599362 141208 606556 141264
rect 599301 141206 606556 141208
rect 599301 141203 599367 141206
rect 581085 140994 581151 140997
rect 576380 140992 581151 140994
rect 576380 140936 581090 140992
rect 581146 140936 581151 140992
rect 576380 140934 581151 140936
rect 581085 140931 581151 140934
rect 599853 140178 599919 140181
rect 599853 140176 606556 140178
rect 599853 140120 599858 140176
rect 599914 140120 606556 140176
rect 599853 140118 606556 140120
rect 599853 140115 599919 140118
rect 666737 139770 666803 139773
rect 666356 139768 666803 139770
rect 666356 139712 666742 139768
rect 666798 139712 666803 139768
rect 666356 139710 666803 139712
rect 666737 139707 666803 139710
rect 581361 139498 581427 139501
rect 576380 139496 581427 139498
rect 576380 139440 581366 139496
rect 581422 139440 581427 139496
rect 576380 139438 581427 139440
rect 581361 139435 581427 139438
rect 600037 139226 600103 139229
rect 600037 139224 606556 139226
rect 600037 139168 600042 139224
rect 600098 139168 606556 139224
rect 600037 139166 606556 139168
rect 600037 139163 600103 139166
rect 672717 138410 672783 138413
rect 670650 138408 672783 138410
rect 670650 138352 672722 138408
rect 672778 138352 672783 138408
rect 670650 138350 672783 138352
rect 670650 138141 670710 138350
rect 672717 138347 672783 138350
rect 599945 138138 600011 138141
rect 670650 138138 670759 138141
rect 599945 138136 606556 138138
rect 599945 138080 599950 138136
rect 600006 138080 606556 138136
rect 599945 138078 606556 138080
rect 666356 138136 670759 138138
rect 666356 138080 670698 138136
rect 670754 138080 670759 138136
rect 666356 138078 670759 138080
rect 599945 138075 600011 138078
rect 670693 138075 670759 138078
rect 580441 138002 580507 138005
rect 576380 138000 580507 138002
rect 576380 137944 580446 138000
rect 580502 137944 580507 138000
rect 576380 137942 580507 137944
rect 580441 137939 580507 137942
rect 599853 137186 599919 137189
rect 599853 137184 606556 137186
rect 599853 137128 599858 137184
rect 599914 137128 606556 137184
rect 599853 137126 606556 137128
rect 599853 137123 599919 137126
rect 580717 136506 580783 136509
rect 576380 136504 580783 136506
rect 576380 136448 580722 136504
rect 580778 136448 580783 136504
rect 576380 136446 580783 136448
rect 580717 136443 580783 136446
rect 599945 136098 600011 136101
rect 599945 136096 606556 136098
rect 599945 136040 599950 136096
rect 600006 136040 606556 136096
rect 599945 136038 606556 136040
rect 599945 136035 600011 136038
rect 600037 135146 600103 135149
rect 600037 135144 606556 135146
rect 600037 135088 600042 135144
rect 600098 135088 606556 135144
rect 600037 135086 606556 135088
rect 600037 135083 600103 135086
rect 581177 135010 581243 135013
rect 576380 135008 581243 135010
rect 576380 134952 581182 135008
rect 581238 134952 581243 135008
rect 576380 134950 581243 134952
rect 581177 134947 581243 134950
rect 670693 134738 670759 134741
rect 666356 134736 670759 134738
rect 666356 134680 670698 134736
rect 670754 134680 670759 134736
rect 666356 134678 670759 134680
rect 670693 134675 670759 134678
rect 599853 134058 599919 134061
rect 599853 134056 606556 134058
rect 599853 134000 599858 134056
rect 599914 134000 606556 134056
rect 599853 133998 606556 134000
rect 599853 133995 599919 133998
rect 580625 133514 580691 133517
rect 576380 133512 580691 133514
rect 576380 133456 580630 133512
rect 580686 133456 580691 133512
rect 576380 133454 580691 133456
rect 580625 133451 580691 133454
rect 599945 133106 600011 133109
rect 676121 133106 676187 133109
rect 676262 133106 676322 133348
rect 599945 133104 606556 133106
rect 599945 133048 599950 133104
rect 600006 133048 606556 133104
rect 599945 133046 606556 133048
rect 676121 133104 676322 133106
rect 676121 133048 676126 133104
rect 676182 133048 676322 133104
rect 676121 133046 676322 133048
rect 599945 133043 600011 133046
rect 676121 133043 676187 133046
rect 666737 132970 666803 132973
rect 672809 132970 672875 132973
rect 666356 132968 672875 132970
rect 666356 132912 666742 132968
rect 666798 132912 672814 132968
rect 672870 132912 672875 132968
rect 666356 132910 672875 132912
rect 666737 132907 666803 132910
rect 672809 132907 672875 132910
rect 676029 132970 676095 132973
rect 676029 132968 676292 132970
rect 676029 132912 676034 132968
rect 676090 132912 676292 132968
rect 676029 132910 676292 132912
rect 676029 132907 676095 132910
rect 676213 132698 676279 132701
rect 676213 132696 676322 132698
rect 676213 132640 676218 132696
rect 676274 132640 676322 132696
rect 676213 132635 676322 132640
rect 676262 132532 676322 132635
rect 676213 132290 676279 132293
rect 676213 132288 676322 132290
rect 676213 132232 676218 132288
rect 676274 132232 676322 132288
rect 676213 132227 676322 132232
rect 676262 132124 676322 132227
rect 580809 132018 580875 132021
rect 576380 132016 580875 132018
rect 576380 131960 580814 132016
rect 580870 131960 580875 132016
rect 576380 131958 580875 131960
rect 580809 131955 580875 131958
rect 598933 132018 598999 132021
rect 598933 132016 606556 132018
rect 598933 131960 598938 132016
rect 598994 131960 606556 132016
rect 598933 131958 606556 131960
rect 598933 131955 598999 131958
rect 676029 131746 676095 131749
rect 676029 131744 676292 131746
rect 676029 131688 676034 131744
rect 676090 131688 676292 131744
rect 676029 131686 676292 131688
rect 676029 131683 676095 131686
rect 676213 131474 676279 131477
rect 676213 131472 676322 131474
rect 676213 131416 676218 131472
rect 676274 131416 676322 131472
rect 676213 131411 676322 131416
rect 676262 131308 676322 131411
rect 599761 131066 599827 131069
rect 599761 131064 606556 131066
rect 599761 131008 599766 131064
rect 599822 131008 606556 131064
rect 599761 131006 606556 131008
rect 599761 131003 599827 131006
rect 676029 130930 676095 130933
rect 676029 130928 676292 130930
rect 676029 130872 676034 130928
rect 676090 130872 676292 130928
rect 676029 130870 676292 130872
rect 676029 130867 676095 130870
rect 676213 130658 676279 130661
rect 676213 130656 676322 130658
rect 676213 130600 676218 130656
rect 676274 130600 676322 130656
rect 676213 130595 676322 130600
rect 582189 130522 582255 130525
rect 576380 130520 582255 130522
rect 576380 130464 582194 130520
rect 582250 130464 582255 130520
rect 676262 130492 676322 130595
rect 576380 130462 582255 130464
rect 582189 130459 582255 130462
rect 676029 130114 676095 130117
rect 676029 130112 676292 130114
rect 676029 130056 676034 130112
rect 676090 130056 676292 130112
rect 676029 130054 676292 130056
rect 676029 130051 676095 130054
rect 599945 129978 600011 129981
rect 599945 129976 606556 129978
rect 599945 129920 599950 129976
rect 600006 129920 606556 129976
rect 599945 129918 606556 129920
rect 599945 129915 600011 129918
rect 676029 129706 676095 129709
rect 676029 129704 676292 129706
rect 676029 129648 676034 129704
rect 676090 129648 676292 129704
rect 676029 129646 676292 129648
rect 676029 129643 676095 129646
rect 666737 129570 666803 129573
rect 666356 129568 666803 129570
rect 666356 129512 666742 129568
rect 666798 129512 666803 129568
rect 666356 129510 666803 129512
rect 666737 129507 666803 129510
rect 676213 129434 676279 129437
rect 676213 129432 676322 129434
rect 676213 129376 676218 129432
rect 676274 129376 676322 129432
rect 676213 129371 676322 129376
rect 676262 129268 676322 129371
rect 582281 129026 582347 129029
rect 576380 129024 582347 129026
rect 576380 128968 582286 129024
rect 582342 128968 582347 129024
rect 576380 128966 582347 128968
rect 582281 128963 582347 128966
rect 599853 129026 599919 129029
rect 599853 129024 606556 129026
rect 599853 128968 599858 129024
rect 599914 128968 606556 129024
rect 599853 128966 606556 128968
rect 599853 128963 599919 128966
rect 676029 128890 676095 128893
rect 676029 128888 676292 128890
rect 676029 128832 676034 128888
rect 676090 128832 676292 128888
rect 676029 128830 676292 128832
rect 676029 128827 676095 128830
rect 675937 128482 676003 128485
rect 675937 128480 676292 128482
rect 675937 128424 675942 128480
rect 675998 128424 676292 128480
rect 675937 128422 676292 128424
rect 675937 128419 676003 128422
rect 675569 128074 675635 128077
rect 675569 128072 676292 128074
rect 675569 128016 675574 128072
rect 675630 128016 676292 128072
rect 675569 128014 676292 128016
rect 675569 128011 675635 128014
rect 599945 127938 600011 127941
rect 666645 127938 666711 127941
rect 672901 127938 672967 127941
rect 599945 127936 606556 127938
rect 599945 127880 599950 127936
rect 600006 127880 606556 127936
rect 599945 127878 606556 127880
rect 666356 127936 672967 127938
rect 666356 127880 666650 127936
rect 666706 127880 672906 127936
rect 672962 127880 672967 127936
rect 666356 127878 672967 127880
rect 599945 127875 600011 127878
rect 666645 127875 666711 127878
rect 672901 127875 672967 127878
rect 676029 127666 676095 127669
rect 676029 127664 676292 127666
rect 676029 127608 676034 127664
rect 676090 127608 676292 127664
rect 676029 127606 676292 127608
rect 676029 127603 676095 127606
rect 580533 127530 580599 127533
rect 576380 127528 580599 127530
rect 576380 127472 580538 127528
rect 580594 127472 580599 127528
rect 576380 127470 580599 127472
rect 580533 127467 580599 127470
rect 675937 127258 676003 127261
rect 675937 127256 676292 127258
rect 675937 127200 675942 127256
rect 675998 127200 676292 127256
rect 675937 127198 676292 127200
rect 675937 127195 676003 127198
rect 600037 126986 600103 126989
rect 600037 126984 606556 126986
rect 600037 126928 600042 126984
rect 600098 126928 606556 126984
rect 600037 126926 606556 126928
rect 600037 126923 600103 126926
rect 676029 126850 676095 126853
rect 676029 126848 676292 126850
rect 676029 126792 676034 126848
rect 676090 126792 676292 126848
rect 676029 126790 676292 126792
rect 676029 126787 676095 126790
rect 675293 126442 675359 126445
rect 675293 126440 676292 126442
rect 675293 126384 675298 126440
rect 675354 126384 676292 126440
rect 675293 126382 676292 126384
rect 675293 126379 675359 126382
rect 581821 126034 581887 126037
rect 576380 126032 581887 126034
rect 576380 125976 581826 126032
rect 581882 125976 581887 126032
rect 576380 125974 581887 125976
rect 581821 125971 581887 125974
rect 676029 126034 676095 126037
rect 676029 126032 676292 126034
rect 676029 125976 676034 126032
rect 676090 125976 676292 126032
rect 676029 125974 676292 125976
rect 676029 125971 676095 125974
rect 599853 125898 599919 125901
rect 599853 125896 606556 125898
rect 599853 125840 599858 125896
rect 599914 125840 606556 125896
rect 599853 125838 606556 125840
rect 599853 125835 599919 125838
rect 675937 125626 676003 125629
rect 675937 125624 676292 125626
rect 675937 125568 675942 125624
rect 675998 125568 676292 125624
rect 675937 125566 676292 125568
rect 675937 125563 676003 125566
rect 599945 124946 600011 124949
rect 676121 124946 676187 124949
rect 676262 124946 676322 125188
rect 599945 124944 606556 124946
rect 599945 124888 599950 124944
rect 600006 124888 606556 124944
rect 599945 124886 606556 124888
rect 676121 124944 676322 124946
rect 676121 124888 676126 124944
rect 676182 124888 676322 124944
rect 676121 124886 676322 124888
rect 599945 124883 600011 124886
rect 676121 124883 676187 124886
rect 582005 124538 582071 124541
rect 666645 124538 666711 124541
rect 576380 124536 582071 124538
rect 576380 124480 582010 124536
rect 582066 124480 582071 124536
rect 576380 124478 582071 124480
rect 666356 124536 666711 124538
rect 666356 124480 666650 124536
rect 666706 124480 666711 124536
rect 666356 124478 666711 124480
rect 582005 124475 582071 124478
rect 666645 124475 666711 124478
rect 676121 124538 676187 124541
rect 676262 124538 676322 124780
rect 676121 124536 676322 124538
rect 676121 124480 676126 124536
rect 676182 124480 676322 124536
rect 676121 124478 676322 124480
rect 676121 124475 676187 124478
rect 676029 124402 676095 124405
rect 676029 124400 676292 124402
rect 676029 124344 676034 124400
rect 676090 124344 676292 124400
rect 676029 124342 676292 124344
rect 676029 124339 676095 124342
rect 676029 123994 676095 123997
rect 676029 123992 676292 123994
rect 676029 123936 676034 123992
rect 676090 123936 676292 123992
rect 676029 123934 676292 123936
rect 676029 123931 676095 123934
rect 599853 123858 599919 123861
rect 599853 123856 606556 123858
rect 599853 123800 599858 123856
rect 599914 123800 606556 123856
rect 599853 123798 606556 123800
rect 599853 123795 599919 123798
rect 676029 123586 676095 123589
rect 676029 123584 676292 123586
rect 676029 123528 676034 123584
rect 676090 123528 676292 123584
rect 676029 123526 676292 123528
rect 676029 123523 676095 123526
rect 673273 123132 673343 123137
rect 673273 123072 673278 123132
rect 673338 123072 676382 123132
rect 673273 123067 673343 123072
rect 581637 122906 581703 122909
rect 576380 122904 581703 122906
rect 576380 122848 581642 122904
rect 581698 122848 581703 122904
rect 576380 122846 581703 122848
rect 581637 122843 581703 122846
rect 599945 122906 600011 122909
rect 666645 122906 666711 122909
rect 672993 122906 673059 122909
rect 599945 122904 606556 122906
rect 599945 122848 599950 122904
rect 600006 122848 606556 122904
rect 599945 122846 606556 122848
rect 666356 122904 673059 122906
rect 666356 122848 666650 122904
rect 666706 122848 672998 122904
rect 673054 122848 673059 122904
rect 666356 122846 673059 122848
rect 599945 122843 600011 122846
rect 666645 122843 666711 122846
rect 672993 122843 673059 122846
rect 673421 122730 673491 122735
rect 673421 122670 673426 122730
rect 673486 122670 676386 122730
rect 673421 122665 673491 122670
rect 599577 121818 599643 121821
rect 599577 121816 606556 121818
rect 599577 121760 599582 121816
rect 599638 121760 606556 121816
rect 599577 121758 606556 121760
rect 599577 121755 599643 121758
rect 676262 121685 676322 121924
rect 676213 121680 676322 121685
rect 676213 121624 676218 121680
rect 676274 121624 676322 121680
rect 676213 121622 676322 121624
rect 676213 121619 676279 121622
rect 582097 121410 582163 121413
rect 576380 121408 582163 121410
rect 576380 121352 582102 121408
rect 582158 121352 582163 121408
rect 576380 121350 582163 121352
rect 582097 121347 582163 121350
rect 600037 120866 600103 120869
rect 600037 120864 606556 120866
rect 600037 120808 600042 120864
rect 600098 120808 606556 120864
rect 600037 120806 606556 120808
rect 600037 120803 600103 120806
rect 581729 119914 581795 119917
rect 576380 119912 581795 119914
rect 576380 119856 581734 119912
rect 581790 119856 581795 119912
rect 576380 119854 581795 119856
rect 581729 119851 581795 119854
rect 599853 119778 599919 119781
rect 599853 119776 606556 119778
rect 599853 119720 599858 119776
rect 599914 119720 606556 119776
rect 599853 119718 606556 119720
rect 599853 119715 599919 119718
rect 666645 119506 666711 119509
rect 666356 119504 666711 119506
rect 666356 119448 666650 119504
rect 666706 119448 666711 119504
rect 666356 119446 666711 119448
rect 666645 119443 666711 119446
rect 599945 118826 600011 118829
rect 599945 118824 606556 118826
rect 599945 118768 599950 118824
rect 600006 118768 606556 118824
rect 599945 118766 606556 118768
rect 599945 118763 600011 118766
rect 581453 118418 581519 118421
rect 576380 118416 581519 118418
rect 576380 118360 581458 118416
rect 581514 118360 581519 118416
rect 576380 118358 581519 118360
rect 581453 118355 581519 118358
rect 670341 117786 670407 117789
rect 666184 117784 670430 117786
rect 599853 117738 599919 117741
rect 599853 117736 606556 117738
rect 599853 117680 599858 117736
rect 599914 117680 606556 117736
rect 666184 117728 670346 117784
rect 670402 117728 670430 117784
rect 666184 117726 670430 117728
rect 670341 117723 670407 117726
rect 599853 117678 606556 117680
rect 599853 117675 599919 117678
rect 581913 116922 581979 116925
rect 576380 116920 581979 116922
rect 576380 116864 581918 116920
rect 581974 116864 581979 116920
rect 576380 116862 581979 116864
rect 581913 116859 581979 116862
rect 599945 116786 600011 116789
rect 599945 116784 606556 116786
rect 599945 116728 599950 116784
rect 600006 116728 606556 116784
rect 599945 116726 606556 116728
rect 599945 116723 600011 116726
rect 670497 116156 670563 116159
rect 666180 116154 670586 116156
rect 666180 116098 670502 116154
rect 670558 116098 670586 116154
rect 666180 116096 670586 116098
rect 670497 116093 670563 116096
rect 599853 115698 599919 115701
rect 599853 115696 606556 115698
rect 599853 115640 599858 115696
rect 599914 115640 606556 115696
rect 599853 115638 606556 115640
rect 599853 115635 599919 115638
rect 581269 115426 581335 115429
rect 576380 115424 581335 115426
rect 576380 115368 581274 115424
rect 581330 115368 581335 115424
rect 576380 115366 581335 115368
rect 581269 115363 581335 115366
rect 600037 114746 600103 114749
rect 600037 114744 606556 114746
rect 600037 114688 600042 114744
rect 600098 114688 606556 114744
rect 600037 114686 606556 114688
rect 600037 114683 600103 114686
rect 671981 114338 672047 114341
rect 666356 114336 672047 114338
rect 666356 114280 671986 114336
rect 672042 114280 672047 114336
rect 666356 114278 672047 114280
rect 671981 114275 672047 114278
rect 580993 113930 581059 113933
rect 576380 113928 581059 113930
rect 576380 113872 580998 113928
rect 581054 113872 581059 113928
rect 576380 113870 581059 113872
rect 580993 113867 581059 113870
rect 599945 113658 600011 113661
rect 599945 113656 606556 113658
rect 599945 113600 599950 113656
rect 600006 113600 606556 113656
rect 599945 113598 606556 113600
rect 599945 113595 600011 113598
rect 673279 112748 673345 112751
rect 666310 112746 673345 112748
rect 598933 112706 598999 112709
rect 598933 112704 606556 112706
rect 598933 112648 598938 112704
rect 598994 112648 606556 112704
rect 666310 112690 673284 112746
rect 673340 112690 673345 112746
rect 666310 112688 673345 112690
rect 673279 112685 673345 112688
rect 598933 112646 606556 112648
rect 598933 112643 598999 112646
rect 581545 112434 581611 112437
rect 576380 112432 581611 112434
rect 576380 112376 581550 112432
rect 581606 112376 581611 112432
rect 576380 112374 581611 112376
rect 581545 112371 581611 112374
rect 599945 111618 600011 111621
rect 599945 111616 606556 111618
rect 599945 111560 599950 111616
rect 600006 111560 606556 111616
rect 599945 111558 606556 111560
rect 599945 111555 600011 111558
rect 673413 110984 673479 110987
rect 666264 110982 673479 110984
rect 579889 110938 579955 110941
rect 576380 110936 579955 110938
rect 576380 110880 579894 110936
rect 579950 110880 579955 110936
rect 666264 110926 673418 110982
rect 673474 110926 673479 110982
rect 666264 110924 673479 110926
rect 673413 110921 673479 110924
rect 576380 110878 579955 110880
rect 579889 110875 579955 110878
rect 593370 110606 606556 110666
rect 580942 110468 580948 110532
rect 581012 110530 581018 110532
rect 593370 110530 593430 110606
rect 581012 110470 593430 110530
rect 581012 110468 581018 110470
rect 599853 109578 599919 109581
rect 599853 109576 606556 109578
rect 599853 109520 599858 109576
rect 599914 109520 606556 109576
rect 599853 109518 606556 109520
rect 599853 109515 599919 109518
rect 581085 109442 581151 109445
rect 576380 109440 581151 109442
rect 576380 109384 581090 109440
rect 581146 109384 581151 109440
rect 576380 109382 581151 109384
rect 581085 109379 581151 109382
rect 672441 109306 672507 109309
rect 666356 109304 672507 109306
rect 666356 109248 672446 109304
rect 672502 109248 672507 109304
rect 666356 109246 672507 109248
rect 672441 109243 672507 109246
rect 599945 108626 600011 108629
rect 599945 108624 606556 108626
rect 599945 108568 599950 108624
rect 600006 108568 606556 108624
rect 599945 108566 606556 108568
rect 599945 108563 600011 108566
rect 581361 107946 581427 107949
rect 576380 107944 581427 107946
rect 576380 107888 581366 107944
rect 581422 107888 581427 107944
rect 576380 107886 581427 107888
rect 581361 107883 581427 107886
rect 599853 107538 599919 107541
rect 670877 107538 670943 107541
rect 599853 107536 606556 107538
rect 599853 107480 599858 107536
rect 599914 107480 606556 107536
rect 599853 107478 606556 107480
rect 666356 107536 670943 107538
rect 666356 107480 670882 107536
rect 670938 107480 670943 107536
rect 666356 107478 670943 107480
rect 599853 107475 599919 107478
rect 670877 107475 670943 107478
rect 599945 106586 600011 106589
rect 599945 106584 606556 106586
rect 599945 106528 599950 106584
rect 600006 106528 606556 106584
rect 599945 106526 606556 106528
rect 599945 106523 600011 106526
rect 579981 106450 580047 106453
rect 576380 106448 580047 106450
rect 576380 106392 579986 106448
rect 580042 106392 580047 106448
rect 576380 106390 580047 106392
rect 579981 106387 580047 106390
rect 672257 105906 672323 105909
rect 666356 105904 672323 105906
rect 666356 105848 672262 105904
rect 672318 105848 672323 105904
rect 666356 105846 672323 105848
rect 672257 105843 672323 105846
rect 600221 105498 600287 105501
rect 600221 105496 606556 105498
rect 600221 105440 600226 105496
rect 600282 105440 606556 105496
rect 600221 105438 606556 105440
rect 600221 105435 600287 105438
rect 579797 104954 579863 104957
rect 576380 104952 579863 104954
rect 576380 104896 579802 104952
rect 579858 104896 579863 104952
rect 576380 104894 579863 104896
rect 579797 104891 579863 104894
rect 600497 104546 600563 104549
rect 600497 104544 606556 104546
rect 600497 104488 600502 104544
rect 600558 104488 606556 104544
rect 600497 104486 606556 104488
rect 600497 104483 600563 104486
rect 672165 104138 672231 104141
rect 666356 104136 672231 104138
rect 666356 104080 672170 104136
rect 672226 104080 672231 104136
rect 666356 104078 672231 104080
rect 672165 104075 672231 104078
rect 580901 103458 580967 103461
rect 576380 103456 580967 103458
rect 576380 103400 580906 103456
rect 580962 103400 580967 103456
rect 576380 103398 580967 103400
rect 580901 103395 580967 103398
rect 600681 103458 600747 103461
rect 600681 103456 606556 103458
rect 600681 103400 600686 103456
rect 600742 103400 606556 103456
rect 600681 103398 606556 103400
rect 600681 103395 600747 103398
rect 600313 102506 600379 102509
rect 672349 102506 672415 102509
rect 600313 102504 606556 102506
rect 600313 102448 600318 102504
rect 600374 102448 606556 102504
rect 600313 102446 606556 102448
rect 666356 102504 672415 102506
rect 666356 102448 672354 102504
rect 672410 102448 672415 102504
rect 666356 102446 672415 102448
rect 600313 102443 600379 102446
rect 672349 102443 672415 102446
rect 580441 101962 580507 101965
rect 576380 101960 580507 101962
rect 576380 101904 580446 101960
rect 580502 101904 580507 101960
rect 576380 101902 580507 101904
rect 580441 101899 580507 101902
rect 600405 101418 600471 101421
rect 600405 101416 606556 101418
rect 600405 101360 600410 101416
rect 600466 101360 606556 101416
rect 600405 101358 606556 101360
rect 600405 101355 600471 101358
rect 672073 100874 672139 100877
rect 666356 100872 672139 100874
rect 666356 100816 672078 100872
rect 672134 100816 672139 100872
rect 666356 100814 672139 100816
rect 672073 100811 672139 100814
rect 599945 100466 600011 100469
rect 599945 100464 606556 100466
rect 599945 100408 599950 100464
rect 600006 100408 606556 100464
rect 599945 100406 606556 100408
rect 599945 100403 600011 100406
rect 580073 100330 580139 100333
rect 576380 100328 580139 100330
rect 576380 100272 580078 100328
rect 580134 100272 580139 100328
rect 576380 100270 580139 100272
rect 580073 100267 580139 100270
rect 580625 98834 580691 98837
rect 576380 98832 580691 98834
rect 576380 98776 580630 98832
rect 580686 98776 580691 98832
rect 576380 98774 580691 98776
rect 580625 98771 580691 98774
rect 581177 97338 581243 97341
rect 576380 97336 581243 97338
rect 576380 97280 581182 97336
rect 581238 97280 581243 97336
rect 576380 97278 581243 97280
rect 581177 97275 581243 97278
rect 628281 95978 628347 95981
rect 628238 95976 628347 95978
rect 628238 95920 628286 95976
rect 628342 95920 628347 95976
rect 628238 95915 628347 95920
rect 633198 95916 633204 95980
rect 633268 95978 633274 95980
rect 642265 95978 642331 95981
rect 633268 95976 642331 95978
rect 633268 95920 642270 95976
rect 642326 95920 642331 95976
rect 633268 95918 642331 95920
rect 633268 95916 633274 95918
rect 642265 95915 642331 95918
rect 582189 95842 582255 95845
rect 576380 95840 582255 95842
rect 576380 95784 582194 95840
rect 582250 95784 582255 95840
rect 576380 95782 582255 95784
rect 582189 95779 582255 95782
rect 628238 95404 628298 95915
rect 662086 95508 662092 95572
rect 662156 95570 662162 95572
rect 662229 95570 662295 95573
rect 662156 95568 662295 95570
rect 662156 95512 662234 95568
rect 662290 95512 662295 95568
rect 662156 95510 662295 95512
rect 662156 95508 662162 95510
rect 662229 95507 662295 95510
rect 642725 95162 642791 95165
rect 642725 95160 642834 95162
rect 642725 95104 642730 95160
rect 642786 95104 642834 95160
rect 642725 95099 642834 95104
rect 642774 94588 642834 95099
rect 657353 94754 657419 94757
rect 657310 94752 657419 94754
rect 657310 94696 657358 94752
rect 657414 94696 657419 94752
rect 657310 94691 657419 94696
rect 627913 94482 627979 94485
rect 627913 94480 628268 94482
rect 627913 94424 627918 94480
rect 627974 94424 628268 94480
rect 627913 94422 628268 94424
rect 627913 94419 627979 94422
rect 580257 94346 580323 94349
rect 576380 94344 580323 94346
rect 576380 94288 580262 94344
rect 580318 94288 580323 94344
rect 576380 94286 580323 94288
rect 580257 94283 580323 94286
rect 657310 94180 657370 94691
rect 663241 93802 663307 93805
rect 663198 93800 663307 93802
rect 663198 93744 663246 93800
rect 663302 93744 663307 93800
rect 663198 93739 663307 93744
rect 627269 93530 627335 93533
rect 627269 93528 628268 93530
rect 627269 93472 627274 93528
rect 627330 93472 628268 93528
rect 627269 93470 628268 93472
rect 627269 93467 627335 93470
rect 655329 93394 655395 93397
rect 655329 93392 656788 93394
rect 655329 93336 655334 93392
rect 655390 93336 656788 93392
rect 663198 93364 663258 93739
rect 655329 93334 656788 93336
rect 655329 93331 655395 93334
rect 663333 93122 663399 93125
rect 663333 93120 663442 93122
rect 663333 93064 663338 93120
rect 663394 93064 663442 93120
rect 663333 93059 663442 93064
rect 580165 92850 580231 92853
rect 576380 92848 580231 92850
rect 576380 92792 580170 92848
rect 580226 92792 580231 92848
rect 576380 92790 580231 92792
rect 580165 92787 580231 92790
rect 642633 92714 642699 92717
rect 642590 92712 642699 92714
rect 642590 92656 642638 92712
rect 642694 92656 642699 92712
rect 642590 92651 642699 92656
rect 626441 92578 626507 92581
rect 626441 92576 628268 92578
rect 626441 92520 626446 92576
rect 626502 92520 628268 92576
rect 626441 92518 628268 92520
rect 626441 92515 626507 92518
rect 642590 92140 642650 92651
rect 651557 92578 651623 92581
rect 651557 92576 656788 92578
rect 651557 92520 651562 92576
rect 651618 92520 656788 92576
rect 663382 92548 663442 93059
rect 651557 92518 656788 92520
rect 651557 92515 651623 92518
rect 663425 92306 663491 92309
rect 663382 92304 663491 92306
rect 663382 92248 663430 92304
rect 663486 92248 663491 92304
rect 663382 92243 663491 92248
rect 663382 91732 663442 92243
rect 625889 91626 625955 91629
rect 625889 91624 628268 91626
rect 625889 91568 625894 91624
rect 625950 91568 628268 91624
rect 625889 91566 628268 91568
rect 625889 91563 625955 91566
rect 654041 91490 654107 91493
rect 654041 91488 656788 91490
rect 654041 91432 654046 91488
rect 654102 91432 656788 91488
rect 654041 91430 656788 91432
rect 654041 91427 654107 91430
rect 580349 91354 580415 91357
rect 576380 91352 580415 91354
rect 576380 91296 580354 91352
rect 580410 91296 580415 91352
rect 576380 91294 580415 91296
rect 580349 91291 580415 91294
rect 663885 91082 663951 91085
rect 663566 91080 663951 91082
rect 663566 91024 663890 91080
rect 663946 91024 663951 91080
rect 663566 91022 663951 91024
rect 623773 90674 623839 90677
rect 652753 90674 652819 90677
rect 623773 90672 628268 90674
rect 623773 90616 623778 90672
rect 623834 90616 628268 90672
rect 623773 90614 628268 90616
rect 652753 90672 656788 90674
rect 652753 90616 652758 90672
rect 652814 90616 656788 90672
rect 663566 90644 663626 91022
rect 663885 91019 663951 91022
rect 652753 90614 656788 90616
rect 623773 90611 623839 90614
rect 652753 90611 652819 90614
rect 656893 90402 656959 90405
rect 663701 90402 663767 90405
rect 656893 90400 657002 90402
rect 656893 90344 656898 90400
rect 656954 90344 657002 90400
rect 656893 90339 657002 90344
rect 580717 89858 580783 89861
rect 576380 89856 580783 89858
rect 576380 89800 580722 89856
rect 580778 89800 580783 89856
rect 656942 89828 657002 90339
rect 663566 90400 663767 90402
rect 663566 90344 663706 90400
rect 663762 90344 663767 90400
rect 663566 90342 663767 90344
rect 663566 89828 663626 90342
rect 663701 90339 663767 90342
rect 576380 89798 580783 89800
rect 580717 89795 580783 89798
rect 623957 89722 624023 89725
rect 646037 89722 646103 89725
rect 623957 89720 628268 89722
rect 623957 89664 623962 89720
rect 624018 89664 628268 89720
rect 623957 89662 628268 89664
rect 642988 89720 646103 89722
rect 642988 89664 646042 89720
rect 646098 89664 646103 89720
rect 642988 89662 646103 89664
rect 623957 89659 624023 89662
rect 646037 89659 646103 89662
rect 663517 89586 663583 89589
rect 663517 89584 663626 89586
rect 663517 89528 663522 89584
rect 663578 89528 663626 89584
rect 663517 89523 663626 89528
rect 663566 89012 663626 89523
rect 622485 88906 622551 88909
rect 622485 88904 628268 88906
rect 622485 88848 622490 88904
rect 622546 88848 628268 88904
rect 622485 88846 628268 88848
rect 622485 88843 622551 88846
rect 662137 88772 662203 88773
rect 662086 88708 662092 88772
rect 662156 88770 662203 88772
rect 662156 88768 662248 88770
rect 662198 88712 662248 88768
rect 662156 88710 662248 88712
rect 662156 88708 662203 88710
rect 662137 88707 662203 88708
rect 580533 88362 580599 88365
rect 576380 88360 580599 88362
rect 576380 88304 580538 88360
rect 580594 88304 580599 88360
rect 576380 88302 580599 88304
rect 580533 88299 580599 88302
rect 623221 87954 623287 87957
rect 623221 87952 628268 87954
rect 623221 87896 623226 87952
rect 623282 87896 628268 87952
rect 623221 87894 628268 87896
rect 623221 87891 623287 87894
rect 645945 87138 646011 87141
rect 642988 87136 646011 87138
rect 642988 87080 645950 87136
rect 646006 87080 646011 87136
rect 642988 87078 646011 87080
rect 645945 87075 646011 87078
rect 623497 87002 623563 87005
rect 623497 87000 628268 87002
rect 623497 86944 623502 87000
rect 623558 86944 628268 87000
rect 623497 86942 628268 86944
rect 623497 86939 623563 86942
rect 580809 86866 580875 86869
rect 576380 86864 580875 86866
rect 576380 86808 580814 86864
rect 580870 86808 580875 86864
rect 576380 86806 580875 86808
rect 580809 86803 580875 86806
rect 621197 86050 621263 86053
rect 621197 86048 628268 86050
rect 621197 85992 621202 86048
rect 621258 85992 628268 86048
rect 621197 85990 628268 85992
rect 621197 85987 621263 85990
rect 582005 85370 582071 85373
rect 576380 85368 582071 85370
rect 576380 85312 582010 85368
rect 582066 85312 582071 85368
rect 576380 85310 582071 85312
rect 582005 85307 582071 85310
rect 623313 85098 623379 85101
rect 623313 85096 628268 85098
rect 623313 85040 623318 85096
rect 623374 85040 628268 85096
rect 623313 85038 628268 85040
rect 623313 85035 623379 85038
rect 646129 84690 646195 84693
rect 642988 84688 646195 84690
rect 642988 84632 646134 84688
rect 646190 84632 646195 84688
rect 642988 84630 646195 84632
rect 646129 84627 646195 84630
rect 623129 84146 623195 84149
rect 623129 84144 628268 84146
rect 623129 84088 623134 84144
rect 623190 84088 628268 84144
rect 623129 84086 628268 84088
rect 623129 84083 623195 84086
rect 582281 83874 582347 83877
rect 576380 83872 582347 83874
rect 576380 83816 582286 83872
rect 582342 83816 582347 83872
rect 576380 83814 582347 83816
rect 582281 83811 582347 83814
rect 621933 83194 621999 83197
rect 621933 83192 628268 83194
rect 621933 83136 621938 83192
rect 621994 83136 628268 83192
rect 621933 83134 628268 83136
rect 621933 83131 621999 83134
rect 579981 82378 580047 82381
rect 576380 82376 580047 82378
rect 576380 82320 579986 82376
rect 580042 82320 580047 82376
rect 576380 82318 580047 82320
rect 579981 82315 580047 82318
rect 645853 82242 645919 82245
rect 642988 82240 645919 82242
rect 628606 81701 628666 82212
rect 642988 82184 645858 82240
rect 645914 82184 645919 82240
rect 642988 82182 645919 82184
rect 645853 82179 645919 82182
rect 628557 81696 628666 81701
rect 628557 81640 628562 81696
rect 628618 81640 628666 81696
rect 628557 81638 628666 81640
rect 628557 81635 628623 81638
rect 579613 80882 579679 80885
rect 576380 80880 579679 80882
rect 576380 80824 579618 80880
rect 579674 80824 579679 80880
rect 576380 80822 579679 80824
rect 628790 80882 628850 81396
rect 629201 80882 629267 80885
rect 628790 80880 629267 80882
rect 628790 80824 629206 80880
rect 629262 80824 629267 80880
rect 628790 80822 629267 80824
rect 579613 80819 579679 80822
rect 629201 80819 629267 80822
rect 626533 80202 626599 80205
rect 628465 80202 628531 80205
rect 626533 80200 628531 80202
rect 626533 80144 626538 80200
rect 626594 80144 628470 80200
rect 628526 80144 628531 80200
rect 626533 80142 628531 80144
rect 626533 80139 626599 80142
rect 628465 80139 628531 80142
rect 633198 80140 633204 80204
rect 633268 80202 633274 80204
rect 634169 80202 634235 80205
rect 633268 80200 634235 80202
rect 633268 80144 634174 80200
rect 634230 80144 634235 80200
rect 633268 80142 634235 80144
rect 633268 80140 633274 80142
rect 634169 80139 634235 80142
rect 582097 79386 582163 79389
rect 576380 79384 582163 79386
rect 576380 79328 582102 79384
rect 582158 79328 582163 79384
rect 576380 79326 582163 79328
rect 582097 79323 582163 79326
rect 581821 77890 581887 77893
rect 576380 77888 581887 77890
rect 576380 77832 581826 77888
rect 581882 77832 581887 77888
rect 576380 77830 581887 77832
rect 581821 77827 581887 77830
rect 581729 76258 581795 76261
rect 576380 76256 581795 76258
rect 576380 76200 581734 76256
rect 581790 76200 581795 76256
rect 576380 76198 581795 76200
rect 581729 76195 581795 76198
rect 626758 75516 626764 75580
rect 626828 75578 626834 75580
rect 628465 75578 628531 75581
rect 626828 75576 628531 75578
rect 626828 75520 628470 75576
rect 628526 75520 628531 75576
rect 626828 75518 628531 75520
rect 626828 75516 626834 75518
rect 628465 75515 628531 75518
rect 633198 75516 633204 75580
rect 633268 75578 633274 75580
rect 634169 75578 634235 75581
rect 633268 75576 634235 75578
rect 633268 75520 634174 75576
rect 634230 75520 634235 75576
rect 633268 75518 634235 75520
rect 633268 75516 633274 75518
rect 634169 75515 634235 75518
rect 640333 75442 640399 75445
rect 640333 75440 640994 75442
rect 640333 75384 640338 75440
rect 640394 75384 640994 75440
rect 640333 75382 640994 75384
rect 640333 75379 640399 75382
rect 640934 74868 640994 75382
rect 581913 74762 581979 74765
rect 576380 74760 581979 74762
rect 576380 74704 581918 74760
rect 581974 74704 581979 74760
rect 576380 74702 581979 74704
rect 581913 74699 581979 74702
rect 642817 73402 642883 73405
rect 641516 73400 642883 73402
rect 641516 73344 642822 73400
rect 642878 73344 642883 73400
rect 641516 73342 642883 73344
rect 642817 73339 642883 73342
rect 581637 73266 581703 73269
rect 576380 73264 581703 73266
rect 576380 73208 581642 73264
rect 581698 73208 581703 73264
rect 576380 73206 581703 73208
rect 581637 73203 581703 73206
rect 640977 72450 641043 72453
rect 640977 72448 641178 72450
rect 640977 72392 640982 72448
rect 641038 72392 641178 72448
rect 640977 72390 641178 72392
rect 640977 72387 641043 72390
rect 641118 71876 641178 72390
rect 581453 71770 581519 71773
rect 576380 71768 581519 71770
rect 576380 71712 581458 71768
rect 581514 71712 581519 71768
rect 576380 71710 581519 71712
rect 581453 71707 581519 71710
rect 641069 70954 641135 70957
rect 641069 70952 641178 70954
rect 641069 70896 641074 70952
rect 641130 70896 641178 70952
rect 641069 70891 641178 70896
rect 641118 70380 641178 70891
rect 581269 70274 581335 70277
rect 576380 70272 581335 70274
rect 576380 70216 581274 70272
rect 581330 70216 581335 70272
rect 576380 70214 581335 70216
rect 581269 70211 581335 70214
rect 576158 69396 576164 69460
rect 576228 69458 576234 69460
rect 591941 69458 592007 69461
rect 576228 69456 592007 69458
rect 576228 69400 591946 69456
rect 592002 69400 592007 69456
rect 576228 69398 592007 69400
rect 576228 69396 576234 69398
rect 591941 69395 592007 69398
rect 642909 68914 642975 68917
rect 641516 68912 642975 68914
rect 641516 68856 642914 68912
rect 642970 68856 642975 68912
rect 641516 68854 642975 68856
rect 642909 68851 642975 68854
rect 580942 68778 580948 68780
rect 576380 68718 580948 68778
rect 580942 68716 580948 68718
rect 581012 68716 581018 68780
rect 643001 67418 643067 67421
rect 641516 67416 643067 67418
rect 641516 67360 643006 67416
rect 643062 67360 643067 67416
rect 641516 67358 643067 67360
rect 643001 67355 643067 67358
rect 581545 67282 581611 67285
rect 576380 67280 581611 67282
rect 576380 67224 581550 67280
rect 581606 67224 581611 67280
rect 576380 67222 581611 67224
rect 581545 67219 581611 67222
rect 642633 65922 642699 65925
rect 641516 65920 642699 65922
rect 641516 65864 642638 65920
rect 642694 65864 642699 65920
rect 641516 65862 642699 65864
rect 642633 65859 642699 65862
rect 580993 65786 581059 65789
rect 576380 65784 581059 65786
rect 576380 65728 580998 65784
rect 581054 65728 581059 65784
rect 576380 65726 581059 65728
rect 580993 65723 581059 65726
rect 643093 64426 643159 64429
rect 641516 64424 643159 64426
rect 641516 64368 643098 64424
rect 643154 64368 643159 64424
rect 641516 64366 643159 64368
rect 643093 64363 643159 64366
rect 581361 64290 581427 64293
rect 576380 64288 581427 64290
rect 576380 64232 581366 64288
rect 581422 64232 581427 64288
rect 576380 64230 581427 64232
rect 581361 64227 581427 64230
rect 581085 62794 581151 62797
rect 576380 62792 581151 62794
rect 576380 62736 581090 62792
rect 581146 62736 581151 62792
rect 576380 62734 581151 62736
rect 581085 62731 581151 62734
rect 580717 61298 580783 61301
rect 576380 61296 580783 61298
rect 576380 61240 580722 61296
rect 580778 61240 580783 61296
rect 576380 61238 580783 61240
rect 580717 61235 580783 61238
rect 579613 59802 579679 59805
rect 576380 59800 579679 59802
rect 576380 59744 579618 59800
rect 579674 59744 579679 59800
rect 576380 59742 579679 59744
rect 579613 59739 579679 59742
rect 579613 58306 579679 58309
rect 576380 58304 579679 58306
rect 576380 58248 579618 58304
rect 579674 58248 579679 58304
rect 576380 58246 579679 58248
rect 579613 58243 579679 58246
rect 580809 56810 580875 56813
rect 576380 56808 580875 56810
rect 576380 56752 580814 56808
rect 580870 56752 580875 56808
rect 576380 56750 580875 56752
rect 580809 56747 580875 56750
rect 580625 55314 580691 55317
rect 576380 55312 580691 55314
rect 576380 55256 580630 55312
rect 580686 55256 580691 55312
rect 576380 55254 580691 55256
rect 580625 55251 580691 55254
rect 580901 53818 580967 53821
rect 576380 53816 580967 53818
rect 576380 53760 580906 53816
rect 580962 53760 580967 53816
rect 576380 53758 580967 53760
rect 580901 53755 580967 53758
rect 339401 52458 339467 52461
rect 346945 52458 347011 52461
rect 626758 52458 626764 52460
rect 339401 52456 626764 52458
rect 339401 52400 339406 52456
rect 339462 52400 346950 52456
rect 347006 52400 626764 52456
rect 339401 52398 626764 52400
rect 339401 52395 339467 52398
rect 346945 52395 347011 52398
rect 626758 52396 626764 52398
rect 626828 52396 626834 52460
rect 184933 51098 184999 51101
rect 633198 51098 633204 51100
rect 184933 51096 633204 51098
rect 184933 51040 184938 51096
rect 184994 51040 633204 51096
rect 184933 51038 633204 51040
rect 184933 51035 184999 51038
rect 633198 51036 633204 51038
rect 633268 51036 633274 51100
rect 590694 49676 590700 49740
rect 590764 49738 590770 49740
rect 597461 49738 597527 49741
rect 590764 49736 597527 49738
rect 590764 49680 597466 49736
rect 597522 49680 597527 49736
rect 590764 49678 597527 49680
rect 590764 49676 590770 49678
rect 597461 49675 597527 49678
rect 666553 49058 666619 49061
rect 661358 49056 666619 49058
rect 661358 49000 666558 49056
rect 666614 49000 666619 49056
rect 661358 48998 666619 49000
rect 661358 48482 661418 48998
rect 666553 48995 666619 48998
rect 216121 48242 216187 48245
rect 521694 48242 521700 48244
rect 216121 48240 521700 48242
rect 216121 48184 216126 48240
rect 216182 48184 521700 48240
rect 216121 48182 521700 48184
rect 216121 48179 216187 48182
rect 521694 48180 521700 48182
rect 521764 48180 521770 48244
rect 470133 43210 470199 43213
rect 600037 43210 600103 43213
rect 470133 43208 600103 43210
rect 470133 43152 470138 43208
rect 470194 43152 600042 43208
rect 600098 43152 600103 43208
rect 470133 43150 600103 43152
rect 470133 43147 470199 43150
rect 600037 43147 600103 43150
rect 521745 42124 521811 42125
rect 521694 42060 521700 42124
rect 521764 42122 521811 42124
rect 521764 42120 521856 42122
rect 521806 42064 521856 42120
rect 521764 42062 521856 42064
rect 521764 42060 521811 42062
rect 521745 42059 521811 42060
rect 194317 41850 194383 41853
rect 307293 41852 307359 41853
rect 194317 41848 194426 41850
rect 194317 41792 194322 41848
rect 194378 41792 194426 41848
rect 194317 41787 194426 41792
rect 307293 41848 307340 41852
rect 307404 41850 307410 41852
rect 361941 41850 362007 41853
rect 415485 41850 415551 41853
rect 416773 41852 416839 41853
rect 307293 41792 307298 41848
rect 307293 41788 307340 41792
rect 307404 41790 307450 41850
rect 361941 41848 362050 41850
rect 361941 41792 361946 41848
rect 362002 41792 362050 41848
rect 307404 41788 307410 41790
rect 307293 41787 307359 41788
rect 361941 41787 362050 41792
rect 415485 41848 415594 41850
rect 415485 41792 415490 41848
rect 415546 41792 415594 41848
rect 415485 41787 415594 41792
rect 416773 41848 416820 41852
rect 416884 41850 416890 41852
rect 419809 41850 419875 41853
rect 471697 41850 471763 41853
rect 520365 41850 520431 41853
rect 416773 41792 416778 41848
rect 416773 41788 416820 41792
rect 416884 41790 416930 41850
rect 419809 41848 420010 41850
rect 419809 41792 419814 41848
rect 419870 41792 420010 41848
rect 419809 41790 420010 41792
rect 416884 41788 416890 41790
rect 416773 41787 416839 41788
rect 419809 41787 419875 41790
rect 194366 41306 194426 41787
rect 223573 41306 223639 41309
rect 194366 41304 223639 41306
rect 194366 41248 223578 41304
rect 223634 41248 223639 41304
rect 194366 41246 223639 41248
rect 361990 41306 362050 41787
rect 390185 41306 390251 41309
rect 361990 41304 390251 41306
rect 361990 41248 390190 41304
rect 390246 41248 390251 41304
rect 361990 41246 390251 41248
rect 223573 41243 223639 41246
rect 390185 41243 390251 41246
rect 415534 41170 415594 41787
rect 419950 41306 420010 41790
rect 471697 41848 477510 41850
rect 471697 41792 471702 41848
rect 471758 41792 477510 41848
rect 471697 41790 477510 41792
rect 471697 41787 471763 41790
rect 477450 41442 477510 41790
rect 516090 41848 520431 41850
rect 516090 41792 520370 41848
rect 520426 41792 520431 41848
rect 516090 41790 520431 41792
rect 513189 41714 513255 41717
rect 516090 41714 516150 41790
rect 520365 41787 520431 41790
rect 513189 41712 516150 41714
rect 513189 41656 513194 41712
rect 513250 41656 516150 41712
rect 513189 41654 516150 41656
rect 513189 41651 513255 41654
rect 568573 41442 568639 41445
rect 477450 41440 568639 41442
rect 477450 41384 568578 41440
rect 568634 41384 568639 41440
rect 477450 41382 568639 41384
rect 568573 41379 568639 41382
rect 543641 41306 543707 41309
rect 419950 41304 543707 41306
rect 419950 41248 543646 41304
rect 543702 41248 543707 41304
rect 419950 41246 543707 41248
rect 543641 41243 543707 41246
rect 530301 41170 530367 41173
rect 415534 41168 530367 41170
rect 415534 41112 530306 41168
rect 530362 41112 530367 41168
rect 415534 41110 530367 41112
rect 530301 41107 530367 41110
rect 475469 41034 475535 41037
rect 530393 41034 530459 41037
rect 475469 41032 530459 41034
rect 475469 40976 475474 41032
rect 475530 40976 530398 41032
rect 530454 40976 530459 41032
rect 475469 40974 530459 40976
rect 475469 40971 475535 40974
rect 530393 40971 530459 40974
<< via3 >>
rect 674420 895460 674484 895524
rect 673868 893828 673932 893892
rect 679204 886620 679268 886684
rect 679204 885804 679268 885868
rect 679204 884988 679268 885052
rect 41828 809100 41892 809164
rect 41828 794472 41892 794476
rect 41828 794416 41878 794472
rect 41878 794416 41892 794472
rect 41828 794412 41892 794416
rect 674972 788292 675036 788356
rect 675156 787128 675220 787132
rect 675156 787072 675206 787128
rect 675206 787072 675220 787128
rect 675156 787068 675220 787072
rect 674052 786796 674116 786860
rect 42012 757012 42076 757076
rect 42748 757012 42812 757076
rect 42748 752932 42812 752996
rect 42012 748716 42076 748780
rect 675340 742928 675404 742932
rect 675340 742872 675390 742928
rect 675390 742872 675404 742928
rect 675340 742868 675404 742872
rect 676648 742732 676712 742796
rect 676812 742596 676876 742660
rect 675708 742520 675772 742524
rect 675708 742464 675722 742520
rect 675722 742464 675772 742520
rect 675708 742460 675772 742464
rect 674236 740284 674300 740348
rect 674604 740148 674668 740212
rect 673500 739604 673564 739668
rect 674788 738652 674852 738716
rect 677180 737972 677244 738036
rect 675524 728996 675588 729060
rect 675524 728180 675588 728244
rect 674052 724644 674116 724708
rect 674052 724236 674116 724300
rect 674420 724236 674484 724300
rect 673868 724100 673932 724164
rect 675156 724100 675220 724164
rect 674420 723964 674484 724028
rect 674972 723964 675036 724028
rect 675892 721516 675956 721580
rect 674052 715260 674116 715324
rect 43116 714368 43180 714372
rect 43116 714312 43130 714368
rect 43130 714312 43180 714368
rect 43116 714308 43180 714312
rect 43668 714172 43732 714236
rect 673684 713628 673748 713692
rect 675892 711996 675956 712060
rect 43116 711452 43180 711516
rect 674420 711180 674484 711244
rect 673868 709548 673932 709612
rect 42748 709412 42812 709476
rect 42748 708868 42812 708932
rect 43668 708460 43732 708524
rect 676076 707236 676140 707300
rect 675892 706692 675956 706756
rect 676996 699620 677060 699684
rect 673868 698124 673932 698188
rect 676076 697172 676140 697236
rect 676812 696628 676876 696692
rect 675892 694724 675956 694788
rect 674052 694316 674116 694380
rect 676648 693500 676712 693564
rect 677180 692956 677244 693020
rect 673684 690508 673748 690572
rect 674420 690100 674484 690164
rect 674236 681124 674300 681188
rect 674236 680308 674300 680372
rect 674604 680308 674668 680372
rect 674604 680172 674668 680236
rect 675340 680172 675404 680236
rect 675892 678464 675956 678468
rect 675892 678408 675942 678464
rect 675942 678408 675956 678464
rect 675892 678404 675956 678408
rect 41460 677724 41524 677788
rect 41460 676908 41524 676972
rect 674604 674732 674668 674796
rect 675340 674732 675404 674796
rect 675892 674792 675956 674796
rect 675892 674736 675942 674792
rect 675942 674736 675956 674792
rect 675892 674732 675956 674736
rect 674236 674596 674300 674660
rect 674604 674596 674668 674660
rect 674236 674052 674300 674116
rect 43300 671060 43364 671124
rect 42932 670652 42996 670716
rect 42932 670516 42996 670580
rect 43852 670516 43916 670580
rect 43300 670380 43364 670444
rect 674236 666844 674300 666908
rect 675340 666028 675404 666092
rect 674604 665620 674668 665684
rect 43852 665212 43916 665276
rect 675708 664396 675772 664460
rect 673500 663988 673564 664052
rect 674788 663580 674852 663644
rect 677364 662492 677428 662556
rect 676996 662084 677060 662148
rect 675708 652624 675772 652628
rect 675708 652568 675722 652624
rect 675722 652568 675772 652624
rect 675708 652564 675772 652568
rect 675156 652156 675220 652220
rect 675340 651672 675404 651676
rect 675340 651616 675390 651672
rect 675390 651616 675404 651672
rect 675340 651612 675404 651616
rect 674972 648892 675036 648956
rect 673500 648620 673564 648684
rect 674788 641684 674852 641748
rect 676076 641684 676140 641748
rect 674604 641548 674668 641612
rect 675892 641548 675956 641612
rect 673868 640188 673932 640252
rect 675708 638208 675772 638212
rect 675708 638152 675758 638208
rect 675758 638152 675772 638208
rect 675708 638148 675772 638152
rect 675340 637604 675404 637668
rect 674788 629308 674852 629372
rect 41828 627464 41892 627468
rect 41828 627408 41842 627464
rect 41842 627408 41892 627464
rect 41828 627404 41892 627408
rect 42380 627464 42444 627468
rect 42380 627408 42430 627464
rect 42430 627408 42444 627464
rect 42380 627404 42444 627408
rect 677548 622780 677612 622844
rect 42380 621964 42444 622028
rect 676812 621964 676876 622028
rect 41828 621480 41892 621484
rect 41828 621424 41878 621480
rect 41878 621424 41892 621480
rect 41828 621420 41892 621424
rect 674420 620604 674484 620668
rect 673684 620196 673748 620260
rect 674604 619380 674668 619444
rect 674052 618972 674116 619036
rect 676648 618700 676712 618764
rect 677180 617476 677244 617540
rect 677364 617068 677428 617132
rect 674236 616932 674300 616996
rect 676668 609180 676732 609244
rect 673684 607820 673748 607884
rect 676076 607276 676140 607340
rect 674236 604964 674300 605028
rect 674604 604420 674668 604484
rect 675340 604480 675404 604484
rect 675340 604424 675354 604480
rect 675354 604424 675404 604480
rect 675340 604420 675404 604424
rect 674420 603740 674484 603804
rect 673868 601836 673932 601900
rect 674052 587964 674116 588028
rect 675156 587964 675220 588028
rect 676076 587752 676140 587756
rect 676076 587696 676090 587752
rect 676090 587696 676140 587752
rect 676076 587692 676140 587696
rect 676076 586256 676140 586260
rect 676076 586200 676090 586256
rect 676090 586200 676140 586256
rect 676076 586196 676140 586200
rect 42196 585244 42260 585308
rect 41828 584216 41892 584220
rect 41828 584160 41842 584216
rect 41842 584160 41892 584216
rect 41828 584156 41892 584160
rect 42932 583884 42996 583948
rect 42932 581844 42996 581908
rect 41828 580620 41892 580684
rect 676996 579260 677060 579324
rect 677548 578444 677612 578508
rect 677180 577628 677244 577692
rect 42196 577008 42260 577012
rect 42196 576952 42210 577008
rect 42210 576952 42260 577008
rect 42196 576948 42260 576952
rect 676812 576812 676876 576876
rect 674788 576540 674852 576604
rect 674052 574092 674116 574156
rect 674972 573684 675036 573748
rect 673500 573276 673564 573340
rect 676668 571916 676732 571980
rect 677364 571508 677428 571572
rect 675156 562396 675220 562460
rect 674052 562260 674116 562324
rect 674972 561172 675036 561236
rect 674788 557500 674852 557564
rect 41644 556684 41708 556748
rect 42380 556004 42444 556068
rect 44036 555188 44100 555252
rect 39988 554236 40052 554300
rect 42564 553964 42628 554028
rect 675524 553828 675588 553892
rect 42748 553148 42812 553212
rect 42196 552740 42260 552804
rect 42932 552332 42996 552396
rect 41828 551516 41892 551580
rect 41460 550972 41524 551036
rect 42012 550700 42076 550764
rect 675524 548040 675588 548044
rect 675524 547984 675538 548040
rect 675538 547984 675588 548040
rect 675524 547980 675588 547984
rect 677180 544036 677244 544100
rect 676812 543900 676876 543964
rect 676996 543764 677060 543828
rect 673684 543084 673748 543148
rect 674420 543084 674484 543148
rect 674604 542676 674668 542740
rect 675340 542676 675404 542740
rect 676076 542736 676140 542740
rect 676076 542680 676126 542736
rect 676126 542680 676140 542736
rect 676076 542676 676140 542680
rect 676076 541240 676140 541244
rect 676076 541184 676126 541240
rect 676126 541184 676140 541240
rect 676076 541180 676140 541184
rect 41644 538460 41708 538524
rect 42932 538324 42996 538388
rect 42380 538188 42444 538252
rect 42012 538052 42076 538116
rect 41460 535332 41524 535396
rect 42564 535332 42628 535396
rect 42196 532748 42260 532812
rect 41828 532612 41892 532676
rect 42748 532612 42812 532676
rect 674420 531796 674484 531860
rect 673500 530980 673564 531044
rect 674236 530572 674300 530636
rect 676076 529348 676140 529412
rect 674604 528940 674668 529004
rect 673684 528532 673748 528596
rect 673868 527036 673932 527100
rect 674972 487596 675036 487660
rect 675156 486780 675220 486844
rect 674052 485148 674116 485212
rect 674788 484740 674852 484804
rect 39988 435916 40052 435980
rect 44036 428028 44100 428092
rect 43116 411436 43180 411500
rect 43116 406872 43180 406876
rect 43116 406816 43166 406872
rect 43166 406816 43180 406872
rect 43116 406812 43180 406816
rect 675156 400556 675220 400620
rect 41644 383012 41708 383076
rect 41460 382196 41524 382260
rect 41644 356900 41708 356964
rect 41460 355676 41524 355740
rect 675156 355812 675220 355876
rect 41460 340172 41524 340236
rect 41644 337316 41708 337380
rect 41828 337180 41892 337244
rect 42564 336772 42628 336836
rect 42196 330108 42260 330172
rect 42012 329972 42076 330036
rect 42380 329836 42444 329900
rect 42564 316372 42628 316436
rect 41828 316296 41892 316300
rect 41828 316240 41842 316296
rect 41842 316240 41892 316296
rect 41828 316236 41892 316240
rect 42380 315420 42444 315484
rect 42012 313848 42076 313852
rect 42012 313792 42026 313848
rect 42026 313792 42076 313848
rect 42012 313788 42076 313792
rect 41644 312972 41708 313036
rect 42196 312352 42260 312356
rect 42196 312296 42210 312352
rect 42210 312296 42260 312352
rect 42196 312292 42260 312296
rect 41828 297604 41892 297668
rect 41828 296788 41892 296852
rect 41828 295972 41892 296036
rect 41828 295564 41892 295628
rect 42012 294340 42076 294404
rect 41828 272368 41892 272372
rect 41828 272312 41842 272368
rect 41842 272312 41892 272368
rect 41828 272308 41892 272312
rect 41460 270404 41524 270468
rect 42012 269784 42076 269788
rect 42012 269728 42026 269784
rect 42026 269728 42076 269784
rect 42012 269724 42076 269728
rect 41644 269316 41708 269380
rect 676076 265236 676140 265300
rect 39988 255444 40052 255508
rect 676076 250140 676140 250204
rect 675156 246256 675220 246260
rect 675156 246200 675206 246256
rect 675206 246200 675220 246256
rect 675156 246196 675220 246200
rect 43852 242252 43916 242316
rect 44036 242116 44100 242180
rect 43668 238036 43732 238100
rect 43852 228788 43916 228852
rect 44036 228652 44100 228716
rect 43668 225660 43732 225724
rect 675156 220628 675220 220692
rect 39988 213012 40052 213076
rect 41460 201316 41524 201380
rect 41644 200228 41708 200292
rect 41828 200092 41892 200156
rect 41828 184240 41892 184244
rect 41828 184184 41878 184240
rect 41878 184184 41892 184240
rect 41828 184180 41892 184184
rect 41460 183364 41524 183428
rect 41644 182956 41708 183020
rect 675892 171124 675956 171188
rect 675892 156980 675956 157044
rect 580948 110468 581012 110532
rect 633204 95916 633268 95980
rect 662092 95508 662156 95572
rect 662092 88768 662156 88772
rect 662092 88712 662142 88768
rect 662142 88712 662156 88768
rect 662092 88708 662156 88712
rect 633204 80140 633268 80204
rect 626764 75516 626828 75580
rect 633204 75516 633268 75580
rect 576164 69396 576228 69460
rect 580948 68716 581012 68780
rect 626764 52396 626828 52460
rect 633204 51036 633268 51100
rect 590700 49676 590764 49740
rect 521700 48180 521764 48244
rect 521700 42120 521764 42124
rect 521700 42064 521750 42120
rect 521750 42064 521764 42120
rect 521700 42060 521764 42064
rect 307340 41848 307404 41852
rect 307340 41792 307354 41848
rect 307354 41792 307404 41848
rect 307340 41788 307404 41792
rect 416820 41848 416884 41852
rect 416820 41792 416834 41848
rect 416834 41792 416884 41848
rect 416820 41788 416884 41792
<< metal4 >>
rect 674419 895524 674485 895525
rect 674419 895460 674420 895524
rect 674484 895460 674485 895524
rect 674419 895459 674485 895460
rect 673867 893892 673933 893893
rect 673867 893828 673868 893892
rect 673932 893828 673933 893892
rect 673867 893827 673933 893828
rect 41827 809164 41893 809165
rect 41827 809100 41828 809164
rect 41892 809100 41893 809164
rect 41827 809099 41893 809100
rect 41830 794477 41890 809099
rect 41827 794476 41893 794477
rect 41827 794412 41828 794476
rect 41892 794412 41893 794476
rect 41827 794411 41893 794412
rect 42011 757076 42077 757077
rect 42011 757012 42012 757076
rect 42076 757012 42077 757076
rect 42011 757011 42077 757012
rect 42747 757076 42813 757077
rect 42747 757012 42748 757076
rect 42812 757012 42813 757076
rect 42747 757011 42813 757012
rect 42014 748781 42074 757011
rect 42750 752997 42810 757011
rect 42747 752996 42813 752997
rect 42747 752932 42748 752996
rect 42812 752932 42813 752996
rect 42747 752931 42813 752932
rect 42011 748780 42077 748781
rect 42011 748716 42012 748780
rect 42076 748716 42077 748780
rect 42011 748715 42077 748716
rect 673499 739668 673565 739669
rect 673499 739604 673500 739668
rect 673564 739604 673565 739668
rect 673499 739603 673565 739604
rect 43115 714372 43181 714373
rect 43115 714308 43116 714372
rect 43180 714308 43181 714372
rect 43115 714307 43181 714308
rect 43118 711517 43178 714307
rect 43667 714236 43733 714237
rect 43667 714172 43668 714236
rect 43732 714172 43733 714236
rect 43667 714171 43733 714172
rect 43115 711516 43181 711517
rect 43115 711452 43116 711516
rect 43180 711452 43181 711516
rect 43115 711451 43181 711452
rect 42747 709476 42813 709477
rect 42747 709412 42748 709476
rect 42812 709412 42813 709476
rect 42747 709411 42813 709412
rect 42750 708933 42810 709411
rect 42747 708932 42813 708933
rect 42747 708868 42748 708932
rect 42812 708868 42813 708932
rect 42747 708867 42813 708868
rect 43670 708525 43730 714171
rect 43667 708524 43733 708525
rect 43667 708460 43668 708524
rect 43732 708460 43733 708524
rect 43667 708459 43733 708460
rect 41459 677788 41525 677789
rect 41459 677724 41460 677788
rect 41524 677724 41525 677788
rect 41459 677723 41525 677724
rect 41462 676973 41522 677723
rect 41459 676972 41525 676973
rect 41459 676908 41460 676972
rect 41524 676908 41525 676972
rect 41459 676907 41525 676908
rect 43299 671124 43365 671125
rect 43299 671060 43300 671124
rect 43364 671060 43365 671124
rect 43299 671059 43365 671060
rect 42931 670716 42997 670717
rect 42931 670652 42932 670716
rect 42996 670652 42997 670716
rect 42931 670651 42997 670652
rect 42934 670581 42994 670651
rect 42931 670580 42997 670581
rect 42931 670516 42932 670580
rect 42996 670516 42997 670580
rect 42931 670515 42997 670516
rect 43302 670445 43362 671059
rect 43851 670580 43917 670581
rect 43851 670516 43852 670580
rect 43916 670516 43917 670580
rect 43851 670515 43917 670516
rect 43299 670444 43365 670445
rect 43299 670380 43300 670444
rect 43364 670380 43365 670444
rect 43299 670379 43365 670380
rect 43854 665277 43914 670515
rect 43851 665276 43917 665277
rect 43851 665212 43852 665276
rect 43916 665212 43917 665276
rect 43851 665211 43917 665212
rect 673502 664053 673562 739603
rect 673870 728670 673930 893827
rect 674051 786860 674117 786861
rect 674051 786796 674052 786860
rect 674116 786796 674117 786860
rect 674051 786795 674117 786796
rect 673686 728610 673930 728670
rect 673686 713693 673746 728610
rect 674054 724709 674114 786795
rect 674235 740348 674301 740349
rect 674235 740284 674236 740348
rect 674300 740284 674301 740348
rect 674235 740283 674301 740284
rect 674051 724708 674117 724709
rect 674051 724644 674052 724708
rect 674116 724644 674117 724708
rect 674051 724643 674117 724644
rect 674051 724300 674117 724301
rect 674051 724236 674052 724300
rect 674116 724236 674117 724300
rect 674051 724235 674117 724236
rect 673867 724164 673933 724165
rect 673867 724100 673868 724164
rect 673932 724100 673933 724164
rect 673867 724099 673933 724100
rect 673683 713692 673749 713693
rect 673683 713628 673684 713692
rect 673748 713628 673749 713692
rect 673683 713627 673749 713628
rect 673870 709613 673930 724099
rect 674054 715325 674114 724235
rect 674051 715324 674117 715325
rect 674051 715260 674052 715324
rect 674116 715260 674117 715324
rect 674051 715259 674117 715260
rect 673867 709612 673933 709613
rect 673867 709548 673868 709612
rect 673932 709548 673933 709612
rect 673867 709547 673933 709548
rect 673867 698188 673933 698189
rect 673867 698124 673868 698188
rect 673932 698124 673933 698188
rect 673867 698123 673933 698124
rect 673683 690572 673749 690573
rect 673683 690508 673684 690572
rect 673748 690508 673749 690572
rect 673683 690507 673749 690508
rect 673499 664052 673565 664053
rect 673499 663988 673500 664052
rect 673564 663988 673565 664052
rect 673499 663987 673565 663988
rect 673499 648684 673565 648685
rect 673499 648620 673500 648684
rect 673564 648620 673565 648684
rect 673499 648619 673565 648620
rect 41827 627468 41893 627469
rect 41827 627404 41828 627468
rect 41892 627404 41893 627468
rect 41827 627403 41893 627404
rect 42379 627468 42445 627469
rect 42379 627404 42380 627468
rect 42444 627404 42445 627468
rect 42379 627403 42445 627404
rect 41830 621485 41890 627403
rect 42382 622029 42442 627403
rect 42379 622028 42445 622029
rect 42379 621964 42380 622028
rect 42444 621964 42445 622028
rect 42379 621963 42445 621964
rect 41827 621484 41893 621485
rect 41827 621420 41828 621484
rect 41892 621420 41893 621484
rect 41827 621419 41893 621420
rect 42195 585308 42261 585309
rect 42195 585244 42196 585308
rect 42260 585244 42261 585308
rect 42195 585243 42261 585244
rect 41827 584220 41893 584221
rect 41827 584156 41828 584220
rect 41892 584156 41893 584220
rect 41827 584155 41893 584156
rect 41830 580685 41890 584155
rect 41827 580684 41893 580685
rect 41827 580620 41828 580684
rect 41892 580620 41893 580684
rect 41827 580619 41893 580620
rect 42198 577013 42258 585243
rect 42931 583948 42997 583949
rect 42931 583884 42932 583948
rect 42996 583884 42997 583948
rect 42931 583883 42997 583884
rect 42934 581909 42994 583883
rect 42931 581908 42997 581909
rect 42931 581844 42932 581908
rect 42996 581844 42997 581908
rect 42931 581843 42997 581844
rect 42195 577012 42261 577013
rect 42195 576948 42196 577012
rect 42260 576948 42261 577012
rect 42195 576947 42261 576948
rect 673502 573341 673562 648619
rect 673686 620261 673746 690507
rect 673870 640253 673930 698123
rect 674051 694380 674117 694381
rect 674051 694316 674052 694380
rect 674116 694316 674117 694380
rect 674051 694315 674117 694316
rect 673867 640252 673933 640253
rect 673867 640188 673868 640252
rect 673932 640188 673933 640252
rect 673867 640187 673933 640188
rect 673683 620260 673749 620261
rect 673683 620196 673684 620260
rect 673748 620196 673749 620260
rect 673683 620195 673749 620196
rect 674054 619037 674114 694315
rect 674238 681189 674298 740283
rect 674422 724301 674482 895459
rect 679203 886684 679269 886685
rect 679203 886620 679204 886684
rect 679268 886620 679269 886684
rect 679203 886619 679269 886620
rect 679206 885869 679266 886619
rect 679203 885868 679269 885869
rect 679203 885804 679204 885868
rect 679268 885804 679269 885868
rect 679203 885803 679269 885804
rect 679206 885053 679266 885803
rect 679203 885052 679269 885053
rect 679203 884988 679204 885052
rect 679268 884988 679269 885052
rect 679203 884987 679269 884988
rect 674971 788356 675037 788357
rect 674971 788292 674972 788356
rect 675036 788292 675037 788356
rect 674971 788291 675037 788292
rect 674603 740212 674669 740213
rect 674603 740148 674604 740212
rect 674668 740148 674669 740212
rect 674603 740147 674669 740148
rect 674419 724300 674485 724301
rect 674419 724236 674420 724300
rect 674484 724236 674485 724300
rect 674419 724235 674485 724236
rect 674419 724028 674485 724029
rect 674419 723964 674420 724028
rect 674484 723964 674485 724028
rect 674419 723963 674485 723964
rect 674422 711245 674482 723963
rect 674419 711244 674485 711245
rect 674419 711180 674420 711244
rect 674484 711180 674485 711244
rect 674419 711179 674485 711180
rect 674419 690164 674485 690165
rect 674419 690100 674420 690164
rect 674484 690100 674485 690164
rect 674419 690099 674485 690100
rect 674235 681188 674301 681189
rect 674235 681124 674236 681188
rect 674300 681124 674301 681188
rect 674235 681123 674301 681124
rect 674235 680372 674301 680373
rect 674235 680308 674236 680372
rect 674300 680308 674301 680372
rect 674235 680307 674301 680308
rect 674238 674661 674298 680307
rect 674235 674660 674301 674661
rect 674235 674596 674236 674660
rect 674300 674596 674301 674660
rect 674235 674595 674301 674596
rect 674235 674116 674301 674117
rect 674235 674052 674236 674116
rect 674300 674052 674301 674116
rect 674235 674051 674301 674052
rect 674238 666909 674298 674051
rect 674235 666908 674301 666909
rect 674235 666844 674236 666908
rect 674300 666844 674301 666908
rect 674235 666843 674301 666844
rect 674422 632070 674482 690099
rect 674606 680373 674666 740147
rect 674787 738716 674853 738717
rect 674787 738652 674788 738716
rect 674852 738652 674853 738716
rect 674787 738651 674853 738652
rect 674603 680372 674669 680373
rect 674603 680308 674604 680372
rect 674668 680308 674669 680372
rect 674603 680307 674669 680308
rect 674603 680236 674669 680237
rect 674603 680172 674604 680236
rect 674668 680172 674669 680236
rect 674603 680171 674669 680172
rect 674606 674797 674666 680171
rect 674603 674796 674669 674797
rect 674603 674732 674604 674796
rect 674668 674732 674669 674796
rect 674603 674731 674669 674732
rect 674603 674660 674669 674661
rect 674603 674596 674604 674660
rect 674668 674596 674669 674660
rect 674603 674595 674669 674596
rect 674606 665685 674666 674595
rect 674603 665684 674669 665685
rect 674603 665620 674604 665684
rect 674668 665620 674669 665684
rect 674603 665619 674669 665620
rect 674790 663645 674850 738651
rect 674974 724029 675034 788291
rect 675155 787132 675221 787133
rect 675155 787068 675156 787132
rect 675220 787068 675221 787132
rect 675155 787067 675221 787068
rect 675158 724165 675218 787067
rect 675339 742932 675405 742933
rect 675339 742868 675340 742932
rect 675404 742868 675405 742932
rect 675339 742867 675405 742868
rect 675155 724164 675221 724165
rect 675155 724100 675156 724164
rect 675220 724100 675221 724164
rect 675155 724099 675221 724100
rect 674971 724028 675037 724029
rect 674971 723964 674972 724028
rect 675036 723964 675037 724028
rect 674971 723963 675037 723964
rect 675342 723890 675402 742867
rect 676647 742796 676713 742797
rect 676647 742732 676648 742796
rect 676712 742732 676713 742796
rect 676647 742731 676713 742732
rect 675707 742524 675773 742525
rect 675707 742460 675708 742524
rect 675772 742460 675773 742524
rect 675707 742459 675773 742460
rect 675523 729060 675589 729061
rect 675523 728996 675524 729060
rect 675588 728996 675589 729060
rect 675523 728995 675589 728996
rect 675526 728245 675586 728995
rect 675523 728244 675589 728245
rect 675523 728180 675524 728244
rect 675588 728180 675589 728244
rect 675523 728179 675589 728180
rect 674974 723830 675402 723890
rect 674974 701070 675034 723830
rect 675710 723210 675770 742459
rect 675158 723150 675770 723210
rect 675158 720390 675218 723150
rect 675891 721580 675957 721581
rect 675891 721516 675892 721580
rect 675956 721516 675957 721580
rect 675891 721515 675957 721516
rect 675158 720330 675770 720390
rect 674974 701010 675402 701070
rect 675342 680237 675402 701010
rect 675710 690030 675770 720330
rect 675894 712061 675954 721515
rect 675891 712060 675957 712061
rect 675891 711996 675892 712060
rect 675956 711996 675957 712060
rect 675891 711995 675957 711996
rect 676650 710290 676710 742731
rect 676811 742660 676877 742661
rect 676811 742596 676812 742660
rect 676876 742596 676877 742660
rect 676811 742595 676877 742596
rect 676814 712058 676874 742595
rect 677179 738036 677245 738037
rect 677179 737972 677180 738036
rect 677244 737972 677245 738036
rect 677179 737971 677245 737972
rect 677182 728670 677242 737971
rect 677182 728610 677426 728670
rect 676814 711998 677058 712058
rect 675894 710230 676710 710290
rect 675894 706757 675954 710230
rect 676998 709610 677058 711998
rect 676262 709550 677058 709610
rect 676075 707300 676141 707301
rect 676075 707236 676076 707300
rect 676140 707298 676141 707300
rect 676262 707298 676322 709550
rect 676140 707238 676322 707298
rect 676140 707236 676141 707238
rect 676075 707235 676141 707236
rect 675891 706756 675957 706757
rect 675891 706692 675892 706756
rect 675956 706692 675957 706756
rect 675891 706691 675957 706692
rect 676995 699684 677061 699685
rect 676995 699620 676996 699684
rect 677060 699620 677061 699684
rect 676995 699619 677061 699620
rect 676075 697236 676141 697237
rect 676075 697172 676076 697236
rect 676140 697172 676141 697236
rect 676075 697171 676141 697172
rect 675891 694788 675957 694789
rect 675891 694724 675892 694788
rect 675956 694724 675957 694788
rect 675891 694723 675957 694724
rect 675526 689970 675770 690030
rect 675339 680236 675405 680237
rect 675339 680172 675340 680236
rect 675404 680172 675405 680236
rect 675339 680171 675405 680172
rect 675526 679010 675586 689970
rect 674974 678950 675586 679010
rect 674974 675610 675034 678950
rect 675894 678469 675954 694723
rect 675891 678468 675957 678469
rect 675891 678404 675892 678468
rect 675956 678404 675957 678468
rect 675891 678403 675957 678404
rect 676078 678330 676138 697171
rect 676811 696692 676877 696693
rect 676811 696628 676812 696692
rect 676876 696628 676877 696692
rect 676811 696627 676877 696628
rect 676647 693564 676713 693565
rect 676647 693500 676648 693564
rect 676712 693500 676713 693564
rect 676647 693499 676713 693500
rect 675158 678270 676138 678330
rect 675158 676290 675218 678270
rect 675158 676230 676138 676290
rect 674974 675550 675770 675610
rect 675339 674796 675405 674797
rect 675339 674732 675340 674796
rect 675404 674732 675405 674796
rect 675339 674731 675405 674732
rect 675342 666093 675402 674731
rect 675339 666092 675405 666093
rect 675339 666028 675340 666092
rect 675404 666028 675405 666092
rect 675339 666027 675405 666028
rect 675710 664461 675770 675550
rect 675891 674796 675957 674797
rect 675891 674732 675892 674796
rect 675956 674732 675957 674796
rect 675891 674731 675957 674732
rect 675707 664460 675773 664461
rect 675707 664396 675708 664460
rect 675772 664396 675773 664460
rect 675707 664395 675773 664396
rect 674787 663644 674853 663645
rect 674787 663580 674788 663644
rect 674852 663580 674853 663644
rect 674787 663579 674853 663580
rect 675707 652628 675773 652629
rect 675707 652564 675708 652628
rect 675772 652564 675773 652628
rect 675707 652563 675773 652564
rect 675155 652220 675221 652221
rect 675155 652156 675156 652220
rect 675220 652156 675221 652220
rect 675155 652155 675221 652156
rect 674971 648956 675037 648957
rect 674971 648892 674972 648956
rect 675036 648892 675037 648956
rect 674971 648891 675037 648892
rect 674787 641748 674853 641749
rect 674787 641684 674788 641748
rect 674852 641684 674853 641748
rect 674787 641683 674853 641684
rect 674603 641612 674669 641613
rect 674603 641548 674604 641612
rect 674668 641548 674669 641612
rect 674603 641547 674669 641548
rect 674238 632010 674482 632070
rect 674051 619036 674117 619037
rect 674051 618972 674052 619036
rect 674116 618972 674117 619036
rect 674051 618971 674117 618972
rect 674238 616997 674298 632010
rect 674606 630730 674666 641547
rect 674422 630670 674666 630730
rect 674422 620669 674482 630670
rect 674790 630050 674850 641683
rect 674606 629990 674850 630050
rect 674419 620668 674485 620669
rect 674419 620604 674420 620668
rect 674484 620604 674485 620668
rect 674419 620603 674485 620604
rect 674606 619445 674666 629990
rect 674787 629372 674853 629373
rect 674787 629308 674788 629372
rect 674852 629308 674853 629372
rect 674787 629307 674853 629308
rect 674603 619444 674669 619445
rect 674603 619380 674604 619444
rect 674668 619380 674669 619444
rect 674603 619379 674669 619380
rect 674235 616996 674301 616997
rect 674235 616932 674236 616996
rect 674300 616932 674301 616996
rect 674235 616931 674301 616932
rect 673683 607884 673749 607885
rect 673683 607820 673684 607884
rect 673748 607820 673749 607884
rect 673683 607819 673749 607820
rect 673499 573340 673565 573341
rect 673499 573276 673500 573340
rect 673564 573276 673565 573340
rect 673499 573275 673565 573276
rect 41643 556748 41709 556749
rect 41643 556684 41644 556748
rect 41708 556684 41709 556748
rect 41643 556683 41709 556684
rect 39987 554300 40053 554301
rect 39987 554236 39988 554300
rect 40052 554236 40053 554300
rect 39987 554235 40053 554236
rect 39990 435981 40050 554235
rect 41459 551036 41525 551037
rect 41459 550972 41460 551036
rect 41524 550972 41525 551036
rect 41459 550971 41525 550972
rect 41462 535397 41522 550971
rect 41646 538525 41706 556683
rect 42379 556068 42445 556069
rect 42379 556004 42380 556068
rect 42444 556004 42445 556068
rect 42379 556003 42445 556004
rect 42195 552804 42261 552805
rect 42195 552740 42196 552804
rect 42260 552740 42261 552804
rect 42195 552739 42261 552740
rect 41827 551580 41893 551581
rect 41827 551516 41828 551580
rect 41892 551516 41893 551580
rect 41827 551515 41893 551516
rect 41643 538524 41709 538525
rect 41643 538460 41644 538524
rect 41708 538460 41709 538524
rect 41643 538459 41709 538460
rect 41459 535396 41525 535397
rect 41459 535332 41460 535396
rect 41524 535332 41525 535396
rect 41459 535331 41525 535332
rect 41830 532677 41890 551515
rect 42011 550764 42077 550765
rect 42011 550700 42012 550764
rect 42076 550700 42077 550764
rect 42011 550699 42077 550700
rect 42014 538117 42074 550699
rect 42011 538116 42077 538117
rect 42011 538052 42012 538116
rect 42076 538052 42077 538116
rect 42011 538051 42077 538052
rect 42198 532813 42258 552739
rect 42382 538253 42442 556003
rect 44035 555252 44101 555253
rect 44035 555188 44036 555252
rect 44100 555188 44101 555252
rect 44035 555187 44101 555188
rect 42563 554028 42629 554029
rect 42563 553964 42564 554028
rect 42628 553964 42629 554028
rect 42563 553963 42629 553964
rect 42379 538252 42445 538253
rect 42379 538188 42380 538252
rect 42444 538188 42445 538252
rect 42379 538187 42445 538188
rect 42566 535397 42626 553963
rect 42747 553212 42813 553213
rect 42747 553148 42748 553212
rect 42812 553148 42813 553212
rect 42747 553147 42813 553148
rect 42563 535396 42629 535397
rect 42563 535332 42564 535396
rect 42628 535332 42629 535396
rect 42563 535331 42629 535332
rect 42195 532812 42261 532813
rect 42195 532748 42196 532812
rect 42260 532748 42261 532812
rect 42195 532747 42261 532748
rect 42750 532677 42810 553147
rect 42931 552396 42997 552397
rect 42931 552332 42932 552396
rect 42996 552332 42997 552396
rect 42931 552331 42997 552332
rect 42934 538389 42994 552331
rect 42931 538388 42997 538389
rect 42931 538324 42932 538388
rect 42996 538324 42997 538388
rect 42931 538323 42997 538324
rect 41827 532676 41893 532677
rect 41827 532612 41828 532676
rect 41892 532612 41893 532676
rect 41827 532611 41893 532612
rect 42747 532676 42813 532677
rect 42747 532612 42748 532676
rect 42812 532612 42813 532676
rect 42747 532611 42813 532612
rect 44038 455970 44098 555187
rect 673686 546510 673746 607819
rect 674235 605028 674301 605029
rect 674235 604964 674236 605028
rect 674300 604964 674301 605028
rect 674235 604963 674301 604964
rect 673867 601900 673933 601901
rect 673867 601836 673868 601900
rect 673932 601836 673933 601900
rect 673867 601835 673933 601836
rect 673502 546450 673746 546510
rect 673502 531045 673562 546450
rect 673683 543148 673749 543149
rect 673683 543084 673684 543148
rect 673748 543084 673749 543148
rect 673683 543083 673749 543084
rect 673499 531044 673565 531045
rect 673499 530980 673500 531044
rect 673564 530980 673565 531044
rect 673499 530979 673565 530980
rect 673686 528597 673746 543083
rect 673683 528596 673749 528597
rect 673683 528532 673684 528596
rect 673748 528532 673749 528596
rect 673683 528531 673749 528532
rect 673870 527101 673930 601835
rect 674051 588028 674117 588029
rect 674051 587964 674052 588028
rect 674116 587964 674117 588028
rect 674051 587963 674117 587964
rect 674054 574157 674114 587963
rect 674051 574156 674117 574157
rect 674051 574092 674052 574156
rect 674116 574092 674117 574156
rect 674051 574091 674117 574092
rect 674051 562324 674117 562325
rect 674051 562260 674052 562324
rect 674116 562260 674117 562324
rect 674051 562259 674117 562260
rect 673867 527100 673933 527101
rect 673867 527036 673868 527100
rect 673932 527036 673933 527100
rect 673867 527035 673933 527036
rect 674054 485213 674114 562259
rect 674238 530637 674298 604963
rect 674603 604484 674669 604485
rect 674603 604420 674604 604484
rect 674668 604420 674669 604484
rect 674603 604419 674669 604420
rect 674419 603804 674485 603805
rect 674419 603740 674420 603804
rect 674484 603740 674485 603804
rect 674419 603739 674485 603740
rect 674422 543149 674482 603739
rect 674419 543148 674485 543149
rect 674419 543084 674420 543148
rect 674484 543084 674485 543148
rect 674419 543083 674485 543084
rect 674606 543010 674666 604419
rect 674790 576605 674850 629307
rect 674787 576604 674853 576605
rect 674787 576540 674788 576604
rect 674852 576540 674853 576604
rect 674787 576539 674853 576540
rect 674974 573749 675034 648891
rect 675158 588029 675218 652155
rect 675339 651676 675405 651677
rect 675339 651612 675340 651676
rect 675404 651612 675405 651676
rect 675339 651611 675405 651612
rect 675342 637669 675402 651611
rect 675710 638213 675770 652563
rect 675894 641613 675954 674731
rect 676078 641749 676138 676230
rect 676075 641748 676141 641749
rect 676075 641684 676076 641748
rect 676140 641684 676141 641748
rect 676075 641683 676141 641684
rect 675891 641612 675957 641613
rect 675891 641548 675892 641612
rect 675956 641548 675957 641612
rect 675891 641547 675957 641548
rect 675707 638212 675773 638213
rect 675707 638148 675708 638212
rect 675772 638148 675773 638212
rect 675707 638147 675773 638148
rect 675339 637668 675405 637669
rect 675339 637604 675340 637668
rect 675404 637604 675405 637668
rect 675339 637603 675405 637604
rect 676650 618765 676710 693499
rect 676814 622029 676874 696627
rect 676998 662149 677058 699619
rect 677179 693020 677245 693021
rect 677179 692956 677180 693020
rect 677244 692956 677245 693020
rect 677179 692955 677245 692956
rect 676995 662148 677061 662149
rect 676995 662084 676996 662148
rect 677060 662084 677061 662148
rect 676995 662083 677061 662084
rect 676811 622028 676877 622029
rect 676811 621964 676812 622028
rect 676876 621964 676877 622028
rect 676811 621963 676877 621964
rect 676647 618764 676713 618765
rect 676647 618700 676648 618764
rect 676712 618700 676713 618764
rect 676647 618699 676713 618700
rect 677182 617541 677242 692955
rect 677366 662557 677426 728610
rect 677363 662556 677429 662557
rect 677363 662492 677364 662556
rect 677428 662492 677429 662556
rect 677363 662491 677429 662492
rect 677547 622844 677613 622845
rect 677547 622780 677548 622844
rect 677612 622780 677613 622844
rect 677547 622779 677613 622780
rect 677179 617540 677245 617541
rect 677179 617476 677180 617540
rect 677244 617476 677245 617540
rect 677179 617475 677245 617476
rect 677363 617132 677429 617133
rect 677363 617068 677364 617132
rect 677428 617068 677429 617132
rect 677363 617067 677429 617068
rect 676667 609244 676733 609245
rect 676667 609180 676668 609244
rect 676732 609180 676733 609244
rect 676667 609179 676733 609180
rect 676075 607340 676141 607341
rect 676075 607276 676076 607340
rect 676140 607276 676141 607340
rect 676075 607275 676141 607276
rect 675339 604484 675405 604485
rect 675339 604420 675340 604484
rect 675404 604420 675405 604484
rect 675339 604419 675405 604420
rect 675155 588028 675221 588029
rect 675155 587964 675156 588028
rect 675220 587964 675221 588028
rect 675155 587963 675221 587964
rect 675342 587890 675402 604419
rect 675158 587830 675402 587890
rect 675158 574110 675218 587830
rect 676078 587757 676138 607275
rect 676075 587756 676141 587757
rect 676075 587692 676076 587756
rect 676140 587692 676141 587756
rect 676075 587691 676141 587692
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675158 574050 675402 574110
rect 674971 573748 675037 573749
rect 674971 573684 674972 573748
rect 675036 573684 675037 573748
rect 674971 573683 675037 573684
rect 675155 562460 675221 562461
rect 675155 562396 675156 562460
rect 675220 562396 675221 562460
rect 675155 562395 675221 562396
rect 674971 561236 675037 561237
rect 674971 561172 674972 561236
rect 675036 561172 675037 561236
rect 674971 561171 675037 561172
rect 674787 557564 674853 557565
rect 674787 557500 674788 557564
rect 674852 557500 674853 557564
rect 674787 557499 674853 557500
rect 674422 542950 674666 543010
rect 674422 531861 674482 542950
rect 674603 542740 674669 542741
rect 674603 542676 674604 542740
rect 674668 542676 674669 542740
rect 674603 542675 674669 542676
rect 674419 531860 674485 531861
rect 674419 531796 674420 531860
rect 674484 531796 674485 531860
rect 674419 531795 674485 531796
rect 674235 530636 674301 530637
rect 674235 530572 674236 530636
rect 674300 530572 674301 530636
rect 674235 530571 674301 530572
rect 674606 529005 674666 542675
rect 674603 529004 674669 529005
rect 674603 528940 674604 529004
rect 674668 528940 674669 529004
rect 674603 528939 674669 528940
rect 674051 485212 674117 485213
rect 674051 485148 674052 485212
rect 674116 485148 674117 485212
rect 674051 485147 674117 485148
rect 674790 484805 674850 557499
rect 674974 487661 675034 561171
rect 674971 487660 675037 487661
rect 674971 487596 674972 487660
rect 675036 487596 675037 487660
rect 674971 487595 675037 487596
rect 675158 486845 675218 562395
rect 675342 542741 675402 574050
rect 675523 553892 675589 553893
rect 675523 553828 675524 553892
rect 675588 553828 675589 553892
rect 675523 553827 675589 553828
rect 675526 548045 675586 553827
rect 675523 548044 675589 548045
rect 675523 547980 675524 548044
rect 675588 547980 675589 548044
rect 675523 547979 675589 547980
rect 676078 542741 676138 586195
rect 676670 571981 676730 609179
rect 676995 579324 677061 579325
rect 676995 579260 676996 579324
rect 677060 579260 677061 579324
rect 676995 579259 677061 579260
rect 676811 576876 676877 576877
rect 676811 576812 676812 576876
rect 676876 576812 676877 576876
rect 676811 576811 676877 576812
rect 676667 571980 676733 571981
rect 676667 571916 676668 571980
rect 676732 571916 676733 571980
rect 676667 571915 676733 571916
rect 676814 543965 676874 576811
rect 676811 543964 676877 543965
rect 676811 543900 676812 543964
rect 676876 543900 676877 543964
rect 676811 543899 676877 543900
rect 676998 543829 677058 579259
rect 677179 577692 677245 577693
rect 677179 577628 677180 577692
rect 677244 577628 677245 577692
rect 677179 577627 677245 577628
rect 677182 544101 677242 577627
rect 677366 571573 677426 617067
rect 677550 578509 677610 622779
rect 677547 578508 677613 578509
rect 677547 578444 677548 578508
rect 677612 578444 677613 578508
rect 677547 578443 677613 578444
rect 677363 571572 677429 571573
rect 677363 571508 677364 571572
rect 677428 571508 677429 571572
rect 677363 571507 677429 571508
rect 677179 544100 677245 544101
rect 677179 544036 677180 544100
rect 677244 544036 677245 544100
rect 677179 544035 677245 544036
rect 676995 543828 677061 543829
rect 676995 543764 676996 543828
rect 677060 543764 677061 543828
rect 676995 543763 677061 543764
rect 675339 542740 675405 542741
rect 675339 542676 675340 542740
rect 675404 542676 675405 542740
rect 675339 542675 675405 542676
rect 676075 542740 676141 542741
rect 676075 542676 676076 542740
rect 676140 542676 676141 542740
rect 676075 542675 676141 542676
rect 676075 541244 676141 541245
rect 676075 541180 676076 541244
rect 676140 541180 676141 541244
rect 676075 541179 676141 541180
rect 676078 529413 676138 541179
rect 676075 529412 676141 529413
rect 676075 529348 676076 529412
rect 676140 529348 676141 529412
rect 676075 529347 676141 529348
rect 675155 486844 675221 486845
rect 675155 486780 675156 486844
rect 675220 486780 675221 486844
rect 675155 486779 675221 486780
rect 674787 484804 674853 484805
rect 674787 484740 674788 484804
rect 674852 484740 674853 484804
rect 674787 484739 674853 484740
rect 44038 455910 44282 455970
rect 44222 450850 44282 455910
rect 44038 450790 44282 450850
rect 44038 445770 44098 450790
rect 44038 445710 44282 445770
rect 44222 440330 44282 445710
rect 44038 440270 44282 440330
rect 39987 435980 40053 435981
rect 39987 435916 39988 435980
rect 40052 435916 40053 435980
rect 39987 435915 40053 435916
rect 44038 428093 44098 440270
rect 44035 428092 44101 428093
rect 44035 428028 44036 428092
rect 44100 428028 44101 428092
rect 44035 428027 44101 428028
rect 43115 411500 43181 411501
rect 43115 411436 43116 411500
rect 43180 411436 43181 411500
rect 43115 411435 43181 411436
rect 43118 406877 43178 411435
rect 43115 406876 43181 406877
rect 43115 406812 43116 406876
rect 43180 406812 43181 406876
rect 43115 406811 43181 406812
rect 675155 400620 675221 400621
rect 675155 400556 675156 400620
rect 675220 400556 675221 400620
rect 675155 400555 675221 400556
rect 41643 383076 41709 383077
rect 41643 383012 41644 383076
rect 41708 383012 41709 383076
rect 41643 383011 41709 383012
rect 41459 382260 41525 382261
rect 41459 382196 41460 382260
rect 41524 382196 41525 382260
rect 41459 382195 41525 382196
rect 41462 355741 41522 382195
rect 41646 356965 41706 383011
rect 41643 356964 41709 356965
rect 41643 356900 41644 356964
rect 41708 356900 41709 356964
rect 41643 356899 41709 356900
rect 675158 355877 675218 400555
rect 675155 355876 675221 355877
rect 675155 355812 675156 355876
rect 675220 355812 675221 355876
rect 675155 355811 675221 355812
rect 41459 355740 41525 355741
rect 41459 355676 41460 355740
rect 41524 355676 41525 355740
rect 41459 355675 41525 355676
rect 41459 340236 41525 340237
rect 41459 340172 41460 340236
rect 41524 340172 41525 340236
rect 41459 340171 41525 340172
rect 41462 298210 41522 340171
rect 41643 337380 41709 337381
rect 41643 337316 41644 337380
rect 41708 337316 41709 337380
rect 41643 337315 41709 337316
rect 41646 313037 41706 337315
rect 41827 337244 41893 337245
rect 41827 337180 41828 337244
rect 41892 337180 41893 337244
rect 41827 337179 41893 337180
rect 41830 316301 41890 337179
rect 42563 336836 42629 336837
rect 42563 336772 42564 336836
rect 42628 336772 42629 336836
rect 42563 336771 42629 336772
rect 42195 330172 42261 330173
rect 42195 330108 42196 330172
rect 42260 330108 42261 330172
rect 42195 330107 42261 330108
rect 42011 330036 42077 330037
rect 42011 329972 42012 330036
rect 42076 329972 42077 330036
rect 42011 329971 42077 329972
rect 41827 316300 41893 316301
rect 41827 316236 41828 316300
rect 41892 316236 41893 316300
rect 41827 316235 41893 316236
rect 42014 313853 42074 329971
rect 42011 313852 42077 313853
rect 42011 313788 42012 313852
rect 42076 313788 42077 313852
rect 42011 313787 42077 313788
rect 41643 313036 41709 313037
rect 41643 312972 41644 313036
rect 41708 312972 41709 313036
rect 41643 312971 41709 312972
rect 42198 312357 42258 330107
rect 42379 329900 42445 329901
rect 42379 329836 42380 329900
rect 42444 329836 42445 329900
rect 42379 329835 42445 329836
rect 42382 315485 42442 329835
rect 42566 316437 42626 336771
rect 42563 316436 42629 316437
rect 42563 316372 42564 316436
rect 42628 316372 42629 316436
rect 42563 316371 42629 316372
rect 42379 315484 42445 315485
rect 42379 315420 42380 315484
rect 42444 315420 42445 315484
rect 42379 315419 42445 315420
rect 42195 312356 42261 312357
rect 42195 312292 42196 312356
rect 42260 312292 42261 312356
rect 42195 312291 42261 312292
rect 41462 298150 41890 298210
rect 41830 297669 41890 298150
rect 41827 297668 41893 297669
rect 41827 297604 41828 297668
rect 41892 297604 41893 297668
rect 41827 297603 41893 297604
rect 41827 296852 41893 296853
rect 41827 296850 41828 296852
rect 41462 296790 41828 296850
rect 41462 270469 41522 296790
rect 41827 296788 41828 296790
rect 41892 296788 41893 296852
rect 41827 296787 41893 296788
rect 41646 296110 41890 296170
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41646 269381 41706 296110
rect 41830 296037 41890 296110
rect 41827 296036 41893 296037
rect 41827 295972 41828 296036
rect 41892 295972 41893 296036
rect 41827 295971 41893 295972
rect 41827 295628 41893 295629
rect 41827 295564 41828 295628
rect 41892 295564 41893 295628
rect 41827 295563 41893 295564
rect 41830 272373 41890 295563
rect 42011 294404 42077 294405
rect 42011 294340 42012 294404
rect 42076 294340 42077 294404
rect 42011 294339 42077 294340
rect 41827 272372 41893 272373
rect 41827 272308 41828 272372
rect 41892 272308 41893 272372
rect 41827 272307 41893 272308
rect 42014 269789 42074 294339
rect 42011 269788 42077 269789
rect 42011 269724 42012 269788
rect 42076 269724 42077 269788
rect 42011 269723 42077 269724
rect 41643 269380 41709 269381
rect 41643 269316 41644 269380
rect 41708 269316 41709 269380
rect 41643 269315 41709 269316
rect 676075 265300 676141 265301
rect 676075 265236 676076 265300
rect 676140 265236 676141 265300
rect 676075 265235 676141 265236
rect 39987 255508 40053 255509
rect 39987 255444 39988 255508
rect 40052 255444 40053 255508
rect 39987 255443 40053 255444
rect 39990 213077 40050 255443
rect 676078 250205 676138 265235
rect 676075 250204 676141 250205
rect 676075 250140 676076 250204
rect 676140 250140 676141 250204
rect 676075 250139 676141 250140
rect 675155 246260 675221 246261
rect 675155 246196 675156 246260
rect 675220 246196 675221 246260
rect 675155 246195 675221 246196
rect 43851 242316 43917 242317
rect 43851 242252 43852 242316
rect 43916 242252 43917 242316
rect 43851 242251 43917 242252
rect 43667 238100 43733 238101
rect 43667 238036 43668 238100
rect 43732 238036 43733 238100
rect 43667 238035 43733 238036
rect 43670 225725 43730 238035
rect 43854 228853 43914 242251
rect 44035 242180 44101 242181
rect 44035 242116 44036 242180
rect 44100 242116 44101 242180
rect 44035 242115 44101 242116
rect 43851 228852 43917 228853
rect 43851 228788 43852 228852
rect 43916 228788 43917 228852
rect 43851 228787 43917 228788
rect 44038 228717 44098 242115
rect 44035 228716 44101 228717
rect 44035 228652 44036 228716
rect 44100 228652 44101 228716
rect 44035 228651 44101 228652
rect 43667 225724 43733 225725
rect 43667 225660 43668 225724
rect 43732 225660 43733 225724
rect 43667 225659 43733 225660
rect 675158 220693 675218 246195
rect 675155 220692 675221 220693
rect 675155 220628 675156 220692
rect 675220 220628 675221 220692
rect 675155 220627 675221 220628
rect 39987 213076 40053 213077
rect 39987 213012 39988 213076
rect 40052 213012 40053 213076
rect 39987 213011 40053 213012
rect 41459 201380 41525 201381
rect 41459 201316 41460 201380
rect 41524 201316 41525 201380
rect 41459 201315 41525 201316
rect 41462 183429 41522 201315
rect 41643 200292 41709 200293
rect 41643 200228 41644 200292
rect 41708 200228 41709 200292
rect 41643 200227 41709 200228
rect 41459 183428 41525 183429
rect 41459 183364 41460 183428
rect 41524 183364 41525 183428
rect 41459 183363 41525 183364
rect 41646 183021 41706 200227
rect 41827 200156 41893 200157
rect 41827 200092 41828 200156
rect 41892 200092 41893 200156
rect 41827 200091 41893 200092
rect 41830 184245 41890 200091
rect 41827 184244 41893 184245
rect 41827 184180 41828 184244
rect 41892 184180 41893 184244
rect 41827 184179 41893 184180
rect 41643 183020 41709 183021
rect 41643 182956 41644 183020
rect 41708 182956 41709 183020
rect 41643 182955 41709 182956
rect 675891 171188 675957 171189
rect 675891 171124 675892 171188
rect 675956 171124 675957 171188
rect 675891 171123 675957 171124
rect 675894 157045 675954 171123
rect 675891 157044 675957 157045
rect 675891 156980 675892 157044
rect 675956 156980 675957 157044
rect 675891 156979 675957 156980
rect 580947 110532 581013 110533
rect 580947 110468 580948 110532
rect 581012 110468 581013 110532
rect 580947 110467 581013 110468
rect 576163 69460 576229 69461
rect 576163 69396 576164 69460
rect 576228 69396 576229 69460
rect 576163 69395 576229 69396
rect 521699 48244 521765 48245
rect 521699 48180 521700 48244
rect 521764 48180 521765 48244
rect 521699 48179 521765 48180
rect 521702 42125 521762 48179
rect 521699 42124 521765 42125
rect 521699 42060 521700 42124
rect 521764 42060 521765 42124
rect 521699 42059 521765 42060
rect 307339 41852 307405 41853
rect 307339 41788 307340 41852
rect 307404 41788 307405 41852
rect 307339 41787 307405 41788
rect 416819 41852 416885 41853
rect 416819 41788 416820 41852
rect 416884 41788 416885 41852
rect 416819 41787 416885 41788
rect 307342 40578 307402 41787
rect 416822 41258 416882 41787
rect 576166 40578 576226 69395
rect 580950 68781 581010 110467
rect 633203 95980 633269 95981
rect 633203 95916 633204 95980
rect 633268 95916 633269 95980
rect 633203 95915 633269 95916
rect 633206 80205 633266 95915
rect 662091 95572 662157 95573
rect 662091 95508 662092 95572
rect 662156 95508 662157 95572
rect 662091 95507 662157 95508
rect 662094 88773 662154 95507
rect 662091 88772 662157 88773
rect 662091 88708 662092 88772
rect 662156 88708 662157 88772
rect 662091 88707 662157 88708
rect 633203 80204 633269 80205
rect 633203 80140 633204 80204
rect 633268 80140 633269 80204
rect 633203 80139 633269 80140
rect 626763 75580 626829 75581
rect 626763 75516 626764 75580
rect 626828 75516 626829 75580
rect 626763 75515 626829 75516
rect 633203 75580 633269 75581
rect 633203 75516 633204 75580
rect 633268 75516 633269 75580
rect 633203 75515 633269 75516
rect 580947 68780 581013 68781
rect 580947 68716 580948 68780
rect 581012 68716 581013 68780
rect 580947 68715 581013 68716
rect 626766 52461 626826 75515
rect 626763 52460 626829 52461
rect 626763 52396 626764 52460
rect 626828 52396 626829 52460
rect 626763 52395 626829 52396
rect 633206 51101 633266 75515
rect 633203 51100 633269 51101
rect 633203 51036 633204 51100
rect 633268 51036 633269 51100
rect 633203 51035 633269 51036
rect 590699 49740 590765 49741
rect 590699 49676 590700 49740
rect 590764 49676 590765 49740
rect 590699 49675 590765 49676
rect 590702 41258 590762 49675
<< via4 >>
rect 416734 41022 416970 41258
rect 590614 41022 590850 41258
rect 307254 40342 307490 40578
rect 576078 40342 576314 40578
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 284410 1018624 296578 1030788
rect 334810 1018624 346978 1030788
rect 386210 1018624 398378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 953022 710788 965190
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 416692 41258 590892 41300
rect 416692 41022 416734 41258
rect 416970 41022 590614 41258
rect 590850 41022 590892 41258
rect 416692 40980 590892 41022
rect 307212 40578 576356 40620
rect 307212 40342 307254 40578
rect 307490 40342 576078 40578
rect 576314 40342 576356 40578
rect 307212 40300 576356 40342
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use caravan_logo  caravan_logo_0
timestamp 1636751500
transform 1 0 255684 0 1 5594
box 2240 2560 37000 11520
use caravan_motto  caravan_motto_0
timestamp 1637698689
transform 1 0 -53810 0 1 -20
box 367960 10204 399802 14768
use caravan_power_routing  caravan_power_routing_0
timestamp 1650915033
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use caravan_signal_routing  caravan_signal_routing_0
timestamp 1649950523
transform 1 0 0 0 1 0
box 39764 415548 677806 997846
use caravel_clocking  clock_ctrl
timestamp 1638876627
transform 1 0 621684 0 1 63608
box -38 -48 20000 12000
use copyright_block_a  copyright_block_a_0
timestamp 1649951985
transform 1 0 149318 0 1 16066
box -262 -10162 35048 2764
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1650900217
transform -1 0 710203 0 1 121000
box 882 416 34000 13000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1650900217
transform -1 0 710203 0 1 166200
box 882 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1650900217
transform 1 0 7631 0 1 289000
box 882 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1650900217
transform 1 0 7631 0 1 245800
box 882 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1650900217
transform 1 0 7631 0 1 202600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1650900217
transform -1 0 710203 0 1 523800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1650900217
transform -1 0 710203 0 1 568800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1650900217
transform -1 0 710203 0 1 614000
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1650900217
transform -1 0 710203 0 1 659000
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1650900217
transform -1 0 710203 0 1 704200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1650900217
transform -1 0 710203 0 1 884800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1650900217
transform -1 0 710203 0 1 211200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1650900217
transform -1 0 710203 0 1 256400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1650900217
transform -1 0 710203 0 1 301400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1650900217
transform -1 0 710203 0 1 346400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1650900217
transform -1 0 710203 0 1 391600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1650900217
transform -1 0 710203 0 1 479800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1650900217
transform 1 0 7631 0 1 805400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1650900217
transform 1 0 7631 0 1 762200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1650900217
transform 1 0 7631 0 1 719000
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1650900217
transform 1 0 7631 0 1 675800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1650900217
transform 1 0 7631 0 1 632600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1650900217
transform 1 0 7631 0 1 589400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1650900217
transform 1 0 7631 0 1 546200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1650900217
transform 1 0 7631 0 1 418600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1650900217
transform 1 0 7631 0 1 375400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1650900217
transform 1 0 7631 0 1 332200
box 882 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0\[0\]
timestamp 1638587925
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_0\[1\]
timestamp 1638587925
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2\[0\]
timestamp 1638587925
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2\[1\]
timestamp 1638587925
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2\[2\]
timestamp 1638587925
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1638587925
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1638587925
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1638587925
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1638587925
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1638587925
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1638587925
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1638587925
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1638587925
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1638587925
transform -1 0 709467 0 1 897800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1638587925
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1638587925
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1638587925
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1638587925
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1638587925
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1638587925
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1638587925
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1638587925
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1638587925
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1638587925
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1638587925
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1638587925
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1638587925
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1638464048
transform 1 0 606434 0 1 100002
box 0 0 60046 110190
use mgmt_protect  mgmt_buffers
timestamp 1649962643
transform 1 0 192180 0 1 232036
box -400 -400 220400 32400
use user_analog_project_wrapper  mprj
timestamp 1632839657
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use open_source  open_source_0 hexdigits
timestamp 1638586442
transform 1 0 206080 0 1 1916
box 752 5164 29030 16242
use chip_io_alt  padframe
timestamp 1638975641
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use digital_pll  pll
timestamp 1638875307
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use simple_por  por
timestamp 1650914729
transform 1 0 650146 0 -1 55282
box -52 -62 11344 8684
use xres_buf  rstb_level
timestamp 1649268499
transform -1 0 145710 0 -1 50488
box 374 -400 3540 3800
use mgmt_core_wrapper  soc
timestamp 1638280046
transform 1 0 52034 0 1 53002
box 382 -400 524400 164400
use spare_logic_block  spare_logic\[0\]
timestamp 1638030917
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1638030917
transform 1 0 168632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1638030917
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1638030917
transform 1 0 428632 0 1 232528
box 0 0 9000 9000
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 96232 0 1 6528
box -656 1508 33720 10344
use user_id_programming  user_id_value
timestamp 1650371074
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 25000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 25000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 25000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 25000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 25000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 25000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 25000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 25000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 25000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 25000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 25000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698624 953022 710788 965190 0 FreeSans 25000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628410 1018624 640578 1030788 0 FreeSans 25000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526610 1018624 538778 1030788 0 FreeSans 25000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475210 1018624 487378 1030788 0 FreeSans 25000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386210 1018624 398378 1030788 0 FreeSans 25000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284410 1018624 296578 1030788 0 FreeSans 25000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 25000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 231810 1018624 243978 1030788 0 FreeSans 25000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181410 1018624 193578 1030788 0 FreeSans 25000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 130010 1018624 142178 1030788 0 FreeSans 25000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78610 1018624 90778 1030788 0 FreeSans 25000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6811 956610 18975 968778 0 FreeSans 25000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 25000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 25000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 25000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 25000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 25000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 25000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 25000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 25000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 25000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 25000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 25000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 25000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 25000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 25000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 25000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 25000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 25000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 25000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 25000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 25000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 25000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144149 18309 0 FreeSans 25000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 25000 0 0 0 vccd1
port 45 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 25000 0 0 0 vccd2
port 46 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 25000 0 0 0 vdda
port 47 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 25000 0 0 0 vdda1
port 48 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 25000 0 0 0 vdda1_2
port 49 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 25000 0 0 0 vdda2
port 50 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 25000 0 0 0 vddio_2
port 51 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 25000 0 0 0 vssa1
port 52 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 25000 0 0 0 vssa1_2
port 53 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 25000 0 0 0 vssa2
port 54 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 25000 0 0 0 vssd1
port 55 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 25000 0 0 0 vssd2
port 56 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 25000 0 0 0 vssio_2
port 57 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 25000 0 0 0 vddio
port 58 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 25000 0 0 0 vssio
port 59 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 25000 0 0 0 vssa
port 60 nsew signal bidirectional
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 25000 0 0 0 vccd
port 61 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 25000 0 0 0 vssd
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
