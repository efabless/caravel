magic
tech sky130A
magscale 1 2
timestamp 1666265755
<< metal1 >>
rect 132494 1001920 132500 1001972
rect 132552 1001960 132558 1001972
rect 133690 1001960 133696 1001972
rect 132552 1001932 133696 1001960
rect 132552 1001920 132558 1001932
rect 133690 1001920 133696 1001932
rect 133748 1001920 133754 1001972
rect 401686 992196 401692 992248
rect 401744 992236 401750 992248
rect 404354 992236 404360 992248
rect 401744 992208 404360 992236
rect 401744 992196 401750 992208
rect 404354 992196 404360 992208
rect 404412 992196 404418 992248
rect 396074 990836 396080 990888
rect 396132 990876 396138 990888
rect 400214 990876 400220 990888
rect 396132 990848 400220 990876
rect 396132 990836 396138 990848
rect 400214 990836 400220 990848
rect 400272 990836 400278 990888
rect 242250 989068 242256 989120
rect 242308 989108 242314 989120
rect 245654 989108 245660 989120
rect 242308 989080 245660 989108
rect 242308 989068 242314 989080
rect 245654 989068 245660 989080
rect 245712 989068 245718 989120
rect 293954 988184 293960 988236
rect 294012 988224 294018 988236
rect 298094 988224 298100 988236
rect 294012 988196 298100 988224
rect 294012 988184 294018 988196
rect 298094 988184 298100 988196
rect 298152 988184 298158 988236
rect 389174 987504 389180 987556
rect 389232 987544 389238 987556
rect 391934 987544 391940 987556
rect 389232 987516 391940 987544
rect 389232 987504 389238 987516
rect 391934 987504 391940 987516
rect 391992 987504 391998 987556
rect 399754 986348 399760 986400
rect 399812 986388 399818 986400
rect 401686 986388 401692 986400
rect 399812 986360 401692 986388
rect 399812 986348 399818 986360
rect 401686 986348 401692 986360
rect 401744 986348 401750 986400
rect 238662 985940 238668 985992
rect 238720 985980 238726 985992
rect 242250 985980 242256 985992
rect 238720 985952 242256 985980
rect 238720 985940 238726 985952
rect 242250 985940 242256 985952
rect 242308 985940 242314 985992
rect 289722 985396 289728 985448
rect 289780 985436 289786 985448
rect 293954 985436 293960 985448
rect 289780 985408 293960 985436
rect 289780 985396 289786 985408
rect 293954 985396 293960 985408
rect 294012 985396 294018 985448
rect 394418 983492 394424 983544
rect 394476 983532 394482 983544
rect 396074 983532 396080 983544
rect 394476 983504 396080 983532
rect 394476 983492 394482 983504
rect 396074 983492 396080 983504
rect 396132 983492 396138 983544
rect 483014 982472 483020 982524
rect 483072 982512 483078 982524
rect 483842 982512 483848 982524
rect 483072 982484 483848 982512
rect 483072 982472 483078 982484
rect 483842 982472 483848 982484
rect 483900 982472 483906 982524
rect 651374 959080 651380 959132
rect 651432 959120 651438 959132
rect 677410 959120 677416 959132
rect 651432 959092 677416 959120
rect 651432 959080 651438 959092
rect 677410 959080 677416 959092
rect 677468 959080 677474 959132
rect 30098 954932 30104 954984
rect 30156 954972 30162 954984
rect 63402 954972 63408 954984
rect 30156 954944 63408 954972
rect 30156 954932 30162 954944
rect 63402 954932 63408 954944
rect 63460 954932 63466 954984
rect 676030 897104 676036 897116
rect 663766 897076 676036 897104
rect 652018 896996 652024 897048
rect 652076 897036 652082 897048
rect 663766 897036 663794 897076
rect 676030 897064 676036 897076
rect 676088 897064 676094 897116
rect 652076 897008 663794 897036
rect 652076 896996 652082 897008
rect 654778 895772 654784 895824
rect 654836 895812 654842 895824
rect 675846 895812 675852 895824
rect 654836 895784 675852 895812
rect 654836 895772 654842 895784
rect 675846 895772 675852 895784
rect 675904 895772 675910 895824
rect 672718 895636 672724 895688
rect 672776 895676 672782 895688
rect 676030 895676 676036 895688
rect 672776 895648 676036 895676
rect 672776 895636 672782 895648
rect 676030 895636 676036 895648
rect 676088 895636 676094 895688
rect 671062 894412 671068 894464
rect 671120 894452 671126 894464
rect 675846 894452 675852 894464
rect 671120 894424 675852 894452
rect 671120 894412 671126 894424
rect 675846 894412 675852 894424
rect 675904 894412 675910 894464
rect 671890 894276 671896 894328
rect 671948 894316 671954 894328
rect 676030 894316 676036 894328
rect 671948 894288 676036 894316
rect 671948 894276 671954 894288
rect 676030 894276 676036 894288
rect 676088 894276 676094 894328
rect 672534 892984 672540 893036
rect 672592 893024 672598 893036
rect 675846 893024 675852 893036
rect 672592 892996 675852 893024
rect 672592 892984 672598 892996
rect 675846 892984 675852 892996
rect 675904 892984 675910 893036
rect 672074 892848 672080 892900
rect 672132 892888 672138 892900
rect 676030 892888 676036 892900
rect 672132 892860 676036 892888
rect 672132 892848 672138 892860
rect 676030 892848 676036 892860
rect 676088 892848 676094 892900
rect 674834 890332 674840 890384
rect 674892 890372 674898 890384
rect 676030 890372 676036 890384
rect 674892 890344 676036 890372
rect 674892 890332 674898 890344
rect 676030 890332 676036 890344
rect 676088 890332 676094 890384
rect 676214 890128 676220 890180
rect 676272 890168 676278 890180
rect 676858 890168 676864 890180
rect 676272 890140 676864 890168
rect 676272 890128 676278 890140
rect 676858 890128 676864 890140
rect 676916 890128 676922 890180
rect 674374 888904 674380 888956
rect 674432 888944 674438 888956
rect 676030 888944 676036 888956
rect 674432 888916 676036 888944
rect 674432 888904 674438 888916
rect 676030 888904 676036 888916
rect 676088 888904 676094 888956
rect 676214 888700 676220 888752
rect 676272 888740 676278 888752
rect 677042 888740 677048 888752
rect 676272 888712 677048 888740
rect 676272 888700 676278 888712
rect 677042 888700 677048 888712
rect 677100 888700 677106 888752
rect 674650 888496 674656 888548
rect 674708 888536 674714 888548
rect 676030 888536 676036 888548
rect 674708 888508 676036 888536
rect 674708 888496 674714 888508
rect 676030 888496 676036 888508
rect 676088 888496 676094 888548
rect 674190 887272 674196 887324
rect 674248 887312 674254 887324
rect 676030 887312 676036 887324
rect 674248 887284 676036 887312
rect 674248 887272 674254 887284
rect 676030 887272 676036 887284
rect 676088 887272 676094 887324
rect 670878 886864 670884 886916
rect 670936 886904 670942 886916
rect 676030 886904 676036 886916
rect 670936 886876 676036 886904
rect 670936 886864 670942 886876
rect 676030 886864 676036 886876
rect 676088 886864 676094 886916
rect 675846 886660 675852 886712
rect 675904 886700 675910 886712
rect 676398 886700 676404 886712
rect 675904 886672 676404 886700
rect 675904 886660 675910 886672
rect 676398 886660 676404 886672
rect 676456 886660 676462 886712
rect 673086 885640 673092 885692
rect 673144 885680 673150 885692
rect 676030 885680 676036 885692
rect 673144 885652 676036 885680
rect 673144 885640 673150 885652
rect 676030 885640 676036 885652
rect 676088 885640 676094 885692
rect 653398 880472 653404 880524
rect 653456 880512 653462 880524
rect 675478 880512 675484 880524
rect 653456 880484 675484 880512
rect 653456 880472 653462 880484
rect 675478 880472 675484 880484
rect 675536 880472 675542 880524
rect 676030 880200 676036 880252
rect 676088 880240 676094 880252
rect 679618 880240 679624 880252
rect 676088 880212 679624 880240
rect 676088 880200 676094 880212
rect 679618 880200 679624 880212
rect 679676 880200 679682 880252
rect 675018 879588 675024 879640
rect 675076 879628 675082 879640
rect 677042 879628 677048 879640
rect 675076 879600 677048 879628
rect 675076 879588 675082 879600
rect 677042 879588 677048 879600
rect 677100 879588 677106 879640
rect 675110 879384 675116 879436
rect 675168 879424 675174 879436
rect 676858 879424 676864 879436
rect 675168 879396 676864 879424
rect 675168 879384 675174 879396
rect 676858 879384 676864 879396
rect 676916 879384 676922 879436
rect 675662 879248 675668 879300
rect 675720 879288 675726 879300
rect 678238 879288 678244 879300
rect 675720 879260 678244 879288
rect 675720 879248 675726 879260
rect 678238 879248 678244 879260
rect 678296 879248 678302 879300
rect 675846 878472 675852 878484
rect 674944 878444 675852 878472
rect 674944 876772 674972 878444
rect 675846 878432 675852 878444
rect 675904 878432 675910 878484
rect 676030 878432 676036 878484
rect 676088 878432 676094 878484
rect 676048 878200 676076 878432
rect 675588 878172 676076 878200
rect 675588 877928 675616 878172
rect 675496 877900 675616 877928
rect 675496 877804 675524 877900
rect 675478 877752 675484 877804
rect 675536 877752 675542 877804
rect 675386 876772 675392 876784
rect 674944 876744 675392 876772
rect 675386 876732 675392 876744
rect 675444 876732 675450 876784
rect 657538 869388 657544 869440
rect 657596 869428 657602 869440
rect 675018 869428 675024 869440
rect 657596 869400 675024 869428
rect 657596 869388 657602 869400
rect 675018 869388 675024 869400
rect 675076 869388 675082 869440
rect 674834 869252 674840 869304
rect 674892 869292 674898 869304
rect 675294 869292 675300 869304
rect 674892 869264 675300 869292
rect 674892 869252 674898 869264
rect 675294 869252 675300 869264
rect 675352 869252 675358 869304
rect 651466 868844 651472 868896
rect 651524 868884 651530 868896
rect 654778 868884 654784 868896
rect 651524 868856 654784 868884
rect 651524 868844 651530 868856
rect 654778 868844 654784 868856
rect 654836 868844 654842 868896
rect 674190 868708 674196 868760
rect 674248 868748 674254 868760
rect 675294 868748 675300 868760
rect 674248 868720 675300 868748
rect 674248 868708 674254 868720
rect 675294 868708 675300 868720
rect 675352 868708 675358 868760
rect 654134 868028 654140 868080
rect 654192 868068 654198 868080
rect 675018 868068 675024 868080
rect 654192 868040 675024 868068
rect 654192 868028 654198 868040
rect 675018 868028 675024 868040
rect 675076 868028 675082 868080
rect 674834 867552 674840 867604
rect 674892 867592 674898 867604
rect 675202 867592 675208 867604
rect 674892 867564 675208 867592
rect 674892 867552 674898 867564
rect 675202 867552 675208 867564
rect 675260 867552 675266 867604
rect 651466 866600 651472 866652
rect 651524 866640 651530 866652
rect 672718 866640 672724 866652
rect 651524 866612 672724 866640
rect 651524 866600 651530 866612
rect 672718 866600 672724 866612
rect 672776 866600 672782 866652
rect 651374 865172 651380 865224
rect 651432 865212 651438 865224
rect 653398 865212 653404 865224
rect 651432 865184 653404 865212
rect 651432 865172 651438 865184
rect 653398 865172 653404 865184
rect 653456 865172 653462 865224
rect 651466 863812 651472 863864
rect 651524 863852 651530 863864
rect 657538 863852 657544 863864
rect 651524 863824 657544 863852
rect 651524 863812 651530 863824
rect 657538 863812 657544 863824
rect 657596 863812 657602 863864
rect 651466 862452 651472 862504
rect 651524 862492 651530 862504
rect 654134 862492 654140 862504
rect 651524 862464 654140 862492
rect 651524 862452 651530 862464
rect 654134 862452 654140 862464
rect 654192 862452 654198 862504
rect 35802 817096 35808 817148
rect 35860 817136 35866 817148
rect 46198 817136 46204 817148
rect 35860 817108 46204 817136
rect 35860 817096 35866 817108
rect 46198 817096 46204 817108
rect 46256 817096 46262 817148
rect 35618 816960 35624 817012
rect 35676 817000 35682 817012
rect 59998 817000 60004 817012
rect 35676 816972 60004 817000
rect 35676 816960 35682 816972
rect 59998 816960 60004 816972
rect 60056 816960 60062 817012
rect 35802 815736 35808 815788
rect 35860 815776 35866 815788
rect 42886 815776 42892 815788
rect 35860 815748 42892 815776
rect 35860 815736 35866 815748
rect 42886 815736 42892 815748
rect 42944 815736 42950 815788
rect 35434 815600 35440 815652
rect 35492 815640 35498 815652
rect 44174 815640 44180 815652
rect 35492 815612 44180 815640
rect 35492 815600 35498 815612
rect 44174 815600 44180 815612
rect 44232 815600 44238 815652
rect 35618 814376 35624 814428
rect 35676 814416 35682 814428
rect 43438 814416 43444 814428
rect 35676 814388 43444 814416
rect 35676 814376 35682 814388
rect 43438 814376 43444 814388
rect 43496 814376 43502 814428
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 45278 814280 45284 814292
rect 35860 814252 45284 814280
rect 35860 814240 35866 814252
rect 45278 814240 45284 814252
rect 45336 814240 45342 814292
rect 41322 812812 41328 812864
rect 41380 812852 41386 812864
rect 44542 812852 44548 812864
rect 41380 812824 44548 812852
rect 41380 812812 41386 812824
rect 44542 812812 44548 812824
rect 44600 812812 44606 812864
rect 41322 811452 41328 811504
rect 41380 811492 41386 811504
rect 43070 811492 43076 811504
rect 41380 811464 43076 811492
rect 41380 811452 41386 811464
rect 43070 811452 43076 811464
rect 43128 811452 43134 811504
rect 40954 810704 40960 810756
rect 41012 810744 41018 810756
rect 42702 810744 42708 810756
rect 41012 810716 42708 810744
rect 41012 810704 41018 810716
rect 42702 810704 42708 810716
rect 42760 810704 42766 810756
rect 44174 810704 44180 810756
rect 44232 810744 44238 810756
rect 62942 810744 62948 810756
rect 44232 810716 62948 810744
rect 44232 810704 44238 810716
rect 62942 810704 62948 810716
rect 63000 810704 63006 810756
rect 41322 808596 41328 808648
rect 41380 808636 41386 808648
rect 42242 808636 42248 808648
rect 41380 808608 42248 808636
rect 41380 808596 41386 808608
rect 42242 808596 42248 808608
rect 42300 808596 42306 808648
rect 41322 807440 41328 807492
rect 41380 807480 41386 807492
rect 43254 807480 43260 807492
rect 41380 807452 43260 807480
rect 41380 807440 41386 807452
rect 43254 807440 43260 807452
rect 43312 807440 43318 807492
rect 41138 807304 41144 807356
rect 41196 807344 41202 807356
rect 44358 807344 44364 807356
rect 41196 807316 44364 807344
rect 41196 807304 41202 807316
rect 44358 807304 44364 807316
rect 44416 807304 44422 807356
rect 41322 806080 41328 806132
rect 41380 806120 41386 806132
rect 50338 806120 50344 806132
rect 41380 806092 50344 806120
rect 41380 806080 41386 806092
rect 50338 806080 50344 806092
rect 50396 806080 50402 806132
rect 41138 805944 41144 805996
rect 41196 805984 41202 805996
rect 62666 805984 62672 805996
rect 41196 805956 62672 805984
rect 41196 805944 41202 805956
rect 62666 805944 62672 805956
rect 62724 805944 62730 805996
rect 34514 802408 34520 802460
rect 34572 802448 34578 802460
rect 41874 802448 41880 802460
rect 34572 802420 41880 802448
rect 34572 802408 34578 802420
rect 41874 802408 41880 802420
rect 41932 802408 41938 802460
rect 37918 801728 37924 801780
rect 37976 801768 37982 801780
rect 39758 801768 39764 801780
rect 37976 801740 39764 801768
rect 37976 801728 37982 801740
rect 39758 801728 39764 801740
rect 39816 801728 39822 801780
rect 31018 801048 31024 801100
rect 31076 801088 31082 801100
rect 42518 801088 42524 801100
rect 31076 801060 42524 801088
rect 31076 801048 31082 801060
rect 42518 801048 42524 801060
rect 42576 801048 42582 801100
rect 36538 800708 36544 800760
rect 36596 800748 36602 800760
rect 40494 800748 40500 800760
rect 36596 800720 40500 800748
rect 36596 800708 36602 800720
rect 40494 800708 40500 800720
rect 40552 800708 40558 800760
rect 42242 799280 42248 799332
rect 42300 799320 42306 799332
rect 42702 799320 42708 799332
rect 42300 799292 42708 799320
rect 42300 799280 42306 799292
rect 42702 799280 42708 799292
rect 42760 799280 42766 799332
rect 43622 799008 43628 799060
rect 43680 799048 43686 799060
rect 53098 799048 53104 799060
rect 43680 799020 53104 799048
rect 43680 799008 43686 799020
rect 53098 799008 53104 799020
rect 53156 799008 53162 799060
rect 43806 797648 43812 797700
rect 43864 797688 43870 797700
rect 57238 797688 57244 797700
rect 43864 797660 57244 797688
rect 43864 797648 43870 797660
rect 57238 797648 57244 797660
rect 57296 797648 57302 797700
rect 42242 795608 42248 795660
rect 42300 795648 42306 795660
rect 43806 795648 43812 795660
rect 42300 795620 43812 795648
rect 42300 795608 42306 795620
rect 43806 795608 43812 795620
rect 43864 795608 43870 795660
rect 42334 793908 42340 793960
rect 42392 793948 42398 793960
rect 44358 793948 44364 793960
rect 42392 793920 44364 793948
rect 42392 793908 42398 793920
rect 44358 793908 44364 793920
rect 44416 793908 44422 793960
rect 653398 790780 653404 790832
rect 653456 790820 653462 790832
rect 675386 790820 675392 790832
rect 653456 790792 675392 790820
rect 653456 790780 653462 790792
rect 675386 790780 675392 790792
rect 675444 790780 675450 790832
rect 53098 790712 53104 790764
rect 53156 790752 53162 790764
rect 62206 790752 62212 790764
rect 53156 790724 62212 790752
rect 53156 790712 53162 790724
rect 62206 790712 62212 790724
rect 62264 790712 62270 790764
rect 42610 789284 42616 789336
rect 42668 789324 42674 789336
rect 43070 789324 43076 789336
rect 42668 789296 43076 789324
rect 42668 789284 42674 789296
rect 43070 789284 43076 789296
rect 43128 789284 43134 789336
rect 57238 789148 57244 789200
rect 57296 789188 57302 789200
rect 62114 789188 62120 789200
rect 57296 789160 62120 789188
rect 57296 789148 57302 789160
rect 62114 789148 62120 789160
rect 62172 789148 62178 789200
rect 42702 786632 42708 786684
rect 42760 786672 42766 786684
rect 62114 786672 62120 786684
rect 42760 786644 62120 786672
rect 42760 786632 42766 786644
rect 62114 786632 62120 786644
rect 62172 786632 62178 786684
rect 59998 786496 60004 786548
rect 60056 786536 60062 786548
rect 62298 786536 62304 786548
rect 60056 786508 62304 786536
rect 60056 786496 60062 786508
rect 62298 786496 62304 786508
rect 62356 786496 62362 786548
rect 46198 785136 46204 785188
rect 46256 785176 46262 785188
rect 62114 785176 62120 785188
rect 46256 785148 62120 785176
rect 46256 785136 46262 785148
rect 62114 785136 62120 785148
rect 62172 785136 62178 785188
rect 670602 784252 670608 784304
rect 670660 784292 670666 784304
rect 675110 784292 675116 784304
rect 670660 784264 675116 784292
rect 670660 784252 670666 784264
rect 675110 784252 675116 784264
rect 675168 784252 675174 784304
rect 669222 784116 669228 784168
rect 669280 784156 669286 784168
rect 675386 784156 675392 784168
rect 669280 784128 675392 784156
rect 669280 784116 669286 784128
rect 675386 784116 675392 784128
rect 675444 784116 675450 784168
rect 673730 782620 673736 782672
rect 673788 782660 673794 782672
rect 675110 782660 675116 782672
rect 673788 782632 675116 782660
rect 673788 782620 673794 782632
rect 675110 782620 675116 782632
rect 675168 782620 675174 782672
rect 669038 782484 669044 782536
rect 669096 782524 669102 782536
rect 675294 782524 675300 782536
rect 669096 782496 675300 782524
rect 669096 782484 669102 782496
rect 675294 782484 675300 782496
rect 675352 782484 675358 782536
rect 655514 781056 655520 781108
rect 655572 781096 655578 781108
rect 675018 781096 675024 781108
rect 655572 781068 675024 781096
rect 655572 781056 655578 781068
rect 675018 781056 675024 781068
rect 675076 781056 675082 781108
rect 673914 779968 673920 780020
rect 673972 780008 673978 780020
rect 675110 780008 675116 780020
rect 673972 779980 675116 780008
rect 673972 779968 673978 779980
rect 675110 779968 675116 779980
rect 675168 779968 675174 780020
rect 655054 778336 655060 778388
rect 655112 778376 655118 778388
rect 674926 778376 674932 778388
rect 655112 778348 674932 778376
rect 655112 778336 655118 778348
rect 674926 778336 674932 778348
rect 674984 778336 674990 778388
rect 651466 777588 651472 777640
rect 651524 777628 651530 777640
rect 660298 777628 660304 777640
rect 651524 777600 660304 777628
rect 651524 777588 651530 777600
rect 660298 777588 660304 777600
rect 660356 777588 660362 777640
rect 670418 776976 670424 777028
rect 670476 777016 670482 777028
rect 675294 777016 675300 777028
rect 670476 776988 675300 777016
rect 670476 776976 670482 776988
rect 675294 776976 675300 776988
rect 675352 776976 675358 777028
rect 672718 775616 672724 775668
rect 672776 775656 672782 775668
rect 674926 775656 674932 775668
rect 672776 775628 674932 775656
rect 672776 775616 672782 775628
rect 674926 775616 674932 775628
rect 674984 775616 674990 775668
rect 651466 775548 651472 775600
rect 651524 775588 651530 775600
rect 669958 775588 669964 775600
rect 651524 775560 669964 775588
rect 651524 775548 651530 775560
rect 669958 775548 669964 775560
rect 670016 775548 670022 775600
rect 651374 775276 651380 775328
rect 651432 775316 651438 775328
rect 653398 775316 653404 775328
rect 651432 775288 653404 775316
rect 651432 775276 651438 775288
rect 653398 775276 653404 775288
rect 653456 775276 653462 775328
rect 35802 774188 35808 774240
rect 35860 774228 35866 774240
rect 41690 774228 41696 774240
rect 35860 774200 41696 774228
rect 35860 774188 35866 774200
rect 41690 774188 41696 774200
rect 41748 774188 41754 774240
rect 42058 774188 42064 774240
rect 42116 774228 42122 774240
rect 58618 774228 58624 774240
rect 42116 774200 58624 774228
rect 42116 774188 42122 774200
rect 58618 774188 58624 774200
rect 58676 774188 58682 774240
rect 651466 774120 651472 774172
rect 651524 774160 651530 774172
rect 655514 774160 655520 774172
rect 651524 774132 655520 774160
rect 651524 774120 651530 774132
rect 655514 774120 655520 774132
rect 655572 774120 655578 774172
rect 651466 773780 651472 773832
rect 651524 773820 651530 773832
rect 655054 773820 655060 773832
rect 651524 773792 655060 773820
rect 651524 773780 651530 773792
rect 655054 773780 655060 773792
rect 655112 773780 655118 773832
rect 35434 773372 35440 773424
rect 35492 773412 35498 773424
rect 41506 773412 41512 773424
rect 35492 773384 41512 773412
rect 35492 773372 35498 773384
rect 41506 773372 41512 773384
rect 41564 773372 41570 773424
rect 671430 773372 671436 773424
rect 671488 773412 671494 773424
rect 675294 773412 675300 773424
rect 671488 773384 675300 773412
rect 671488 773372 671494 773384
rect 675294 773372 675300 773384
rect 675352 773372 675358 773424
rect 41690 773208 41696 773220
rect 41386 773180 41696 773208
rect 35802 773100 35808 773152
rect 35860 773140 35866 773152
rect 41386 773140 41414 773180
rect 41690 773168 41696 773180
rect 41748 773168 41754 773220
rect 42058 773168 42064 773220
rect 42116 773208 42122 773220
rect 42886 773208 42892 773220
rect 42116 773180 42892 773208
rect 42116 773168 42122 773180
rect 42886 773168 42892 773180
rect 42944 773168 42950 773220
rect 35860 773112 41414 773140
rect 35860 773100 35866 773112
rect 41690 773072 41696 773084
rect 41524 773044 41696 773072
rect 35618 772964 35624 773016
rect 35676 773004 35682 773016
rect 41524 773004 41552 773044
rect 41690 773032 41696 773044
rect 41748 773032 41754 773084
rect 42058 773032 42064 773084
rect 42116 773072 42122 773084
rect 46198 773072 46204 773084
rect 42116 773044 46204 773072
rect 42116 773032 42122 773044
rect 46198 773032 46204 773044
rect 46256 773032 46262 773084
rect 35676 772976 41552 773004
rect 35676 772964 35682 772976
rect 35250 772828 35256 772880
rect 35308 772868 35314 772880
rect 41690 772868 41696 772880
rect 35308 772840 41696 772868
rect 35308 772828 35314 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 42058 772828 42064 772880
rect 42116 772868 42122 772880
rect 61378 772868 61384 772880
rect 42116 772840 61384 772868
rect 42116 772828 42122 772840
rect 61378 772828 61384 772840
rect 61436 772828 61442 772880
rect 35802 771808 35808 771860
rect 35860 771848 35866 771860
rect 39942 771848 39948 771860
rect 35860 771820 39948 771848
rect 35860 771808 35866 771820
rect 39942 771808 39948 771820
rect 40000 771808 40006 771860
rect 40310 771644 40316 771656
rect 36004 771616 40316 771644
rect 35618 771536 35624 771588
rect 35676 771576 35682 771588
rect 36004 771576 36032 771616
rect 40310 771604 40316 771616
rect 40368 771604 40374 771656
rect 35676 771548 36032 771576
rect 35676 771536 35682 771548
rect 42058 771468 42064 771520
rect 42116 771508 42122 771520
rect 45278 771508 45284 771520
rect 42116 771480 45284 771508
rect 42116 771468 42122 771480
rect 45278 771468 45284 771480
rect 45336 771468 45342 771520
rect 35802 771400 35808 771452
rect 35860 771440 35866 771452
rect 41690 771440 41696 771452
rect 35860 771412 41696 771440
rect 35860 771400 35866 771412
rect 41690 771400 41696 771412
rect 41748 771400 41754 771452
rect 35802 770448 35808 770500
rect 35860 770488 35866 770500
rect 40310 770488 40316 770500
rect 35860 770460 40316 770488
rect 35860 770448 35866 770460
rect 40310 770448 40316 770460
rect 40368 770448 40374 770500
rect 41690 770284 41696 770296
rect 41386 770256 41696 770284
rect 35434 770176 35440 770228
rect 35492 770216 35498 770228
rect 41386 770216 41414 770256
rect 41690 770244 41696 770256
rect 41748 770244 41754 770296
rect 42058 770244 42064 770296
rect 42116 770284 42122 770296
rect 43070 770284 43076 770296
rect 42116 770256 43076 770284
rect 42116 770244 42122 770256
rect 43070 770244 43076 770256
rect 43128 770244 43134 770296
rect 35492 770188 41414 770216
rect 35492 770176 35498 770188
rect 42058 770108 42064 770160
rect 42116 770148 42122 770160
rect 44542 770148 44548 770160
rect 42116 770120 44548 770148
rect 42116 770108 42122 770120
rect 44542 770108 44548 770120
rect 44600 770108 44606 770160
rect 35618 770040 35624 770092
rect 35676 770080 35682 770092
rect 41690 770080 41696 770092
rect 35676 770052 41696 770080
rect 35676 770040 35682 770052
rect 41690 770040 41696 770052
rect 41748 770040 41754 770092
rect 35802 768816 35808 768868
rect 35860 768856 35866 768868
rect 40034 768856 40040 768868
rect 35860 768828 40040 768856
rect 35860 768816 35866 768828
rect 40034 768816 40040 768828
rect 40092 768816 40098 768868
rect 35618 768680 35624 768732
rect 35676 768720 35682 768732
rect 41690 768720 41696 768732
rect 35676 768692 41696 768720
rect 35676 768680 35682 768692
rect 41690 768680 41696 768692
rect 41748 768680 41754 768732
rect 35802 767592 35808 767644
rect 35860 767632 35866 767644
rect 36538 767632 36544 767644
rect 35860 767604 36544 767632
rect 35860 767592 35866 767604
rect 36538 767592 36544 767604
rect 36596 767592 36602 767644
rect 35802 766028 35808 766080
rect 35860 766068 35866 766080
rect 39390 766068 39396 766080
rect 35860 766040 39396 766068
rect 35860 766028 35866 766040
rect 39390 766028 39396 766040
rect 39448 766028 39454 766080
rect 40034 765280 40040 765332
rect 40092 765320 40098 765332
rect 41690 765320 41696 765332
rect 40092 765292 41696 765320
rect 40092 765280 40098 765292
rect 41690 765280 41696 765292
rect 41748 765280 41754 765332
rect 42058 765144 42064 765196
rect 42116 765184 42122 765196
rect 42426 765184 42432 765196
rect 42116 765156 42432 765184
rect 42116 765144 42122 765156
rect 42426 765144 42432 765156
rect 42484 765144 42490 765196
rect 35802 764804 35808 764856
rect 35860 764844 35866 764856
rect 39942 764844 39948 764856
rect 35860 764816 39948 764844
rect 35860 764804 35866 764816
rect 39942 764804 39948 764816
rect 40000 764804 40006 764856
rect 41690 764640 41696 764652
rect 36004 764612 41696 764640
rect 35618 764532 35624 764584
rect 35676 764572 35682 764584
rect 36004 764572 36032 764612
rect 41690 764600 41696 764612
rect 41748 764600 41754 764652
rect 42058 764600 42064 764652
rect 42116 764640 42122 764652
rect 43438 764640 43444 764652
rect 42116 764612 43444 764640
rect 42116 764600 42122 764612
rect 43438 764600 43444 764612
rect 43496 764600 43502 764652
rect 35676 764544 36032 764572
rect 35676 764532 35682 764544
rect 35618 763444 35624 763496
rect 35676 763484 35682 763496
rect 39942 763484 39948 763496
rect 35676 763456 39948 763484
rect 35676 763444 35682 763456
rect 39942 763444 39948 763456
rect 40000 763444 40006 763496
rect 42058 763376 42064 763428
rect 42116 763376 42122 763428
rect 42076 763280 42104 763376
rect 38626 763252 41736 763280
rect 35802 763172 35808 763224
rect 35860 763212 35866 763224
rect 38626 763212 38654 763252
rect 35860 763184 38654 763212
rect 35860 763172 35866 763184
rect 41708 763156 41736 763252
rect 41984 763252 48314 763280
rect 41690 763104 41696 763156
rect 41748 763104 41754 763156
rect 41984 763144 42012 763252
rect 42076 763144 42104 763252
rect 48286 763212 48314 763252
rect 59998 763212 60004 763224
rect 48286 763184 60004 763212
rect 59998 763172 60004 763184
rect 60056 763172 60062 763224
rect 41984 763116 42104 763144
rect 42058 761880 42064 761932
rect 42116 761920 42122 761932
rect 48958 761920 48964 761932
rect 42116 761892 48964 761920
rect 42116 761880 42122 761892
rect 48958 761880 48964 761892
rect 49016 761880 49022 761932
rect 35802 761812 35808 761864
rect 35860 761852 35866 761864
rect 41690 761852 41696 761864
rect 35860 761824 41696 761852
rect 35860 761812 35866 761824
rect 41690 761812 41696 761824
rect 41748 761812 41754 761864
rect 35158 759772 35164 759824
rect 35216 759812 35222 759824
rect 39666 759812 39672 759824
rect 35216 759784 39672 759812
rect 35216 759772 35222 759784
rect 39666 759772 39672 759784
rect 39724 759772 39730 759824
rect 32398 759636 32404 759688
rect 32456 759676 32462 759688
rect 41598 759676 41604 759688
rect 32456 759648 41604 759676
rect 32456 759636 32462 759648
rect 41598 759636 41604 759648
rect 41656 759636 41662 759688
rect 33778 758276 33784 758328
rect 33836 758316 33842 758328
rect 39942 758316 39948 758328
rect 33836 758288 39948 758316
rect 33836 758276 33842 758288
rect 39942 758276 39948 758288
rect 40000 758276 40006 758328
rect 43898 755488 43904 755540
rect 43956 755528 43962 755540
rect 62942 755528 62948 755540
rect 43956 755500 62948 755528
rect 43956 755488 43962 755500
rect 62942 755488 62948 755500
rect 63000 755488 63006 755540
rect 42610 753720 42616 753772
rect 42668 753720 42674 753772
rect 42628 753636 42656 753720
rect 42610 753584 42616 753636
rect 42668 753584 42674 753636
rect 42242 749708 42248 749760
rect 42300 749708 42306 749760
rect 42260 749216 42288 749708
rect 42242 749164 42248 749216
rect 42300 749164 42306 749216
rect 61378 747260 61384 747312
rect 61436 747300 61442 747312
rect 63034 747300 63040 747312
rect 61436 747272 63040 747300
rect 61436 747260 61442 747272
rect 63034 747260 63040 747272
rect 63092 747260 63098 747312
rect 653398 746580 653404 746632
rect 653456 746620 653462 746632
rect 675386 746620 675392 746632
rect 653456 746592 675392 746620
rect 653456 746580 653462 746592
rect 675386 746580 675392 746592
rect 675444 746580 675450 746632
rect 45278 746512 45284 746564
rect 45336 746552 45342 746564
rect 62114 746552 62120 746564
rect 45336 746524 62120 746552
rect 45336 746512 45342 746524
rect 62114 746512 62120 746524
rect 62172 746512 62178 746564
rect 42242 745288 42248 745340
rect 42300 745288 42306 745340
rect 42260 745136 42288 745288
rect 42242 745084 42248 745136
rect 42300 745084 42306 745136
rect 42794 743996 42800 744048
rect 42852 744036 42858 744048
rect 42852 744008 45554 744036
rect 42852 743996 42858 744008
rect 45526 743900 45554 744008
rect 62114 743900 62120 743912
rect 45526 743872 62120 743900
rect 62114 743860 62120 743872
rect 62172 743860 62178 743912
rect 46198 743724 46204 743776
rect 46256 743764 46262 743776
rect 62114 743764 62120 743776
rect 46256 743736 62120 743764
rect 46256 743724 46262 743736
rect 62114 743724 62120 743736
rect 62172 743724 62178 743776
rect 671798 742432 671804 742484
rect 671856 742472 671862 742484
rect 675386 742472 675392 742484
rect 671856 742444 675392 742472
rect 671856 742432 671862 742444
rect 675386 742432 675392 742444
rect 675444 742432 675450 742484
rect 58618 742364 58624 742416
rect 58676 742404 58682 742416
rect 62114 742404 62120 742416
rect 58676 742376 62120 742404
rect 58676 742364 58682 742376
rect 62114 742364 62120 742376
rect 62172 742364 62178 742416
rect 671614 741140 671620 741192
rect 671672 741180 671678 741192
rect 675202 741180 675208 741192
rect 671672 741152 675208 741180
rect 671672 741140 671678 741152
rect 675202 741140 675208 741152
rect 675260 741140 675266 741192
rect 672258 739100 672264 739152
rect 672316 739140 672322 739152
rect 675386 739140 675392 739152
rect 672316 739112 675392 739140
rect 672316 739100 672322 739112
rect 675386 739100 675392 739112
rect 675444 739100 675450 739152
rect 673546 738692 673552 738744
rect 673604 738732 673610 738744
rect 675386 738732 675392 738744
rect 673604 738704 675392 738732
rect 673604 738692 673610 738704
rect 675386 738692 675392 738704
rect 675444 738692 675450 738744
rect 674834 738556 674840 738608
rect 674892 738596 674898 738608
rect 675202 738596 675208 738608
rect 674892 738568 675208 738596
rect 674892 738556 674898 738568
rect 675202 738556 675208 738568
rect 675260 738556 675266 738608
rect 652018 736856 652024 736908
rect 652076 736896 652082 736908
rect 656158 736896 656164 736908
rect 652076 736868 656164 736896
rect 652076 736856 652082 736868
rect 656158 736856 656164 736868
rect 656216 736856 656222 736908
rect 675110 736012 675116 736024
rect 663766 735984 675116 736012
rect 657538 735564 657544 735616
rect 657596 735604 657602 735616
rect 663766 735604 663794 735984
rect 675110 735972 675116 735984
rect 675168 735972 675174 736024
rect 657596 735576 663794 735604
rect 657596 735564 657602 735576
rect 674006 735088 674012 735140
rect 674064 735128 674070 735140
rect 675294 735128 675300 735140
rect 674064 735100 675300 735128
rect 674064 735088 674070 735100
rect 675294 735088 675300 735100
rect 675352 735088 675358 735140
rect 675110 734584 675116 734596
rect 663766 734556 675116 734584
rect 654778 734136 654784 734188
rect 654836 734176 654842 734188
rect 663766 734176 663794 734556
rect 675110 734544 675116 734556
rect 675168 734544 675174 734596
rect 654836 734148 663794 734176
rect 654836 734136 654842 734148
rect 651466 733388 651472 733440
rect 651524 733428 651530 733440
rect 668578 733428 668584 733440
rect 651524 733400 668584 733428
rect 651524 733388 651530 733400
rect 668578 733388 668584 733400
rect 668636 733388 668642 733440
rect 672902 732708 672908 732760
rect 672960 732748 672966 732760
rect 675294 732748 675300 732760
rect 672960 732720 675300 732748
rect 672960 732708 672966 732720
rect 675294 732708 675300 732720
rect 675352 732708 675358 732760
rect 651466 731416 651472 731468
rect 651524 731456 651530 731468
rect 658918 731456 658924 731468
rect 651524 731428 658924 731456
rect 651524 731416 651530 731428
rect 658918 731416 658924 731428
rect 658976 731416 658982 731468
rect 35802 731144 35808 731196
rect 35860 731184 35866 731196
rect 35860 731156 38654 731184
rect 35860 731144 35866 731156
rect 38626 731116 38654 731156
rect 41690 731116 41696 731128
rect 38626 731088 41696 731116
rect 41690 731076 41696 731088
rect 41748 731076 41754 731128
rect 651374 731076 651380 731128
rect 651432 731116 651438 731128
rect 653398 731116 653404 731128
rect 651432 731088 653404 731116
rect 651432 731076 651438 731088
rect 653398 731076 653404 731088
rect 653456 731076 653462 731128
rect 652662 730668 652668 730720
rect 652720 730708 652726 730720
rect 661678 730708 661684 730720
rect 652720 730680 661684 730708
rect 652720 730668 652726 730680
rect 661678 730668 661684 730680
rect 661736 730668 661742 730720
rect 35802 730328 35808 730380
rect 35860 730368 35866 730380
rect 40402 730368 40408 730380
rect 35860 730340 40408 730368
rect 35860 730328 35866 730340
rect 40402 730328 40408 730340
rect 40460 730328 40466 730380
rect 35434 730056 35440 730108
rect 35492 730096 35498 730108
rect 41690 730096 41696 730108
rect 35492 730068 41696 730096
rect 35492 730056 35498 730068
rect 41690 730056 41696 730068
rect 41748 730056 41754 730108
rect 42058 730056 42064 730108
rect 42116 730096 42122 730108
rect 61378 730096 61384 730108
rect 42116 730068 61384 730096
rect 42116 730056 42122 730068
rect 61378 730056 61384 730068
rect 61436 730056 61442 730108
rect 651466 729988 651472 730040
rect 651524 730028 651530 730040
rect 657538 730028 657544 730040
rect 651524 730000 657544 730028
rect 651524 729988 651530 730000
rect 657538 729988 657544 730000
rect 657596 729988 657602 730040
rect 35618 729444 35624 729496
rect 35676 729484 35682 729496
rect 35676 729456 35894 729484
rect 35676 729444 35682 729456
rect 35866 729280 35894 729456
rect 42058 729308 42064 729360
rect 42116 729348 42122 729360
rect 62942 729348 62948 729360
rect 42116 729320 62948 729348
rect 42116 729308 42122 729320
rect 62942 729308 62948 729320
rect 63000 729308 63006 729360
rect 41690 729280 41696 729292
rect 35866 729252 41696 729280
rect 41690 729240 41696 729252
rect 41748 729240 41754 729292
rect 675294 729240 675300 729292
rect 675352 729240 675358 729292
rect 675312 729088 675340 729240
rect 35802 729036 35808 729088
rect 35860 729076 35866 729088
rect 41506 729076 41512 729088
rect 35860 729048 41512 729076
rect 35860 729036 35866 729048
rect 41506 729036 41512 729048
rect 41564 729036 41570 729088
rect 675294 729036 675300 729088
rect 675352 729036 675358 729088
rect 42058 728832 42064 728884
rect 42116 728872 42122 728884
rect 44266 728872 44272 728884
rect 42116 728844 44272 728872
rect 42116 728832 42122 728844
rect 44266 728832 44272 728844
rect 44324 728832 44330 728884
rect 35618 728764 35624 728816
rect 35676 728804 35682 728816
rect 41690 728804 41696 728816
rect 35676 728776 41696 728804
rect 35676 728764 35682 728776
rect 41690 728764 41696 728776
rect 41748 728764 41754 728816
rect 35434 728628 35440 728680
rect 35492 728668 35498 728680
rect 41690 728668 41696 728680
rect 35492 728640 41696 728668
rect 35492 728628 35498 728640
rect 41690 728628 41696 728640
rect 41748 728628 41754 728680
rect 42058 728628 42064 728680
rect 42116 728668 42122 728680
rect 44542 728668 44548 728680
rect 42116 728640 44548 728668
rect 42116 728628 42122 728640
rect 44542 728628 44548 728640
rect 44600 728628 44606 728680
rect 651466 728492 651472 728544
rect 651524 728532 651530 728544
rect 654778 728532 654784 728544
rect 651524 728504 654784 728532
rect 651524 728492 651530 728504
rect 654778 728492 654784 728504
rect 654836 728492 654842 728544
rect 673086 728288 673092 728340
rect 673144 728328 673150 728340
rect 673144 728300 674176 728328
rect 673144 728288 673150 728300
rect 670878 728084 670884 728136
rect 670936 728124 670942 728136
rect 670936 728096 674058 728124
rect 670936 728084 670942 728096
rect 35802 727812 35808 727864
rect 35860 727852 35866 727864
rect 40034 727852 40040 727864
rect 35860 727824 40040 727852
rect 35860 727812 35866 727824
rect 40034 727812 40040 727824
rect 40092 727812 40098 727864
rect 41690 727648 41696 727660
rect 36004 727620 41696 727648
rect 35434 727540 35440 727592
rect 35492 727580 35498 727592
rect 36004 727580 36032 727620
rect 41690 727608 41696 727620
rect 41748 727608 41754 727660
rect 35492 727552 36032 727580
rect 35492 727540 35498 727552
rect 35802 727404 35808 727456
rect 35860 727444 35866 727456
rect 41690 727444 41696 727456
rect 35860 727416 41696 727444
rect 35860 727404 35866 727416
rect 41690 727404 41696 727416
rect 41748 727404 41754 727456
rect 42058 727404 42064 727456
rect 42116 727444 42122 727456
rect 43438 727444 43444 727456
rect 42116 727416 43444 727444
rect 42116 727404 42122 727416
rect 43438 727404 43444 727416
rect 43496 727404 43502 727456
rect 35618 727268 35624 727320
rect 35676 727308 35682 727320
rect 41690 727308 41696 727320
rect 35676 727280 41696 727308
rect 35676 727268 35682 727280
rect 41690 727268 41696 727280
rect 41748 727268 41754 727320
rect 42058 727268 42064 727320
rect 42116 727308 42122 727320
rect 43622 727308 43628 727320
rect 42116 727280 43628 727308
rect 42116 727268 42122 727280
rect 43622 727268 43628 727280
rect 43680 727268 43686 727320
rect 674834 727200 674840 727252
rect 674892 727240 674898 727252
rect 680998 727240 681004 727252
rect 674892 727212 681004 727240
rect 674892 727200 674898 727212
rect 680998 727200 681004 727212
rect 681056 727200 681062 727252
rect 674558 726724 674564 726776
rect 674616 726764 674622 726776
rect 683390 726764 683396 726776
rect 674616 726736 683396 726764
rect 674616 726724 674622 726736
rect 683390 726724 683396 726736
rect 683448 726724 683454 726776
rect 674374 726588 674380 726640
rect 674432 726628 674438 726640
rect 684034 726628 684040 726640
rect 674432 726600 684040 726628
rect 674432 726588 674438 726600
rect 684034 726588 684040 726600
rect 684092 726588 684098 726640
rect 41322 726044 41328 726096
rect 41380 726084 41386 726096
rect 41690 726084 41696 726096
rect 41380 726056 41696 726084
rect 41380 726044 41386 726056
rect 41690 726044 41696 726056
rect 41748 726044 41754 726096
rect 42058 726044 42064 726096
rect 42116 726084 42122 726096
rect 42518 726084 42524 726096
rect 42116 726056 42524 726084
rect 42116 726044 42122 726056
rect 42518 726044 42524 726056
rect 42576 726044 42582 726096
rect 41138 725908 41144 725960
rect 41196 725948 41202 725960
rect 41598 725948 41604 725960
rect 41196 725920 41604 725948
rect 41196 725908 41202 725920
rect 41598 725908 41604 725920
rect 41656 725908 41662 725960
rect 675294 721692 675300 721744
rect 675352 721692 675358 721744
rect 675312 721268 675340 721692
rect 675294 721216 675300 721268
rect 675352 721216 675358 721268
rect 675294 720808 675300 720860
rect 675352 720808 675358 720860
rect 675312 720520 675340 720808
rect 675294 720468 675300 720520
rect 675352 720468 675358 720520
rect 43622 718972 43628 719024
rect 43680 719012 43686 719024
rect 53098 719012 53104 719024
rect 43680 718984 53104 719012
rect 43680 718972 43686 718984
rect 53098 718972 53104 718984
rect 53156 718972 53162 719024
rect 672810 717476 672816 717528
rect 672868 717516 672874 717528
rect 673270 717516 673276 717528
rect 672868 717488 673276 717516
rect 672868 717476 672874 717488
rect 673270 717476 673276 717488
rect 673328 717476 673334 717528
rect 32398 716864 32404 716916
rect 32456 716904 32462 716916
rect 41690 716904 41696 716916
rect 32456 716876 41696 716904
rect 32456 716864 32462 716876
rect 41690 716864 41696 716876
rect 41748 716864 41754 716916
rect 42058 716728 42064 716780
rect 42116 716768 42122 716780
rect 42702 716768 42708 716780
rect 42116 716740 42708 716768
rect 42116 716728 42122 716740
rect 42702 716728 42708 716740
rect 42760 716728 42766 716780
rect 42058 716592 42064 716644
rect 42116 716632 42122 716644
rect 42518 716632 42524 716644
rect 42116 716604 42524 716632
rect 42116 716592 42122 716604
rect 42518 716592 42524 716604
rect 42576 716592 42582 716644
rect 656158 716252 656164 716304
rect 656216 716292 656222 716304
rect 673270 716292 673276 716304
rect 656216 716264 673276 716292
rect 656216 716252 656222 716264
rect 673270 716252 673276 716264
rect 673328 716252 673334 716304
rect 35158 715708 35164 715760
rect 35216 715748 35222 715760
rect 41322 715748 41328 715760
rect 35216 715720 41328 715748
rect 35216 715708 35222 715720
rect 41322 715708 41328 715720
rect 41380 715708 41386 715760
rect 669958 715708 669964 715760
rect 670016 715748 670022 715760
rect 673086 715748 673092 715760
rect 670016 715720 673092 715748
rect 670016 715708 670022 715720
rect 673086 715708 673092 715720
rect 673144 715708 673150 715760
rect 31662 715504 31668 715556
rect 31720 715544 31726 715556
rect 40586 715544 40592 715556
rect 31720 715516 40592 715544
rect 31720 715504 31726 715516
rect 40586 715504 40592 715516
rect 40644 715504 40650 715556
rect 671062 715300 671068 715352
rect 671120 715340 671126 715352
rect 673086 715340 673092 715352
rect 671120 715312 673092 715340
rect 671120 715300 671126 715312
rect 673086 715300 673092 715312
rect 673144 715300 673150 715352
rect 660298 714960 660304 715012
rect 660356 715000 660362 715012
rect 673270 715000 673276 715012
rect 660356 714972 673276 715000
rect 660356 714960 660362 714972
rect 673270 714960 673276 714972
rect 673328 714960 673334 715012
rect 671890 714484 671896 714536
rect 671948 714524 671954 714536
rect 673270 714524 673276 714536
rect 671948 714496 673276 714524
rect 671948 714484 671954 714496
rect 673270 714484 673276 714496
rect 673328 714484 673334 714536
rect 673270 713532 673276 713584
rect 673328 713572 673334 713584
rect 673328 713544 673500 713572
rect 673328 713532 673334 713544
rect 672074 713396 672080 713448
rect 672132 713436 672138 713448
rect 673270 713436 673276 713448
rect 672132 713408 673276 713436
rect 672132 713396 672138 713408
rect 673270 713396 673276 713408
rect 673328 713396 673334 713448
rect 672626 713260 672632 713312
rect 672684 713300 672690 713312
rect 673472 713300 673500 713544
rect 672684 713272 673500 713300
rect 672684 713260 672690 713272
rect 671062 712580 671068 712632
rect 671120 712620 671126 712632
rect 671982 712620 671988 712632
rect 671120 712592 671988 712620
rect 671120 712580 671126 712592
rect 671982 712580 671988 712592
rect 672040 712580 672046 712632
rect 43622 712104 43628 712156
rect 43680 712144 43686 712156
rect 51718 712144 51724 712156
rect 43680 712116 51724 712144
rect 43680 712104 43686 712116
rect 51718 712104 51724 712116
rect 51776 712104 51782 712156
rect 672442 712036 672448 712088
rect 672500 712076 672506 712088
rect 673270 712076 673276 712088
rect 672500 712048 673276 712076
rect 672500 712036 672506 712048
rect 673270 712036 673276 712048
rect 673328 712036 673334 712088
rect 672442 711764 672448 711816
rect 672500 711804 672506 711816
rect 673086 711804 673092 711816
rect 672500 711776 673092 711804
rect 672500 711764 672506 711776
rect 673086 711764 673092 711776
rect 673144 711764 673150 711816
rect 42242 710404 42248 710456
rect 42300 710444 42306 710456
rect 44726 710444 44732 710456
rect 42300 710416 44732 710444
rect 42300 710404 42306 710416
rect 44726 710404 44732 710416
rect 44784 710404 44790 710456
rect 671430 709996 671436 710048
rect 671488 710036 671494 710048
rect 673086 710036 673092 710048
rect 671488 710008 673092 710036
rect 671488 709996 671494 710008
rect 673086 709996 673092 710008
rect 673144 709996 673150 710048
rect 43622 709316 43628 709368
rect 43680 709356 43686 709368
rect 45094 709356 45100 709368
rect 43680 709328 45100 709356
rect 43680 709316 43686 709328
rect 45094 709316 45100 709328
rect 45152 709316 45158 709368
rect 669038 709316 669044 709368
rect 669096 709356 669102 709368
rect 673270 709356 673276 709368
rect 669096 709328 673276 709356
rect 669096 709316 669102 709328
rect 673270 709316 673276 709328
rect 673328 709316 673334 709368
rect 670602 709180 670608 709232
rect 670660 709220 670666 709232
rect 673270 709220 673276 709232
rect 670660 709192 673276 709220
rect 670660 709180 670666 709192
rect 673270 709180 673276 709192
rect 673328 709180 673334 709232
rect 669222 708228 669228 708280
rect 669280 708268 669286 708280
rect 673270 708268 673276 708280
rect 669280 708240 673276 708268
rect 669280 708228 669286 708240
rect 673270 708228 673276 708240
rect 673328 708228 673334 708280
rect 42242 707820 42248 707872
rect 42300 707860 42306 707872
rect 43622 707860 43628 707872
rect 42300 707832 43628 707860
rect 42300 707820 42306 707832
rect 43622 707820 43628 707832
rect 43680 707820 43686 707872
rect 42242 707412 42248 707464
rect 42300 707452 42306 707464
rect 42702 707452 42708 707464
rect 42300 707424 42708 707452
rect 42300 707412 42306 707424
rect 42702 707412 42708 707424
rect 42760 707412 42766 707464
rect 674650 707140 674656 707192
rect 674708 707180 674714 707192
rect 676030 707180 676036 707192
rect 674708 707152 676036 707180
rect 674708 707140 674714 707152
rect 676030 707140 676036 707152
rect 676088 707140 676094 707192
rect 42518 706664 42524 706716
rect 42576 706664 42582 706716
rect 42536 706500 42564 706664
rect 42702 706500 42708 706512
rect 42536 706472 42708 706500
rect 42702 706460 42708 706472
rect 42760 706460 42766 706512
rect 42242 705508 42248 705560
rect 42300 705548 42306 705560
rect 43806 705548 43812 705560
rect 42300 705520 43812 705548
rect 42300 705508 42306 705520
rect 43806 705508 43812 705520
rect 43864 705508 43870 705560
rect 670418 705372 670424 705424
rect 670476 705412 670482 705424
rect 673270 705412 673276 705424
rect 670476 705384 673276 705412
rect 670476 705372 670482 705384
rect 673270 705372 673276 705384
rect 673328 705372 673334 705424
rect 674282 705304 674288 705356
rect 674340 705344 674346 705356
rect 683114 705344 683120 705356
rect 674340 705316 683120 705344
rect 674340 705304 674346 705316
rect 683114 705304 683120 705316
rect 683172 705304 683178 705356
rect 673730 705276 673736 705288
rect 669286 705248 673736 705276
rect 667842 705168 667848 705220
rect 667900 705208 667906 705220
rect 669286 705208 669314 705248
rect 673730 705236 673736 705248
rect 673788 705236 673794 705288
rect 667900 705180 669314 705208
rect 667900 705168 667906 705180
rect 51718 705100 51724 705152
rect 51776 705140 51782 705152
rect 62114 705140 62120 705152
rect 51776 705112 62120 705140
rect 51776 705100 51782 705112
rect 62114 705100 62120 705112
rect 62172 705100 62178 705152
rect 667014 703808 667020 703860
rect 667072 703848 667078 703860
rect 673730 703848 673736 703860
rect 667072 703820 673736 703848
rect 667072 703808 667078 703820
rect 673730 703808 673736 703820
rect 673788 703808 673794 703860
rect 44726 703740 44732 703792
rect 44784 703780 44790 703792
rect 62114 703780 62120 703792
rect 44784 703752 62120 703780
rect 44784 703740 44790 703752
rect 62114 703740 62120 703752
rect 62172 703740 62178 703792
rect 654778 701156 654784 701208
rect 654836 701196 654842 701208
rect 673730 701196 673736 701208
rect 654836 701168 673736 701196
rect 654836 701156 654842 701168
rect 673730 701156 673736 701168
rect 673788 701156 673794 701208
rect 42702 701088 42708 701140
rect 42760 701128 42766 701140
rect 42760 701100 51074 701128
rect 42760 701088 42766 701100
rect 51046 701060 51074 701100
rect 62942 701060 62948 701072
rect 51046 701032 62948 701060
rect 62942 701020 62948 701032
rect 63000 701020 63006 701072
rect 46198 698232 46204 698284
rect 46256 698272 46262 698284
rect 62206 698272 62212 698284
rect 46256 698244 62212 698272
rect 46256 698232 46262 698244
rect 62206 698232 62212 698244
rect 62264 698232 62270 698284
rect 674282 692996 674288 693048
rect 674340 693036 674346 693048
rect 675386 693036 675392 693048
rect 674340 693008 675392 693036
rect 674340 692996 674346 693008
rect 675386 692996 675392 693008
rect 675444 692996 675450 693048
rect 668394 692792 668400 692844
rect 668452 692832 668458 692844
rect 673730 692832 673736 692844
rect 668452 692804 673736 692832
rect 668452 692792 668458 692804
rect 673730 692792 673736 692804
rect 673788 692792 673794 692844
rect 656434 690072 656440 690124
rect 656492 690112 656498 690124
rect 673730 690112 673736 690124
rect 656492 690084 673736 690112
rect 656492 690072 656498 690084
rect 673730 690072 673736 690084
rect 673788 690072 673794 690124
rect 674834 688984 674840 689036
rect 674892 689024 674898 689036
rect 675202 689024 675208 689036
rect 674892 688996 675208 689024
rect 674892 688984 674898 688996
rect 675202 688984 675208 688996
rect 675260 688984 675266 689036
rect 652754 688780 652760 688832
rect 652812 688820 652818 688832
rect 673730 688820 673736 688832
rect 652812 688792 673736 688820
rect 652812 688780 652818 688792
rect 673730 688780 673736 688792
rect 673788 688780 673794 688832
rect 651466 688644 651472 688696
rect 651524 688684 651530 688696
rect 657538 688684 657544 688696
rect 651524 688656 657544 688684
rect 651524 688644 651530 688656
rect 657538 688644 657544 688656
rect 657596 688644 657602 688696
rect 35802 687488 35808 687540
rect 35860 687528 35866 687540
rect 41690 687528 41696 687540
rect 35860 687500 41696 687528
rect 35860 687488 35866 687500
rect 41690 687488 41696 687500
rect 41748 687488 41754 687540
rect 35434 687216 35440 687268
rect 35492 687256 35498 687268
rect 35492 687228 38654 687256
rect 35492 687216 35498 687228
rect 38626 687188 38654 687228
rect 651466 687216 651472 687268
rect 651524 687256 651530 687268
rect 669958 687256 669964 687268
rect 651524 687228 669964 687256
rect 651524 687216 651530 687228
rect 669958 687216 669964 687228
rect 670016 687216 670022 687268
rect 41690 687188 41696 687200
rect 38626 687160 41696 687188
rect 41690 687148 41696 687160
rect 41748 687148 41754 687200
rect 651466 687012 651472 687064
rect 651524 687052 651530 687064
rect 654778 687052 654784 687064
rect 651524 687024 654784 687052
rect 651524 687012 651530 687024
rect 654778 687012 654784 687024
rect 654836 687012 654842 687064
rect 42058 686468 42064 686520
rect 42116 686508 42122 686520
rect 62942 686508 62948 686520
rect 42116 686480 62948 686508
rect 42116 686468 42122 686480
rect 62942 686468 62948 686480
rect 63000 686468 63006 686520
rect 651650 686468 651656 686520
rect 651708 686508 651714 686520
rect 667198 686508 667204 686520
rect 651708 686480 667204 686508
rect 651708 686468 651714 686480
rect 667198 686468 667204 686480
rect 667256 686468 667262 686520
rect 35618 686400 35624 686452
rect 35676 686440 35682 686452
rect 41690 686440 41696 686452
rect 35676 686412 41696 686440
rect 35676 686400 35682 686412
rect 41690 686400 41696 686412
rect 41748 686400 41754 686452
rect 35802 686264 35808 686316
rect 35860 686304 35866 686316
rect 41690 686304 41696 686316
rect 35860 686276 41696 686304
rect 35860 686264 35866 686276
rect 41690 686264 41696 686276
rect 41748 686264 41754 686316
rect 42058 686264 42064 686316
rect 42116 686304 42122 686316
rect 43622 686304 43628 686316
rect 42116 686276 43628 686304
rect 42116 686264 42122 686276
rect 43622 686264 43628 686276
rect 43680 686264 43686 686316
rect 42058 686060 42064 686112
rect 42116 686100 42122 686112
rect 44542 686100 44548 686112
rect 42116 686072 44548 686100
rect 42116 686060 42122 686072
rect 44542 686060 44548 686072
rect 44600 686060 44606 686112
rect 35434 685992 35440 686044
rect 35492 686032 35498 686044
rect 41690 686032 41696 686044
rect 35492 686004 41696 686032
rect 35492 685992 35498 686004
rect 41690 685992 41696 686004
rect 41748 685992 41754 686044
rect 35802 685856 35808 685908
rect 35860 685896 35866 685908
rect 41690 685896 41696 685908
rect 35860 685868 41696 685896
rect 35860 685856 35866 685868
rect 41690 685856 41696 685868
rect 41748 685856 41754 685908
rect 42058 685856 42064 685908
rect 42116 685896 42122 685908
rect 44266 685896 44272 685908
rect 42116 685868 44272 685896
rect 42116 685856 42122 685868
rect 44266 685856 44272 685868
rect 44324 685856 44330 685908
rect 651466 685516 651472 685568
rect 651524 685556 651530 685568
rect 656434 685556 656440 685568
rect 651524 685528 656440 685556
rect 651524 685516 651530 685528
rect 656434 685516 656440 685528
rect 656492 685516 656498 685568
rect 35802 684972 35808 685024
rect 35860 685012 35866 685024
rect 35860 684972 35894 685012
rect 35866 684944 35894 684972
rect 41690 684944 41696 684956
rect 35866 684916 41696 684944
rect 41690 684904 41696 684916
rect 41748 684904 41754 684956
rect 42242 684768 42248 684820
rect 42300 684808 42306 684820
rect 45278 684808 45284 684820
rect 42300 684780 45284 684808
rect 42300 684768 42306 684780
rect 45278 684768 45284 684780
rect 45336 684768 45342 684820
rect 35618 684632 35624 684684
rect 35676 684672 35682 684684
rect 41690 684672 41696 684684
rect 35676 684644 41696 684672
rect 35676 684632 35682 684644
rect 41690 684632 41696 684644
rect 41748 684632 41754 684684
rect 35802 684496 35808 684548
rect 35860 684536 35866 684548
rect 41690 684536 41696 684548
rect 35860 684508 41696 684536
rect 35860 684496 35866 684508
rect 41690 684496 41696 684508
rect 41748 684496 41754 684548
rect 42058 684496 42064 684548
rect 42116 684536 42122 684548
rect 43070 684536 43076 684548
rect 42116 684508 43076 684536
rect 42116 684496 42122 684508
rect 43070 684496 43076 684508
rect 43128 684496 43134 684548
rect 35802 683408 35808 683460
rect 35860 683448 35866 683460
rect 41690 683448 41696 683460
rect 35860 683420 41696 683448
rect 35860 683408 35866 683420
rect 41690 683408 41696 683420
rect 41748 683408 41754 683460
rect 35618 683272 35624 683324
rect 35676 683312 35682 683324
rect 41506 683312 41512 683324
rect 35676 683284 41512 683312
rect 35676 683272 35682 683284
rect 41506 683272 41512 683284
rect 41564 683272 41570 683324
rect 35434 683136 35440 683188
rect 35492 683176 35498 683188
rect 35492 683148 38654 683176
rect 35492 683136 35498 683148
rect 38626 683108 38654 683148
rect 41690 683108 41696 683120
rect 38626 683080 41696 683108
rect 41690 683068 41696 683080
rect 41748 683068 41754 683120
rect 675478 682524 675484 682576
rect 675536 682564 675542 682576
rect 683206 682564 683212 682576
rect 675536 682536 683212 682564
rect 675536 682524 675542 682536
rect 683206 682524 683212 682536
rect 683264 682524 683270 682576
rect 674834 682388 674840 682440
rect 674892 682428 674898 682440
rect 683482 682428 683488 682440
rect 674892 682400 683488 682428
rect 674892 682388 674898 682400
rect 683482 682388 683488 682400
rect 683540 682388 683546 682440
rect 35618 681844 35624 681896
rect 35676 681884 35682 681896
rect 41690 681884 41696 681896
rect 35676 681856 41696 681884
rect 35676 681844 35682 681856
rect 41690 681844 41696 681856
rect 41748 681844 41754 681896
rect 35802 681708 35808 681760
rect 35860 681748 35866 681760
rect 41506 681748 41512 681760
rect 35860 681720 41512 681748
rect 35860 681708 35866 681720
rect 41506 681708 41512 681720
rect 41564 681708 41570 681760
rect 35802 680484 35808 680536
rect 35860 680524 35866 680536
rect 41690 680524 41696 680536
rect 35860 680496 41696 680524
rect 35860 680484 35866 680496
rect 41690 680484 41696 680496
rect 41748 680484 41754 680536
rect 35802 679396 35808 679448
rect 35860 679436 35866 679448
rect 41690 679436 41696 679448
rect 35860 679408 41696 679436
rect 35860 679396 35866 679408
rect 41690 679396 41696 679408
rect 41748 679396 41754 679448
rect 35802 679124 35808 679176
rect 35860 679164 35866 679176
rect 41506 679164 41512 679176
rect 35860 679136 41512 679164
rect 35860 679124 35866 679136
rect 41506 679124 41512 679136
rect 41564 679124 41570 679176
rect 35618 678988 35624 679040
rect 35676 679028 35682 679040
rect 41690 679028 41696 679040
rect 35676 679000 41696 679028
rect 35676 678988 35682 679000
rect 41690 678988 41696 679000
rect 41748 678988 41754 679040
rect 43990 676200 43996 676252
rect 44048 676240 44054 676252
rect 57238 676240 57244 676252
rect 44048 676212 57244 676240
rect 44048 676200 44054 676212
rect 57238 676200 57244 676212
rect 57296 676200 57302 676252
rect 33042 674092 33048 674144
rect 33100 674132 33106 674144
rect 41506 674132 41512 674144
rect 33100 674104 41512 674132
rect 33100 674092 33106 674104
rect 41506 674092 41512 674104
rect 41564 674092 41570 674144
rect 35158 672800 35164 672852
rect 35216 672840 35222 672852
rect 41690 672840 41696 672852
rect 35216 672812 41696 672840
rect 35216 672800 35222 672812
rect 41690 672800 41696 672812
rect 41748 672800 41754 672852
rect 42058 672664 42064 672716
rect 42116 672704 42122 672716
rect 42518 672704 42524 672716
rect 42116 672676 42524 672704
rect 42116 672664 42122 672676
rect 42518 672664 42524 672676
rect 42576 672664 42582 672716
rect 31018 672460 31024 672512
rect 31076 672500 31082 672512
rect 41690 672500 41696 672512
rect 31076 672472 41696 672500
rect 31076 672460 31082 672472
rect 41690 672460 41696 672472
rect 41748 672460 41754 672512
rect 673546 671304 673552 671356
rect 673604 671344 673610 671356
rect 673604 671316 673776 671344
rect 673604 671304 673610 671316
rect 668578 671100 668584 671152
rect 668636 671140 668642 671152
rect 673546 671140 673552 671152
rect 668636 671112 673552 671140
rect 668636 671100 668642 671112
rect 673546 671100 673552 671112
rect 673604 671100 673610 671152
rect 661678 670692 661684 670744
rect 661736 670732 661742 670744
rect 673748 670732 673776 671316
rect 661736 670704 673776 670732
rect 661736 670692 661742 670704
rect 673546 670352 673552 670404
rect 673604 670392 673610 670404
rect 673604 670364 673776 670392
rect 673604 670352 673610 670364
rect 670234 670216 670240 670268
rect 670292 670256 670298 670268
rect 673546 670256 673552 670268
rect 670292 670228 673552 670256
rect 670292 670216 670298 670228
rect 673546 670216 673552 670228
rect 673604 670216 673610 670268
rect 44082 669400 44088 669452
rect 44140 669440 44146 669452
rect 44140 669412 51074 669440
rect 44140 669400 44146 669412
rect 51046 669372 51074 669412
rect 58618 669372 58624 669384
rect 51046 669344 58624 669372
rect 58618 669332 58624 669344
rect 58676 669332 58682 669384
rect 658918 669332 658924 669384
rect 658976 669372 658982 669384
rect 673748 669372 673776 670364
rect 658976 669344 673776 669372
rect 658976 669332 658982 669344
rect 673546 668652 673552 668704
rect 673604 668692 673610 668704
rect 673604 668664 673776 668692
rect 673604 668652 673610 668664
rect 671062 668516 671068 668568
rect 671120 668556 671126 668568
rect 673546 668556 673552 668568
rect 671120 668528 673552 668556
rect 671120 668516 671126 668528
rect 673546 668516 673552 668528
rect 673604 668516 673610 668568
rect 671430 668176 671436 668228
rect 671488 668216 671494 668228
rect 673748 668216 673776 668664
rect 671488 668188 673776 668216
rect 671488 668176 671494 668188
rect 45646 667904 45652 667956
rect 45704 667944 45710 667956
rect 61378 667944 61384 667956
rect 45704 667916 61384 667944
rect 45704 667904 45710 667916
rect 61378 667904 61384 667916
rect 61436 667904 61442 667956
rect 671062 667904 671068 667956
rect 671120 667944 671126 667956
rect 673546 667944 673552 667956
rect 671120 667916 673552 667944
rect 671120 667904 671126 667916
rect 673546 667904 673552 667916
rect 673604 667904 673610 667956
rect 673546 667292 673552 667344
rect 673604 667332 673610 667344
rect 673604 667304 673776 667332
rect 673604 667292 673610 667304
rect 671614 667156 671620 667208
rect 671672 667196 671678 667208
rect 673546 667196 673552 667208
rect 671672 667168 673552 667196
rect 671672 667156 671678 667168
rect 673546 667156 673552 667168
rect 673604 667156 673610 667208
rect 42242 667020 42248 667072
rect 42300 667060 42306 667072
rect 45646 667060 45652 667072
rect 42300 667032 45652 667060
rect 42300 667020 42306 667032
rect 45646 667020 45652 667032
rect 45704 667020 45710 667072
rect 671982 666884 671988 666936
rect 672040 666924 672046 666936
rect 673748 666924 673776 667304
rect 672040 666896 673776 666924
rect 672040 666884 672046 666896
rect 674834 666612 674840 666664
rect 674892 666652 674898 666664
rect 676030 666652 676036 666664
rect 674892 666624 676036 666652
rect 674892 666612 674898 666624
rect 676030 666612 676036 666624
rect 676088 666612 676094 666664
rect 671890 666544 671896 666596
rect 671948 666584 671954 666596
rect 673546 666584 673552 666596
rect 671948 666556 673552 666584
rect 671948 666544 671954 666556
rect 673546 666544 673552 666556
rect 673604 666544 673610 666596
rect 669590 665252 669596 665304
rect 669648 665292 669654 665304
rect 673546 665292 673552 665304
rect 669648 665264 673552 665292
rect 669648 665252 669654 665264
rect 673546 665252 673552 665264
rect 673604 665252 673610 665304
rect 671706 664368 671712 664420
rect 671764 664408 671770 664420
rect 673546 664408 673552 664420
rect 671764 664380 673552 664408
rect 671764 664368 671770 664380
rect 673546 664368 673552 664380
rect 673604 664368 673610 664420
rect 669406 663892 669412 663944
rect 669464 663932 669470 663944
rect 673546 663932 673552 663944
rect 669464 663904 673552 663932
rect 669464 663892 669470 663904
rect 673546 663892 673552 663904
rect 673604 663892 673610 663944
rect 674834 663756 674840 663808
rect 674892 663796 674898 663808
rect 676030 663796 676036 663808
rect 674892 663768 676036 663796
rect 674892 663756 674898 663768
rect 676030 663756 676036 663768
rect 676088 663756 676094 663808
rect 42242 663280 42248 663332
rect 42300 663320 42306 663332
rect 42300 663292 42564 663320
rect 42300 663280 42306 663292
rect 42536 663128 42564 663292
rect 42518 663076 42524 663128
rect 42576 663076 42582 663128
rect 42242 662940 42248 662992
rect 42300 662980 42306 662992
rect 44450 662980 44456 662992
rect 42300 662952 44456 662980
rect 42300 662940 42306 662952
rect 44450 662940 44456 662952
rect 44508 662940 44514 662992
rect 671246 661580 671252 661632
rect 671304 661620 671310 661632
rect 674006 661620 674012 661632
rect 671304 661592 674012 661620
rect 671304 661580 671310 661592
rect 674006 661580 674012 661592
rect 674064 661580 674070 661632
rect 669222 661104 669228 661156
rect 669280 661144 669286 661156
rect 674006 661144 674012 661156
rect 669280 661116 674012 661144
rect 669280 661104 669286 661116
rect 674006 661104 674012 661116
rect 674064 661104 674070 661156
rect 42150 661036 42156 661088
rect 42208 661076 42214 661088
rect 43806 661076 43812 661088
rect 42208 661048 43812 661076
rect 42208 661036 42214 661048
rect 43806 661036 43812 661048
rect 43864 661036 43870 661088
rect 58618 660900 58624 660952
rect 58676 660940 58682 660952
rect 62114 660940 62120 660952
rect 58676 660912 62120 660940
rect 58676 660900 58682 660912
rect 62114 660900 62120 660912
rect 62172 660900 62178 660952
rect 668854 660152 668860 660204
rect 668912 660192 668918 660204
rect 674006 660192 674012 660204
rect 668912 660164 674012 660192
rect 668912 660152 668918 660164
rect 674006 660152 674012 660164
rect 674064 660152 674070 660204
rect 674834 659812 674840 659864
rect 674892 659852 674898 659864
rect 683114 659852 683120 659864
rect 674892 659824 683120 659852
rect 674892 659812 674898 659824
rect 683114 659812 683120 659824
rect 683172 659812 683178 659864
rect 672166 659676 672172 659728
rect 672224 659716 672230 659728
rect 674006 659716 674012 659728
rect 672224 659688 674012 659716
rect 672224 659676 672230 659688
rect 674006 659676 674012 659688
rect 674064 659676 674070 659728
rect 42518 657500 42524 657552
rect 42576 657540 42582 657552
rect 62114 657540 62120 657552
rect 42576 657512 62120 657540
rect 42576 657500 42582 657512
rect 62114 657500 62120 657512
rect 62172 657500 62178 657552
rect 46198 656820 46204 656872
rect 46256 656860 46262 656872
rect 62114 656860 62120 656872
rect 46256 656832 62120 656860
rect 46256 656820 46262 656832
rect 62114 656820 62120 656832
rect 62172 656820 62178 656872
rect 653398 655528 653404 655580
rect 653456 655568 653462 655580
rect 674006 655568 674012 655580
rect 653456 655540 674012 655568
rect 653456 655528 653462 655540
rect 674006 655528 674012 655540
rect 674064 655528 674070 655580
rect 45462 655460 45468 655512
rect 45520 655500 45526 655512
rect 62114 655500 62120 655512
rect 45520 655472 62120 655500
rect 45520 655460 45526 655472
rect 62114 655460 62120 655472
rect 62172 655460 62178 655512
rect 655514 645872 655520 645924
rect 655572 645912 655578 645924
rect 671246 645912 671252 645924
rect 655572 645884 671252 645912
rect 655572 645872 655578 645884
rect 671246 645872 671252 645884
rect 671304 645872 671310 645924
rect 35802 644444 35808 644496
rect 35860 644484 35866 644496
rect 41690 644484 41696 644496
rect 35860 644456 41696 644484
rect 35860 644444 35866 644456
rect 41690 644444 41696 644456
rect 41748 644444 41754 644496
rect 42058 644444 42064 644496
rect 42116 644484 42122 644496
rect 58618 644484 58624 644496
rect 42116 644456 58624 644484
rect 42116 644444 42122 644456
rect 58618 644444 58624 644456
rect 58676 644444 58682 644496
rect 674788 643764 674794 643816
rect 674846 643764 674852 643816
rect 35802 643492 35808 643544
rect 35860 643532 35866 643544
rect 41138 643532 41144 643544
rect 35860 643504 41144 643532
rect 35860 643492 35866 643504
rect 41138 643492 41144 643504
rect 41196 643492 41202 643544
rect 674806 643396 674834 643764
rect 674926 643396 674932 643408
rect 674806 643368 674932 643396
rect 674926 643356 674932 643368
rect 674984 643356 674990 643408
rect 41690 643328 41696 643340
rect 41386 643300 41696 643328
rect 35526 643220 35532 643272
rect 35584 643260 35590 643272
rect 41386 643260 41414 643300
rect 41690 643288 41696 643300
rect 41748 643288 41754 643340
rect 42058 643288 42064 643340
rect 42116 643328 42122 643340
rect 43622 643328 43628 643340
rect 42116 643300 43628 643328
rect 42116 643288 42122 643300
rect 43622 643288 43628 643300
rect 43680 643288 43686 643340
rect 35584 643232 41414 643260
rect 35584 643220 35590 643232
rect 35342 643084 35348 643136
rect 35400 643124 35406 643136
rect 41690 643124 41696 643136
rect 35400 643096 41696 643124
rect 35400 643084 35406 643096
rect 41690 643084 41696 643096
rect 41748 643084 41754 643136
rect 42058 643084 42064 643136
rect 42116 643124 42122 643136
rect 61378 643124 61384 643136
rect 42116 643096 61384 643124
rect 42116 643084 42122 643096
rect 61378 643084 61384 643096
rect 61436 643084 61442 643136
rect 655330 643084 655336 643136
rect 655388 643124 655394 643136
rect 671246 643124 671252 643136
rect 655388 643096 671252 643124
rect 655388 643084 655394 643096
rect 671246 643084 671252 643096
rect 671304 643084 671310 643136
rect 38562 642472 38568 642524
rect 38620 642512 38626 642524
rect 41690 642512 41696 642524
rect 38620 642484 41696 642512
rect 38620 642472 38626 642484
rect 41690 642472 41696 642484
rect 41748 642472 41754 642524
rect 42058 642336 42064 642388
rect 42116 642376 42122 642388
rect 62942 642376 62948 642388
rect 42116 642348 62948 642376
rect 42116 642336 42122 642348
rect 62942 642336 62948 642348
rect 63000 642336 63006 642388
rect 651466 642336 651472 642388
rect 651524 642376 651530 642388
rect 658918 642376 658924 642388
rect 651524 642348 658924 642376
rect 651524 642336 651530 642348
rect 658918 642336 658924 642348
rect 658976 642336 658982 642388
rect 35802 642132 35808 642184
rect 35860 642172 35866 642184
rect 39390 642172 39396 642184
rect 35860 642144 39396 642172
rect 35860 642132 35866 642144
rect 39390 642132 39396 642144
rect 39448 642132 39454 642184
rect 41690 641968 41696 641980
rect 41386 641940 41696 641968
rect 35434 641860 35440 641912
rect 35492 641900 35498 641912
rect 41386 641900 41414 641940
rect 41690 641928 41696 641940
rect 41748 641928 41754 641980
rect 42058 641928 42064 641980
rect 42116 641968 42122 641980
rect 43070 641968 43076 641980
rect 42116 641940 43076 641968
rect 42116 641928 42122 641940
rect 43070 641928 43076 641940
rect 43128 641928 43134 641980
rect 35492 641872 41414 641900
rect 35492 641860 35498 641872
rect 35618 641724 35624 641776
rect 35676 641764 35682 641776
rect 41690 641764 41696 641776
rect 35676 641736 41696 641764
rect 35676 641724 35682 641736
rect 41690 641724 41696 641736
rect 41748 641724 41754 641776
rect 42058 641724 42064 641776
rect 42116 641764 42122 641776
rect 45278 641764 45284 641776
rect 42116 641736 45284 641764
rect 42116 641724 42122 641736
rect 45278 641724 45284 641736
rect 45336 641724 45342 641776
rect 42058 640908 42064 640960
rect 42116 640948 42122 640960
rect 45094 640948 45100 640960
rect 42116 640920 45100 640948
rect 42116 640908 42122 640920
rect 45094 640908 45100 640920
rect 45152 640908 45158 640960
rect 35802 640772 35808 640824
rect 35860 640812 35866 640824
rect 35860 640772 35894 640812
rect 35866 640608 35894 640772
rect 40862 640608 40868 640620
rect 35866 640580 40868 640608
rect 40862 640568 40868 640580
rect 40920 640568 40926 640620
rect 35618 640432 35624 640484
rect 35676 640472 35682 640484
rect 41690 640472 41696 640484
rect 35676 640444 41696 640472
rect 35676 640432 35682 640444
rect 41690 640432 41696 640444
rect 41748 640432 41754 640484
rect 675202 640472 675208 640484
rect 675036 640444 675208 640472
rect 35802 640296 35808 640348
rect 35860 640336 35866 640348
rect 41690 640336 41696 640348
rect 35860 640308 41696 640336
rect 35860 640296 35866 640308
rect 41690 640296 41696 640308
rect 41748 640296 41754 640348
rect 42058 640296 42064 640348
rect 42116 640336 42122 640348
rect 45370 640336 45376 640348
rect 42116 640308 45376 640336
rect 42116 640296 42122 640308
rect 45370 640296 45376 640308
rect 45428 640296 45434 640348
rect 651466 640296 651472 640348
rect 651524 640336 651530 640348
rect 668578 640336 668584 640348
rect 651524 640308 668584 640336
rect 651524 640296 651530 640308
rect 668578 640296 668584 640308
rect 668636 640296 668642 640348
rect 675036 640144 675064 640444
rect 675202 640432 675208 640444
rect 675260 640432 675266 640484
rect 651374 640092 651380 640144
rect 651432 640132 651438 640144
rect 653398 640132 653404 640144
rect 651432 640104 653404 640132
rect 651432 640092 651438 640104
rect 653398 640092 653404 640104
rect 653456 640092 653462 640144
rect 675018 640092 675024 640144
rect 675076 640092 675082 640144
rect 35802 639208 35808 639260
rect 35860 639248 35866 639260
rect 41690 639248 41696 639260
rect 35860 639220 41696 639248
rect 35860 639208 35866 639220
rect 41690 639208 41696 639220
rect 41748 639208 41754 639260
rect 35526 639072 35532 639124
rect 35584 639112 35590 639124
rect 39298 639112 39304 639124
rect 35584 639084 39304 639112
rect 35584 639072 35590 639084
rect 39298 639072 39304 639084
rect 39356 639072 39362 639124
rect 651650 638868 651656 638920
rect 651708 638908 651714 638920
rect 655330 638908 655336 638920
rect 651708 638880 655336 638908
rect 651708 638868 651714 638880
rect 655330 638868 655336 638880
rect 655388 638868 655394 638920
rect 651466 638732 651472 638784
rect 651524 638772 651530 638784
rect 655514 638772 655520 638784
rect 651524 638744 655520 638772
rect 651524 638732 651530 638744
rect 655514 638732 655520 638744
rect 655572 638732 655578 638784
rect 34422 638188 34428 638240
rect 34480 638228 34486 638240
rect 41690 638228 41696 638240
rect 34480 638200 41696 638228
rect 34480 638188 34486 638200
rect 41690 638188 41696 638200
rect 41748 638188 41754 638240
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 36538 637616 36544 637628
rect 35860 637588 36544 637616
rect 35860 637576 35866 637588
rect 36538 637576 36544 637588
rect 36596 637576 36602 637628
rect 674466 636964 674472 637016
rect 674524 637004 674530 637016
rect 683206 637004 683212 637016
rect 674524 636976 683212 637004
rect 674524 636964 674530 636976
rect 683206 636964 683212 636976
rect 683264 636964 683270 637016
rect 35618 636896 35624 636948
rect 35676 636936 35682 636948
rect 40586 636936 40592 636948
rect 35676 636908 40592 636936
rect 35676 636896 35682 636908
rect 40586 636896 40592 636908
rect 40644 636896 40650 636948
rect 674282 636828 674288 636880
rect 674340 636868 674346 636880
rect 683390 636868 683396 636880
rect 674340 636840 683396 636868
rect 674340 636828 674346 636840
rect 683390 636828 683396 636840
rect 683448 636828 683454 636880
rect 35802 636692 35808 636744
rect 35860 636732 35866 636744
rect 35860 636692 35894 636732
rect 35866 636664 35894 636692
rect 35866 636636 38654 636664
rect 38626 636596 38654 636636
rect 40034 636596 40040 636608
rect 38626 636568 40040 636596
rect 40034 636556 40040 636568
rect 40092 636556 40098 636608
rect 39574 636460 39580 636472
rect 36004 636432 39580 636460
rect 35802 636352 35808 636404
rect 35860 636392 35866 636404
rect 36004 636392 36032 636432
rect 39574 636420 39580 636432
rect 39632 636420 39638 636472
rect 35860 636364 36032 636392
rect 35860 636352 35866 636364
rect 35526 636216 35532 636268
rect 35584 636256 35590 636268
rect 35584 636228 38654 636256
rect 35584 636216 35590 636228
rect 38626 636188 38654 636228
rect 39114 636188 39120 636200
rect 38626 636160 39120 636188
rect 39114 636148 39120 636160
rect 39172 636148 39178 636200
rect 674926 635468 674932 635520
rect 674984 635508 674990 635520
rect 675662 635508 675668 635520
rect 674984 635480 675668 635508
rect 674984 635468 674990 635480
rect 675662 635468 675668 635480
rect 675720 635468 675726 635520
rect 35802 634924 35808 634976
rect 35860 634964 35866 634976
rect 40126 634964 40132 634976
rect 35860 634936 40132 634964
rect 35860 634924 35866 634936
rect 40126 634924 40132 634936
rect 40184 634924 40190 634976
rect 652018 634040 652024 634092
rect 652076 634080 652082 634092
rect 660298 634080 660304 634092
rect 652076 634052 660304 634080
rect 652076 634040 652082 634052
rect 660298 634040 660304 634052
rect 660356 634040 660362 634092
rect 35802 633836 35808 633888
rect 35860 633876 35866 633888
rect 35860 633836 35894 633876
rect 35866 633740 35894 633836
rect 40034 633740 40040 633752
rect 35866 633712 40040 633740
rect 40034 633700 40040 633712
rect 40092 633700 40098 633752
rect 35802 633428 35808 633480
rect 35860 633468 35866 633480
rect 41598 633468 41604 633480
rect 35860 633440 41604 633468
rect 35860 633428 35866 633440
rect 41598 633428 41604 633440
rect 41656 633428 41662 633480
rect 42058 633428 42064 633480
rect 42116 633468 42122 633480
rect 60182 633468 60188 633480
rect 42116 633440 60188 633468
rect 42116 633428 42122 633440
rect 60182 633428 60188 633440
rect 60240 633428 60246 633480
rect 671522 632952 671528 633004
rect 671580 632952 671586 633004
rect 671338 632924 671344 632936
rect 671172 632896 671344 632924
rect 671172 632652 671200 632896
rect 671338 632884 671344 632896
rect 671396 632884 671402 632936
rect 671338 632748 671344 632800
rect 671396 632788 671402 632800
rect 671540 632788 671568 632952
rect 671396 632760 671568 632788
rect 671396 632748 671402 632760
rect 671522 632652 671528 632664
rect 671172 632624 671528 632652
rect 671522 632612 671528 632624
rect 671580 632612 671586 632664
rect 36538 630572 36544 630624
rect 36596 630612 36602 630624
rect 41598 630612 41604 630624
rect 36596 630584 41604 630612
rect 36596 630572 36602 630584
rect 41598 630572 41604 630584
rect 41656 630572 41662 630624
rect 672442 629688 672448 629740
rect 672500 629728 672506 629740
rect 673270 629728 673276 629740
rect 672500 629700 673276 629728
rect 672500 629688 672506 629700
rect 673270 629688 673276 629700
rect 673328 629688 673334 629740
rect 35158 628668 35164 628720
rect 35216 628708 35222 628720
rect 39390 628708 39396 628720
rect 35216 628680 39396 628708
rect 35216 628668 35222 628680
rect 39390 628668 39396 628680
rect 39448 628668 39454 628720
rect 667198 626084 667204 626136
rect 667256 626124 667262 626136
rect 673270 626124 673276 626136
rect 667256 626096 673276 626124
rect 667256 626084 667262 626096
rect 673270 626084 673276 626096
rect 673328 626084 673334 626136
rect 44174 625988 44180 626000
rect 42352 625960 44180 625988
rect 42352 625184 42380 625960
rect 44174 625948 44180 625960
rect 44232 625948 44238 626000
rect 44174 625812 44180 625864
rect 44232 625852 44238 625864
rect 63126 625852 63132 625864
rect 44232 625824 63132 625852
rect 44232 625812 44238 625824
rect 63126 625812 63132 625824
rect 63184 625812 63190 625864
rect 669958 625404 669964 625456
rect 670016 625444 670022 625456
rect 673270 625444 673276 625456
rect 670016 625416 673276 625444
rect 670016 625404 670022 625416
rect 673270 625404 673276 625416
rect 673328 625404 673334 625456
rect 42334 625132 42340 625184
rect 42392 625132 42398 625184
rect 657538 625132 657544 625184
rect 657596 625172 657602 625184
rect 673270 625172 673276 625184
rect 657596 625144 673276 625172
rect 657596 625132 657602 625144
rect 673270 625132 673276 625144
rect 673328 625132 673334 625184
rect 674282 625132 674288 625184
rect 674340 625172 674346 625184
rect 676214 625172 676220 625184
rect 674340 625144 676220 625172
rect 674340 625132 674346 625144
rect 676214 625132 676220 625144
rect 676272 625132 676278 625184
rect 670234 624452 670240 624504
rect 670292 624492 670298 624504
rect 672626 624492 672632 624504
rect 670292 624464 672632 624492
rect 670292 624452 670298 624464
rect 672626 624452 672632 624464
rect 672684 624452 672690 624504
rect 669406 623908 669412 623960
rect 669464 623948 669470 623960
rect 674006 623948 674012 623960
rect 669464 623920 674012 623948
rect 669464 623908 669470 623920
rect 674006 623908 674012 623920
rect 674064 623908 674070 623960
rect 674282 623840 674288 623892
rect 674340 623880 674346 623892
rect 676214 623880 676220 623892
rect 674340 623852 676220 623880
rect 674340 623840 674346 623852
rect 676214 623840 676220 623852
rect 676272 623840 676278 623892
rect 43990 623812 43996 623824
rect 42260 623784 43996 623812
rect 42260 622872 42288 623784
rect 43990 623772 43996 623784
rect 44048 623772 44054 623824
rect 670234 623772 670240 623824
rect 670292 623812 670298 623824
rect 672626 623812 672632 623824
rect 670292 623784 672632 623812
rect 670292 623772 670298 623784
rect 672626 623772 672632 623784
rect 672684 623772 672690 623824
rect 671062 623228 671068 623280
rect 671120 623268 671126 623280
rect 672626 623268 672632 623280
rect 671120 623240 672632 623268
rect 671120 623228 671126 623240
rect 672626 623228 672632 623240
rect 672684 623228 672690 623280
rect 674650 623024 674656 623076
rect 674708 623064 674714 623076
rect 683390 623064 683396 623076
rect 674708 623036 683396 623064
rect 674708 623024 674714 623036
rect 683390 623024 683396 623036
rect 683448 623024 683454 623076
rect 42242 622820 42248 622872
rect 42300 622820 42306 622872
rect 671890 622616 671896 622668
rect 671948 622656 671954 622668
rect 671948 622628 673454 622656
rect 671948 622616 671954 622628
rect 673426 622588 673454 622628
rect 674282 622616 674288 622668
rect 674340 622656 674346 622668
rect 676030 622656 676036 622668
rect 674340 622628 676036 622656
rect 674340 622616 674346 622628
rect 676030 622616 676036 622628
rect 676088 622616 676094 622668
rect 674006 622588 674012 622600
rect 673426 622560 674012 622588
rect 674006 622548 674012 622560
rect 674064 622548 674070 622600
rect 670418 622412 670424 622464
rect 670476 622452 670482 622464
rect 672626 622452 672632 622464
rect 670476 622424 672632 622452
rect 670476 622412 670482 622424
rect 672626 622412 672632 622424
rect 672684 622412 672690 622464
rect 674282 622412 674288 622464
rect 674340 622452 674346 622464
rect 676398 622452 676404 622464
rect 674340 622424 676404 622452
rect 674340 622412 674346 622424
rect 676398 622412 676404 622424
rect 676456 622412 676462 622464
rect 674282 621392 674288 621444
rect 674340 621432 674346 621444
rect 676030 621432 676036 621444
rect 674340 621404 676036 621432
rect 674340 621392 674346 621404
rect 676030 621392 676036 621404
rect 676088 621392 676094 621444
rect 673178 621324 673184 621376
rect 673236 621364 673242 621376
rect 674006 621364 674012 621376
rect 673236 621336 674012 621364
rect 673236 621324 673242 621336
rect 674006 621324 674012 621336
rect 674064 621324 674070 621376
rect 671430 621120 671436 621172
rect 671488 621160 671494 621172
rect 673270 621160 673276 621172
rect 671488 621132 673276 621160
rect 671488 621120 671494 621132
rect 673270 621120 673276 621132
rect 673328 621120 673334 621172
rect 667658 620984 667664 621036
rect 667716 621024 667722 621036
rect 674006 621024 674012 621036
rect 667716 620996 674012 621024
rect 667716 620984 667722 620996
rect 674006 620984 674012 620996
rect 674064 620984 674070 621036
rect 670878 620780 670884 620832
rect 670936 620820 670942 620832
rect 674006 620820 674012 620832
rect 670936 620792 674012 620820
rect 670936 620780 670942 620792
rect 674006 620780 674012 620792
rect 674064 620780 674070 620832
rect 674282 620780 674288 620832
rect 674340 620820 674346 620832
rect 676214 620820 676220 620832
rect 674340 620792 676220 620820
rect 674340 620780 674346 620792
rect 676214 620780 676220 620792
rect 676272 620780 676278 620832
rect 42242 620236 42248 620288
rect 42300 620276 42306 620288
rect 42702 620276 42708 620288
rect 42300 620248 42708 620276
rect 42300 620236 42306 620248
rect 42702 620236 42708 620248
rect 42760 620236 42766 620288
rect 669774 620236 669780 620288
rect 669832 620276 669838 620288
rect 674006 620276 674012 620288
rect 669832 620248 674012 620276
rect 669832 620236 669838 620248
rect 674006 620236 674012 620248
rect 674064 620236 674070 620288
rect 674282 620100 674288 620152
rect 674340 620140 674346 620152
rect 676490 620140 676496 620152
rect 674340 620112 676496 620140
rect 674340 620100 674346 620112
rect 676490 620100 676496 620112
rect 676548 620100 676554 620152
rect 674282 619896 674288 619948
rect 674340 619936 674346 619948
rect 676214 619936 676220 619948
rect 674340 619908 676220 619936
rect 674340 619896 674346 619908
rect 676214 619896 676220 619908
rect 676272 619896 676278 619948
rect 668394 619692 668400 619744
rect 668452 619732 668458 619744
rect 674006 619732 674012 619744
rect 668452 619704 674012 619732
rect 668452 619692 668458 619704
rect 674006 619692 674012 619704
rect 674064 619692 674070 619744
rect 42242 619624 42248 619676
rect 42300 619664 42306 619676
rect 43070 619664 43076 619676
rect 42300 619636 43076 619664
rect 42300 619624 42306 619636
rect 43070 619624 43076 619636
rect 43128 619624 43134 619676
rect 672442 619556 672448 619608
rect 672500 619596 672506 619608
rect 674006 619596 674012 619608
rect 672500 619568 674012 619596
rect 672500 619556 672506 619568
rect 674006 619556 674012 619568
rect 674064 619556 674070 619608
rect 674282 619488 674288 619540
rect 674340 619528 674346 619540
rect 676214 619528 676220 619540
rect 674340 619500 676220 619528
rect 674340 619488 674346 619500
rect 676214 619488 676220 619500
rect 676272 619488 676278 619540
rect 43806 618304 43812 618316
rect 42260 618276 43812 618304
rect 42260 617364 42288 618276
rect 43806 618264 43812 618276
rect 43864 618264 43870 618316
rect 668210 617448 668216 617500
rect 668268 617488 668274 617500
rect 673270 617488 673276 617500
rect 668268 617460 673276 617488
rect 668268 617448 668274 617460
rect 673270 617448 673276 617460
rect 673328 617448 673334 617500
rect 42242 617312 42248 617364
rect 42300 617312 42306 617364
rect 674282 617108 674288 617160
rect 674340 617148 674346 617160
rect 676030 617148 676036 617160
rect 674340 617120 676036 617148
rect 674340 617108 674346 617120
rect 676030 617108 676036 617120
rect 676088 617108 676094 617160
rect 669038 616836 669044 616888
rect 669096 616876 669102 616888
rect 674006 616876 674012 616888
rect 669096 616848 674012 616876
rect 669096 616836 669102 616848
rect 674006 616836 674012 616848
rect 674064 616836 674070 616888
rect 44174 616768 44180 616820
rect 44232 616808 44238 616820
rect 62114 616808 62120 616820
rect 44232 616780 62120 616808
rect 44232 616768 44238 616780
rect 62114 616768 62120 616780
rect 62172 616768 62178 616820
rect 42150 616292 42156 616344
rect 42208 616332 42214 616344
rect 42518 616332 42524 616344
rect 42208 616304 42524 616332
rect 42208 616292 42214 616304
rect 42518 616292 42524 616304
rect 42576 616292 42582 616344
rect 670602 615612 670608 615664
rect 670660 615652 670666 615664
rect 674006 615652 674012 615664
rect 670660 615624 674012 615652
rect 670660 615612 670666 615624
rect 674006 615612 674012 615624
rect 674064 615612 674070 615664
rect 674282 615476 674288 615528
rect 674340 615516 674346 615528
rect 683114 615516 683120 615528
rect 674340 615488 683120 615516
rect 674340 615476 674346 615488
rect 683114 615476 683120 615488
rect 683172 615476 683178 615528
rect 670602 614864 670608 614916
rect 670660 614904 670666 614916
rect 674006 614904 674012 614916
rect 670660 614876 674012 614904
rect 670660 614864 670666 614876
rect 674006 614864 674012 614876
rect 674064 614864 674070 614916
rect 42702 614116 42708 614168
rect 42760 614156 42766 614168
rect 62114 614156 62120 614168
rect 42760 614128 62120 614156
rect 42760 614116 42766 614128
rect 62114 614116 62120 614128
rect 62172 614116 62178 614168
rect 43254 612620 43260 612672
rect 43312 612660 43318 612672
rect 43312 612632 43691 612660
rect 43312 612620 43318 612632
rect 42242 612348 42248 612400
rect 42300 612388 42306 612400
rect 42300 612360 43562 612388
rect 42300 612348 42306 612360
rect 43663 612306 43691 612632
rect 58618 612620 58624 612672
rect 58676 612660 58682 612672
rect 62114 612660 62120 612672
rect 58676 612632 62120 612660
rect 58676 612620 58682 612632
rect 62114 612620 62120 612632
rect 62172 612620 62178 612672
rect 43766 611992 43818 611998
rect 44910 611980 44916 611992
rect 43901 611952 44916 611980
rect 44910 611940 44916 611952
rect 44968 611940 44974 611992
rect 43766 611934 43818 611940
rect 43996 611652 44048 611658
rect 43996 611594 44048 611600
rect 44205 611572 44211 611584
rect 44114 611544 44211 611572
rect 44205 611532 44211 611544
rect 44263 611532 44269 611584
rect 653398 611328 653404 611380
rect 653456 611368 653462 611380
rect 674006 611368 674012 611380
rect 653456 611340 674012 611368
rect 653456 611328 653462 611340
rect 674006 611328 674012 611340
rect 674064 611328 674070 611380
rect 674282 611328 674288 611380
rect 674340 611368 674346 611380
rect 675386 611368 675392 611380
rect 674340 611340 675392 611368
rect 674340 611328 674346 611340
rect 675386 611328 675392 611340
rect 675444 611328 675450 611380
rect 50154 611300 50160 611312
rect 44237 611272 50160 611300
rect 50154 611260 50160 611272
rect 50212 611260 50218 611312
rect 44726 611096 44732 611108
rect 44344 611068 44732 611096
rect 44726 611056 44732 611068
rect 44784 611056 44790 611108
rect 46198 610892 46204 610904
rect 44461 610864 46204 610892
rect 46198 610852 46204 610864
rect 46256 610852 46262 610904
rect 44726 610756 44732 610768
rect 44574 610728 44732 610756
rect 44726 610716 44732 610728
rect 44784 610716 44790 610768
rect 50154 609968 50160 610020
rect 50212 610008 50218 610020
rect 61378 610008 61384 610020
rect 50212 609980 61384 610008
rect 50212 609968 50218 609980
rect 61378 609968 61384 609980
rect 61436 609968 61442 610020
rect 667658 608608 667664 608660
rect 667716 608648 667722 608660
rect 674006 608648 674012 608660
rect 667716 608620 674012 608648
rect 667716 608608 667722 608620
rect 674006 608608 674012 608620
rect 674064 608608 674070 608660
rect 674282 608608 674288 608660
rect 674340 608648 674346 608660
rect 675110 608648 675116 608660
rect 674340 608620 675116 608648
rect 674340 608608 674346 608620
rect 675110 608608 675116 608620
rect 675168 608608 675174 608660
rect 674466 603236 674472 603288
rect 674524 603276 674530 603288
rect 675110 603276 675116 603288
rect 674524 603248 675116 603276
rect 674524 603236 674530 603248
rect 675110 603236 675116 603248
rect 675168 603236 675174 603288
rect 35802 601672 35808 601724
rect 35860 601712 35866 601724
rect 36538 601712 36544 601724
rect 35860 601684 36544 601712
rect 35860 601672 35866 601684
rect 36538 601672 36544 601684
rect 36596 601672 36602 601724
rect 674006 600488 674012 600500
rect 663766 600460 674012 600488
rect 657538 600312 657544 600364
rect 657596 600352 657602 600364
rect 663766 600352 663794 600460
rect 674006 600448 674012 600460
rect 674064 600448 674070 600500
rect 657596 600324 663794 600352
rect 657596 600312 657602 600324
rect 674282 600312 674288 600364
rect 674340 600352 674346 600364
rect 675110 600352 675116 600364
rect 674340 600324 675116 600352
rect 674340 600312 674346 600324
rect 675110 600312 675116 600324
rect 675168 600312 675174 600364
rect 674650 599564 674656 599616
rect 674708 599604 674714 599616
rect 675294 599604 675300 599616
rect 674708 599576 675300 599604
rect 674708 599564 674714 599576
rect 675294 599564 675300 599576
rect 675352 599564 675358 599616
rect 674006 599536 674012 599548
rect 663766 599508 674012 599536
rect 654778 598952 654784 599004
rect 654836 598992 654842 599004
rect 663766 598992 663794 599508
rect 674006 599496 674012 599508
rect 674064 599496 674070 599548
rect 674282 599360 674288 599412
rect 674340 599400 674346 599412
rect 675294 599400 675300 599412
rect 674340 599372 675300 599400
rect 674340 599360 674346 599372
rect 675294 599360 675300 599372
rect 675352 599360 675358 599412
rect 654836 598964 663794 598992
rect 654836 598952 654842 598964
rect 675294 598408 675300 598460
rect 675352 598408 675358 598460
rect 675312 598188 675340 598408
rect 675294 598136 675300 598188
rect 675352 598136 675358 598188
rect 651466 597524 651472 597576
rect 651524 597564 651530 597576
rect 669958 597564 669964 597576
rect 651524 597536 669964 597564
rect 651524 597524 651530 597536
rect 669958 597524 669964 597536
rect 670016 597524 670022 597576
rect 42886 597388 42892 597440
rect 42944 597388 42950 597440
rect 42904 597032 42932 597388
rect 42886 596980 42892 597032
rect 42944 596980 42950 597032
rect 651466 596164 651472 596216
rect 651524 596204 651530 596216
rect 664438 596204 664444 596216
rect 651524 596176 664444 596204
rect 651524 596164 651530 596176
rect 664438 596164 664444 596176
rect 664496 596164 664502 596216
rect 40126 595756 40132 595808
rect 40184 595796 40190 595808
rect 41690 595796 41696 595808
rect 40184 595768 41696 595796
rect 40184 595756 40190 595768
rect 41690 595756 41696 595768
rect 41748 595756 41754 595808
rect 651650 595484 651656 595536
rect 651708 595524 651714 595536
rect 653398 595524 653404 595536
rect 651708 595496 653404 595524
rect 651708 595484 651714 595496
rect 653398 595484 653404 595496
rect 653456 595484 653462 595536
rect 651466 594804 651472 594856
rect 651524 594844 651530 594856
rect 661678 594844 661684 594856
rect 651524 594816 661684 594844
rect 651524 594804 651530 594816
rect 661678 594804 661684 594816
rect 661736 594804 661742 594856
rect 41322 594736 41328 594788
rect 41380 594776 41386 594788
rect 41506 594776 41512 594788
rect 41380 594748 41512 594776
rect 41380 594736 41386 594748
rect 41506 594736 41512 594748
rect 41564 594736 41570 594788
rect 651466 594668 651472 594720
rect 651524 594708 651530 594720
rect 657538 594708 657544 594720
rect 651524 594680 657544 594708
rect 651524 594668 651530 594680
rect 657538 594668 657544 594680
rect 657596 594668 657602 594720
rect 39942 594532 39948 594584
rect 40000 594572 40006 594584
rect 41690 594572 41696 594584
rect 40000 594544 41696 594572
rect 40000 594532 40006 594544
rect 41690 594532 41696 594544
rect 41748 594532 41754 594584
rect 651466 593240 651472 593292
rect 651524 593280 651530 593292
rect 654778 593280 654784 593292
rect 651524 593252 654784 593280
rect 651524 593240 651530 593252
rect 654778 593240 654784 593252
rect 654836 593240 654842 593292
rect 675294 592628 675300 592680
rect 675352 592668 675358 592680
rect 683390 592668 683396 592680
rect 675352 592640 683396 592668
rect 675352 592628 675358 592640
rect 683390 592628 683396 592640
rect 683448 592628 683454 592680
rect 40954 592492 40960 592544
rect 41012 592532 41018 592544
rect 41690 592532 41696 592544
rect 41012 592504 41696 592532
rect 41012 592492 41018 592504
rect 41690 592492 41696 592504
rect 41748 592492 41754 592544
rect 35618 590928 35624 590980
rect 35676 590968 35682 590980
rect 41690 590968 41696 590980
rect 35676 590940 41696 590968
rect 35676 590928 35682 590940
rect 41690 590928 41696 590940
rect 41748 590928 41754 590980
rect 35802 590656 35808 590708
rect 35860 590696 35866 590708
rect 39758 590696 39764 590708
rect 35860 590668 39764 590696
rect 35860 590656 35866 590668
rect 39758 590656 39764 590668
rect 39816 590656 39822 590708
rect 674834 590588 674840 590640
rect 674892 590628 674898 590640
rect 682378 590628 682384 590640
rect 674892 590600 682384 590628
rect 674892 590588 674898 590600
rect 682378 590588 682384 590600
rect 682436 590588 682442 590640
rect 674282 588548 674288 588600
rect 674340 588588 674346 588600
rect 684034 588588 684040 588600
rect 674340 588560 684040 588588
rect 674340 588548 674346 588560
rect 684034 588548 684040 588560
rect 684092 588548 684098 588600
rect 33042 587120 33048 587172
rect 33100 587160 33106 587172
rect 41506 587160 41512 587172
rect 33100 587132 41512 587160
rect 33100 587120 33106 587132
rect 41506 587120 41512 587132
rect 41564 587120 41570 587172
rect 42058 587120 42064 587172
rect 42116 587160 42122 587172
rect 42610 587160 42616 587172
rect 42116 587132 42616 587160
rect 42116 587120 42122 587132
rect 42610 587120 42616 587132
rect 42668 587120 42674 587172
rect 42058 586236 42064 586288
rect 42116 586276 42122 586288
rect 42116 586248 42472 586276
rect 42116 586236 42122 586248
rect 35158 586168 35164 586220
rect 35216 586208 35222 586220
rect 41690 586208 41696 586220
rect 35216 586180 41696 586208
rect 35216 586168 35222 586180
rect 41690 586168 41696 586180
rect 41748 586168 41754 586220
rect 42444 586140 42472 586248
rect 42794 586140 42800 586152
rect 42444 586112 42800 586140
rect 42794 586100 42800 586112
rect 42852 586100 42858 586152
rect 42242 586032 42248 586084
rect 42300 586032 42306 586084
rect 33778 585896 33784 585948
rect 33836 585936 33842 585948
rect 39850 585936 39856 585948
rect 33836 585908 39856 585936
rect 33836 585896 33842 585908
rect 39850 585896 39856 585908
rect 39908 585896 39914 585948
rect 31018 585760 31024 585812
rect 31076 585800 31082 585812
rect 40586 585800 40592 585812
rect 31076 585772 40592 585800
rect 31076 585760 31082 585772
rect 40586 585760 40592 585772
rect 40644 585760 40650 585812
rect 42260 585608 42288 586032
rect 42242 585556 42248 585608
rect 42300 585556 42306 585608
rect 660298 581000 660304 581052
rect 660356 581040 660362 581052
rect 674006 581040 674012 581052
rect 660356 581012 674012 581040
rect 660356 581000 660362 581012
rect 674006 581000 674012 581012
rect 674064 581000 674070 581052
rect 668578 579980 668584 580032
rect 668636 580020 668642 580032
rect 674006 580020 674012 580032
rect 668636 579992 674012 580020
rect 668636 579980 668642 579992
rect 674006 579980 674012 579992
rect 674064 579980 674070 580032
rect 670234 579844 670240 579896
rect 670292 579884 670298 579896
rect 674006 579884 674012 579896
rect 670292 579856 674012 579884
rect 670292 579844 670298 579856
rect 674006 579844 674012 579856
rect 674064 579844 674070 579896
rect 658918 579640 658924 579692
rect 658976 579680 658982 579692
rect 673546 579680 673552 579692
rect 658976 579652 673552 579680
rect 658976 579640 658982 579652
rect 673546 579640 673552 579652
rect 673604 579640 673610 579692
rect 670786 579368 670792 579420
rect 670844 579408 670850 579420
rect 674006 579408 674012 579420
rect 670844 579380 674012 579408
rect 670844 579368 670850 579380
rect 674006 579368 674012 579380
rect 674064 579368 674070 579420
rect 669406 579028 669412 579080
rect 669464 579068 669470 579080
rect 674006 579068 674012 579080
rect 669464 579040 674012 579068
rect 669464 579028 669470 579040
rect 674006 579028 674012 579040
rect 674064 579028 674070 579080
rect 42242 578960 42248 579012
rect 42300 579000 42306 579012
rect 43254 579000 43260 579012
rect 42300 578972 43260 579000
rect 42300 578960 42306 578972
rect 43254 578960 43260 578972
rect 43312 578960 43318 579012
rect 671154 578552 671160 578604
rect 671212 578592 671218 578604
rect 674006 578592 674012 578604
rect 671212 578564 674012 578592
rect 671212 578552 671218 578564
rect 674006 578552 674012 578564
rect 674064 578552 674070 578604
rect 670418 578144 670424 578196
rect 670476 578184 670482 578196
rect 674006 578184 674012 578196
rect 670476 578156 674012 578184
rect 670476 578144 670482 578156
rect 674006 578144 674012 578156
rect 674064 578144 674070 578196
rect 42242 577736 42248 577788
rect 42300 577776 42306 577788
rect 42794 577776 42800 577788
rect 42300 577748 42800 577776
rect 42300 577736 42306 577748
rect 42794 577736 42800 577748
rect 42852 577736 42858 577788
rect 670234 577736 670240 577788
rect 670292 577776 670298 577788
rect 674006 577776 674012 577788
rect 670292 577748 674012 577776
rect 670292 577736 670298 577748
rect 674006 577736 674012 577748
rect 674064 577736 674070 577788
rect 671430 577396 671436 577448
rect 671488 577436 671494 577448
rect 674006 577436 674012 577448
rect 671488 577408 674012 577436
rect 671488 577396 671494 577408
rect 674006 577396 674012 577408
rect 674064 577396 674070 577448
rect 669406 576920 669412 576972
rect 669464 576960 669470 576972
rect 674006 576960 674012 576972
rect 669464 576932 674012 576960
rect 669464 576920 669470 576932
rect 674006 576920 674012 576932
rect 674064 576920 674070 576972
rect 45094 575424 45100 575476
rect 45152 575464 45158 575476
rect 62114 575464 62120 575476
rect 45152 575436 62120 575464
rect 45152 575424 45158 575436
rect 62114 575424 62120 575436
rect 62172 575424 62178 575476
rect 671614 574540 671620 574592
rect 671672 574580 671678 574592
rect 673546 574580 673552 574592
rect 671672 574552 673552 574580
rect 671672 574540 671678 574552
rect 673546 574540 673552 574552
rect 673604 574540 673610 574592
rect 671982 574268 671988 574320
rect 672040 574308 672046 574320
rect 673546 574308 673552 574320
rect 672040 574280 673552 574308
rect 672040 574268 672046 574280
rect 673546 574268 673552 574280
rect 673604 574268 673610 574320
rect 667474 574064 667480 574116
rect 667532 574104 667538 574116
rect 674006 574104 674012 574116
rect 667532 574076 674012 574104
rect 667532 574064 667538 574076
rect 674006 574064 674012 574076
rect 674064 574064 674070 574116
rect 46934 573996 46940 574048
rect 46992 574036 46998 574048
rect 62114 574036 62120 574048
rect 46992 574008 62120 574036
rect 46992 573996 46998 574008
rect 62114 573996 62120 574008
rect 62172 573996 62178 574048
rect 669590 572228 669596 572280
rect 669648 572268 669654 572280
rect 674006 572268 674012 572280
rect 669648 572240 674012 572268
rect 669648 572228 669654 572240
rect 674006 572228 674012 572240
rect 674064 572228 674070 572280
rect 671798 571548 671804 571600
rect 671856 571588 671862 571600
rect 674006 571588 674012 571600
rect 671856 571560 674012 571588
rect 671856 571548 671862 571560
rect 674006 571548 674012 571560
rect 674064 571548 674070 571600
rect 674466 571548 674472 571600
rect 674524 571588 674530 571600
rect 676214 571588 676220 571600
rect 674524 571560 676220 571588
rect 674524 571548 674530 571560
rect 676214 571548 676220 571560
rect 676272 571548 676278 571600
rect 42058 570936 42064 570988
rect 42116 570976 42122 570988
rect 42610 570976 42616 570988
rect 42116 570948 42616 570976
rect 42116 570936 42122 570948
rect 42610 570936 42616 570948
rect 42668 570936 42674 570988
rect 674834 570460 674840 570512
rect 674892 570500 674898 570512
rect 675478 570500 675484 570512
rect 674892 570472 675484 570500
rect 674892 570460 674898 570472
rect 675478 570460 675484 570472
rect 675536 570500 675542 570512
rect 683114 570500 683120 570512
rect 675536 570472 683120 570500
rect 675536 570460 675542 570472
rect 683114 570460 683120 570472
rect 683172 570460 683178 570512
rect 671338 570392 671344 570444
rect 671396 570432 671402 570444
rect 673546 570432 673552 570444
rect 671396 570404 673552 570432
rect 671396 570392 671402 570404
rect 673546 570392 673552 570404
rect 673604 570392 673610 570444
rect 671982 570120 671988 570172
rect 672040 570160 672046 570172
rect 674006 570160 674012 570172
rect 672040 570132 674012 570160
rect 672040 570120 672046 570132
rect 674006 570120 674012 570132
rect 674064 570120 674070 570172
rect 669774 568556 669780 568608
rect 669832 568596 669838 568608
rect 674006 568596 674012 568608
rect 669832 568568 674012 568596
rect 669832 568556 669838 568568
rect 674006 568556 674012 568568
rect 674064 568556 674070 568608
rect 653398 565836 653404 565888
rect 653456 565876 653462 565888
rect 673546 565876 673552 565888
rect 653456 565848 673552 565876
rect 653456 565836 653462 565848
rect 673546 565836 673552 565848
rect 673604 565836 673610 565888
rect 665082 564408 665088 564460
rect 665140 564448 665146 564460
rect 673546 564448 673552 564460
rect 665140 564420 673552 564448
rect 665140 564408 665146 564420
rect 673546 564408 673552 564420
rect 673604 564408 673610 564460
rect 35802 557540 35808 557592
rect 35860 557580 35866 557592
rect 40954 557580 40960 557592
rect 35860 557552 40960 557580
rect 35860 557540 35866 557552
rect 40954 557540 40960 557552
rect 41012 557540 41018 557592
rect 35802 555024 35808 555076
rect 35860 555064 35866 555076
rect 40494 555064 40500 555076
rect 35860 555036 40500 555064
rect 35860 555024 35866 555036
rect 40494 555024 40500 555036
rect 40552 555024 40558 555076
rect 35802 554752 35808 554804
rect 35860 554792 35866 554804
rect 39850 554792 39856 554804
rect 35860 554764 39856 554792
rect 35860 554752 35866 554764
rect 39850 554752 39856 554764
rect 39908 554752 39914 554804
rect 657814 554752 657820 554804
rect 657872 554792 657878 554804
rect 673546 554792 673552 554804
rect 657872 554764 673552 554792
rect 657872 554752 657878 554764
rect 673546 554752 673552 554764
rect 673604 554752 673610 554804
rect 35618 553528 35624 553580
rect 35676 553568 35682 553580
rect 41690 553568 41696 553580
rect 35676 553540 41696 553568
rect 35676 553528 35682 553540
rect 41690 553528 41696 553540
rect 41748 553528 41754 553580
rect 35802 553392 35808 553444
rect 35860 553432 35866 553444
rect 41322 553432 41328 553444
rect 35860 553404 41328 553432
rect 35860 553392 35866 553404
rect 41322 553392 41328 553404
rect 41380 553392 41386 553444
rect 655146 553392 655152 553444
rect 655204 553432 655210 553444
rect 670418 553432 670424 553444
rect 655204 553404 670424 553432
rect 655204 553392 655210 553404
rect 670418 553392 670424 553404
rect 670476 553392 670482 553444
rect 651466 552644 651472 552696
rect 651524 552684 651530 552696
rect 665818 552684 665824 552696
rect 651524 552656 665824 552684
rect 651524 552644 651530 552656
rect 665818 552644 665824 552656
rect 665876 552644 665882 552696
rect 41322 552032 41328 552084
rect 41380 552072 41386 552084
rect 41690 552072 41696 552084
rect 41380 552044 41696 552072
rect 41380 552032 41386 552044
rect 41690 552032 41696 552044
rect 41748 552032 41754 552084
rect 675202 551760 675208 551812
rect 675260 551760 675266 551812
rect 675220 551608 675248 551760
rect 675202 551556 675208 551608
rect 675260 551556 675266 551608
rect 41138 550604 41144 550656
rect 41196 550644 41202 550656
rect 41690 550644 41696 550656
rect 41196 550616 41696 550644
rect 41196 550604 41202 550616
rect 41690 550604 41696 550616
rect 41748 550604 41754 550656
rect 42058 550604 42064 550656
rect 42116 550644 42122 550656
rect 42978 550644 42984 550656
rect 42116 550616 42984 550644
rect 42116 550604 42122 550616
rect 42978 550604 42984 550616
rect 43036 550604 43042 550656
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 660298 550644 660304 550656
rect 651524 550616 660304 550644
rect 651524 550604 651530 550616
rect 660298 550604 660304 550616
rect 660356 550604 660362 550656
rect 651374 550332 651380 550384
rect 651432 550372 651438 550384
rect 653398 550372 653404 550384
rect 651432 550344 653404 550372
rect 651432 550332 651438 550344
rect 653398 550332 653404 550344
rect 653456 550332 653462 550384
rect 40862 550196 40868 550248
rect 40920 550236 40926 550248
rect 41690 550236 41696 550248
rect 40920 550208 41696 550236
rect 40920 550196 40926 550208
rect 41690 550196 41696 550208
rect 41748 550196 41754 550248
rect 651650 549856 651656 549908
rect 651708 549896 651714 549908
rect 663058 549896 663064 549908
rect 651708 549868 663064 549896
rect 651708 549856 651714 549868
rect 663058 549856 663064 549868
rect 663116 549856 663122 549908
rect 675294 549488 675300 549500
rect 675128 549460 675300 549488
rect 651466 549176 651472 549228
rect 651524 549216 651530 549228
rect 657814 549216 657820 549228
rect 651524 549188 657820 549216
rect 651524 549176 651530 549188
rect 657814 549176 657820 549188
rect 657872 549176 657878 549228
rect 675128 548944 675156 549460
rect 675294 549448 675300 549460
rect 675352 549448 675358 549500
rect 675036 548916 675156 548944
rect 675036 548820 675064 548916
rect 651466 548768 651472 548820
rect 651524 548808 651530 548820
rect 655146 548808 655152 548820
rect 651524 548780 655152 548808
rect 651524 548768 651530 548780
rect 655146 548768 655152 548780
rect 655204 548768 655210 548820
rect 675018 548768 675024 548820
rect 675076 548768 675082 548820
rect 41322 547884 41328 547936
rect 41380 547924 41386 547936
rect 41690 547924 41696 547936
rect 41380 547896 41696 547924
rect 41380 547884 41386 547896
rect 41690 547884 41696 547896
rect 41748 547884 41754 547936
rect 29638 547136 29644 547188
rect 29696 547176 29702 547188
rect 41690 547176 41696 547188
rect 29696 547148 41696 547176
rect 29696 547136 29702 547148
rect 41690 547136 41696 547148
rect 41748 547136 41754 547188
rect 675570 547136 675576 547188
rect 675628 547176 675634 547188
rect 683206 547176 683212 547188
rect 675628 547148 683212 547176
rect 675628 547136 675634 547148
rect 683206 547136 683212 547148
rect 683264 547136 683270 547188
rect 674834 545844 674840 545896
rect 674892 545884 674898 545896
rect 682378 545884 682384 545896
rect 674892 545856 682384 545884
rect 674892 545844 674898 545856
rect 682378 545844 682384 545856
rect 682436 545844 682442 545896
rect 673914 540880 673920 540932
rect 673972 540880 673978 540932
rect 673730 540608 673736 540660
rect 673788 540648 673794 540660
rect 673932 540648 673960 540880
rect 673788 540620 673960 540648
rect 673788 540608 673794 540620
rect 669958 535780 669964 535832
rect 670016 535820 670022 535832
rect 674006 535820 674012 535832
rect 670016 535792 674012 535820
rect 670016 535780 670022 535792
rect 674006 535780 674012 535792
rect 674064 535780 674070 535832
rect 674282 535712 674288 535764
rect 674340 535752 674346 535764
rect 676030 535752 676036 535764
rect 674340 535724 676036 535752
rect 674340 535712 674346 535724
rect 676030 535712 676036 535724
rect 676088 535712 676094 535764
rect 674282 535508 674288 535560
rect 674340 535548 674346 535560
rect 676214 535548 676220 535560
rect 674340 535520 676220 535548
rect 674340 535508 674346 535520
rect 676214 535508 676220 535520
rect 676272 535508 676278 535560
rect 664438 535440 664444 535492
rect 664496 535480 664502 535492
rect 674006 535480 674012 535492
rect 664496 535452 674012 535480
rect 664496 535440 664502 535452
rect 674006 535440 674012 535452
rect 674064 535440 674070 535492
rect 670786 534964 670792 535016
rect 670844 535004 670850 535016
rect 674006 535004 674012 535016
rect 670844 534976 674012 535004
rect 670844 534964 670850 534976
rect 674006 534964 674012 534976
rect 674064 534964 674070 535016
rect 674282 534896 674288 534948
rect 674340 534936 674346 534948
rect 676030 534936 676036 534948
rect 674340 534908 676036 534936
rect 674340 534896 674346 534908
rect 676030 534896 676036 534908
rect 676088 534896 676094 534948
rect 674282 534420 674288 534472
rect 674340 534460 674346 534472
rect 676030 534460 676036 534472
rect 674340 534432 676036 534460
rect 674340 534420 674346 534432
rect 676030 534420 676036 534432
rect 676088 534420 676094 534472
rect 670786 534352 670792 534404
rect 670844 534392 670850 534404
rect 674006 534392 674012 534404
rect 670844 534364 674012 534392
rect 670844 534352 670850 534364
rect 674006 534352 674012 534364
rect 674064 534352 674070 534404
rect 674282 534284 674288 534336
rect 674340 534324 674346 534336
rect 676214 534324 676220 534336
rect 674340 534296 676220 534324
rect 674340 534284 674346 534296
rect 676214 534284 676220 534296
rect 676272 534284 676278 534336
rect 661678 534216 661684 534268
rect 661736 534256 661742 534268
rect 674006 534256 674012 534268
rect 661736 534228 674012 534256
rect 661736 534216 661742 534228
rect 674006 534216 674012 534228
rect 674064 534216 674070 534268
rect 671154 534080 671160 534132
rect 671212 534120 671218 534132
rect 674006 534120 674012 534132
rect 671212 534092 674012 534120
rect 671212 534080 671218 534092
rect 674006 534080 674012 534092
rect 674064 534080 674070 534132
rect 674282 534080 674288 534132
rect 674340 534120 674346 534132
rect 676030 534120 676036 534132
rect 674340 534092 676036 534120
rect 674340 534080 674346 534092
rect 676030 534080 676036 534092
rect 676088 534080 676094 534132
rect 674282 533332 674288 533384
rect 674340 533372 674346 533384
rect 683574 533372 683580 533384
rect 674340 533344 683580 533372
rect 674340 533332 674346 533344
rect 683574 533332 683580 533344
rect 683632 533332 683638 533384
rect 671614 533060 671620 533112
rect 671672 533100 671678 533112
rect 674006 533100 674012 533112
rect 671672 533072 674012 533100
rect 671672 533060 671678 533072
rect 674006 533060 674012 533072
rect 674064 533060 674070 533112
rect 674282 533060 674288 533112
rect 674340 533100 674346 533112
rect 676214 533100 676220 533112
rect 674340 533072 676220 533100
rect 674340 533060 674346 533072
rect 676214 533060 676220 533072
rect 676272 533060 676278 533112
rect 674282 532924 674288 532976
rect 674340 532964 674346 532976
rect 676030 532964 676036 532976
rect 674340 532936 676036 532964
rect 674340 532924 674346 532936
rect 676030 532924 676036 532936
rect 676088 532924 676094 532976
rect 670234 532856 670240 532908
rect 670292 532896 670298 532908
rect 674006 532896 674012 532908
rect 670292 532868 674012 532896
rect 670292 532856 670298 532868
rect 674006 532856 674012 532868
rect 674064 532856 674070 532908
rect 674282 532788 674288 532840
rect 674340 532828 674346 532840
rect 676398 532828 676404 532840
rect 674340 532800 676404 532828
rect 674340 532788 674346 532800
rect 676398 532788 676404 532800
rect 676456 532788 676462 532840
rect 672718 532720 672724 532772
rect 672776 532760 672782 532772
rect 674006 532760 674012 532772
rect 672776 532732 674012 532760
rect 672776 532720 672782 532732
rect 674006 532720 674012 532732
rect 674064 532720 674070 532772
rect 674282 532176 674288 532228
rect 674340 532216 674346 532228
rect 676398 532216 676404 532228
rect 674340 532188 676404 532216
rect 674340 532176 674346 532188
rect 676398 532176 676404 532188
rect 676456 532176 676462 532228
rect 667658 532108 667664 532160
rect 667716 532148 667722 532160
rect 674006 532148 674012 532160
rect 667716 532120 674012 532148
rect 667716 532108 667722 532120
rect 674006 532108 674012 532120
rect 674064 532108 674070 532160
rect 674282 532040 674288 532092
rect 674340 532080 674346 532092
rect 676214 532080 676220 532092
rect 674340 532052 676220 532080
rect 674340 532040 674346 532052
rect 676214 532040 676220 532052
rect 676272 532040 676278 532092
rect 44726 531972 44732 532024
rect 44784 532012 44790 532024
rect 62114 532012 62120 532024
rect 44784 531984 62120 532012
rect 44784 531972 44790 531984
rect 62114 531972 62120 531984
rect 62172 531972 62178 532024
rect 674006 531972 674012 532024
rect 674064 531972 674070 532024
rect 669406 531564 669412 531616
rect 669464 531604 669470 531616
rect 674024 531604 674052 531972
rect 674282 531700 674288 531752
rect 674340 531740 674346 531752
rect 676030 531740 676036 531752
rect 674340 531712 676036 531740
rect 674340 531700 674346 531712
rect 676030 531700 676036 531712
rect 676088 531700 676094 531752
rect 669464 531576 674052 531604
rect 669464 531564 669470 531576
rect 671154 531428 671160 531480
rect 671212 531468 671218 531480
rect 674006 531468 674012 531480
rect 671212 531440 674012 531468
rect 671212 531428 671218 531440
rect 674006 531428 674012 531440
rect 674064 531428 674070 531480
rect 51718 531224 51724 531276
rect 51776 531264 51782 531276
rect 62298 531264 62304 531276
rect 51776 531236 62304 531264
rect 51776 531224 51782 531236
rect 62298 531224 62304 531236
rect 62356 531224 62362 531276
rect 42150 530680 42156 530732
rect 42208 530720 42214 530732
rect 42702 530720 42708 530732
rect 42208 530692 42708 530720
rect 42208 530680 42214 530692
rect 42702 530680 42708 530692
rect 42760 530680 42766 530732
rect 42242 530272 42248 530324
rect 42300 530312 42306 530324
rect 42702 530312 42708 530324
rect 42300 530284 42708 530312
rect 42300 530272 42306 530284
rect 42702 530272 42708 530284
rect 42760 530272 42766 530324
rect 667290 529932 667296 529984
rect 667348 529972 667354 529984
rect 674006 529972 674012 529984
rect 667348 529944 674012 529972
rect 667348 529932 667354 529944
rect 674006 529932 674012 529944
rect 674064 529932 674070 529984
rect 674282 529932 674288 529984
rect 674340 529972 674346 529984
rect 676030 529972 676036 529984
rect 674340 529944 676036 529972
rect 674340 529932 674346 529944
rect 676030 529932 676036 529944
rect 676088 529932 676094 529984
rect 674282 529320 674288 529372
rect 674340 529360 674346 529372
rect 676214 529360 676220 529372
rect 674340 529332 676220 529360
rect 674340 529320 674346 529332
rect 676214 529320 676220 529332
rect 676272 529320 676278 529372
rect 668946 529116 668952 529168
rect 669004 529156 669010 529168
rect 674006 529156 674012 529168
rect 669004 529128 674012 529156
rect 669004 529116 669010 529128
rect 674006 529116 674012 529128
rect 674064 529116 674070 529168
rect 674282 528980 674288 529032
rect 674340 529020 674346 529032
rect 676214 529020 676220 529032
rect 674340 528992 676220 529020
rect 674340 528980 674346 528992
rect 676214 528980 676220 528992
rect 676272 528980 676278 529032
rect 670970 528912 670976 528964
rect 671028 528952 671034 528964
rect 674006 528952 674012 528964
rect 671028 528924 674012 528952
rect 671028 528912 671034 528924
rect 674006 528912 674012 528924
rect 674064 528912 674070 528964
rect 672350 528708 672356 528760
rect 672408 528748 672414 528760
rect 674006 528748 674012 528760
rect 672408 528720 674012 528748
rect 672408 528708 672414 528720
rect 674006 528708 674012 528720
rect 674064 528708 674070 528760
rect 674282 528708 674288 528760
rect 674340 528748 674346 528760
rect 676030 528748 676036 528760
rect 674340 528720 676036 528748
rect 674340 528708 674346 528720
rect 676030 528708 676036 528720
rect 676088 528708 676094 528760
rect 44818 528572 44824 528624
rect 44876 528612 44882 528624
rect 62114 528612 62120 528624
rect 44876 528584 62120 528612
rect 44876 528572 44882 528584
rect 62114 528572 62120 528584
rect 62172 528572 62178 528624
rect 672534 528096 672540 528148
rect 672592 528136 672598 528148
rect 673362 528136 673368 528148
rect 672592 528108 673368 528136
rect 672592 528096 672598 528108
rect 673362 528096 673368 528108
rect 673420 528096 673426 528148
rect 47578 527076 47584 527128
rect 47636 527116 47642 527128
rect 62114 527116 62120 527128
rect 47636 527088 62120 527116
rect 47636 527076 47642 527088
rect 62114 527076 62120 527088
rect 62172 527076 62178 527128
rect 674650 526736 674656 526788
rect 674708 526776 674714 526788
rect 676030 526776 676036 526788
rect 674708 526748 676036 526776
rect 674708 526736 674714 526748
rect 676030 526736 676036 526748
rect 676088 526736 676094 526788
rect 674282 526328 674288 526380
rect 674340 526368 674346 526380
rect 676030 526368 676036 526380
rect 674340 526340 676036 526368
rect 674340 526328 674346 526340
rect 676030 526328 676036 526340
rect 676088 526328 676094 526380
rect 662414 525036 662420 525088
rect 662472 525076 662478 525088
rect 668762 525076 668768 525088
rect 662472 525048 668768 525076
rect 662472 525036 662478 525048
rect 668762 525036 668768 525048
rect 668820 525076 668826 525088
rect 674006 525076 674012 525088
rect 668820 525048 674012 525076
rect 668820 525036 668826 525048
rect 674006 525036 674012 525048
rect 674064 525036 674070 525088
rect 674282 524560 674288 524612
rect 674340 524600 674346 524612
rect 683114 524600 683120 524612
rect 674340 524572 683120 524600
rect 674340 524560 674346 524572
rect 683114 524560 683120 524572
rect 683172 524560 683178 524612
rect 658918 521976 658924 522028
rect 658976 522016 658982 522028
rect 662414 522016 662420 522028
rect 658976 521988 662420 522016
rect 658976 521976 658982 521988
rect 662414 521976 662420 521988
rect 662472 521976 662478 522028
rect 675478 520208 675484 520260
rect 675536 520248 675542 520260
rect 678974 520248 678980 520260
rect 675536 520220 678980 520248
rect 675536 520208 675542 520220
rect 678974 520208 678980 520220
rect 679032 520208 679038 520260
rect 675662 518780 675668 518832
rect 675720 518820 675726 518832
rect 677870 518820 677876 518832
rect 675720 518792 677876 518820
rect 675720 518780 675726 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 656158 512864 656164 512916
rect 656216 512904 656222 512916
rect 658918 512904 658924 512916
rect 656216 512876 658924 512904
rect 656216 512864 656222 512876
rect 658918 512864 658924 512876
rect 658976 512864 658982 512916
rect 675110 503616 675116 503668
rect 675168 503656 675174 503668
rect 679618 503656 679624 503668
rect 675168 503628 679624 503656
rect 675168 503616 675174 503628
rect 679618 503616 679624 503628
rect 679676 503616 679682 503668
rect 675294 503480 675300 503532
rect 675352 503520 675358 503532
rect 680998 503520 681004 503532
rect 675352 503492 681004 503520
rect 675352 503480 675358 503492
rect 680998 503480 681004 503492
rect 681056 503480 681062 503532
rect 674926 500896 674932 500948
rect 674984 500936 674990 500948
rect 681182 500936 681188 500948
rect 674984 500908 681188 500936
rect 674984 500896 674990 500908
rect 681182 500896 681188 500908
rect 681240 500896 681246 500948
rect 650638 499536 650644 499588
rect 650696 499576 650702 499588
rect 656158 499576 656164 499588
rect 650696 499548 656164 499576
rect 650696 499536 650702 499548
rect 656158 499536 656164 499548
rect 656216 499536 656222 499588
rect 674282 494980 674288 495032
rect 674340 495020 674346 495032
rect 674650 495020 674656 495032
rect 674340 494992 674656 495020
rect 674340 494980 674346 494992
rect 674650 494980 674656 494992
rect 674708 494980 674714 495032
rect 674282 491648 674288 491700
rect 674340 491688 674346 491700
rect 676030 491688 676036 491700
rect 674340 491660 676036 491688
rect 674340 491648 674346 491660
rect 676030 491648 676036 491660
rect 676088 491648 676094 491700
rect 665818 491580 665824 491632
rect 665876 491620 665882 491632
rect 674006 491620 674012 491632
rect 665876 491592 674012 491620
rect 665876 491580 665882 491592
rect 674006 491580 674012 491592
rect 674064 491580 674070 491632
rect 663058 491444 663064 491496
rect 663116 491484 663122 491496
rect 673822 491484 673828 491496
rect 663116 491456 673828 491484
rect 663116 491444 663122 491456
rect 673822 491444 673828 491456
rect 673880 491444 673886 491496
rect 660298 491308 660304 491360
rect 660356 491348 660362 491360
rect 674006 491348 674012 491360
rect 660356 491320 674012 491348
rect 660356 491308 660362 491320
rect 674006 491308 674012 491320
rect 674064 491308 674070 491360
rect 670786 490900 670792 490952
rect 670844 490940 670850 490952
rect 674006 490940 674012 490952
rect 670844 490912 674012 490940
rect 670844 490900 670850 490912
rect 674006 490900 674012 490912
rect 674064 490900 674070 490952
rect 672626 489880 672632 489932
rect 672684 489920 672690 489932
rect 673362 489920 673368 489932
rect 672684 489892 673368 489920
rect 672684 489880 672690 489892
rect 673362 489880 673368 489892
rect 673420 489880 673426 489932
rect 672442 489608 672448 489660
rect 672500 489648 672506 489660
rect 674006 489648 674012 489660
rect 672500 489620 674012 489648
rect 672500 489608 672506 489620
rect 674006 489608 674012 489620
rect 674064 489608 674070 489660
rect 671614 489268 671620 489320
rect 671672 489308 671678 489320
rect 674006 489308 674012 489320
rect 671672 489280 674012 489308
rect 671672 489268 671678 489280
rect 674006 489268 674012 489280
rect 674064 489268 674070 489320
rect 671154 488452 671160 488504
rect 671212 488492 671218 488504
rect 674006 488492 674012 488504
rect 671212 488464 674012 488492
rect 671212 488452 671218 488464
rect 674006 488452 674012 488464
rect 674064 488452 674070 488504
rect 674282 486752 674288 486804
rect 674340 486792 674346 486804
rect 676030 486792 676036 486804
rect 674340 486764 676036 486792
rect 674340 486752 674346 486764
rect 676030 486752 676036 486764
rect 676088 486752 676094 486804
rect 665082 485800 665088 485852
rect 665140 485840 665146 485852
rect 674006 485840 674012 485852
rect 665140 485812 674012 485840
rect 665140 485800 665146 485812
rect 674006 485800 674012 485812
rect 674064 485800 674070 485852
rect 674282 485120 674288 485172
rect 674340 485160 674346 485172
rect 676030 485160 676036 485172
rect 674340 485132 676036 485160
rect 674340 485120 674346 485132
rect 676030 485120 676036 485132
rect 676088 485120 676094 485172
rect 668578 484372 668584 484424
rect 668636 484412 668642 484424
rect 674006 484412 674012 484424
rect 668636 484384 674012 484412
rect 668636 484372 668642 484384
rect 674006 484372 674012 484384
rect 674064 484372 674070 484424
rect 674466 483964 674472 484016
rect 674524 484004 674530 484016
rect 676030 484004 676036 484016
rect 674524 483976 676036 484004
rect 674524 483964 674530 483976
rect 676030 483964 676036 483976
rect 676088 483964 676094 484016
rect 671798 483148 671804 483200
rect 671856 483188 671862 483200
rect 674006 483188 674012 483200
rect 671856 483160 674012 483188
rect 671856 483148 671862 483160
rect 674006 483148 674012 483160
rect 674064 483148 674070 483200
rect 676214 482944 676220 482996
rect 676272 482984 676278 482996
rect 677410 482984 677416 482996
rect 676272 482956 677416 482984
rect 676272 482944 676278 482956
rect 677410 482944 677416 482956
rect 677468 482944 677474 482996
rect 670418 480360 670424 480412
rect 670476 480400 670482 480412
rect 674006 480400 674012 480412
rect 670476 480372 674012 480400
rect 670476 480360 670482 480372
rect 674006 480360 674012 480372
rect 674064 480360 674070 480412
rect 674282 480360 674288 480412
rect 674340 480400 674346 480412
rect 683114 480400 683120 480412
rect 674340 480372 683120 480400
rect 674340 480360 674346 480372
rect 683114 480360 683120 480372
rect 683172 480360 683178 480412
rect 667474 477504 667480 477556
rect 667532 477544 667538 477556
rect 670418 477544 670424 477556
rect 667532 477516 670424 477544
rect 667532 477504 667538 477516
rect 670418 477504 670424 477516
rect 670476 477504 670482 477556
rect 676030 476076 676036 476128
rect 676088 476116 676094 476128
rect 680354 476116 680360 476128
rect 676088 476088 680360 476116
rect 676088 476076 676094 476088
rect 680354 476076 680360 476088
rect 680412 476076 680418 476128
rect 664438 474240 664444 474292
rect 664496 474280 664502 474292
rect 667474 474280 667480 474292
rect 664496 474252 667480 474280
rect 664496 474240 664502 474252
rect 667474 474240 667480 474252
rect 667532 474240 667538 474292
rect 652754 467100 652760 467152
rect 652812 467140 652818 467152
rect 664438 467140 664444 467152
rect 652812 467112 664444 467140
rect 652812 467100 652818 467112
rect 664438 467100 664444 467112
rect 664496 467100 664502 467152
rect 650822 461320 650828 461372
rect 650880 461360 650886 461372
rect 652754 461360 652760 461372
rect 650880 461332 652760 461360
rect 650880 461320 650886 461332
rect 652754 461320 652760 461332
rect 652812 461320 652818 461372
rect 667014 456560 667020 456612
rect 667072 456600 667078 456612
rect 667072 456572 673988 456600
rect 667072 456560 667078 456572
rect 673960 456246 673988 456572
rect 667842 455948 667848 456000
rect 667900 455988 667906 456000
rect 667900 455960 673854 455988
rect 667900 455948 667906 455960
rect 672166 455812 672172 455864
rect 672224 455852 672230 455864
rect 672224 455824 673762 455852
rect 672224 455812 672230 455824
rect 669222 455608 669228 455660
rect 669280 455648 669286 455660
rect 669280 455620 673624 455648
rect 669280 455608 669286 455620
rect 673270 455336 673276 455388
rect 673328 455336 673334 455388
rect 673288 455022 673316 455336
rect 673388 455252 673440 455258
rect 673388 455194 673440 455200
rect 673506 455252 673558 455258
rect 673506 455194 673558 455200
rect 674282 454860 674288 454912
rect 674340 454900 674346 454912
rect 675846 454900 675852 454912
rect 674340 454872 675852 454900
rect 674340 454860 674346 454872
rect 675846 454860 675852 454872
rect 675904 454860 675910 454912
rect 672074 454792 672080 454844
rect 672132 454832 672138 454844
rect 672132 454804 673190 454832
rect 672132 454792 672138 454804
rect 673046 454640 673098 454646
rect 674282 454588 674288 454640
rect 674340 454628 674346 454640
rect 675478 454628 675484 454640
rect 674340 454600 675484 454628
rect 674340 454588 674346 454600
rect 675478 454588 675484 454600
rect 675536 454588 675542 454640
rect 673046 454582 673098 454588
rect 672810 454452 672816 454504
rect 672868 454452 672874 454504
rect 672828 454206 672856 454452
rect 672954 454368 673006 454374
rect 674282 454316 674288 454368
rect 674340 454356 674346 454368
rect 675662 454356 675668 454368
rect 674340 454328 675668 454356
rect 674340 454316 674346 454328
rect 675662 454316 675668 454328
rect 675720 454316 675726 454368
rect 672954 454310 673006 454316
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 674282 453908 674288 453960
rect 674340 453948 674346 453960
rect 676030 453948 676036 453960
rect 674340 453920 676036 453948
rect 674340 453908 674346 453920
rect 676030 453908 676036 453920
rect 676088 453908 676094 453960
rect 35802 429156 35808 429208
rect 35860 429196 35866 429208
rect 41690 429196 41696 429208
rect 35860 429168 41696 429196
rect 35860 429156 35866 429168
rect 41690 429156 41696 429168
rect 41748 429156 41754 429208
rect 35802 427932 35808 427984
rect 35860 427972 35866 427984
rect 41690 427972 41696 427984
rect 35860 427944 41696 427972
rect 35860 427932 35866 427944
rect 41690 427932 41696 427944
rect 41748 427932 41754 427984
rect 41138 424328 41144 424380
rect 41196 424368 41202 424380
rect 41690 424368 41696 424380
rect 41196 424340 41696 424368
rect 41196 424328 41202 424340
rect 41690 424328 41696 424340
rect 41748 424328 41754 424380
rect 32766 417392 32772 417444
rect 32824 417432 32830 417444
rect 41690 417432 41696 417444
rect 32824 417404 41696 417432
rect 32824 417392 32830 417404
rect 41690 417392 41696 417404
rect 41748 417392 41754 417444
rect 42058 417256 42064 417308
rect 42116 417296 42122 417308
rect 42610 417296 42616 417308
rect 42116 417268 42616 417296
rect 42116 417256 42122 417268
rect 42610 417256 42616 417268
rect 42668 417256 42674 417308
rect 34514 416032 34520 416084
rect 34572 416072 34578 416084
rect 41598 416072 41604 416084
rect 34572 416044 41604 416072
rect 34572 416032 34578 416044
rect 41598 416032 41604 416044
rect 41656 416032 41662 416084
rect 42242 406988 42248 407040
rect 42300 407028 42306 407040
rect 42610 407028 42616 407040
rect 42300 407000 42616 407028
rect 42300 406988 42306 407000
rect 42610 406988 42616 407000
rect 42668 406988 42674 407040
rect 45278 404268 45284 404320
rect 45336 404308 45342 404320
rect 62114 404308 62120 404320
rect 45336 404280 62120 404308
rect 45336 404268 45342 404280
rect 62114 404268 62120 404280
rect 62172 404268 62178 404320
rect 674558 403248 674564 403300
rect 674616 403288 674622 403300
rect 676214 403288 676220 403300
rect 674616 403260 676220 403288
rect 674616 403248 674622 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 51442 402908 51448 402960
rect 51500 402948 51506 402960
rect 62114 402948 62120 402960
rect 51500 402920 62120 402948
rect 51500 402908 51506 402920
rect 62114 402908 62120 402920
rect 62172 402908 62178 402960
rect 42426 402500 42432 402552
rect 42484 402540 42490 402552
rect 42978 402540 42984 402552
rect 42484 402512 42984 402540
rect 42484 402500 42490 402512
rect 42978 402500 42984 402512
rect 43036 402500 43042 402552
rect 42426 402024 42432 402076
rect 42484 402064 42490 402076
rect 43254 402064 43260 402076
rect 42484 402036 43260 402064
rect 42484 402024 42490 402036
rect 43254 402024 43260 402036
rect 43312 402024 43318 402076
rect 51074 400188 51080 400240
rect 51132 400228 51138 400240
rect 62114 400228 62120 400240
rect 51132 400200 62120 400228
rect 51132 400188 51138 400200
rect 62114 400188 62120 400200
rect 62172 400188 62178 400240
rect 44818 400052 44824 400104
rect 44876 400092 44882 400104
rect 62114 400092 62120 400104
rect 44876 400064 62120 400092
rect 44876 400052 44882 400064
rect 62114 400052 62120 400064
rect 62172 400052 62178 400104
rect 674926 398828 674932 398880
rect 674984 398868 674990 398880
rect 676030 398868 676036 398880
rect 674984 398840 676036 398868
rect 674984 398828 674990 398840
rect 676030 398828 676036 398840
rect 676088 398828 676094 398880
rect 47762 398760 47768 398812
rect 47820 398800 47826 398812
rect 62114 398800 62120 398812
rect 47820 398772 62120 398800
rect 47820 398760 47826 398772
rect 62114 398760 62120 398772
rect 62172 398760 62178 398812
rect 674558 396040 674564 396092
rect 674616 396080 674622 396092
rect 676030 396080 676036 396092
rect 674616 396052 676036 396080
rect 674616 396040 674622 396052
rect 676030 396040 676036 396052
rect 676088 396040 676094 396092
rect 675202 395700 675208 395752
rect 675260 395740 675266 395752
rect 676214 395740 676220 395752
rect 675260 395712 676220 395740
rect 675260 395700 675266 395712
rect 676214 395700 676220 395712
rect 676272 395700 676278 395752
rect 674374 394272 674380 394324
rect 674432 394312 674438 394324
rect 676214 394312 676220 394324
rect 674432 394284 676220 394312
rect 674432 394272 674438 394284
rect 676214 394272 676220 394284
rect 676272 394272 676278 394324
rect 679618 386764 679624 386776
rect 675588 386736 679624 386764
rect 41322 386384 41328 386436
rect 41380 386424 41386 386436
rect 41690 386424 41696 386436
rect 41380 386396 41696 386424
rect 41380 386384 41386 386396
rect 41690 386384 41696 386396
rect 41748 386384 41754 386436
rect 675588 386424 675616 386736
rect 679618 386724 679624 386736
rect 679676 386724 679682 386776
rect 675496 386396 675616 386424
rect 675496 386028 675524 386396
rect 675478 385976 675484 386028
rect 675536 385976 675542 386028
rect 674834 384752 674840 384804
rect 674892 384792 674898 384804
rect 675386 384792 675392 384804
rect 674892 384764 675392 384792
rect 674892 384752 674898 384764
rect 675386 384752 675392 384764
rect 675444 384752 675450 384804
rect 41322 382372 41328 382424
rect 41380 382412 41386 382424
rect 41690 382412 41696 382424
rect 41380 382384 41696 382412
rect 41380 382372 41386 382384
rect 41690 382372 41696 382384
rect 41748 382372 41754 382424
rect 674374 382168 674380 382220
rect 674432 382208 674438 382220
rect 675110 382208 675116 382220
rect 674432 382180 675116 382208
rect 674432 382168 674438 382180
rect 675110 382168 675116 382180
rect 675168 382168 675174 382220
rect 41322 379720 41328 379772
rect 41380 379760 41386 379772
rect 41506 379760 41512 379772
rect 41380 379732 41512 379760
rect 41380 379720 41386 379732
rect 41506 379720 41512 379732
rect 41564 379720 41570 379772
rect 35802 379584 35808 379636
rect 35860 379624 35866 379636
rect 40402 379624 40408 379636
rect 35860 379596 36032 379624
rect 35860 379584 35866 379596
rect 36004 379488 36032 379596
rect 36096 379596 40408 379624
rect 36096 379488 36124 379596
rect 40402 379584 40408 379596
rect 40460 379584 40466 379636
rect 36004 379460 36124 379488
rect 35802 378156 35808 378208
rect 35860 378196 35866 378208
rect 41690 378196 41696 378208
rect 35860 378168 41696 378196
rect 35860 378156 35866 378168
rect 41690 378156 41696 378168
rect 41748 378156 41754 378208
rect 674374 378088 674380 378140
rect 674432 378128 674438 378140
rect 675110 378128 675116 378140
rect 674432 378100 675116 378128
rect 674432 378088 674438 378100
rect 675110 378088 675116 378100
rect 675168 378088 675174 378140
rect 651466 373940 651472 373992
rect 651524 373980 651530 373992
rect 657538 373980 657544 373992
rect 651524 373952 657544 373980
rect 651524 373940 651530 373952
rect 657538 373940 657544 373952
rect 657596 373940 657602 373992
rect 33962 373260 33968 373312
rect 34020 373300 34026 373312
rect 41690 373300 41696 373312
rect 34020 373272 41696 373300
rect 34020 373260 34026 373272
rect 41690 373260 41696 373272
rect 41748 373260 41754 373312
rect 39298 371832 39304 371884
rect 39356 371872 39362 371884
rect 41690 371872 41696 371884
rect 39356 371844 41696 371872
rect 39356 371832 39362 371844
rect 41690 371832 41696 371844
rect 41748 371832 41754 371884
rect 42058 371696 42064 371748
rect 42116 371736 42122 371748
rect 42702 371736 42708 371748
rect 42116 371708 42708 371736
rect 42116 371696 42122 371708
rect 42702 371696 42708 371708
rect 42760 371696 42766 371748
rect 651466 370948 651472 371000
rect 651524 370988 651530 371000
rect 654778 370988 654784 371000
rect 651524 370960 654784 370988
rect 651524 370948 651530 370960
rect 654778 370948 654784 370960
rect 654836 370948 654842 371000
rect 42334 366800 42340 366852
rect 42392 366840 42398 366852
rect 43070 366840 43076 366852
rect 42392 366812 43076 366840
rect 42392 366800 42398 366812
rect 43070 366800 43076 366812
rect 43128 366800 43134 366852
rect 42242 364964 42248 365016
rect 42300 365004 42306 365016
rect 42702 365004 42708 365016
rect 42300 364976 42708 365004
rect 42300 364964 42306 364976
rect 42702 364964 42708 364976
rect 42760 364964 42766 365016
rect 651006 362924 651012 362976
rect 651064 362964 651070 362976
rect 655514 362964 655520 362976
rect 651064 362936 655520 362964
rect 651064 362924 651070 362936
rect 655514 362924 655520 362936
rect 655572 362924 655578 362976
rect 45646 361496 45652 361548
rect 45704 361536 45710 361548
rect 62114 361536 62120 361548
rect 45704 361508 62120 361536
rect 45704 361496 45710 361508
rect 62114 361496 62120 361508
rect 62172 361496 62178 361548
rect 51074 360136 51080 360188
rect 51132 360176 51138 360188
rect 62114 360176 62120 360188
rect 51132 360148 62120 360176
rect 51132 360136 51138 360148
rect 62114 360136 62120 360148
rect 62172 360136 62178 360188
rect 44634 357416 44640 357468
rect 44692 357456 44698 357468
rect 62114 357456 62120 357468
rect 44692 357428 62120 357456
rect 44692 357416 44698 357428
rect 62114 357416 62120 357428
rect 62172 357416 62178 357468
rect 42242 355988 42248 356040
rect 42300 356028 42306 356040
rect 42886 356028 42892 356040
rect 42300 356000 42892 356028
rect 42300 355988 42306 356000
rect 42886 355988 42892 356000
rect 42944 355988 42950 356040
rect 47762 355988 47768 356040
rect 47820 356028 47826 356040
rect 62114 356028 62120 356040
rect 47820 356000 62120 356028
rect 47820 355988 47826 356000
rect 62114 355988 62120 356000
rect 62172 355988 62178 356040
rect 44640 354544 44692 354550
rect 44640 354486 44692 354492
rect 44732 354408 44784 354414
rect 44732 354350 44784 354356
rect 45646 354328 45652 354340
rect 44881 354300 45652 354328
rect 45646 354288 45652 354300
rect 45704 354288 45710 354340
rect 45830 354192 45836 354204
rect 45091 354164 45836 354192
rect 45091 354056 45119 354164
rect 45830 354152 45836 354164
rect 45888 354152 45894 354204
rect 44988 354028 45119 354056
rect 45462 354016 45468 354068
rect 45520 354056 45526 354068
rect 45520 354028 45692 354056
rect 45520 354016 45526 354028
rect 45462 353920 45468 353932
rect 45105 353892 45468 353920
rect 45462 353880 45468 353892
rect 45520 353880 45526 353932
rect 45664 353784 45692 354028
rect 45204 353756 45692 353784
rect 45204 353702 45232 353756
rect 45462 353444 45468 353456
rect 45329 353416 45468 353444
rect 45462 353404 45468 353416
rect 45520 353404 45526 353456
rect 45422 353184 45474 353190
rect 45422 353126 45474 353132
rect 35802 344564 35808 344616
rect 35860 344604 35866 344616
rect 39850 344604 39856 344616
rect 35860 344576 39856 344604
rect 35860 344564 35866 344576
rect 39850 344564 39856 344576
rect 39908 344564 39914 344616
rect 35618 343612 35624 343664
rect 35676 343652 35682 343664
rect 40034 343652 40040 343664
rect 35676 343624 40040 343652
rect 35676 343612 35682 343624
rect 40034 343612 40040 343624
rect 40092 343612 40098 343664
rect 35802 342252 35808 342304
rect 35860 342292 35866 342304
rect 40218 342292 40224 342304
rect 35860 342264 40224 342292
rect 35860 342252 35866 342264
rect 40218 342252 40224 342264
rect 40276 342252 40282 342304
rect 33042 341368 33048 341420
rect 33100 341408 33106 341420
rect 40218 341408 40224 341420
rect 33100 341380 40224 341408
rect 33100 341368 33106 341380
rect 40218 341368 40224 341380
rect 40276 341368 40282 341420
rect 45462 341368 45468 341420
rect 45520 341408 45526 341420
rect 62298 341408 62304 341420
rect 45520 341380 62304 341408
rect 45520 341368 45526 341380
rect 62298 341368 62304 341380
rect 62356 341368 62362 341420
rect 35802 341164 35808 341216
rect 35860 341204 35866 341216
rect 40218 341204 40224 341216
rect 35860 341176 40224 341204
rect 35860 341164 35866 341176
rect 40218 341164 40224 341176
rect 40276 341164 40282 341216
rect 35802 341028 35808 341080
rect 35860 341068 35866 341080
rect 40034 341068 40040 341080
rect 35860 341040 40040 341068
rect 35860 341028 35866 341040
rect 40034 341028 40040 341040
rect 40092 341028 40098 341080
rect 35802 339600 35808 339652
rect 35860 339640 35866 339652
rect 37918 339640 37924 339652
rect 35860 339612 37924 339640
rect 35860 339600 35866 339612
rect 37918 339600 37924 339612
rect 37976 339600 37982 339652
rect 35526 339464 35532 339516
rect 35584 339504 35590 339516
rect 38654 339504 38660 339516
rect 35584 339476 38660 339504
rect 35584 339464 35590 339476
rect 38654 339464 38660 339476
rect 38712 339464 38718 339516
rect 35802 335316 35808 335368
rect 35860 335356 35866 335368
rect 40218 335356 40224 335368
rect 35860 335328 40224 335356
rect 35860 335316 35866 335328
rect 40218 335316 40224 335328
rect 40276 335316 40282 335368
rect 35802 334092 35808 334144
rect 35860 334132 35866 334144
rect 39758 334132 39764 334144
rect 35860 334104 39764 334132
rect 35860 334092 35866 334104
rect 39758 334092 39764 334104
rect 39816 334092 39822 334144
rect 674466 331032 674472 331084
rect 674524 331072 674530 331084
rect 675110 331072 675116 331084
rect 674524 331044 675116 331072
rect 674524 331032 674530 331044
rect 675110 331032 675116 331044
rect 675168 331032 675174 331084
rect 651374 328244 651380 328296
rect 651432 328284 651438 328296
rect 654778 328284 654784 328296
rect 651432 328256 654784 328284
rect 651432 328244 651438 328256
rect 654778 328244 654784 328256
rect 654836 328244 654842 328296
rect 651374 325592 651380 325644
rect 651432 325632 651438 325644
rect 653398 325632 653404 325644
rect 651432 325604 653404 325632
rect 651432 325592 651438 325604
rect 653398 325592 653404 325604
rect 653456 325592 653462 325644
rect 42426 322872 42432 322924
rect 42484 322912 42490 322924
rect 43070 322912 43076 322924
rect 42484 322884 43076 322912
rect 42484 322872 42490 322884
rect 43070 322872 43076 322884
rect 43128 322872 43134 322924
rect 42242 321512 42248 321564
rect 42300 321552 42306 321564
rect 42886 321552 42892 321564
rect 42300 321524 42892 321552
rect 42300 321512 42306 321524
rect 42886 321512 42892 321524
rect 42944 321512 42950 321564
rect 45462 317364 45468 317416
rect 45520 317404 45526 317416
rect 62114 317404 62120 317416
rect 45520 317376 62120 317404
rect 45520 317364 45526 317376
rect 62114 317364 62120 317376
rect 62172 317364 62178 317416
rect 62114 314752 62120 314764
rect 45526 314724 62120 314752
rect 45526 314696 45554 314724
rect 62114 314712 62120 314724
rect 62172 314712 62178 314764
rect 45462 314644 45468 314696
rect 45520 314656 45554 314696
rect 45520 314644 45526 314656
rect 674374 311992 674380 312044
rect 674432 312032 674438 312044
rect 675478 312032 675484 312044
rect 674432 312004 675484 312032
rect 674432 311992 674438 312004
rect 675478 311992 675484 312004
rect 675536 311992 675542 312044
rect 674742 309816 674748 309868
rect 674800 309856 674806 309868
rect 675478 309856 675484 309868
rect 674800 309828 675484 309856
rect 674800 309816 674806 309828
rect 675478 309816 675484 309828
rect 675536 309816 675542 309868
rect 676214 306348 676220 306400
rect 676272 306388 676278 306400
rect 676858 306388 676864 306400
rect 676272 306360 676864 306388
rect 676272 306348 676278 306360
rect 676858 306348 676864 306360
rect 676916 306348 676922 306400
rect 675846 304852 675852 304904
rect 675904 304892 675910 304904
rect 676398 304892 676404 304904
rect 675904 304864 676404 304892
rect 675904 304852 675910 304864
rect 676398 304852 676404 304864
rect 676456 304852 676462 304904
rect 651374 303492 651380 303544
rect 651432 303532 651438 303544
rect 653398 303532 653404 303544
rect 651432 303504 653404 303532
rect 651432 303492 651438 303504
rect 653398 303492 653404 303504
rect 653456 303492 653462 303544
rect 41322 300840 41328 300892
rect 41380 300880 41386 300892
rect 41690 300880 41696 300892
rect 41380 300852 41696 300880
rect 41380 300840 41386 300852
rect 41690 300840 41696 300852
rect 41748 300840 41754 300892
rect 46382 300772 46388 300824
rect 46440 300812 46446 300824
rect 52086 300812 52092 300824
rect 46440 300784 52092 300812
rect 46440 300772 46446 300784
rect 52086 300772 52092 300784
rect 52144 300772 52150 300824
rect 651466 300772 651472 300824
rect 651524 300812 651530 300824
rect 658918 300812 658924 300824
rect 651524 300784 658924 300812
rect 651524 300772 651530 300784
rect 658918 300772 658924 300784
rect 658976 300772 658982 300824
rect 47578 299412 47584 299464
rect 47636 299452 47642 299464
rect 54478 299452 54484 299464
rect 47636 299424 54484 299452
rect 47636 299412 47642 299424
rect 54478 299412 54484 299424
rect 54536 299412 54542 299464
rect 41138 299072 41144 299124
rect 41196 299112 41202 299124
rect 41690 299112 41696 299124
rect 41196 299084 41696 299112
rect 41196 299072 41202 299084
rect 41690 299072 41696 299084
rect 41748 299072 41754 299124
rect 651466 298120 651472 298172
rect 651524 298160 651530 298172
rect 660574 298160 660580 298172
rect 651524 298132 660580 298160
rect 651524 298120 651530 298132
rect 660574 298120 660580 298132
rect 660632 298120 660638 298172
rect 674742 297780 674748 297832
rect 674800 297820 674806 297832
rect 675478 297820 675484 297832
rect 674800 297792 675484 297820
rect 674800 297780 674806 297792
rect 675478 297780 675484 297792
rect 675536 297780 675542 297832
rect 676030 297576 676036 297628
rect 676088 297616 676094 297628
rect 678974 297616 678980 297628
rect 676088 297588 678980 297616
rect 676088 297576 676094 297588
rect 678974 297576 678980 297588
rect 679032 297576 679038 297628
rect 675846 297440 675852 297492
rect 675904 297480 675910 297492
rect 678238 297480 678244 297492
rect 675904 297452 678244 297480
rect 675904 297440 675910 297452
rect 678238 297440 678244 297452
rect 678296 297440 678302 297492
rect 652202 296760 652208 296812
rect 652260 296800 652266 296812
rect 652260 296772 654134 296800
rect 652260 296760 652266 296772
rect 654106 296732 654134 296772
rect 658918 296732 658924 296744
rect 654106 296704 658924 296732
rect 658918 296692 658924 296704
rect 658976 296692 658982 296744
rect 675294 296148 675300 296200
rect 675352 296148 675358 296200
rect 41138 295468 41144 295520
rect 41196 295508 41202 295520
rect 41690 295508 41696 295520
rect 41196 295480 41696 295508
rect 41196 295468 41202 295480
rect 41690 295468 41696 295480
rect 41748 295468 41754 295520
rect 675312 295452 675340 296148
rect 675294 295400 675300 295452
rect 675352 295400 675358 295452
rect 45462 295332 45468 295384
rect 45520 295372 45526 295384
rect 62114 295372 62120 295384
rect 45520 295344 62120 295372
rect 45520 295332 45526 295344
rect 62114 295332 62120 295344
rect 62172 295332 62178 295384
rect 41322 294244 41328 294296
rect 41380 294284 41386 294296
rect 41690 294284 41696 294296
rect 41380 294256 41696 294284
rect 41380 294244 41386 294256
rect 41690 294244 41696 294256
rect 41748 294244 41754 294296
rect 42058 294244 42064 294296
rect 42116 294284 42122 294296
rect 42610 294284 42616 294296
rect 42116 294256 42616 294284
rect 42116 294244 42122 294256
rect 42610 294244 42616 294256
rect 42668 294244 42674 294296
rect 57422 294040 57428 294092
rect 57480 294080 57486 294092
rect 62114 294080 62120 294092
rect 57480 294052 62120 294080
rect 57480 294040 57486 294052
rect 62114 294040 62120 294052
rect 62172 294040 62178 294092
rect 651466 293972 651472 294024
rect 651524 294012 651530 294024
rect 664438 294012 664444 294024
rect 651524 293984 664444 294012
rect 651524 293972 651530 293984
rect 664438 293972 664444 293984
rect 664496 293972 664502 294024
rect 42058 293020 42064 293072
rect 42116 293060 42122 293072
rect 43346 293060 43352 293072
rect 42116 293032 43352 293060
rect 42116 293020 42122 293032
rect 43346 293020 43352 293032
rect 43404 293020 43410 293072
rect 41690 292788 41696 292800
rect 41386 292760 41696 292788
rect 41386 292732 41414 292760
rect 41690 292748 41696 292760
rect 41748 292748 41754 292800
rect 41322 292680 41328 292732
rect 41380 292692 41414 292732
rect 41380 292680 41386 292692
rect 60366 292544 60372 292596
rect 60424 292584 60430 292596
rect 62298 292584 62304 292596
rect 60424 292556 62304 292584
rect 60424 292544 60430 292556
rect 62298 292544 62304 292556
rect 62356 292544 62362 292596
rect 651466 292544 651472 292596
rect 651524 292584 651530 292596
rect 660298 292584 660304 292596
rect 651524 292556 660304 292584
rect 651524 292544 651530 292556
rect 660298 292544 660304 292556
rect 660356 292544 660362 292596
rect 45462 292408 45468 292460
rect 45520 292448 45526 292460
rect 62114 292448 62120 292460
rect 45520 292420 62120 292448
rect 45520 292408 45526 292420
rect 62114 292408 62120 292420
rect 62172 292408 62178 292460
rect 651466 289824 651472 289876
rect 651524 289864 651530 289876
rect 663058 289864 663064 289876
rect 651524 289836 663064 289864
rect 651524 289824 651530 289836
rect 663058 289824 663064 289836
rect 663116 289824 663122 289876
rect 54478 288396 54484 288448
rect 54536 288436 54542 288448
rect 57606 288436 57612 288448
rect 54536 288408 57612 288436
rect 54536 288396 54542 288408
rect 57606 288396 57612 288408
rect 57664 288396 57670 288448
rect 651466 288396 651472 288448
rect 651524 288436 651530 288448
rect 672166 288436 672172 288448
rect 651524 288408 672172 288436
rect 651524 288396 651530 288408
rect 672166 288396 672172 288408
rect 672224 288396 672230 288448
rect 651466 287036 651472 287088
rect 651524 287076 651530 287088
rect 667566 287076 667572 287088
rect 651524 287048 667572 287076
rect 651524 287036 651530 287048
rect 667566 287036 667572 287048
rect 667624 287036 667630 287088
rect 33778 286288 33784 286340
rect 33836 286328 33842 286340
rect 41506 286328 41512 286340
rect 33836 286300 41512 286328
rect 33836 286288 33842 286300
rect 41506 286288 41512 286300
rect 41564 286288 41570 286340
rect 45462 285676 45468 285728
rect 45520 285716 45526 285728
rect 62114 285716 62120 285728
rect 45520 285688 62120 285716
rect 45520 285676 45526 285688
rect 62114 285676 62120 285688
rect 62172 285676 62178 285728
rect 651466 285676 651472 285728
rect 651524 285716 651530 285728
rect 667382 285716 667388 285728
rect 651524 285688 667388 285716
rect 651524 285676 651530 285688
rect 667382 285676 667388 285688
rect 667440 285676 667446 285728
rect 39942 284452 39948 284504
rect 40000 284492 40006 284504
rect 41690 284492 41696 284504
rect 40000 284464 41696 284492
rect 40000 284452 40006 284464
rect 41690 284452 41696 284464
rect 41748 284452 41754 284504
rect 46382 284316 46388 284368
rect 46440 284356 46446 284368
rect 63218 284356 63224 284368
rect 46440 284328 63224 284356
rect 46440 284316 46446 284328
rect 63218 284316 63224 284328
rect 63276 284316 63282 284368
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 672350 284356 672356 284368
rect 651524 284328 672356 284356
rect 651524 284316 651530 284328
rect 672350 284316 672356 284328
rect 672408 284316 672414 284368
rect 51718 282888 51724 282940
rect 51776 282928 51782 282940
rect 62114 282928 62120 282940
rect 51776 282900 62120 282928
rect 51776 282888 51782 282900
rect 62114 282888 62120 282900
rect 62172 282888 62178 282940
rect 651466 282888 651472 282940
rect 651524 282928 651530 282940
rect 666554 282928 666560 282940
rect 651524 282900 666560 282928
rect 651524 282888 651530 282900
rect 666554 282888 666560 282900
rect 666612 282888 666618 282940
rect 56042 281528 56048 281580
rect 56100 281568 56106 281580
rect 62850 281568 62856 281580
rect 56100 281540 62856 281568
rect 56100 281528 56106 281540
rect 62850 281528 62856 281540
rect 62908 281528 62914 281580
rect 651466 280168 651472 280220
rect 651524 280208 651530 280220
rect 667198 280208 667204 280220
rect 651524 280180 667204 280208
rect 651524 280168 651530 280180
rect 667198 280168 667204 280180
rect 667256 280168 667262 280220
rect 42426 280100 42432 280152
rect 42484 280140 42490 280152
rect 43070 280140 43076 280152
rect 42484 280112 43076 280140
rect 42484 280100 42490 280112
rect 43070 280100 43076 280112
rect 43128 280100 43134 280152
rect 58618 280032 58624 280084
rect 58676 280072 58682 280084
rect 61930 280072 61936 280084
rect 58676 280044 61936 280072
rect 58676 280032 58682 280044
rect 61930 280032 61936 280044
rect 61988 280032 61994 280084
rect 57606 278672 57612 278724
rect 57664 278712 57670 278724
rect 61746 278712 61752 278724
rect 57664 278684 61752 278712
rect 57664 278672 57670 278684
rect 61746 278672 61752 278684
rect 61804 278672 61810 278724
rect 63494 278672 63500 278724
rect 63552 278712 63558 278724
rect 671338 278712 671344 278724
rect 63552 278684 671344 278712
rect 63552 278672 63558 278684
rect 671338 278672 671344 278684
rect 671396 278672 671402 278724
rect 49326 278536 49332 278588
rect 49384 278576 49390 278588
rect 49384 278548 60044 278576
rect 49384 278536 49390 278548
rect 60016 278440 60044 278548
rect 60550 278536 60556 278588
rect 60608 278576 60614 278588
rect 61930 278576 61936 278588
rect 60608 278548 61936 278576
rect 60608 278536 60614 278548
rect 61930 278536 61936 278548
rect 61988 278536 61994 278588
rect 63310 278536 63316 278588
rect 63368 278576 63374 278588
rect 671706 278576 671712 278588
rect 63368 278548 671712 278576
rect 63368 278536 63374 278548
rect 671706 278536 671712 278548
rect 671764 278536 671770 278588
rect 650822 278440 650828 278452
rect 60016 278412 650828 278440
rect 650822 278400 650828 278412
rect 650880 278400 650886 278452
rect 52086 278264 52092 278316
rect 52144 278304 52150 278316
rect 60550 278304 60556 278316
rect 52144 278276 60556 278304
rect 52144 278264 52150 278276
rect 60550 278264 60556 278276
rect 60608 278264 60614 278316
rect 61746 278264 61752 278316
rect 61804 278304 61810 278316
rect 651006 278304 651012 278316
rect 61804 278276 651012 278304
rect 61804 278264 61810 278276
rect 651006 278264 651012 278276
rect 651064 278264 651070 278316
rect 51902 278128 51908 278180
rect 51960 278168 51966 278180
rect 629938 278168 629944 278180
rect 51960 278140 629944 278168
rect 51960 278128 51966 278140
rect 629938 278128 629944 278140
rect 629996 278128 630002 278180
rect 630122 278128 630128 278180
rect 630180 278168 630186 278180
rect 650638 278168 650644 278180
rect 630180 278140 650644 278168
rect 630180 278128 630186 278140
rect 650638 278128 650644 278140
rect 650696 278128 650702 278180
rect 47762 277992 47768 278044
rect 47820 278032 47826 278044
rect 635090 278032 635096 278044
rect 47820 278004 635096 278032
rect 47820 277992 47826 278004
rect 635090 277992 635096 278004
rect 635148 277992 635154 278044
rect 64322 277856 64328 277908
rect 64380 277896 64386 277908
rect 637758 277896 637764 277908
rect 64380 277868 637764 277896
rect 64380 277856 64386 277868
rect 637758 277856 637764 277868
rect 637816 277856 637822 277908
rect 74506 277732 625154 277760
rect 61930 277584 61936 277636
rect 61988 277624 61994 277636
rect 74506 277624 74534 277732
rect 61988 277596 74534 277624
rect 625126 277624 625154 277732
rect 629938 277720 629944 277772
rect 629996 277760 630002 277772
rect 636286 277760 636292 277772
rect 629996 277732 636292 277760
rect 629996 277720 630002 277732
rect 636286 277720 636292 277732
rect 636344 277720 636350 277772
rect 630122 277624 630128 277636
rect 625126 277596 630128 277624
rect 61988 277584 61994 277596
rect 630122 277584 630128 277596
rect 630180 277584 630186 277636
rect 479978 277312 479984 277364
rect 480036 277352 480042 277364
rect 555234 277352 555240 277364
rect 480036 277324 555240 277352
rect 480036 277312 480042 277324
rect 555234 277312 555240 277324
rect 555292 277312 555298 277364
rect 487982 277176 487988 277228
rect 488040 277216 488046 277228
rect 565814 277216 565820 277228
rect 488040 277188 565820 277216
rect 488040 277176 488046 277188
rect 565814 277176 565820 277188
rect 565872 277176 565878 277228
rect 497918 277040 497924 277092
rect 497976 277080 497982 277092
rect 579982 277080 579988 277092
rect 497976 277052 579988 277080
rect 497976 277040 497982 277052
rect 579982 277040 579988 277052
rect 580040 277040 580046 277092
rect 511626 276904 511632 276956
rect 511684 276944 511690 276956
rect 600130 276944 600136 276956
rect 511684 276916 600136 276944
rect 511684 276904 511690 276916
rect 600130 276904 600136 276916
rect 600188 276904 600194 276956
rect 42242 276768 42248 276820
rect 42300 276808 42306 276820
rect 42610 276808 42616 276820
rect 42300 276780 42616 276808
rect 42300 276768 42306 276780
rect 42610 276768 42616 276780
rect 42668 276768 42674 276820
rect 514478 276768 514484 276820
rect 514536 276808 514542 276820
rect 603626 276808 603632 276820
rect 514536 276780 603632 276808
rect 514536 276768 514542 276780
rect 603626 276768 603632 276780
rect 603684 276768 603690 276820
rect 53282 276632 53288 276684
rect 53340 276672 53346 276684
rect 62114 276672 62120 276684
rect 53340 276644 62120 276672
rect 53340 276632 53346 276644
rect 62114 276632 62120 276644
rect 62172 276632 62178 276684
rect 518710 276632 518716 276684
rect 518768 276672 518774 276684
rect 609606 276672 609612 276684
rect 518768 276644 609612 276672
rect 518768 276632 518774 276644
rect 609606 276632 609612 276644
rect 609664 276632 609670 276684
rect 482830 276496 482836 276548
rect 482888 276536 482894 276548
rect 557534 276536 557540 276548
rect 482888 276508 557540 276536
rect 482888 276496 482894 276508
rect 557534 276496 557540 276508
rect 557592 276496 557598 276548
rect 477034 276360 477040 276412
rect 477092 276400 477098 276412
rect 550450 276400 550456 276412
rect 477092 276372 550456 276400
rect 477092 276360 477098 276372
rect 550450 276360 550456 276372
rect 550508 276360 550514 276412
rect 471606 276224 471612 276276
rect 471664 276264 471670 276276
rect 543366 276264 543372 276276
rect 471664 276236 543372 276264
rect 471664 276224 471670 276236
rect 543366 276224 543372 276236
rect 543424 276224 543430 276276
rect 107194 275952 107200 276004
rect 107252 275992 107258 276004
rect 163498 275992 163504 276004
rect 107252 275964 163504 275992
rect 107252 275952 107258 275964
rect 163498 275952 163504 275964
rect 163556 275952 163562 276004
rect 167546 275952 167552 276004
rect 167604 275992 167610 276004
rect 178678 275992 178684 276004
rect 167604 275964 178684 275992
rect 167604 275952 167610 275964
rect 178678 275952 178684 275964
rect 178736 275952 178742 276004
rect 185210 275952 185216 276004
rect 185268 275992 185274 276004
rect 221274 275992 221280 276004
rect 185268 275964 221280 275992
rect 185268 275952 185274 275964
rect 221274 275952 221280 275964
rect 221332 275952 221338 276004
rect 232498 275952 232504 276004
rect 232556 275992 232562 276004
rect 239214 275992 239220 276004
rect 232556 275964 239220 275992
rect 232556 275952 232562 275964
rect 239214 275952 239220 275964
rect 239272 275952 239278 276004
rect 410794 275952 410800 276004
rect 410852 275992 410858 276004
rect 455874 275992 455880 276004
rect 410852 275964 455880 275992
rect 410852 275952 410858 275964
rect 455874 275952 455880 275964
rect 455932 275952 455938 276004
rect 456058 275952 456064 276004
rect 456116 275992 456122 276004
rect 509050 275992 509056 276004
rect 456116 275964 509056 275992
rect 456116 275952 456122 275964
rect 509050 275952 509056 275964
rect 509108 275952 509114 276004
rect 513190 275952 513196 276004
rect 513248 275992 513254 276004
rect 601326 275992 601332 276004
rect 513248 275964 601332 275992
rect 513248 275952 513254 275964
rect 601326 275952 601332 275964
rect 601384 275952 601390 276004
rect 139118 275816 139124 275868
rect 139176 275856 139182 275868
rect 174262 275856 174268 275868
rect 139176 275828 174268 275856
rect 139176 275816 139182 275828
rect 174262 275816 174268 275828
rect 174320 275816 174326 275868
rect 178126 275816 178132 275868
rect 178184 275856 178190 275868
rect 216674 275856 216680 275868
rect 178184 275828 216680 275856
rect 178184 275816 178190 275828
rect 216674 275816 216680 275828
rect 216732 275816 216738 275868
rect 224218 275816 224224 275868
rect 224276 275856 224282 275868
rect 232682 275856 232688 275868
rect 224276 275828 232688 275856
rect 224276 275816 224282 275828
rect 232682 275816 232688 275828
rect 232740 275816 232746 275868
rect 236086 275816 236092 275868
rect 236144 275856 236150 275868
rect 250438 275856 250444 275868
rect 236144 275828 250444 275856
rect 236144 275816 236150 275828
rect 250438 275816 250444 275828
rect 250496 275816 250502 275868
rect 286870 275816 286876 275868
rect 286928 275856 286934 275868
rect 291838 275856 291844 275868
rect 286928 275828 291844 275856
rect 286928 275816 286934 275828
rect 291838 275816 291844 275828
rect 291896 275816 291902 275868
rect 430206 275816 430212 275868
rect 430264 275856 430270 275868
rect 484302 275856 484308 275868
rect 430264 275828 484308 275856
rect 430264 275816 430270 275828
rect 484302 275816 484308 275828
rect 484360 275816 484366 275868
rect 490558 275816 490564 275868
rect 490616 275856 490622 275868
rect 505554 275856 505560 275868
rect 490616 275828 505560 275856
rect 490616 275816 490622 275828
rect 505554 275816 505560 275828
rect 505612 275816 505618 275868
rect 522758 275816 522764 275868
rect 522816 275856 522822 275868
rect 615494 275856 615500 275868
rect 522816 275828 615500 275856
rect 522816 275816 522822 275828
rect 615494 275816 615500 275828
rect 615552 275816 615558 275868
rect 260926 275748 260932 275800
rect 260984 275788 260990 275800
rect 266354 275788 266360 275800
rect 260984 275760 266360 275788
rect 260984 275748 260990 275760
rect 266354 275748 266360 275760
rect 266412 275748 266418 275800
rect 100110 275680 100116 275732
rect 100168 275720 100174 275732
rect 159450 275720 159456 275732
rect 100168 275692 159456 275720
rect 100168 275680 100174 275692
rect 159450 275680 159456 275692
rect 159508 275680 159514 275732
rect 160462 275680 160468 275732
rect 160520 275720 160526 275732
rect 199562 275720 199568 275732
rect 160520 275692 199568 275720
rect 160520 275680 160526 275692
rect 199562 275680 199568 275692
rect 199620 275680 199626 275732
rect 217134 275680 217140 275732
rect 217192 275720 217198 275732
rect 224218 275720 224224 275732
rect 217192 275692 224224 275720
rect 217192 275680 217198 275692
rect 224218 275680 224224 275692
rect 224276 275680 224282 275732
rect 229002 275680 229008 275732
rect 229060 275720 229066 275732
rect 243538 275720 243544 275732
rect 229060 275692 243544 275720
rect 229060 275680 229066 275692
rect 243538 275680 243544 275692
rect 243596 275680 243602 275732
rect 250254 275680 250260 275732
rect 250312 275720 250318 275732
rect 259362 275720 259368 275732
rect 250312 275692 259368 275720
rect 250312 275680 250318 275692
rect 259362 275680 259368 275692
rect 259420 275680 259426 275732
rect 284570 275680 284576 275732
rect 284628 275720 284634 275732
rect 290090 275720 290096 275732
rect 284628 275692 290096 275720
rect 284628 275680 284634 275692
rect 290090 275680 290096 275692
rect 290148 275680 290154 275732
rect 445018 275680 445024 275732
rect 445076 275720 445082 275732
rect 498470 275720 498476 275732
rect 445076 275692 498476 275720
rect 445076 275680 445082 275692
rect 498470 275680 498476 275692
rect 498528 275680 498534 275732
rect 498838 275680 498844 275732
rect 498896 275720 498902 275732
rect 512638 275720 512644 275732
rect 498896 275692 512644 275720
rect 498896 275680 498902 275692
rect 512638 275680 512644 275692
rect 512696 275680 512702 275732
rect 528186 275680 528192 275732
rect 528244 275720 528250 275732
rect 622578 275720 622584 275732
rect 528244 275692 622584 275720
rect 528244 275680 528250 275692
rect 622578 275680 622584 275692
rect 622636 275680 622642 275732
rect 291654 275612 291660 275664
rect 291712 275652 291718 275664
rect 295334 275652 295340 275664
rect 291712 275624 295340 275652
rect 291712 275612 291718 275624
rect 295334 275612 295340 275624
rect 295392 275612 295398 275664
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86218 275584 86224 275596
rect 76524 275556 86224 275584
rect 76524 275544 76530 275556
rect 86218 275544 86224 275556
rect 86276 275544 86282 275596
rect 90726 275544 90732 275596
rect 90784 275584 90790 275596
rect 154758 275584 154764 275596
rect 90784 275556 154764 275584
rect 90784 275544 90790 275556
rect 154758 275544 154764 275556
rect 154816 275544 154822 275596
rect 171042 275544 171048 275596
rect 171100 275584 171106 275596
rect 211614 275584 211620 275596
rect 171100 275556 211620 275584
rect 171100 275544 171106 275556
rect 211614 275544 211620 275556
rect 211672 275544 211678 275596
rect 218330 275544 218336 275596
rect 218388 275584 218394 275596
rect 233878 275584 233884 275596
rect 218388 275556 233884 275584
rect 218388 275544 218394 275556
rect 233878 275544 233884 275556
rect 233936 275544 233942 275596
rect 239582 275544 239588 275596
rect 239640 275584 239646 275596
rect 255958 275584 255964 275596
rect 239640 275556 255964 275584
rect 239640 275544 239646 275556
rect 255958 275544 255964 275556
rect 256016 275544 256022 275596
rect 257338 275544 257344 275596
rect 257396 275584 257402 275596
rect 262306 275584 262312 275596
rect 257396 275556 262312 275584
rect 257396 275544 257402 275556
rect 262306 275544 262312 275556
rect 262364 275544 262370 275596
rect 266814 275544 266820 275596
rect 266872 275584 266878 275596
rect 276474 275584 276480 275596
rect 266872 275556 276480 275584
rect 266872 275544 266878 275556
rect 276474 275544 276480 275556
rect 276532 275544 276538 275596
rect 363874 275544 363880 275596
rect 363932 275584 363938 275596
rect 388530 275584 388536 275596
rect 363932 275556 388536 275584
rect 363932 275544 363938 275556
rect 388530 275544 388536 275556
rect 388588 275544 388594 275596
rect 416406 275544 416412 275596
rect 416464 275584 416470 275596
rect 462958 275584 462964 275596
rect 416464 275556 462964 275584
rect 416464 275544 416470 275556
rect 462958 275544 462964 275556
rect 463016 275544 463022 275596
rect 463142 275544 463148 275596
rect 463200 275584 463206 275596
rect 516226 275584 516232 275596
rect 463200 275556 516232 275584
rect 463200 275544 463206 275556
rect 516226 275544 516232 275556
rect 516284 275544 516290 275596
rect 516778 275544 516784 275596
rect 516836 275584 516842 275596
rect 526806 275584 526812 275596
rect 516836 275556 526812 275584
rect 516836 275544 516842 275556
rect 526806 275544 526812 275556
rect 526864 275544 526870 275596
rect 532326 275544 532332 275596
rect 532384 275584 532390 275596
rect 629662 275584 629668 275596
rect 532384 275556 629668 275584
rect 532384 275544 532390 275556
rect 629662 275544 629668 275556
rect 629720 275544 629726 275596
rect 277486 275476 277492 275528
rect 277544 275516 277550 275528
rect 285122 275516 285128 275528
rect 277544 275488 285128 275516
rect 277544 275476 277550 275488
rect 285122 275476 285128 275488
rect 285180 275476 285186 275528
rect 81250 275408 81256 275460
rect 81308 275448 81314 275460
rect 144914 275448 144920 275460
rect 81308 275420 144920 275448
rect 81308 275408 81314 275420
rect 144914 275408 144920 275420
rect 144972 275408 144978 275460
rect 156874 275408 156880 275460
rect 156932 275448 156938 275460
rect 156932 275420 161474 275448
rect 156932 275408 156938 275420
rect 96614 275272 96620 275324
rect 96672 275312 96678 275324
rect 149606 275312 149612 275324
rect 96672 275284 149612 275312
rect 96672 275272 96678 275284
rect 149606 275272 149612 275284
rect 149664 275272 149670 275324
rect 161446 275312 161474 275420
rect 163958 275408 163964 275460
rect 164016 275448 164022 275460
rect 206370 275448 206376 275460
rect 164016 275420 206376 275448
rect 164016 275408 164022 275420
rect 206370 275408 206376 275420
rect 206428 275408 206434 275460
rect 221918 275408 221924 275460
rect 221976 275448 221982 275460
rect 243722 275448 243728 275460
rect 221976 275420 243728 275448
rect 221976 275408 221982 275420
rect 243722 275408 243728 275420
rect 243780 275408 243786 275460
rect 256142 275408 256148 275460
rect 256200 275448 256206 275460
rect 256200 275420 268976 275448
rect 256200 275408 256206 275420
rect 200758 275312 200764 275324
rect 161446 275284 200764 275312
rect 200758 275272 200764 275284
rect 200816 275272 200822 275324
rect 214834 275272 214840 275324
rect 214892 275312 214898 275324
rect 239398 275312 239404 275324
rect 214892 275284 239404 275312
rect 214892 275272 214898 275284
rect 239398 275272 239404 275284
rect 239456 275272 239462 275324
rect 243170 275272 243176 275324
rect 243228 275312 243234 275324
rect 256694 275312 256700 275324
rect 243228 275284 256700 275312
rect 243228 275272 243234 275284
rect 256694 275272 256700 275284
rect 256752 275272 256758 275324
rect 268948 275244 268976 275420
rect 285674 275408 285680 275460
rect 285732 275448 285738 275460
rect 291286 275448 291292 275460
rect 285732 275420 291292 275448
rect 285732 275408 285738 275420
rect 291286 275408 291292 275420
rect 291344 275408 291350 275460
rect 358630 275408 358636 275460
rect 358688 275448 358694 275460
rect 381446 275448 381452 275460
rect 358688 275420 381452 275448
rect 358688 275408 358694 275420
rect 381446 275408 381452 275420
rect 381504 275408 381510 275460
rect 386046 275408 386052 275460
rect 386104 275448 386110 275460
rect 420454 275448 420460 275460
rect 386104 275420 420460 275448
rect 386104 275408 386110 275420
rect 420454 275408 420460 275420
rect 420512 275408 420518 275460
rect 435634 275408 435640 275460
rect 435692 275448 435698 275460
rect 485038 275448 485044 275460
rect 435692 275420 485044 275448
rect 435692 275408 435698 275420
rect 485038 275408 485044 275420
rect 485096 275408 485102 275460
rect 485222 275408 485228 275460
rect 485280 275448 485286 275460
rect 530394 275448 530400 275460
rect 485280 275420 530400 275448
rect 485280 275408 485286 275420
rect 530394 275408 530400 275420
rect 530452 275408 530458 275460
rect 537662 275408 537668 275460
rect 537720 275448 537726 275460
rect 636746 275448 636752 275460
rect 537720 275420 636752 275448
rect 537720 275408 537726 275420
rect 636746 275408 636752 275420
rect 636804 275408 636810 275460
rect 269206 275340 269212 275392
rect 269264 275380 269270 275392
rect 274634 275380 274640 275392
rect 269264 275352 274640 275380
rect 269264 275340 269270 275352
rect 274634 275340 274640 275352
rect 274692 275340 274698 275392
rect 297542 275340 297548 275392
rect 297600 275380 297606 275392
rect 299566 275380 299572 275392
rect 297600 275352 299572 275380
rect 297600 275340 297606 275352
rect 299566 275340 299572 275352
rect 299624 275340 299630 275392
rect 299934 275340 299940 275392
rect 299992 275380 299998 275392
rect 301130 275380 301136 275392
rect 299992 275352 301136 275380
rect 299992 275340 299998 275352
rect 301130 275340 301136 275352
rect 301188 275340 301194 275392
rect 276290 275272 276296 275324
rect 276348 275312 276354 275324
rect 283098 275312 283104 275324
rect 276348 275284 283104 275312
rect 276348 275272 276354 275284
rect 283098 275272 283104 275284
rect 283156 275272 283162 275324
rect 290458 275272 290464 275324
rect 290516 275312 290522 275324
rect 294138 275312 294144 275324
rect 290516 275284 294144 275312
rect 290516 275272 290522 275284
rect 294138 275272 294144 275284
rect 294196 275272 294202 275324
rect 326430 275272 326436 275324
rect 326488 275312 326494 275324
rect 335354 275312 335360 275324
rect 326488 275284 335360 275312
rect 326488 275272 326494 275284
rect 335354 275272 335360 275284
rect 335412 275272 335418 275324
rect 371050 275272 371056 275324
rect 371108 275312 371114 275324
rect 399202 275312 399208 275324
rect 371108 275284 399208 275312
rect 371108 275272 371114 275284
rect 399202 275272 399208 275284
rect 399260 275272 399266 275324
rect 418798 275272 418804 275324
rect 418856 275312 418862 275324
rect 466546 275312 466552 275324
rect 418856 275284 466552 275312
rect 418856 275272 418862 275284
rect 466546 275272 466552 275284
rect 466604 275272 466610 275324
rect 467558 275272 467564 275324
rect 467616 275312 467622 275324
rect 537478 275312 537484 275324
rect 467616 275284 537484 275312
rect 467616 275272 467622 275284
rect 537478 275272 537484 275284
rect 537536 275272 537542 275324
rect 542262 275272 542268 275324
rect 542320 275312 542326 275324
rect 643830 275312 643836 275324
rect 542320 275284 643836 275312
rect 542320 275272 542326 275284
rect 643830 275272 643836 275284
rect 643888 275272 643894 275324
rect 269114 275244 269120 275256
rect 268948 275216 269120 275244
rect 269114 275204 269120 275216
rect 269172 275204 269178 275256
rect 298738 275204 298744 275256
rect 298796 275244 298802 275256
rect 300026 275244 300032 275256
rect 298796 275216 300032 275244
rect 298796 275204 298802 275216
rect 300026 275204 300032 275216
rect 300084 275204 300090 275256
rect 93026 275136 93032 275188
rect 93084 275176 93090 275188
rect 152826 275176 152832 275188
rect 93084 275148 152832 275176
rect 93084 275136 93090 275148
rect 152826 275136 152832 275148
rect 152884 275136 152890 275188
rect 153378 275136 153384 275188
rect 153436 275176 153442 275188
rect 169018 275176 169024 275188
rect 153436 275148 169024 275176
rect 153436 275136 153442 275148
rect 169018 275136 169024 275148
rect 169076 275136 169082 275188
rect 189994 275136 190000 275188
rect 190052 275176 190058 275188
rect 222930 275176 222936 275188
rect 190052 275148 222936 275176
rect 190052 275136 190058 275148
rect 222930 275136 222936 275148
rect 222988 275136 222994 275188
rect 292850 275136 292856 275188
rect 292908 275176 292914 275188
rect 295794 275176 295800 275188
rect 292908 275148 295800 275176
rect 292908 275136 292914 275148
rect 295794 275136 295800 275148
rect 295852 275136 295858 275188
rect 427078 275136 427084 275188
rect 427136 275176 427142 275188
rect 477218 275176 477224 275188
rect 427136 275148 477224 275176
rect 427136 275136 427142 275148
rect 477218 275136 477224 275148
rect 477276 275136 477282 275188
rect 485038 275136 485044 275188
rect 485096 275176 485102 275188
rect 491386 275176 491392 275188
rect 485096 275148 491392 275176
rect 485096 275136 485102 275148
rect 491386 275136 491392 275148
rect 491444 275136 491450 275188
rect 507486 275136 507492 275188
rect 507544 275176 507550 275188
rect 594242 275176 594248 275188
rect 507544 275148 594248 275176
rect 507544 275136 507550 275148
rect 594242 275136 594248 275148
rect 594300 275136 594306 275188
rect 263226 275068 263232 275120
rect 263284 275108 263290 275120
rect 273254 275108 273260 275120
rect 263284 275080 273260 275108
rect 263284 275068 263290 275080
rect 273254 275068 273260 275080
rect 273312 275068 273318 275120
rect 71774 275000 71780 275052
rect 71832 275040 71838 275052
rect 141050 275040 141056 275052
rect 71832 275012 141056 275040
rect 71832 275000 71838 275012
rect 141050 275000 141056 275012
rect 141108 275000 141114 275052
rect 149790 275000 149796 275052
rect 149848 275040 149854 275052
rect 189074 275040 189080 275052
rect 149848 275012 189080 275040
rect 149848 275000 149854 275012
rect 189074 275000 189080 275012
rect 189132 275000 189138 275052
rect 288066 275000 288072 275052
rect 288124 275040 288130 275052
rect 292666 275040 292672 275052
rect 288124 275012 292672 275040
rect 288124 275000 288130 275012
rect 292666 275000 292672 275012
rect 292724 275000 292730 275052
rect 420546 275000 420552 275052
rect 420604 275040 420610 275052
rect 470134 275040 470140 275052
rect 420604 275012 470140 275040
rect 420604 275000 420610 275012
rect 470134 275000 470140 275012
rect 470192 275000 470198 275052
rect 484302 275000 484308 275052
rect 484360 275040 484366 275052
rect 485222 275040 485228 275052
rect 484360 275012 485228 275040
rect 484360 275000 484366 275012
rect 485222 275000 485228 275012
rect 485280 275000 485286 275052
rect 503438 275000 503444 275052
rect 503496 275040 503502 275052
rect 587066 275040 587072 275052
rect 503496 275012 587072 275040
rect 503496 275000 503502 275012
rect 587066 275000 587072 275012
rect 587124 275000 587130 275052
rect 293954 274932 293960 274984
rect 294012 274972 294018 274984
rect 296806 274972 296812 274984
rect 294012 274944 296812 274972
rect 294012 274932 294018 274944
rect 296806 274932 296812 274944
rect 296864 274932 296870 274984
rect 146202 274864 146208 274916
rect 146260 274904 146266 274916
rect 185578 274904 185584 274916
rect 146260 274876 185584 274904
rect 146260 274864 146266 274876
rect 185578 274864 185584 274876
rect 185636 274864 185642 274916
rect 473078 274864 473084 274916
rect 473136 274904 473142 274916
rect 544562 274904 544568 274916
rect 473136 274876 544568 274904
rect 473136 274864 473142 274876
rect 544562 274864 544568 274876
rect 544620 274864 544626 274916
rect 289262 274796 289268 274848
rect 289320 274836 289326 274848
rect 293402 274836 293408 274848
rect 289320 274808 293408 274836
rect 289320 274796 289326 274808
rect 293402 274796 293408 274808
rect 293460 274796 293466 274848
rect 295150 274796 295156 274848
rect 295208 274836 295214 274848
rect 297450 274836 297456 274848
rect 295208 274808 297456 274836
rect 295208 274796 295214 274808
rect 297450 274796 297456 274808
rect 297508 274796 297514 274848
rect 128538 274728 128544 274780
rect 128596 274768 128602 274780
rect 168282 274768 168288 274780
rect 128596 274740 168288 274768
rect 128596 274728 128602 274740
rect 168282 274728 168288 274740
rect 168340 274728 168346 274780
rect 207750 274728 207756 274780
rect 207808 274768 207814 274780
rect 210694 274768 210700 274780
rect 207808 274740 210700 274768
rect 207808 274728 207814 274740
rect 210694 274728 210700 274740
rect 210752 274728 210758 274780
rect 476758 274728 476764 274780
rect 476816 274768 476822 274780
rect 523310 274768 523316 274780
rect 476816 274740 523316 274768
rect 476816 274728 476822 274740
rect 523310 274728 523316 274740
rect 523368 274728 523374 274780
rect 523678 274728 523684 274780
rect 523736 274768 523742 274780
rect 533890 274768 533896 274780
rect 523736 274740 533896 274768
rect 523736 274728 523742 274740
rect 533890 274728 533896 274740
rect 533948 274728 533954 274780
rect 534718 274728 534724 274780
rect 534776 274768 534782 274780
rect 540974 274768 540980 274780
rect 534776 274740 540980 274768
rect 534776 274728 534782 274740
rect 540974 274728 540980 274740
rect 541032 274728 541038 274780
rect 74166 274660 74172 274712
rect 74224 274700 74230 274712
rect 76834 274700 76840 274712
rect 74224 274672 76840 274700
rect 74224 274660 74230 274672
rect 76834 274660 76840 274672
rect 76892 274660 76898 274712
rect 85942 274660 85948 274712
rect 86000 274700 86006 274712
rect 90358 274700 90364 274712
rect 86000 274672 90364 274700
rect 86000 274660 86006 274672
rect 90358 274660 90364 274672
rect 90416 274660 90422 274712
rect 103698 274660 103704 274712
rect 103756 274700 103762 274712
rect 104802 274700 104808 274712
rect 103756 274672 104808 274700
rect 103756 274660 103762 274672
rect 104802 274660 104808 274672
rect 104860 274660 104866 274712
rect 110782 274660 110788 274712
rect 110840 274700 110846 274712
rect 111702 274700 111708 274712
rect 110840 274672 111708 274700
rect 110840 274660 110846 274672
rect 111702 274660 111708 274672
rect 111760 274660 111766 274712
rect 253842 274660 253848 274712
rect 253900 274700 253906 274712
rect 256878 274700 256884 274712
rect 253900 274672 256884 274700
rect 253900 274660 253906 274672
rect 256878 274660 256884 274672
rect 256936 274660 256942 274712
rect 275094 274660 275100 274712
rect 275152 274700 275158 274712
rect 278038 274700 278044 274712
rect 275152 274672 278044 274700
rect 275152 274660 275158 274672
rect 278038 274660 278044 274672
rect 278096 274660 278102 274712
rect 283374 274660 283380 274712
rect 283432 274700 283438 274712
rect 289170 274700 289176 274712
rect 283432 274672 289176 274700
rect 283432 274660 283438 274672
rect 289170 274660 289176 274672
rect 289228 274660 289234 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 303430 274660 303436 274712
rect 303488 274700 303494 274712
rect 303982 274700 303988 274712
rect 303488 274672 303988 274700
rect 303488 274660 303494 274672
rect 303982 274660 303988 274672
rect 304040 274660 304046 274712
rect 321186 274660 321192 274712
rect 321244 274700 321250 274712
rect 328270 274700 328276 274712
rect 321244 274672 328276 274700
rect 321244 274660 321250 274672
rect 328270 274660 328276 274672
rect 328328 274660 328334 274712
rect 114370 274592 114376 274644
rect 114428 274632 114434 274644
rect 171594 274632 171600 274644
rect 114428 274604 171600 274632
rect 114428 274592 114434 274604
rect 171594 274592 171600 274604
rect 171652 274592 171658 274644
rect 179322 274592 179328 274644
rect 179380 274632 179386 274644
rect 214558 274632 214564 274644
rect 179380 274604 214564 274632
rect 179380 274592 179386 274604
rect 214558 274592 214564 274604
rect 214616 274592 214622 274644
rect 409782 274592 409788 274644
rect 409840 274632 409846 274644
rect 453574 274632 453580 274644
rect 409840 274604 453580 274632
rect 409840 274592 409846 274604
rect 453574 274592 453580 274604
rect 453632 274592 453638 274644
rect 457438 274592 457444 274644
rect 457496 274632 457502 274644
rect 480714 274632 480720 274644
rect 457496 274604 480720 274632
rect 457496 274592 457502 274604
rect 480714 274592 480720 274604
rect 480772 274592 480778 274644
rect 486786 274592 486792 274644
rect 486844 274632 486850 274644
rect 563422 274632 563428 274644
rect 486844 274604 563428 274632
rect 486844 274592 486850 274604
rect 563422 274592 563428 274604
rect 563480 274592 563486 274644
rect 101306 274456 101312 274508
rect 101364 274496 101370 274508
rect 160922 274496 160928 274508
rect 101364 274468 160928 274496
rect 101364 274456 101370 274468
rect 160922 274456 160928 274468
rect 160980 274456 160986 274508
rect 168742 274456 168748 274508
rect 168800 274496 168806 274508
rect 208394 274496 208400 274508
rect 168800 274468 208400 274496
rect 168800 274456 168806 274468
rect 208394 274456 208400 274468
rect 208452 274456 208458 274508
rect 381538 274456 381544 274508
rect 381596 274496 381602 274508
rect 392118 274496 392124 274508
rect 381596 274468 392124 274496
rect 381596 274456 381602 274468
rect 392118 274456 392124 274468
rect 392176 274456 392182 274508
rect 413830 274456 413836 274508
rect 413888 274496 413894 274508
rect 460658 274496 460664 274508
rect 413888 274468 460664 274496
rect 413888 274456 413894 274468
rect 460658 274456 460664 274468
rect 460716 274456 460722 274508
rect 463234 274456 463240 274508
rect 463292 274496 463298 274508
rect 484302 274496 484308 274508
rect 463292 274468 484308 274496
rect 463292 274456 463298 274468
rect 484302 274456 484308 274468
rect 484360 274456 484366 274508
rect 488350 274456 488356 274508
rect 488408 274496 488414 274508
rect 567010 274496 567016 274508
rect 488408 274468 567016 274496
rect 488408 274456 488414 274468
rect 567010 274456 567016 274468
rect 567068 274456 567074 274508
rect 95418 274320 95424 274372
rect 95476 274360 95482 274372
rect 157610 274360 157616 274372
rect 95476 274332 157616 274360
rect 95476 274320 95482 274332
rect 157610 274320 157616 274332
rect 157668 274320 157674 274372
rect 159266 274320 159272 274372
rect 159324 274360 159330 274372
rect 202322 274360 202328 274372
rect 159324 274332 202328 274360
rect 159324 274320 159330 274332
rect 202322 274320 202328 274332
rect 202380 274320 202386 274372
rect 223114 274320 223120 274372
rect 223172 274360 223178 274372
rect 247218 274360 247224 274372
rect 223172 274332 247224 274360
rect 223172 274320 223178 274332
rect 247218 274320 247224 274332
rect 247276 274320 247282 274372
rect 369118 274320 369124 274372
rect 369176 274360 369182 274372
rect 387334 274360 387340 274372
rect 369176 274332 387340 274360
rect 369176 274320 369182 274332
rect 387334 274320 387340 274332
rect 387392 274320 387398 274372
rect 419074 274320 419080 274372
rect 419132 274360 419138 274372
rect 467742 274360 467748 274372
rect 419132 274332 467748 274360
rect 419132 274320 419138 274332
rect 467742 274320 467748 274332
rect 467800 274320 467806 274372
rect 506198 274320 506204 274372
rect 506256 274360 506262 274372
rect 591850 274360 591856 274372
rect 506256 274332 591856 274360
rect 506256 274320 506262 274332
rect 591850 274320 591856 274332
rect 591908 274320 591914 274372
rect 67082 274184 67088 274236
rect 67140 274224 67146 274236
rect 130378 274224 130384 274236
rect 67140 274196 130384 274224
rect 67140 274184 67146 274196
rect 130378 274184 130384 274196
rect 130436 274184 130442 274236
rect 130838 274184 130844 274236
rect 130896 274224 130902 274236
rect 182450 274224 182456 274236
rect 130896 274196 182456 274224
rect 130896 274184 130902 274196
rect 182450 274184 182456 274196
rect 182508 274184 182514 274236
rect 192386 274184 192392 274236
rect 192444 274224 192450 274236
rect 224954 274224 224960 274236
rect 192444 274196 224960 274224
rect 192444 274184 192450 274196
rect 224954 274184 224960 274196
rect 225012 274184 225018 274236
rect 239214 274184 239220 274236
rect 239272 274224 239278 274236
rect 253934 274224 253940 274236
rect 239272 274196 253940 274224
rect 239272 274184 239278 274196
rect 253934 274184 253940 274196
rect 253992 274184 253998 274236
rect 331858 274184 331864 274236
rect 331916 274224 331922 274236
rect 337746 274224 337752 274236
rect 331916 274196 337752 274224
rect 331916 274184 331922 274196
rect 337746 274184 337752 274196
rect 337804 274184 337810 274236
rect 359458 274184 359464 274236
rect 359516 274224 359522 274236
rect 380250 274224 380256 274236
rect 359516 274196 380256 274224
rect 359516 274184 359522 274196
rect 380250 274184 380256 274196
rect 380308 274184 380314 274236
rect 388990 274184 388996 274236
rect 389048 274224 389054 274236
rect 425238 274224 425244 274236
rect 389048 274196 425244 274224
rect 389048 274184 389054 274196
rect 425238 274184 425244 274196
rect 425296 274184 425302 274236
rect 425698 274184 425704 274236
rect 425756 274224 425762 274236
rect 474826 274224 474832 274236
rect 425756 274196 474832 274224
rect 425756 274184 425762 274196
rect 474826 274184 474832 274196
rect 474884 274184 474890 274236
rect 511810 274184 511816 274236
rect 511868 274224 511874 274236
rect 598934 274224 598940 274236
rect 511868 274196 598940 274224
rect 511868 274184 511874 274196
rect 598934 274184 598940 274196
rect 598992 274184 598998 274236
rect 77662 274048 77668 274100
rect 77720 274088 77726 274100
rect 145098 274088 145104 274100
rect 77720 274060 145104 274088
rect 77720 274048 77726 274060
rect 145098 274048 145104 274060
rect 145156 274048 145162 274100
rect 154482 274048 154488 274100
rect 154540 274088 154546 274100
rect 198090 274088 198096 274100
rect 154540 274060 198096 274088
rect 154540 274048 154546 274060
rect 198090 274048 198096 274060
rect 198148 274048 198154 274100
rect 210050 274048 210056 274100
rect 210108 274088 210114 274100
rect 237834 274088 237840 274100
rect 210108 274060 237840 274088
rect 210108 274048 210114 274060
rect 237834 274048 237840 274060
rect 237892 274048 237898 274100
rect 249058 274048 249064 274100
rect 249116 274088 249122 274100
rect 265250 274088 265256 274100
rect 249116 274060 265256 274088
rect 249116 274048 249122 274060
rect 265250 274048 265256 274060
rect 265308 274048 265314 274100
rect 266354 274048 266360 274100
rect 266412 274088 266418 274100
rect 273530 274088 273536 274100
rect 266412 274060 273536 274088
rect 266412 274048 266418 274060
rect 273530 274048 273536 274060
rect 273588 274048 273594 274100
rect 278590 274048 278596 274100
rect 278648 274088 278654 274100
rect 285858 274088 285864 274100
rect 278648 274060 285864 274088
rect 278648 274048 278654 274060
rect 285858 274048 285864 274060
rect 285916 274048 285922 274100
rect 337746 274048 337752 274100
rect 337804 274088 337810 274100
rect 351914 274088 351920 274100
rect 337804 274060 351920 274088
rect 337804 274048 337810 274060
rect 351914 274048 351920 274060
rect 351972 274048 351978 274100
rect 353938 274048 353944 274100
rect 353996 274088 354002 274100
rect 369578 274088 369584 274100
rect 353996 274060 369584 274088
rect 353996 274048 354002 274060
rect 369578 274048 369584 274060
rect 369636 274048 369642 274100
rect 373258 274048 373264 274100
rect 373316 274088 373322 274100
rect 400306 274088 400312 274100
rect 373316 274060 400312 274088
rect 373316 274048 373322 274060
rect 400306 274048 400312 274060
rect 400364 274048 400370 274100
rect 401502 274048 401508 274100
rect 401560 274088 401566 274100
rect 442902 274088 442908 274100
rect 401560 274060 442908 274088
rect 401560 274048 401566 274060
rect 442902 274048 442908 274060
rect 442960 274048 442966 274100
rect 451182 274048 451188 274100
rect 451240 274088 451246 274100
rect 513834 274088 513840 274100
rect 451240 274060 513840 274088
rect 451240 274048 451246 274060
rect 513834 274048 513840 274060
rect 513892 274048 513898 274100
rect 536742 274048 536748 274100
rect 536800 274088 536806 274100
rect 634354 274088 634360 274100
rect 536800 274060 634360 274088
rect 536800 274048 536806 274060
rect 634354 274048 634360 274060
rect 634412 274048 634418 274100
rect 69382 273912 69388 273964
rect 69440 273952 69446 273964
rect 139394 273952 139400 273964
rect 69440 273924 139400 273952
rect 69440 273912 69446 273924
rect 139394 273912 139400 273924
rect 139452 273912 139458 273964
rect 144914 273912 144920 273964
rect 144972 273952 144978 273964
rect 147858 273952 147864 273964
rect 144972 273924 147864 273952
rect 144972 273912 144978 273924
rect 147858 273912 147864 273924
rect 147916 273912 147922 273964
rect 148594 273912 148600 273964
rect 148652 273952 148658 273964
rect 194778 273952 194784 273964
rect 148652 273924 194784 273952
rect 148652 273912 148658 273924
rect 194778 273912 194784 273924
rect 194836 273912 194842 273964
rect 208854 273912 208860 273964
rect 208912 273952 208918 273964
rect 237374 273952 237380 273964
rect 208912 273924 237380 273952
rect 208912 273912 208918 273924
rect 237374 273912 237380 273924
rect 237432 273912 237438 273964
rect 238478 273912 238484 273964
rect 238536 273952 238542 273964
rect 238536 273924 238754 273952
rect 238536 273912 238542 273924
rect 88334 273776 88340 273828
rect 88392 273816 88398 273828
rect 119338 273816 119344 273828
rect 88392 273788 119344 273816
rect 88392 273776 88398 273788
rect 119338 273776 119344 273788
rect 119396 273776 119402 273828
rect 120258 273776 120264 273828
rect 120316 273816 120322 273828
rect 175274 273816 175280 273828
rect 120316 273788 175280 273816
rect 120316 273776 120322 273788
rect 175274 273776 175280 273788
rect 175332 273776 175338 273828
rect 193490 273776 193496 273828
rect 193548 273816 193554 273828
rect 226426 273816 226432 273828
rect 193548 273788 226432 273816
rect 193548 273776 193554 273788
rect 226426 273776 226432 273788
rect 226484 273776 226490 273828
rect 238726 273816 238754 273924
rect 271506 273912 271512 273964
rect 271564 273952 271570 273964
rect 280338 273952 280344 273964
rect 271564 273924 280344 273952
rect 271564 273912 271570 273924
rect 280338 273912 280344 273924
rect 280396 273912 280402 273964
rect 322750 273912 322756 273964
rect 322808 273952 322814 273964
rect 330570 273952 330576 273964
rect 322808 273924 330576 273952
rect 322808 273912 322814 273924
rect 330570 273912 330576 273924
rect 330628 273912 330634 273964
rect 335262 273912 335268 273964
rect 335320 273952 335326 273964
rect 348326 273952 348332 273964
rect 335320 273924 348332 273952
rect 335320 273912 335326 273924
rect 348326 273912 348332 273924
rect 348384 273912 348390 273964
rect 350350 273912 350356 273964
rect 350408 273952 350414 273964
rect 368474 273952 368480 273964
rect 350408 273924 368480 273952
rect 350408 273912 350414 273924
rect 368474 273912 368480 273924
rect 368532 273912 368538 273964
rect 377674 273912 377680 273964
rect 377732 273952 377738 273964
rect 408586 273952 408592 273964
rect 377732 273924 408592 273952
rect 377732 273912 377738 273924
rect 408586 273912 408592 273924
rect 408644 273912 408650 273964
rect 422110 273912 422116 273964
rect 422168 273952 422174 273964
rect 472434 273952 472440 273964
rect 422168 273924 472440 273952
rect 422168 273912 422174 273924
rect 472434 273912 472440 273924
rect 472492 273912 472498 273964
rect 474642 273912 474648 273964
rect 474700 273952 474706 273964
rect 545758 273952 545764 273964
rect 474700 273924 545764 273952
rect 474700 273912 474706 273924
rect 545758 273912 545764 273924
rect 545816 273912 545822 273964
rect 545942 273912 545948 273964
rect 546000 273952 546006 273964
rect 639138 273952 639144 273964
rect 546000 273924 639144 273952
rect 546000 273912 546006 273924
rect 639138 273912 639144 273924
rect 639196 273912 639202 273964
rect 258074 273816 258080 273828
rect 238726 273788 258080 273816
rect 258074 273776 258080 273788
rect 258132 273776 258138 273828
rect 259362 273776 259368 273828
rect 259420 273816 259426 273828
rect 266354 273816 266360 273828
rect 259420 273788 266360 273816
rect 259420 273776 259426 273788
rect 266354 273776 266360 273788
rect 266412 273776 266418 273828
rect 396994 273776 397000 273828
rect 397052 273816 397058 273828
rect 435818 273816 435824 273828
rect 397052 273788 435824 273816
rect 397052 273776 397058 273788
rect 435818 273776 435824 273788
rect 435876 273776 435882 273828
rect 438118 273776 438124 273828
rect 438176 273816 438182 273828
rect 473630 273816 473636 273828
rect 438176 273788 473636 273816
rect 438176 273776 438182 273788
rect 473630 273776 473636 273788
rect 473688 273776 473694 273828
rect 481358 273776 481364 273828
rect 481416 273816 481422 273828
rect 556338 273816 556344 273828
rect 481416 273788 556344 273816
rect 481416 273776 481422 273788
rect 556338 273776 556344 273788
rect 556396 273776 556402 273828
rect 556798 273776 556804 273828
rect 556856 273816 556862 273828
rect 590654 273816 590660 273828
rect 556856 273788 590660 273816
rect 556856 273776 556862 273788
rect 590654 273776 590660 273788
rect 590712 273776 590718 273828
rect 119062 273640 119068 273692
rect 119120 273680 119126 273692
rect 173250 273680 173256 273692
rect 119120 273652 173256 273680
rect 119120 273640 119126 273652
rect 173250 273640 173256 273652
rect 173308 273640 173314 273692
rect 447778 273640 447784 273692
rect 447836 273680 447842 273692
rect 481910 273680 481916 273692
rect 447836 273652 481916 273680
rect 447836 273640 447842 273652
rect 481910 273640 481916 273652
rect 481968 273640 481974 273692
rect 484210 273640 484216 273692
rect 484268 273680 484274 273692
rect 559926 273680 559932 273692
rect 484268 273652 559932 273680
rect 484268 273640 484274 273652
rect 559926 273640 559932 273652
rect 559984 273640 559990 273692
rect 132034 273504 132040 273556
rect 132092 273544 132098 273556
rect 153838 273544 153844 273556
rect 132092 273516 153844 273544
rect 132092 273504 132098 273516
rect 153838 273504 153844 273516
rect 153896 273504 153902 273556
rect 440878 273504 440884 273556
rect 440936 273544 440942 273556
rect 471238 273544 471244 273556
rect 440936 273516 471244 273544
rect 440936 273504 440942 273516
rect 471238 273504 471244 273516
rect 471296 273504 471302 273556
rect 476022 273504 476028 273556
rect 476080 273544 476086 273556
rect 549254 273544 549260 273556
rect 476080 273516 549260 273544
rect 476080 273504 476086 273516
rect 549254 273504 549260 273516
rect 549312 273504 549318 273556
rect 549898 273504 549904 273556
rect 549956 273544 549962 273556
rect 583570 273544 583576 273556
rect 549956 273516 583576 273544
rect 549956 273504 549962 273516
rect 583570 273504 583576 273516
rect 583628 273504 583634 273556
rect 478690 273368 478696 273420
rect 478748 273408 478754 273420
rect 552842 273408 552848 273420
rect 478748 273380 552848 273408
rect 478748 273368 478754 273380
rect 552842 273368 552848 273380
rect 552900 273368 552906 273420
rect 460566 273300 460572 273352
rect 460624 273340 460630 273352
rect 461394 273340 461400 273352
rect 460624 273312 461400 273340
rect 460624 273300 460630 273312
rect 461394 273300 461400 273312
rect 461452 273300 461458 273352
rect 327718 273232 327724 273284
rect 327776 273272 327782 273284
rect 329466 273272 329472 273284
rect 327776 273244 329472 273272
rect 327776 273232 327782 273244
rect 329466 273232 329472 273244
rect 329524 273232 329530 273284
rect 108390 273164 108396 273216
rect 108448 273204 108454 273216
rect 165890 273204 165896 273216
rect 108448 273176 165896 273204
rect 108448 273164 108454 273176
rect 165890 273164 165896 273176
rect 165948 273164 165954 273216
rect 186406 273164 186412 273216
rect 186464 273204 186470 273216
rect 218698 273204 218704 273216
rect 186464 273176 218704 273204
rect 186464 273164 186470 273176
rect 218698 273164 218704 273176
rect 218756 273164 218762 273216
rect 362770 273164 362776 273216
rect 362828 273204 362834 273216
rect 385862 273204 385868 273216
rect 362828 273176 385868 273204
rect 362828 273164 362834 273176
rect 385862 273164 385868 273176
rect 385920 273164 385926 273216
rect 400030 273164 400036 273216
rect 400088 273204 400094 273216
rect 439314 273204 439320 273216
rect 400088 273176 439320 273204
rect 400088 273164 400094 273176
rect 439314 273164 439320 273176
rect 439372 273164 439378 273216
rect 444006 273164 444012 273216
rect 444064 273204 444070 273216
rect 503162 273204 503168 273216
rect 444064 273176 503168 273204
rect 444064 273164 444070 273176
rect 503162 273164 503168 273176
rect 503220 273164 503226 273216
rect 504174 273164 504180 273216
rect 504232 273204 504238 273216
rect 511442 273204 511448 273216
rect 504232 273176 511448 273204
rect 504232 273164 504238 273176
rect 511442 273164 511448 273176
rect 511500 273164 511506 273216
rect 518526 273204 518532 273216
rect 512012 273176 518532 273204
rect 102502 273028 102508 273080
rect 102560 273068 102566 273080
rect 162854 273068 162860 273080
rect 102560 273040 162860 273068
rect 102560 273028 102566 273040
rect 162854 273028 162860 273040
rect 162912 273028 162918 273080
rect 172238 273028 172244 273080
rect 172296 273068 172302 273080
rect 209774 273068 209780 273080
rect 172296 273040 209780 273068
rect 172296 273028 172302 273040
rect 209774 273028 209780 273040
rect 209832 273028 209838 273080
rect 219526 273028 219532 273080
rect 219584 273068 219590 273080
rect 244550 273068 244556 273080
rect 219584 273040 244556 273068
rect 219584 273028 219590 273040
rect 244550 273028 244556 273040
rect 244608 273028 244614 273080
rect 280982 273028 280988 273080
rect 281040 273068 281046 273080
rect 286318 273068 286324 273080
rect 281040 273040 286324 273068
rect 281040 273028 281046 273040
rect 286318 273028 286324 273040
rect 286376 273028 286382 273080
rect 361206 273028 361212 273080
rect 361264 273068 361270 273080
rect 384942 273068 384948 273080
rect 361264 273040 384948 273068
rect 361264 273028 361270 273040
rect 384942 273028 384948 273040
rect 385000 273028 385006 273080
rect 385678 273028 385684 273080
rect 385736 273068 385742 273080
rect 395614 273068 395620 273080
rect 385736 273040 395620 273068
rect 385736 273028 385742 273040
rect 395614 273028 395620 273040
rect 395672 273028 395678 273080
rect 404170 273028 404176 273080
rect 404228 273068 404234 273080
rect 446490 273068 446496 273080
rect 404228 273040 446496 273068
rect 404228 273028 404234 273040
rect 446490 273028 446496 273040
rect 446548 273028 446554 273080
rect 452286 273028 452292 273080
rect 452344 273068 452350 273080
rect 452344 273040 461624 273068
rect 452344 273028 452350 273040
rect 94222 272892 94228 272944
rect 94280 272932 94286 272944
rect 156138 272932 156144 272944
rect 94280 272904 156144 272932
rect 94280 272892 94286 272904
rect 156138 272892 156144 272904
rect 156196 272892 156202 272944
rect 166350 272892 166356 272944
rect 166408 272932 166414 272944
rect 207290 272932 207296 272944
rect 166408 272904 207296 272932
rect 166408 272892 166414 272904
rect 207290 272892 207296 272904
rect 207348 272892 207354 272944
rect 211246 272892 211252 272944
rect 211304 272932 211310 272944
rect 220078 272932 220084 272944
rect 211304 272904 220084 272932
rect 211304 272892 211310 272904
rect 220078 272892 220084 272904
rect 220136 272892 220142 272944
rect 220722 272892 220728 272944
rect 220780 272932 220786 272944
rect 245746 272932 245752 272944
rect 220780 272904 245752 272932
rect 220780 272892 220786 272904
rect 245746 272892 245752 272904
rect 245804 272892 245810 272944
rect 247862 272892 247868 272944
rect 247920 272932 247926 272944
rect 264238 272932 264244 272944
rect 247920 272904 264244 272932
rect 247920 272892 247926 272904
rect 264238 272892 264244 272904
rect 264296 272892 264302 272944
rect 333790 272892 333796 272944
rect 333848 272932 333854 272944
rect 345934 272932 345940 272944
rect 333848 272904 345940 272932
rect 333848 272892 333854 272904
rect 345934 272892 345940 272904
rect 345992 272892 345998 272944
rect 348418 272892 348424 272944
rect 348476 272932 348482 272944
rect 362494 272932 362500 272944
rect 348476 272904 362500 272932
rect 348476 272892 348482 272904
rect 362494 272892 362500 272904
rect 362552 272892 362558 272944
rect 365438 272892 365444 272944
rect 365496 272932 365502 272944
rect 390922 272932 390928 272944
rect 365496 272904 390928 272932
rect 365496 272892 365502 272904
rect 390922 272892 390928 272904
rect 390980 272892 390986 272944
rect 405550 272892 405556 272944
rect 405608 272932 405614 272944
rect 448790 272932 448796 272944
rect 405608 272904 448796 272932
rect 405608 272892 405614 272904
rect 448790 272892 448796 272904
rect 448848 272892 448854 272944
rect 455322 272892 455328 272944
rect 455380 272932 455386 272944
rect 460566 272932 460572 272944
rect 455380 272904 460572 272932
rect 455380 272892 455386 272904
rect 460566 272892 460572 272904
rect 460624 272892 460630 272944
rect 461596 272932 461624 273040
rect 461762 273028 461768 273080
rect 461820 273068 461826 273080
rect 512012 273068 512040 273176
rect 518526 273164 518532 273176
rect 518584 273164 518590 273216
rect 519722 273204 519728 273216
rect 518866 273176 519728 273204
rect 515030 273068 515036 273080
rect 461820 273040 512040 273068
rect 512104 273040 515036 273068
rect 461820 273028 461826 273040
rect 512104 272932 512132 273040
rect 515030 273028 515036 273040
rect 515088 273028 515094 273080
rect 515398 273028 515404 273080
rect 515456 273068 515462 273080
rect 518866 273068 518894 273176
rect 519722 273164 519728 273176
rect 519780 273164 519786 273216
rect 521470 273164 521476 273216
rect 521528 273204 521534 273216
rect 614298 273204 614304 273216
rect 521528 273176 614304 273204
rect 521528 273164 521534 273176
rect 614298 273164 614304 273176
rect 614356 273164 614362 273216
rect 515456 273040 518894 273068
rect 515456 273028 515462 273040
rect 526806 273028 526812 273080
rect 526864 273068 526870 273080
rect 621382 273068 621388 273080
rect 526864 273040 621388 273068
rect 526864 273028 526870 273040
rect 621382 273028 621388 273040
rect 621440 273028 621446 273080
rect 525610 272932 525616 272944
rect 461596 272904 512132 272932
rect 514036 272904 525616 272932
rect 82446 272756 82452 272808
rect 82504 272796 82510 272808
rect 148410 272796 148416 272808
rect 82504 272768 148416 272796
rect 82504 272756 82510 272768
rect 148410 272756 148416 272768
rect 148468 272756 148474 272808
rect 155678 272756 155684 272808
rect 155736 272796 155742 272808
rect 200114 272796 200120 272808
rect 155736 272768 200120 272796
rect 155736 272756 155742 272768
rect 200114 272756 200120 272768
rect 200172 272756 200178 272808
rect 205358 272756 205364 272808
rect 205416 272796 205422 272808
rect 234798 272796 234804 272808
rect 205416 272768 234804 272796
rect 205416 272756 205422 272768
rect 234798 272756 234804 272768
rect 234856 272756 234862 272808
rect 245378 272756 245384 272808
rect 245436 272796 245442 272808
rect 245436 272768 258074 272796
rect 245436 272756 245442 272768
rect 72970 272620 72976 272672
rect 73028 272660 73034 272672
rect 142154 272660 142160 272672
rect 73028 272632 142160 272660
rect 73028 272620 73034 272632
rect 142154 272620 142160 272632
rect 142212 272620 142218 272672
rect 142706 272620 142712 272672
rect 142764 272660 142770 272672
rect 145558 272660 145564 272672
rect 142764 272632 145564 272660
rect 142764 272620 142770 272632
rect 145558 272620 145564 272632
rect 145616 272620 145622 272672
rect 145742 272620 145748 272672
rect 145800 272660 145806 272672
rect 192386 272660 192392 272672
rect 145800 272632 192392 272660
rect 145800 272620 145806 272632
rect 192386 272620 192392 272632
rect 192444 272620 192450 272672
rect 197078 272620 197084 272672
rect 197136 272660 197142 272672
rect 229094 272660 229100 272672
rect 197136 272632 229100 272660
rect 197136 272620 197142 272632
rect 229094 272620 229100 272632
rect 229152 272620 229158 272672
rect 233694 272620 233700 272672
rect 233752 272660 233758 272672
rect 254394 272660 254400 272672
rect 233752 272632 254400 272660
rect 233752 272620 233758 272632
rect 254394 272620 254400 272632
rect 254452 272620 254458 272672
rect 258046 272660 258074 272768
rect 262306 272756 262312 272808
rect 262364 272796 262370 272808
rect 270954 272796 270960 272808
rect 262364 272768 270960 272796
rect 262364 272756 262370 272768
rect 270954 272756 270960 272768
rect 271012 272756 271018 272808
rect 274266 272756 274272 272808
rect 274324 272796 274330 272808
rect 282914 272796 282920 272808
rect 274324 272768 282920 272796
rect 274324 272756 274330 272768
rect 282914 272756 282920 272768
rect 282972 272756 282978 272808
rect 325326 272756 325332 272808
rect 325384 272796 325390 272808
rect 332962 272796 332968 272808
rect 325384 272768 332968 272796
rect 325384 272756 325390 272768
rect 332962 272756 332968 272768
rect 333020 272756 333026 272808
rect 344646 272756 344652 272808
rect 344704 272796 344710 272808
rect 361390 272796 361396 272808
rect 344704 272768 361396 272796
rect 344704 272756 344710 272768
rect 361390 272756 361396 272768
rect 361448 272756 361454 272808
rect 362218 272756 362224 272808
rect 362276 272796 362282 272808
rect 370314 272796 370320 272808
rect 362276 272768 370320 272796
rect 362276 272756 362282 272768
rect 370314 272756 370320 272768
rect 370372 272756 370378 272808
rect 370498 272756 370504 272808
rect 370556 272796 370562 272808
rect 396810 272796 396816 272808
rect 370556 272768 396816 272796
rect 370556 272756 370562 272768
rect 396810 272756 396816 272768
rect 396868 272756 396874 272808
rect 406838 272756 406844 272808
rect 406896 272796 406902 272808
rect 449986 272796 449992 272808
rect 406896 272768 449992 272796
rect 406896 272756 406902 272768
rect 449986 272756 449992 272768
rect 450044 272756 450050 272808
rect 450538 272756 450544 272808
rect 450596 272796 450602 272808
rect 501046 272796 501052 272808
rect 450596 272768 501052 272796
rect 450596 272756 450602 272768
rect 501046 272756 501052 272768
rect 501104 272756 501110 272808
rect 504358 272756 504364 272808
rect 504416 272796 504422 272808
rect 514036 272796 514064 272904
rect 525610 272892 525616 272904
rect 525668 272892 525674 272944
rect 532510 272892 532516 272944
rect 532568 272932 532574 272944
rect 537938 272932 537944 272944
rect 532568 272904 537944 272932
rect 532568 272892 532574 272904
rect 537938 272892 537944 272904
rect 537996 272892 538002 272944
rect 538122 272892 538128 272944
rect 538180 272932 538186 272944
rect 624970 272932 624976 272944
rect 538180 272904 624976 272932
rect 538180 272892 538186 272904
rect 624970 272892 624976 272904
rect 625028 272892 625034 272944
rect 504416 272768 514064 272796
rect 504416 272756 504422 272768
rect 514202 272756 514208 272808
rect 514260 272796 514266 272808
rect 562134 272796 562140 272808
rect 514260 272768 562140 272796
rect 514260 272756 514266 272768
rect 562134 272756 562140 272768
rect 562192 272756 562198 272808
rect 562318 272756 562324 272808
rect 562376 272796 562382 272808
rect 601142 272796 601148 272808
rect 562376 272768 601148 272796
rect 562376 272756 562382 272768
rect 601142 272756 601148 272768
rect 601200 272756 601206 272808
rect 262674 272660 262680 272672
rect 258046 272632 262680 272660
rect 262674 272620 262680 272632
rect 262732 272620 262738 272672
rect 264422 272620 264428 272672
rect 264480 272660 264486 272672
rect 276014 272660 276020 272672
rect 264480 272632 276020 272660
rect 264480 272620 264486 272632
rect 276014 272620 276020 272632
rect 276072 272620 276078 272672
rect 324038 272620 324044 272672
rect 324096 272660 324102 272672
rect 331398 272660 331404 272672
rect 324096 272632 331404 272660
rect 324096 272620 324102 272632
rect 331398 272620 331404 272632
rect 331456 272620 331462 272672
rect 332318 272620 332324 272672
rect 332376 272660 332382 272672
rect 343634 272660 343640 272672
rect 332376 272632 343640 272660
rect 332376 272620 332382 272632
rect 343634 272620 343640 272632
rect 343692 272620 343698 272672
rect 346210 272620 346216 272672
rect 346268 272660 346274 272672
rect 363690 272660 363696 272672
rect 346268 272632 363696 272660
rect 346268 272620 346274 272632
rect 363690 272620 363696 272632
rect 363748 272620 363754 272672
rect 376110 272620 376116 272672
rect 376168 272660 376174 272672
rect 406286 272660 406292 272672
rect 376168 272632 406292 272660
rect 376168 272620 376174 272632
rect 406286 272620 406292 272632
rect 406344 272620 406350 272672
rect 412266 272620 412272 272672
rect 412324 272660 412330 272672
rect 457070 272660 457076 272672
rect 412324 272632 457076 272660
rect 412324 272620 412330 272632
rect 457070 272620 457076 272632
rect 457128 272620 457134 272672
rect 457254 272620 457260 272672
rect 457312 272660 457318 272672
rect 459370 272660 459376 272672
rect 457312 272632 459376 272660
rect 457312 272620 457318 272632
rect 459370 272620 459376 272632
rect 459428 272620 459434 272672
rect 459554 272620 459560 272672
rect 459612 272660 459618 272672
rect 459612 272632 464108 272660
rect 459612 272620 459618 272632
rect 464080 272592 464108 272632
rect 466408 272620 466414 272672
rect 466466 272660 466472 272672
rect 522114 272660 522120 272672
rect 466466 272632 522120 272660
rect 466466 272620 466472 272632
rect 522114 272620 522120 272632
rect 522172 272620 522178 272672
rect 529842 272620 529848 272672
rect 529900 272660 529906 272672
rect 529900 272632 532924 272660
rect 529900 272620 529906 272632
rect 464080 272564 466316 272592
rect 65886 272484 65892 272536
rect 65944 272524 65950 272536
rect 136818 272524 136824 272536
rect 65944 272496 136824 272524
rect 65944 272484 65950 272496
rect 136818 272484 136824 272496
rect 136876 272484 136882 272536
rect 137922 272484 137928 272536
rect 137980 272524 137986 272536
rect 137980 272496 180794 272524
rect 137980 272484 137986 272496
rect 116670 272348 116676 272400
rect 116728 272388 116734 272400
rect 172514 272388 172520 272400
rect 116728 272360 172520 272388
rect 116728 272348 116734 272360
rect 172514 272348 172520 272360
rect 172572 272348 172578 272400
rect 180766 272388 180794 272496
rect 181714 272484 181720 272536
rect 181772 272524 181778 272536
rect 186958 272524 186964 272536
rect 181772 272496 186964 272524
rect 181772 272484 181778 272496
rect 186958 272484 186964 272496
rect 187016 272484 187022 272536
rect 195882 272484 195888 272536
rect 195940 272524 195946 272536
rect 227898 272524 227904 272536
rect 195940 272496 227904 272524
rect 195940 272484 195946 272496
rect 227898 272484 227904 272496
rect 227956 272484 227962 272536
rect 228082 272484 228088 272536
rect 228140 272524 228146 272536
rect 249058 272524 249064 272536
rect 228140 272496 249064 272524
rect 228140 272484 228146 272496
rect 249058 272484 249064 272496
rect 249116 272484 249122 272536
rect 254946 272484 254952 272536
rect 255004 272524 255010 272536
rect 269298 272524 269304 272536
rect 255004 272496 269304 272524
rect 255004 272484 255010 272496
rect 269298 272484 269304 272496
rect 269356 272484 269362 272536
rect 270310 272484 270316 272536
rect 270368 272524 270374 272536
rect 280522 272524 280528 272536
rect 270368 272496 280528 272524
rect 270368 272484 270374 272496
rect 280522 272484 280528 272496
rect 280580 272484 280586 272536
rect 329742 272484 329748 272536
rect 329800 272524 329806 272536
rect 338850 272524 338856 272536
rect 329800 272496 338856 272524
rect 329800 272484 329806 272496
rect 338850 272484 338856 272496
rect 338908 272484 338914 272536
rect 339218 272484 339224 272536
rect 339276 272524 339282 272536
rect 354214 272524 354220 272536
rect 339276 272496 354220 272524
rect 339276 272484 339282 272496
rect 354214 272484 354220 272496
rect 354272 272484 354278 272536
rect 354490 272484 354496 272536
rect 354548 272524 354554 272536
rect 375558 272524 375564 272536
rect 354548 272496 375564 272524
rect 354548 272484 354554 272496
rect 375558 272484 375564 272496
rect 375616 272484 375622 272536
rect 379422 272484 379428 272536
rect 379480 272524 379486 272536
rect 410978 272524 410984 272536
rect 379480 272496 410984 272524
rect 379480 272484 379486 272496
rect 410978 272484 410984 272496
rect 411036 272484 411042 272536
rect 416590 272484 416596 272536
rect 416648 272524 416654 272536
rect 463878 272524 463884 272536
rect 416648 272496 463884 272524
rect 416648 272484 416654 272496
rect 463878 272484 463884 272496
rect 463936 272484 463942 272536
rect 466288 272524 466316 272564
rect 470548 272524 470554 272536
rect 466288 272496 470554 272524
rect 470548 272484 470554 272496
rect 470606 272484 470612 272536
rect 470686 272484 470692 272536
rect 470744 272524 470750 272536
rect 532694 272524 532700 272536
rect 470744 272496 532700 272524
rect 470744 272484 470750 272496
rect 532694 272484 532700 272496
rect 532752 272484 532758 272536
rect 532896 272524 532924 272632
rect 533706 272620 533712 272672
rect 533764 272660 533770 272672
rect 533764 272632 538444 272660
rect 533764 272620 533770 272632
rect 536374 272524 536380 272536
rect 532896 272496 536380 272524
rect 536374 272484 536380 272496
rect 536432 272484 536438 272536
rect 536558 272484 536564 272536
rect 536616 272524 536622 272536
rect 538122 272524 538128 272536
rect 536616 272496 538128 272524
rect 536616 272484 536622 272496
rect 538122 272484 538128 272496
rect 538180 272484 538186 272536
rect 538416 272524 538444 272632
rect 538674 272620 538680 272672
rect 538732 272660 538738 272672
rect 628466 272660 628472 272672
rect 538732 272632 628472 272660
rect 538732 272620 538738 272632
rect 628466 272620 628472 272632
rect 628524 272620 628530 272672
rect 634078 272620 634084 272672
rect 634136 272660 634142 272672
rect 640334 272660 640340 272672
rect 634136 272632 640340 272660
rect 634136 272620 634142 272632
rect 640334 272620 640340 272632
rect 640392 272620 640398 272672
rect 632054 272524 632060 272536
rect 538416 272496 632060 272524
rect 632054 272484 632060 272496
rect 632112 272484 632118 272536
rect 187694 272388 187700 272400
rect 180766 272360 187700 272388
rect 187694 272348 187700 272360
rect 187752 272348 187758 272400
rect 194962 272348 194968 272400
rect 195020 272388 195026 272400
rect 227162 272388 227168 272400
rect 195020 272360 227168 272388
rect 195020 272348 195026 272360
rect 227162 272348 227168 272360
rect 227220 272348 227226 272400
rect 318702 272348 318708 272400
rect 318760 272388 318766 272400
rect 324682 272388 324688 272400
rect 318760 272360 324688 272388
rect 318760 272348 318766 272360
rect 324682 272348 324688 272360
rect 324740 272348 324746 272400
rect 395982 272348 395988 272400
rect 396040 272388 396046 272400
rect 434622 272388 434628 272400
rect 396040 272360 434628 272388
rect 396040 272348 396046 272360
rect 434622 272348 434628 272360
rect 434680 272348 434686 272400
rect 446858 272348 446864 272400
rect 446916 272388 446922 272400
rect 500862 272388 500868 272400
rect 446916 272360 500868 272388
rect 446916 272348 446922 272360
rect 500862 272348 500868 272360
rect 500920 272348 500926 272400
rect 501046 272348 501052 272400
rect 501104 272388 501110 272400
rect 509694 272388 509700 272400
rect 501104 272360 509700 272388
rect 501104 272348 501110 272360
rect 509694 272348 509700 272360
rect 509752 272348 509758 272400
rect 517422 272348 517428 272400
rect 517480 272388 517486 272400
rect 600958 272388 600964 272400
rect 517480 272360 600964 272388
rect 517480 272348 517486 272360
rect 600958 272348 600964 272360
rect 601016 272348 601022 272400
rect 601142 272348 601148 272400
rect 601200 272388 601206 272400
rect 635550 272388 635556 272400
rect 601200 272360 635556 272388
rect 601200 272348 601206 272360
rect 635550 272348 635556 272360
rect 635608 272348 635614 272400
rect 269114 272280 269120 272332
rect 269172 272320 269178 272332
rect 270586 272320 270592 272332
rect 269172 272292 270592 272320
rect 269172 272280 269178 272292
rect 270586 272280 270592 272292
rect 270644 272280 270650 272332
rect 127342 272212 127348 272264
rect 127400 272252 127406 272264
rect 179874 272252 179880 272264
rect 127400 272224 179880 272252
rect 127400 272212 127406 272224
rect 179874 272212 179880 272224
rect 179932 272212 179938 272264
rect 189074 272212 189080 272264
rect 189132 272252 189138 272264
rect 196434 272252 196440 272264
rect 189132 272224 196440 272252
rect 189132 272212 189138 272224
rect 196434 272212 196440 272224
rect 196492 272212 196498 272264
rect 391842 272212 391848 272264
rect 391900 272252 391906 272264
rect 428734 272252 428740 272264
rect 391900 272224 428740 272252
rect 391900 272212 391906 272224
rect 428734 272212 428740 272224
rect 428792 272212 428798 272264
rect 449710 272212 449716 272264
rect 449768 272252 449774 272264
rect 504174 272252 504180 272264
rect 449768 272224 504180 272252
rect 449768 272212 449774 272224
rect 504174 272212 504180 272224
rect 504232 272212 504238 272264
rect 504542 272212 504548 272264
rect 504600 272252 504606 272264
rect 507946 272252 507952 272264
rect 504600 272224 507952 272252
rect 504600 272212 504606 272224
rect 507946 272212 507952 272224
rect 508004 272212 508010 272264
rect 509694 272212 509700 272264
rect 509752 272252 509758 272264
rect 514202 272252 514208 272264
rect 509752 272224 514208 272252
rect 509752 272212 509758 272224
rect 514202 272212 514208 272224
rect 514260 272212 514266 272264
rect 520090 272212 520096 272264
rect 520148 272252 520154 272264
rect 610710 272252 610716 272264
rect 520148 272224 610716 272252
rect 520148 272212 520154 272224
rect 610710 272212 610716 272224
rect 610768 272212 610774 272264
rect 147398 272076 147404 272128
rect 147456 272116 147462 272128
rect 193214 272116 193220 272128
rect 147456 272088 193220 272116
rect 147456 272076 147462 272088
rect 193214 272076 193220 272088
rect 193272 272076 193278 272128
rect 384942 272076 384948 272128
rect 385000 272116 385006 272128
rect 418062 272116 418068 272128
rect 385000 272088 418068 272116
rect 385000 272076 385006 272088
rect 418062 272076 418068 272088
rect 418120 272076 418126 272128
rect 428458 272076 428464 272128
rect 428516 272116 428522 272128
rect 470548 272116 470554 272128
rect 428516 272088 470554 272116
rect 428516 272076 428522 272088
rect 470548 272076 470554 272088
rect 470606 272076 470612 272128
rect 470778 272076 470784 272128
rect 470836 272116 470842 272128
rect 470836 272088 482600 272116
rect 470836 272076 470842 272088
rect 124950 271940 124956 271992
rect 125008 271980 125014 271992
rect 151078 271980 151084 271992
rect 125008 271952 151084 271980
rect 125008 271940 125014 271952
rect 151078 271940 151084 271952
rect 151136 271940 151142 271992
rect 431678 271940 431684 271992
rect 431736 271980 431742 271992
rect 482572 271980 482600 272088
rect 483014 272076 483020 272128
rect 483072 272116 483078 272128
rect 547506 272116 547512 272128
rect 483072 272088 547512 272116
rect 483072 272076 483078 272088
rect 547506 272076 547512 272088
rect 547564 272076 547570 272128
rect 547690 272076 547696 272128
rect 547748 272116 547754 272128
rect 562318 272116 562324 272128
rect 547748 272088 562324 272116
rect 547748 272076 547754 272088
rect 562318 272076 562324 272088
rect 562376 272076 562382 272128
rect 600958 272076 600964 272128
rect 601016 272116 601022 272128
rect 607214 272116 607220 272128
rect 601016 272088 607220 272116
rect 601016 272076 601022 272088
rect 607214 272076 607220 272088
rect 607272 272076 607278 272128
rect 504358 271980 504364 271992
rect 431736 271952 480484 271980
rect 482572 271952 504364 271980
rect 431736 271940 431742 271952
rect 105998 271804 106004 271856
rect 106056 271844 106062 271856
rect 164970 271844 164976 271856
rect 106056 271816 164976 271844
rect 106056 271804 106062 271816
rect 164970 271804 164976 271816
rect 165028 271804 165034 271856
rect 174262 271804 174268 271856
rect 174320 271844 174326 271856
rect 189166 271844 189172 271856
rect 174320 271816 189172 271844
rect 174320 271804 174326 271816
rect 189166 271804 189172 271816
rect 189224 271804 189230 271856
rect 202966 271804 202972 271856
rect 203024 271844 203030 271856
rect 233234 271844 233240 271856
rect 203024 271816 233240 271844
rect 203024 271804 203030 271816
rect 233234 271804 233240 271816
rect 233292 271804 233298 271856
rect 274634 271804 274640 271856
rect 274692 271844 274698 271856
rect 279234 271844 279240 271856
rect 274692 271816 279240 271844
rect 274692 271804 274698 271816
rect 279234 271804 279240 271816
rect 279292 271804 279298 271856
rect 355318 271804 355324 271856
rect 355376 271844 355382 271856
rect 356606 271844 356612 271856
rect 355376 271816 356612 271844
rect 355376 271804 355382 271816
rect 356606 271804 356612 271816
rect 356664 271804 356670 271856
rect 375282 271804 375288 271856
rect 375340 271844 375346 271856
rect 403894 271844 403900 271856
rect 375340 271816 403900 271844
rect 375340 271804 375346 271816
rect 403894 271804 403900 271816
rect 403952 271804 403958 271856
rect 433150 271804 433156 271856
rect 433208 271844 433214 271856
rect 480162 271844 480168 271856
rect 433208 271816 480168 271844
rect 433208 271804 433214 271816
rect 480162 271804 480168 271816
rect 480220 271804 480226 271856
rect 480456 271844 480484 271952
rect 504358 271940 504364 271952
rect 504416 271940 504422 271992
rect 504542 271940 504548 271992
rect 504600 271980 504606 271992
rect 561950 271980 561956 271992
rect 504600 271952 561956 271980
rect 504600 271940 504606 271952
rect 561950 271940 561956 271952
rect 562008 271940 562014 271992
rect 562134 271940 562140 271992
rect 562192 271980 562198 271992
rect 569402 271980 569408 271992
rect 562192 271952 569408 271980
rect 562192 271940 562198 271952
rect 569402 271940 569408 271952
rect 569460 271940 569466 271992
rect 484854 271844 484860 271856
rect 480456 271816 484860 271844
rect 484854 271804 484860 271816
rect 484912 271804 484918 271856
rect 494698 271804 494704 271856
rect 494756 271844 494762 271856
rect 501414 271844 501420 271856
rect 494756 271816 501420 271844
rect 494756 271804 494762 271816
rect 501414 271804 501420 271816
rect 501472 271804 501478 271856
rect 504358 271804 504364 271856
rect 504416 271844 504422 271856
rect 578510 271844 578516 271856
rect 504416 271816 578516 271844
rect 504416 271804 504422 271816
rect 578510 271804 578516 271816
rect 578568 271804 578574 271856
rect 578878 271804 578884 271856
rect 578936 271844 578942 271856
rect 604822 271844 604828 271856
rect 578936 271816 604828 271844
rect 578936 271804 578942 271816
rect 604822 271804 604828 271816
rect 604880 271804 604886 271856
rect 97810 271668 97816 271720
rect 97868 271708 97874 271720
rect 158806 271708 158812 271720
rect 97868 271680 158812 271708
rect 97868 271668 97874 271680
rect 158806 271668 158812 271680
rect 158864 271668 158870 271720
rect 169846 271668 169852 271720
rect 169904 271708 169910 271720
rect 209958 271708 209964 271720
rect 169904 271680 209964 271708
rect 169904 271668 169910 271680
rect 209958 271668 209964 271680
rect 210016 271668 210022 271720
rect 225414 271668 225420 271720
rect 225472 271708 225478 271720
rect 228358 271708 228364 271720
rect 225472 271680 228364 271708
rect 225472 271668 225478 271680
rect 228358 271668 228364 271680
rect 228416 271668 228422 271720
rect 351178 271668 351184 271720
rect 351236 271708 351242 271720
rect 366082 271708 366088 271720
rect 351236 271680 366088 271708
rect 351236 271668 351242 271680
rect 366082 271668 366088 271680
rect 366140 271668 366146 271720
rect 381998 271668 382004 271720
rect 382056 271708 382062 271720
rect 414566 271708 414572 271720
rect 382056 271680 414572 271708
rect 382056 271668 382062 271680
rect 414566 271668 414572 271680
rect 414624 271668 414630 271720
rect 421650 271708 421656 271720
rect 417160 271680 421656 271708
rect 87138 271532 87144 271584
rect 87196 271572 87202 271584
rect 151998 271572 152004 271584
rect 87196 271544 152004 271572
rect 87196 271532 87202 271544
rect 151998 271532 152004 271544
rect 152056 271532 152062 271584
rect 165154 271532 165160 271584
rect 165212 271572 165218 271584
rect 205634 271572 205640 271584
rect 165212 271544 205640 271572
rect 165212 271532 165218 271544
rect 205634 271532 205640 271544
rect 205692 271532 205698 271584
rect 215938 271532 215944 271584
rect 215996 271572 216002 271584
rect 242066 271572 242072 271584
rect 215996 271544 242072 271572
rect 215996 271532 216002 271544
rect 242066 271532 242072 271544
rect 242124 271532 242130 271584
rect 337930 271532 337936 271584
rect 337988 271572 337994 271584
rect 350718 271572 350724 271584
rect 337988 271544 350724 271572
rect 337988 271532 337994 271544
rect 350718 271532 350724 271544
rect 350776 271532 350782 271584
rect 360838 271532 360844 271584
rect 360896 271572 360902 271584
rect 377858 271572 377864 271584
rect 360896 271544 377864 271572
rect 360896 271532 360902 271544
rect 377858 271532 377864 271544
rect 377916 271532 377922 271584
rect 387702 271532 387708 271584
rect 387760 271572 387766 271584
rect 417160 271572 417188 271680
rect 421650 271668 421656 271680
rect 421708 271668 421714 271720
rect 430390 271668 430396 271720
rect 430448 271708 430454 271720
rect 483198 271708 483204 271720
rect 430448 271680 483204 271708
rect 430448 271668 430454 271680
rect 483198 271668 483204 271680
rect 483256 271668 483262 271720
rect 499298 271668 499304 271720
rect 499356 271708 499362 271720
rect 582374 271708 582380 271720
rect 499356 271680 582380 271708
rect 499356 271668 499362 271680
rect 582374 271668 582380 271680
rect 582432 271668 582438 271720
rect 583018 271668 583024 271720
rect 583076 271708 583082 271720
rect 611906 271708 611912 271720
rect 583076 271680 611912 271708
rect 583076 271668 583082 271680
rect 611906 271668 611912 271680
rect 611964 271668 611970 271720
rect 387760 271544 417188 271572
rect 387760 271532 387766 271544
rect 420178 271532 420184 271584
rect 420236 271572 420242 271584
rect 431126 271572 431132 271584
rect 420236 271544 431132 271572
rect 420236 271532 420242 271544
rect 431126 271532 431132 271544
rect 431184 271532 431190 271584
rect 437198 271532 437204 271584
rect 437256 271572 437262 271584
rect 493686 271572 493692 271584
rect 437256 271544 493692 271572
rect 437256 271532 437262 271544
rect 493686 271532 493692 271544
rect 493744 271532 493750 271584
rect 497274 271572 497280 271584
rect 493888 271544 497280 271572
rect 75362 271396 75368 271448
rect 75420 271436 75426 271448
rect 142706 271436 142712 271448
rect 75420 271408 142712 271436
rect 75420 271396 75426 271408
rect 142706 271396 142712 271408
rect 142764 271396 142770 271448
rect 162670 271396 162676 271448
rect 162728 271436 162734 271448
rect 204714 271436 204720 271448
rect 162728 271408 204720 271436
rect 162728 271396 162734 271408
rect 204714 271396 204720 271408
rect 204772 271396 204778 271448
rect 213638 271396 213644 271448
rect 213696 271436 213702 271448
rect 240410 271436 240416 271448
rect 213696 271408 240416 271436
rect 213696 271396 213702 271408
rect 240410 271396 240416 271408
rect 240468 271396 240474 271448
rect 240778 271396 240784 271448
rect 240836 271436 240842 271448
rect 259638 271436 259644 271448
rect 240836 271408 259644 271436
rect 240836 271396 240842 271408
rect 259638 271396 259644 271408
rect 259696 271396 259702 271448
rect 259822 271396 259828 271448
rect 259880 271436 259886 271448
rect 272610 271436 272616 271448
rect 259880 271408 272616 271436
rect 259880 271396 259886 271408
rect 272610 271396 272616 271408
rect 272668 271396 272674 271448
rect 325510 271396 325516 271448
rect 325568 271436 325574 271448
rect 334158 271436 334164 271448
rect 325568 271408 334164 271436
rect 325568 271396 325574 271408
rect 334158 271396 334164 271408
rect 334216 271396 334222 271448
rect 347682 271396 347688 271448
rect 347740 271436 347746 271448
rect 364886 271436 364892 271448
rect 347740 271408 364892 271436
rect 347740 271396 347746 271408
rect 364886 271396 364892 271408
rect 364944 271396 364950 271448
rect 366358 271396 366364 271448
rect 366416 271436 366422 271448
rect 383838 271436 383844 271448
rect 366416 271408 383844 271436
rect 366416 271396 366422 271408
rect 383838 271396 383844 271408
rect 383896 271396 383902 271448
rect 384758 271396 384764 271448
rect 384816 271436 384822 271448
rect 419258 271436 419264 271448
rect 384816 271408 419264 271436
rect 384816 271396 384822 271408
rect 419258 271396 419264 271408
rect 419316 271396 419322 271448
rect 426342 271436 426348 271448
rect 424336 271408 426348 271436
rect 76834 271260 76840 271312
rect 76892 271300 76898 271312
rect 143534 271300 143540 271312
rect 76892 271272 143540 271300
rect 76892 271260 76898 271272
rect 143534 271260 143540 271272
rect 143592 271260 143598 271312
rect 152182 271260 152188 271312
rect 152240 271300 152246 271312
rect 197354 271300 197360 271312
rect 152240 271272 197360 271300
rect 152240 271260 152246 271272
rect 197354 271260 197360 271272
rect 197412 271260 197418 271312
rect 198274 271260 198280 271312
rect 198332 271300 198338 271312
rect 229554 271300 229560 271312
rect 198332 271272 229560 271300
rect 198332 271260 198338 271272
rect 229554 271260 229560 271272
rect 229612 271260 229618 271312
rect 235258 271260 235264 271312
rect 235316 271300 235322 271312
rect 255314 271300 255320 271312
rect 235316 271272 255320 271300
rect 235316 271260 235322 271272
rect 255314 271260 255320 271272
rect 255372 271260 255378 271312
rect 256694 271260 256700 271312
rect 256752 271300 256758 271312
rect 261018 271300 261024 271312
rect 256752 271272 261024 271300
rect 256752 271260 256758 271272
rect 261018 271260 261024 271272
rect 261076 271260 261082 271312
rect 262030 271260 262036 271312
rect 262088 271300 262094 271312
rect 274634 271300 274640 271312
rect 262088 271272 274640 271300
rect 262088 271260 262094 271272
rect 274634 271260 274640 271272
rect 274692 271260 274698 271312
rect 329558 271260 329564 271312
rect 329616 271300 329622 271312
rect 340046 271300 340052 271312
rect 329616 271272 340052 271300
rect 329616 271260 329622 271272
rect 340046 271260 340052 271272
rect 340104 271260 340110 271312
rect 340598 271260 340604 271312
rect 340656 271300 340662 271312
rect 355134 271300 355140 271312
rect 340656 271272 355140 271300
rect 340656 271260 340662 271272
rect 355134 271260 355140 271272
rect 355192 271260 355198 271312
rect 357158 271260 357164 271312
rect 357216 271300 357222 271312
rect 379054 271300 379060 271312
rect 357216 271272 379060 271300
rect 357216 271260 357222 271272
rect 379054 271260 379060 271272
rect 379112 271260 379118 271312
rect 390278 271260 390284 271312
rect 390336 271300 390342 271312
rect 424336 271300 424364 271408
rect 426342 271396 426348 271408
rect 426400 271396 426406 271448
rect 439958 271396 439964 271448
rect 440016 271436 440022 271448
rect 493888 271436 493916 271544
rect 497274 271532 497280 271544
rect 497332 271532 497338 271584
rect 501966 271532 501972 271584
rect 502024 271572 502030 271584
rect 585962 271572 585968 271584
rect 502024 271544 585968 271572
rect 502024 271532 502030 271544
rect 585962 271532 585968 271544
rect 586020 271532 586026 271584
rect 611998 271532 612004 271584
rect 612056 271572 612062 271584
rect 618990 271572 618996 271584
rect 612056 271544 618996 271572
rect 612056 271532 612062 271544
rect 618990 271532 618996 271544
rect 619048 271532 619054 271584
rect 440016 271408 493916 271436
rect 440016 271396 440022 271408
rect 496538 271396 496544 271448
rect 496596 271436 496602 271448
rect 504358 271436 504364 271448
rect 496596 271408 504364 271436
rect 496596 271396 496602 271408
rect 504358 271396 504364 271408
rect 504416 271396 504422 271448
rect 505002 271396 505008 271448
rect 505060 271436 505066 271448
rect 589458 271436 589464 271448
rect 505060 271408 589464 271436
rect 505060 271396 505066 271408
rect 589458 271396 589464 271408
rect 589516 271396 589522 271448
rect 589918 271396 589924 271448
rect 589976 271436 589982 271448
rect 633250 271436 633256 271448
rect 589976 271408 633256 271436
rect 589976 271396 589982 271408
rect 633250 271396 633256 271408
rect 633308 271396 633314 271448
rect 432230 271300 432236 271312
rect 390336 271272 424364 271300
rect 425992 271272 432236 271300
rect 390336 271260 390342 271272
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 138474 271164 138480 271176
rect 68244 271136 138480 271164
rect 68244 271124 68250 271136
rect 138474 271124 138480 271136
rect 138532 271124 138538 271176
rect 141510 271124 141516 271176
rect 141568 271164 141574 271176
rect 189810 271164 189816 271176
rect 141568 271136 189816 271164
rect 141568 271124 141574 271136
rect 189810 271124 189816 271136
rect 189868 271124 189874 271176
rect 191190 271124 191196 271176
rect 191248 271164 191254 271176
rect 225138 271164 225144 271176
rect 191248 271136 225144 271164
rect 191248 271124 191254 271136
rect 225138 271124 225144 271136
rect 225196 271124 225202 271176
rect 230198 271124 230204 271176
rect 230256 271164 230262 271176
rect 252002 271164 252008 271176
rect 230256 271136 252008 271164
rect 230256 271124 230262 271136
rect 252002 271124 252008 271136
rect 252060 271124 252066 271176
rect 268010 271124 268016 271176
rect 268068 271164 268074 271176
rect 278774 271164 278780 271176
rect 268068 271136 278780 271164
rect 268068 271124 268074 271136
rect 278774 271124 278780 271136
rect 278832 271124 278838 271176
rect 279786 271124 279792 271176
rect 279844 271164 279850 271176
rect 287054 271164 287060 271176
rect 279844 271136 287060 271164
rect 279844 271124 279850 271136
rect 287054 271124 287060 271136
rect 287112 271124 287118 271176
rect 331122 271124 331128 271176
rect 331180 271164 331186 271176
rect 342438 271164 342444 271176
rect 331180 271136 342444 271164
rect 331180 271124 331186 271136
rect 342438 271124 342444 271136
rect 342496 271124 342502 271176
rect 343542 271124 343548 271176
rect 343600 271164 343606 271176
rect 360194 271164 360200 271176
rect 343600 271136 360200 271164
rect 343600 271124 343606 271136
rect 360194 271124 360200 271136
rect 360252 271124 360258 271176
rect 364150 271124 364156 271176
rect 364208 271164 364214 271176
rect 389726 271164 389732 271176
rect 364208 271136 389732 271164
rect 364208 271124 364214 271136
rect 389726 271124 389732 271136
rect 389784 271124 389790 271176
rect 394326 271124 394332 271176
rect 394384 271164 394390 271176
rect 425992 271164 426020 271272
rect 432230 271260 432236 271272
rect 432288 271260 432294 271312
rect 442902 271260 442908 271312
rect 442960 271300 442966 271312
rect 500678 271300 500684 271312
rect 442960 271272 500684 271300
rect 442960 271260 442966 271272
rect 500678 271260 500684 271272
rect 500736 271260 500742 271312
rect 507670 271260 507676 271312
rect 507728 271300 507734 271312
rect 593046 271300 593052 271312
rect 507728 271272 593052 271300
rect 507728 271260 507734 271272
rect 593046 271260 593052 271272
rect 593104 271260 593110 271312
rect 598198 271260 598204 271312
rect 598256 271300 598262 271312
rect 645026 271300 645032 271312
rect 598256 271272 645032 271300
rect 598256 271260 598262 271272
rect 645026 271260 645032 271272
rect 645084 271260 645090 271312
rect 437934 271164 437940 271176
rect 394384 271136 426020 271164
rect 427096 271136 437940 271164
rect 394384 271124 394390 271136
rect 113450 270988 113456 271040
rect 113508 271028 113514 271040
rect 169938 271028 169944 271040
rect 113508 271000 169944 271028
rect 113508 270988 113514 271000
rect 169938 270988 169944 271000
rect 169996 270988 170002 271040
rect 187418 270988 187424 271040
rect 187476 271028 187482 271040
rect 215938 271028 215944 271040
rect 187476 271000 215944 271028
rect 187476 270988 187482 271000
rect 215938 270988 215944 271000
rect 215996 270988 216002 271040
rect 251450 270988 251456 271040
rect 251508 271028 251514 271040
rect 266906 271028 266912 271040
rect 251508 271000 266912 271028
rect 251508 270988 251514 271000
rect 266906 270988 266912 271000
rect 266964 270988 266970 271040
rect 417418 270988 417424 271040
rect 417476 271028 417482 271040
rect 427096 271028 427124 271136
rect 437934 271124 437940 271136
rect 437992 271124 437998 271176
rect 441338 271124 441344 271176
rect 441396 271164 441402 271176
rect 445018 271164 445024 271176
rect 441396 271136 445024 271164
rect 441396 271124 441402 271136
rect 445018 271124 445024 271136
rect 445076 271124 445082 271176
rect 445662 271124 445668 271176
rect 445720 271164 445726 271176
rect 503990 271164 503996 271176
rect 445720 271136 503996 271164
rect 445720 271124 445726 271136
rect 503990 271124 503996 271136
rect 504048 271124 504054 271176
rect 524046 271124 524052 271176
rect 524104 271164 524110 271176
rect 617334 271164 617340 271176
rect 524104 271136 617340 271164
rect 524104 271124 524110 271136
rect 617334 271124 617340 271136
rect 617392 271124 617398 271176
rect 617518 271124 617524 271176
rect 617576 271164 617582 271176
rect 626074 271164 626080 271176
rect 617576 271136 626080 271164
rect 617576 271124 617582 271136
rect 626074 271124 626080 271136
rect 626132 271124 626138 271176
rect 417476 271000 427124 271028
rect 417476 270988 417482 271000
rect 427446 270988 427452 271040
rect 427504 271028 427510 271040
rect 479150 271028 479156 271040
rect 427504 271000 479156 271028
rect 427504 270988 427510 271000
rect 479150 270988 479156 271000
rect 479208 270988 479214 271040
rect 485038 270988 485044 271040
rect 485096 271028 485102 271040
rect 494698 271028 494704 271040
rect 485096 271000 494704 271028
rect 485096 270988 485102 271000
rect 494698 270988 494704 271000
rect 494756 270988 494762 271040
rect 495066 270988 495072 271040
rect 495124 271028 495130 271040
rect 575290 271028 575296 271040
rect 495124 271000 575296 271028
rect 495124 270988 495130 271000
rect 575290 270988 575296 271000
rect 575348 270988 575354 271040
rect 123754 270852 123760 270904
rect 123812 270892 123818 270904
rect 177482 270892 177488 270904
rect 123812 270864 177488 270892
rect 123812 270852 123818 270864
rect 177482 270852 177488 270864
rect 177540 270852 177546 270904
rect 407758 270852 407764 270904
rect 407816 270892 407822 270904
rect 440510 270892 440516 270904
rect 407816 270864 440516 270892
rect 407816 270852 407822 270864
rect 440510 270852 440516 270864
rect 440568 270852 440574 270904
rect 449158 270852 449164 270904
rect 449216 270892 449222 270904
rect 490190 270892 490196 270904
rect 449216 270864 490196 270892
rect 449216 270852 449222 270864
rect 490190 270852 490196 270864
rect 490248 270852 490254 270904
rect 492582 270852 492588 270904
rect 492640 270892 492646 270904
rect 571702 270892 571708 270904
rect 492640 270864 571708 270892
rect 492640 270852 492646 270864
rect 571702 270852 571708 270864
rect 571760 270852 571766 270904
rect 134426 270716 134432 270768
rect 134484 270756 134490 270768
rect 185118 270756 185124 270768
rect 134484 270728 185124 270756
rect 134484 270716 134490 270728
rect 185118 270716 185124 270728
rect 185176 270716 185182 270768
rect 321370 270716 321376 270768
rect 321428 270756 321434 270768
rect 327074 270756 327080 270768
rect 321428 270728 327080 270756
rect 321428 270716 321434 270728
rect 327074 270716 327080 270728
rect 327132 270716 327138 270768
rect 414658 270716 414664 270768
rect 414716 270756 414722 270768
rect 450814 270756 450820 270768
rect 414716 270728 450820 270756
rect 414716 270716 414722 270728
rect 450814 270716 450820 270728
rect 450872 270716 450878 270768
rect 480254 270716 480260 270768
rect 480312 270756 480318 270768
rect 486602 270756 486608 270768
rect 480312 270728 486608 270756
rect 480312 270716 480318 270728
rect 486602 270716 486608 270728
rect 486660 270716 486666 270768
rect 486970 270716 486976 270768
rect 487028 270756 487034 270768
rect 564618 270756 564624 270768
rect 487028 270728 564624 270756
rect 487028 270716 487034 270728
rect 564618 270716 564624 270728
rect 564676 270716 564682 270768
rect 567838 270716 567844 270768
rect 567896 270756 567902 270768
rect 597738 270756 597744 270768
rect 567896 270728 597744 270756
rect 567896 270716 567902 270728
rect 597738 270716 597744 270728
rect 597796 270716 597802 270768
rect 121454 270580 121460 270632
rect 121512 270620 121518 270632
rect 168098 270620 168104 270632
rect 121512 270592 168104 270620
rect 121512 270580 121518 270592
rect 168098 270580 168104 270592
rect 168156 270580 168162 270632
rect 403618 270580 403624 270632
rect 403676 270620 403682 270632
rect 433426 270620 433432 270632
rect 403676 270592 433432 270620
rect 403676 270580 403682 270592
rect 433426 270580 433432 270592
rect 433484 270580 433490 270632
rect 453298 270580 453304 270632
rect 453356 270620 453362 270632
rect 487798 270620 487804 270632
rect 453356 270592 487804 270620
rect 453356 270580 453362 270592
rect 487798 270580 487804 270592
rect 487856 270580 487862 270632
rect 489638 270580 489644 270632
rect 489696 270620 489702 270632
rect 568206 270620 568212 270632
rect 489696 270592 568212 270620
rect 489696 270580 489702 270592
rect 568206 270580 568212 270592
rect 568264 270580 568270 270632
rect 78858 270444 78864 270496
rect 78916 270484 78922 270496
rect 132494 270484 132500 270496
rect 78916 270456 132500 270484
rect 78916 270444 78922 270456
rect 132494 270444 132500 270456
rect 132552 270444 132558 270496
rect 133782 270444 133788 270496
rect 133840 270484 133846 270496
rect 136634 270484 136640 270496
rect 133840 270456 136640 270484
rect 133840 270444 133846 270456
rect 136634 270444 136640 270456
rect 136692 270444 136698 270496
rect 137002 270444 137008 270496
rect 137060 270484 137066 270496
rect 137060 270456 137692 270484
rect 137060 270444 137066 270456
rect 84102 270308 84108 270360
rect 84160 270348 84166 270360
rect 137462 270348 137468 270360
rect 84160 270320 137468 270348
rect 84160 270308 84166 270320
rect 137462 270308 137468 270320
rect 137520 270308 137526 270360
rect 137664 270348 137692 270456
rect 137830 270444 137836 270496
rect 137888 270484 137894 270496
rect 183646 270484 183652 270496
rect 137888 270456 183652 270484
rect 137888 270444 137894 270456
rect 183646 270444 183652 270456
rect 183704 270444 183710 270496
rect 185578 270444 185584 270496
rect 185636 270484 185642 270496
rect 194410 270484 194416 270496
rect 185636 270456 194416 270484
rect 185636 270444 185642 270456
rect 194410 270444 194416 270456
rect 194468 270444 194474 270496
rect 200758 270444 200764 270496
rect 200816 270484 200822 270496
rect 201862 270484 201868 270496
rect 200816 270456 201868 270484
rect 200816 270444 200822 270456
rect 201862 270444 201868 270456
rect 201920 270444 201926 270496
rect 206830 270444 206836 270496
rect 206888 270484 206894 270496
rect 235810 270484 235816 270496
rect 206888 270456 235816 270484
rect 206888 270444 206894 270456
rect 235810 270444 235816 270456
rect 235868 270444 235874 270496
rect 278038 270444 278044 270496
rect 278096 270484 278102 270496
rect 283834 270484 283840 270496
rect 278096 270456 283840 270484
rect 278096 270444 278102 270456
rect 283834 270444 283840 270456
rect 283892 270444 283898 270496
rect 400858 270444 400864 270496
rect 400916 270484 400922 270496
rect 441614 270484 441620 270496
rect 400916 270456 441620 270484
rect 400916 270444 400922 270456
rect 441614 270444 441620 270456
rect 441672 270444 441678 270496
rect 456426 270444 456432 270496
rect 456484 270484 456490 270496
rect 520274 270484 520280 270496
rect 456484 270456 520280 270484
rect 456484 270444 456490 270456
rect 520274 270444 520280 270456
rect 520332 270444 520338 270496
rect 523126 270444 523132 270496
rect 523184 270484 523190 270496
rect 532878 270484 532884 270496
rect 523184 270456 532884 270484
rect 523184 270444 523190 270456
rect 532878 270444 532884 270456
rect 532936 270444 532942 270496
rect 619634 270484 619640 270496
rect 533356 270456 619640 270484
rect 186130 270348 186136 270360
rect 137664 270320 186136 270348
rect 186130 270308 186136 270320
rect 186188 270308 186194 270360
rect 199930 270308 199936 270360
rect 199988 270348 199994 270360
rect 230842 270348 230848 270360
rect 199988 270320 230848 270348
rect 199988 270308 199994 270320
rect 230842 270308 230848 270320
rect 230900 270308 230906 270360
rect 232682 270308 232688 270360
rect 232740 270348 232746 270360
rect 248230 270348 248236 270360
rect 232740 270320 248236 270348
rect 232740 270308 232746 270320
rect 248230 270308 248236 270320
rect 248288 270308 248294 270360
rect 283098 270308 283104 270360
rect 283156 270348 283162 270360
rect 284662 270348 284668 270360
rect 283156 270320 284668 270348
rect 283156 270308 283162 270320
rect 284662 270308 284668 270320
rect 284720 270308 284726 270360
rect 355042 270308 355048 270360
rect 355100 270348 355106 270360
rect 376938 270348 376944 270360
rect 355100 270320 376944 270348
rect 355100 270308 355106 270320
rect 376938 270308 376944 270320
rect 376996 270308 377002 270360
rect 380526 270308 380532 270360
rect 380584 270348 380590 270360
rect 404354 270348 404360 270360
rect 380584 270320 404360 270348
rect 380584 270308 380590 270320
rect 404354 270308 404360 270320
rect 404412 270308 404418 270360
rect 409598 270308 409604 270360
rect 409656 270348 409662 270360
rect 454310 270348 454316 270360
rect 409656 270320 454316 270348
rect 409656 270308 409662 270320
rect 454310 270308 454316 270320
rect 454368 270308 454374 270360
rect 458818 270308 458824 270360
rect 458876 270348 458882 270360
rect 524414 270348 524420 270360
rect 458876 270320 524420 270348
rect 458876 270308 458882 270320
rect 524414 270308 524420 270320
rect 524472 270308 524478 270360
rect 525610 270308 525616 270360
rect 525668 270348 525674 270360
rect 533356 270348 533384 270456
rect 619634 270444 619640 270456
rect 619692 270444 619698 270496
rect 525668 270320 533384 270348
rect 525668 270308 525674 270320
rect 533522 270308 533528 270360
rect 533580 270348 533586 270360
rect 626534 270348 626540 270360
rect 533580 270320 626540 270348
rect 533580 270308 533586 270320
rect 626534 270308 626540 270320
rect 626592 270308 626598 270360
rect 111978 270172 111984 270224
rect 112036 270212 112042 270224
rect 168742 270212 168748 270224
rect 112036 270184 168748 270212
rect 112036 270172 112042 270184
rect 168742 270172 168748 270184
rect 168800 270172 168806 270224
rect 184842 270172 184848 270224
rect 184900 270212 184906 270224
rect 219342 270212 219348 270224
rect 184900 270184 219348 270212
rect 184900 270172 184906 270184
rect 219342 270172 219348 270184
rect 219400 270172 219406 270224
rect 244366 270172 244372 270224
rect 244424 270212 244430 270224
rect 262306 270212 262312 270224
rect 244424 270184 262312 270212
rect 244424 270172 244430 270184
rect 262306 270172 262312 270184
rect 262364 270172 262370 270224
rect 334342 270172 334348 270224
rect 334400 270212 334406 270224
rect 346394 270212 346400 270224
rect 334400 270184 346400 270212
rect 334400 270172 334406 270184
rect 346394 270172 346400 270184
rect 346452 270172 346458 270224
rect 372246 270172 372252 270224
rect 372304 270212 372310 270224
rect 397454 270212 397460 270224
rect 372304 270184 397460 270212
rect 372304 270172 372310 270184
rect 397454 270172 397460 270184
rect 397512 270172 397518 270224
rect 398742 270172 398748 270224
rect 398800 270212 398806 270224
rect 412634 270212 412640 270224
rect 398800 270184 412640 270212
rect 398800 270172 398806 270184
rect 412634 270172 412640 270184
rect 412692 270172 412698 270224
rect 415026 270172 415032 270224
rect 415084 270212 415090 270224
rect 460934 270212 460940 270224
rect 415084 270184 460940 270212
rect 415084 270172 415090 270184
rect 460934 270172 460940 270184
rect 460992 270172 460998 270224
rect 461394 270172 461400 270224
rect 461452 270212 461458 270224
rect 527174 270212 527180 270224
rect 461452 270184 527180 270212
rect 461452 270172 461458 270184
rect 527174 270172 527180 270184
rect 527232 270172 527238 270224
rect 528370 270172 528376 270224
rect 528428 270212 528434 270224
rect 623958 270212 623964 270224
rect 528428 270184 623964 270212
rect 528428 270172 528434 270184
rect 623958 270172 623964 270184
rect 624016 270172 624022 270224
rect 89622 270036 89628 270088
rect 89680 270076 89686 270088
rect 153010 270076 153016 270088
rect 89680 270048 153016 270076
rect 89680 270036 89686 270048
rect 153010 270036 153016 270048
rect 153068 270036 153074 270088
rect 176562 270036 176568 270088
rect 176620 270076 176626 270088
rect 211154 270076 211160 270088
rect 176620 270048 211160 270076
rect 176620 270036 176626 270048
rect 211154 270036 211160 270048
rect 211212 270036 211218 270088
rect 212442 270036 212448 270088
rect 212500 270076 212506 270088
rect 239950 270076 239956 270088
rect 212500 270048 239956 270076
rect 212500 270036 212506 270048
rect 239950 270036 239956 270048
rect 240008 270036 240014 270088
rect 241882 270036 241888 270088
rect 241940 270076 241946 270088
rect 260650 270076 260656 270088
rect 241940 270048 260656 270076
rect 241940 270036 241946 270048
rect 260650 270036 260656 270048
rect 260708 270036 260714 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 277210 270076 277216 270088
rect 266228 270048 277216 270076
rect 266228 270036 266234 270048
rect 277210 270036 277216 270048
rect 277268 270036 277274 270088
rect 345290 270036 345296 270088
rect 345348 270076 345354 270088
rect 358814 270076 358820 270088
rect 345348 270048 358820 270076
rect 345348 270036 345354 270048
rect 358814 270036 358820 270048
rect 358872 270036 358878 270088
rect 366634 270036 366640 270088
rect 366692 270076 366698 270088
rect 393314 270076 393320 270088
rect 366692 270048 393320 270076
rect 366692 270036 366698 270048
rect 393314 270036 393320 270048
rect 393372 270036 393378 270088
rect 394970 270036 394976 270088
rect 395028 270076 395034 270088
rect 408770 270076 408776 270088
rect 395028 270048 408776 270076
rect 395028 270036 395034 270048
rect 408770 270036 408776 270048
rect 408828 270036 408834 270088
rect 412450 270036 412456 270088
rect 412508 270076 412514 270088
rect 458266 270076 458272 270088
rect 412508 270048 458272 270076
rect 412508 270036 412514 270048
rect 458266 270036 458272 270048
rect 458324 270036 458330 270088
rect 463510 270036 463516 270088
rect 463568 270076 463574 270088
rect 530762 270076 530768 270088
rect 463568 270048 530768 270076
rect 463568 270036 463574 270048
rect 530762 270036 530768 270048
rect 530820 270036 530826 270088
rect 530946 270036 530952 270088
rect 531004 270076 531010 270088
rect 533154 270076 533160 270088
rect 531004 270048 533160 270076
rect 531004 270036 531010 270048
rect 533154 270036 533160 270048
rect 533212 270036 533218 270088
rect 538122 270076 538128 270088
rect 533356 270048 538128 270076
rect 85482 269900 85488 269952
rect 85540 269940 85546 269952
rect 149422 269940 149428 269952
rect 85540 269912 149428 269940
rect 85540 269900 85546 269912
rect 149422 269900 149428 269912
rect 149480 269900 149486 269952
rect 152826 269900 152832 269952
rect 152884 269940 152890 269952
rect 157150 269940 157156 269952
rect 152884 269912 157156 269940
rect 152884 269900 152890 269912
rect 157150 269900 157156 269912
rect 157208 269900 157214 269952
rect 173710 269900 173716 269952
rect 173768 269940 173774 269952
rect 212626 269940 212632 269952
rect 173768 269912 212632 269940
rect 173768 269900 173774 269912
rect 212626 269900 212632 269912
rect 212684 269900 212690 269952
rect 226610 269900 226616 269952
rect 226668 269940 226674 269952
rect 249886 269940 249892 269952
rect 226668 269912 249892 269940
rect 226668 269900 226674 269912
rect 249886 269900 249892 269912
rect 249944 269900 249950 269952
rect 256878 269900 256884 269952
rect 256936 269940 256942 269952
rect 268930 269940 268936 269952
rect 256936 269912 268936 269940
rect 256936 269900 256942 269912
rect 268930 269900 268936 269912
rect 268988 269900 268994 269952
rect 330202 269900 330208 269952
rect 330260 269940 330266 269952
rect 340874 269940 340880 269952
rect 330260 269912 340880 269940
rect 330260 269900 330266 269912
rect 340874 269900 340880 269912
rect 340932 269900 340938 269952
rect 341794 269900 341800 269952
rect 341852 269940 341858 269952
rect 357526 269940 357532 269952
rect 341852 269912 357532 269940
rect 341852 269900 341858 269912
rect 357526 269900 357532 269912
rect 357584 269900 357590 269952
rect 359182 269900 359188 269952
rect 359240 269940 359246 269952
rect 382274 269940 382280 269952
rect 359240 269912 382280 269940
rect 359240 269900 359246 269912
rect 382274 269900 382280 269912
rect 382332 269900 382338 269952
rect 383010 269900 383016 269952
rect 383068 269940 383074 269952
rect 411254 269940 411260 269952
rect 383068 269912 411260 269940
rect 383068 269900 383074 269912
rect 411254 269900 411260 269912
rect 411312 269900 411318 269952
rect 419626 269900 419632 269952
rect 419684 269940 419690 269952
rect 468110 269940 468116 269952
rect 419684 269912 468116 269940
rect 419684 269900 419690 269912
rect 468110 269900 468116 269912
rect 468168 269900 468174 269952
rect 468478 269900 468484 269952
rect 468536 269940 468542 269952
rect 533356 269940 533384 270048
rect 538122 270036 538128 270048
rect 538180 270036 538186 270088
rect 538306 270036 538312 270088
rect 538364 270076 538370 270088
rect 630674 270076 630680 270088
rect 538364 270048 630680 270076
rect 538364 270036 538370 270048
rect 630674 270036 630680 270048
rect 630732 270036 630738 270088
rect 468536 269912 533384 269940
rect 468536 269900 468542 269912
rect 533982 269900 533988 269952
rect 534040 269940 534046 269952
rect 537846 269940 537852 269952
rect 534040 269912 537852 269940
rect 534040 269900 534046 269912
rect 537846 269900 537852 269912
rect 537904 269900 537910 269952
rect 538030 269900 538036 269952
rect 538088 269940 538094 269952
rect 538088 269912 543044 269940
rect 538088 269900 538094 269912
rect 70578 269764 70584 269816
rect 70636 269804 70642 269816
rect 79318 269804 79324 269816
rect 70636 269776 79324 269804
rect 70636 269764 70642 269776
rect 79318 269764 79324 269776
rect 79376 269764 79382 269816
rect 80054 269764 80060 269816
rect 80112 269804 80118 269816
rect 146386 269804 146392 269816
rect 80112 269776 146392 269804
rect 80112 269764 80118 269776
rect 146386 269764 146392 269776
rect 146444 269764 146450 269816
rect 158622 269764 158628 269816
rect 158680 269804 158686 269816
rect 201034 269804 201040 269816
rect 158680 269776 201040 269804
rect 158680 269764 158686 269776
rect 201034 269764 201040 269776
rect 201092 269764 201098 269816
rect 201678 269764 201684 269816
rect 201736 269804 201742 269816
rect 232498 269804 232504 269816
rect 201736 269776 232504 269804
rect 201736 269764 201742 269776
rect 232498 269764 232504 269776
rect 232556 269764 232562 269816
rect 237190 269764 237196 269816
rect 237248 269804 237254 269816
rect 257338 269804 257344 269816
rect 237248 269776 257344 269804
rect 237248 269764 237254 269776
rect 257338 269764 257344 269776
rect 257396 269764 257402 269816
rect 258534 269764 258540 269816
rect 258592 269804 258598 269816
rect 272242 269804 272248 269816
rect 258592 269776 272248 269804
rect 258592 269764 258598 269776
rect 272242 269764 272248 269776
rect 272300 269764 272306 269816
rect 273070 269764 273076 269816
rect 273128 269804 273134 269816
rect 282178 269804 282184 269816
rect 273128 269776 282184 269804
rect 273128 269764 273134 269776
rect 282178 269764 282184 269776
rect 282236 269764 282242 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335538 269804 335544 269816
rect 326948 269776 335544 269804
rect 326948 269764 326954 269776
rect 335538 269764 335544 269776
rect 335596 269764 335602 269816
rect 335998 269764 336004 269816
rect 336056 269804 336062 269816
rect 349154 269804 349160 269816
rect 336056 269776 349160 269804
rect 336056 269764 336062 269776
rect 349154 269764 349160 269776
rect 349212 269764 349218 269816
rect 351730 269764 351736 269816
rect 351788 269804 351794 269816
rect 371234 269804 371240 269816
rect 351788 269776 371240 269804
rect 351788 269764 351794 269776
rect 371234 269764 371240 269776
rect 371292 269764 371298 269816
rect 376570 269764 376576 269816
rect 376628 269804 376634 269816
rect 407114 269804 407120 269816
rect 376628 269776 407120 269804
rect 376628 269764 376634 269776
rect 407114 269764 407120 269776
rect 407172 269764 407178 269816
rect 417142 269764 417148 269816
rect 417200 269804 417206 269816
rect 465074 269804 465080 269816
rect 417200 269776 465080 269804
rect 417200 269764 417206 269776
rect 465074 269764 465080 269776
rect 465132 269764 465138 269816
rect 465994 269764 466000 269816
rect 466052 269804 466058 269816
rect 530394 269804 530400 269816
rect 466052 269776 530400 269804
rect 466052 269764 466058 269776
rect 530394 269764 530400 269776
rect 530452 269764 530458 269816
rect 538582 269804 538588 269816
rect 530596 269776 538588 269804
rect 122742 269628 122748 269680
rect 122800 269668 122806 269680
rect 176194 269668 176200 269680
rect 122800 269640 176200 269668
rect 122800 269628 122806 269640
rect 176194 269628 176200 269640
rect 176252 269628 176258 269680
rect 183462 269628 183468 269680
rect 183520 269668 183526 269680
rect 205450 269668 205456 269680
rect 183520 269640 205456 269668
rect 183520 269628 183526 269640
rect 205450 269628 205456 269640
rect 205508 269628 205514 269680
rect 392026 269628 392032 269680
rect 392084 269668 392090 269680
rect 401686 269668 401692 269680
rect 392084 269640 401692 269668
rect 392084 269628 392090 269640
rect 401686 269628 401692 269640
rect 401744 269628 401750 269680
rect 404354 269628 404360 269680
rect 404412 269668 404418 269680
rect 423674 269668 423680 269680
rect 404412 269640 423680 269668
rect 404412 269628 404418 269640
rect 423674 269628 423680 269640
rect 423732 269628 423738 269680
rect 423950 269628 423956 269680
rect 424008 269668 424014 269680
rect 451366 269668 451372 269680
rect 424008 269640 451372 269668
rect 424008 269628 424014 269640
rect 451366 269628 451372 269640
rect 451424 269628 451430 269680
rect 453574 269628 453580 269680
rect 453632 269668 453638 269680
rect 509234 269668 509240 269680
rect 453632 269640 509240 269668
rect 453632 269628 453638 269640
rect 509234 269628 509240 269640
rect 509292 269628 509298 269680
rect 530596 269668 530624 269776
rect 538582 269764 538588 269776
rect 538640 269764 538646 269816
rect 538766 269764 538772 269816
rect 538824 269804 538830 269816
rect 542814 269804 542820 269816
rect 538824 269776 542820 269804
rect 538824 269764 538830 269776
rect 542814 269764 542820 269776
rect 542872 269764 542878 269816
rect 543016 269804 543044 269912
rect 543182 269900 543188 269952
rect 543240 269940 543246 269952
rect 640518 269940 640524 269952
rect 543240 269912 640524 269940
rect 543240 269900 543246 269912
rect 640518 269900 640524 269912
rect 640576 269900 640582 269952
rect 637574 269804 637580 269816
rect 543016 269776 637580 269804
rect 637574 269764 637580 269776
rect 637632 269764 637638 269816
rect 509712 269640 530624 269668
rect 129642 269492 129648 269544
rect 129700 269532 129706 269544
rect 181162 269532 181168 269544
rect 129700 269504 181168 269532
rect 129700 269492 129706 269504
rect 181162 269492 181168 269504
rect 181220 269492 181226 269544
rect 204162 269492 204168 269544
rect 204220 269532 204226 269544
rect 223482 269532 223488 269544
rect 204220 269504 223488 269532
rect 204220 269492 204226 269504
rect 223482 269492 223488 269504
rect 223540 269492 223546 269544
rect 401686 269492 401692 269544
rect 401744 269532 401750 269544
rect 416774 269532 416780 269544
rect 401744 269504 416780 269532
rect 401744 269492 401750 269504
rect 416774 269492 416780 269504
rect 416832 269492 416838 269544
rect 424594 269492 424600 269544
rect 424652 269532 424658 269544
rect 475010 269532 475016 269544
rect 424652 269504 475016 269532
rect 424652 269492 424658 269504
rect 475010 269492 475016 269504
rect 475068 269492 475074 269544
rect 495250 269492 495256 269544
rect 495308 269532 495314 269544
rect 509712 269532 509740 269640
rect 532878 269628 532884 269680
rect 532936 269668 532942 269680
rect 616230 269668 616236 269680
rect 532936 269640 616236 269668
rect 532936 269628 532942 269640
rect 616230 269628 616236 269640
rect 616288 269628 616294 269680
rect 495308 269504 509740 269532
rect 495308 269492 495314 269504
rect 509878 269492 509884 269544
rect 509936 269532 509942 269544
rect 596174 269532 596180 269544
rect 509936 269504 596180 269532
rect 509936 269492 509942 269504
rect 596174 269492 596180 269504
rect 596232 269492 596238 269544
rect 126882 269356 126888 269408
rect 126940 269396 126946 269408
rect 178310 269396 178316 269408
rect 126940 269368 178316 269396
rect 126940 269356 126946 269368
rect 178310 269356 178316 269368
rect 178368 269356 178374 269408
rect 408402 269356 408408 269408
rect 408460 269396 408466 269408
rect 426526 269396 426532 269408
rect 408460 269368 426532 269396
rect 408460 269356 408466 269368
rect 426526 269356 426532 269368
rect 426584 269356 426590 269408
rect 441614 269356 441620 269408
rect 441672 269396 441678 269408
rect 458450 269396 458456 269408
rect 441672 269368 458456 269396
rect 441672 269356 441678 269368
rect 458450 269356 458456 269368
rect 458508 269356 458514 269408
rect 470962 269356 470968 269408
rect 471020 269396 471026 269408
rect 471020 269368 538444 269396
rect 471020 269356 471026 269368
rect 143902 269220 143908 269272
rect 143960 269260 143966 269272
rect 191098 269260 191104 269272
rect 143960 269232 191104 269260
rect 143960 269220 143966 269232
rect 191098 269220 191104 269232
rect 191156 269220 191162 269272
rect 282730 269220 282736 269272
rect 282788 269260 282794 269272
rect 288802 269260 288808 269272
rect 282788 269232 288808 269260
rect 282788 269220 282794 269232
rect 288802 269220 288808 269232
rect 288860 269220 288866 269272
rect 474274 269220 474280 269272
rect 474332 269260 474338 269272
rect 538214 269260 538220 269272
rect 474332 269232 538220 269260
rect 474332 269220 474338 269232
rect 538214 269220 538220 269232
rect 538272 269220 538278 269272
rect 538416 269260 538444 269368
rect 538582 269356 538588 269408
rect 538640 269396 538646 269408
rect 575474 269396 575480 269408
rect 538640 269368 575480 269396
rect 538640 269356 538646 269368
rect 575474 269356 575480 269368
rect 575532 269356 575538 269408
rect 540606 269260 540612 269272
rect 538416 269232 540612 269260
rect 540606 269220 540612 269232
rect 540664 269220 540670 269272
rect 540790 269220 540796 269272
rect 540848 269260 540854 269272
rect 543182 269260 543188 269272
rect 540848 269232 543188 269260
rect 540848 269220 540854 269232
rect 543182 269220 543188 269232
rect 543240 269220 543246 269272
rect 543366 269152 543372 269204
rect 543424 269192 543430 269204
rect 546494 269192 546500 269204
rect 543424 269164 546500 269192
rect 543424 269152 543430 269164
rect 546494 269152 546500 269164
rect 546552 269152 546558 269204
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 42150 269016 42156 269068
rect 42208 269056 42214 269068
rect 42886 269056 42892 269068
rect 42208 269028 42892 269056
rect 42208 269016 42214 269028
rect 42886 269016 42892 269028
rect 42944 269016 42950 269068
rect 118602 269016 118608 269068
rect 118660 269056 118666 269068
rect 174538 269056 174544 269068
rect 118660 269028 174544 269056
rect 118660 269016 118666 269028
rect 174538 269016 174544 269028
rect 174596 269016 174602 269068
rect 175090 269016 175096 269068
rect 175148 269056 175154 269068
rect 177666 269056 177672 269068
rect 175148 269028 177672 269056
rect 175148 269016 175154 269028
rect 177666 269016 177672 269028
rect 177724 269016 177730 269068
rect 273254 269016 273260 269068
rect 273312 269056 273318 269068
rect 275554 269056 275560 269068
rect 273312 269028 275560 269056
rect 273312 269016 273318 269028
rect 275554 269016 275560 269028
rect 275612 269016 275618 269068
rect 436554 269016 436560 269068
rect 436612 269056 436618 269068
rect 491662 269056 491668 269068
rect 436612 269028 491668 269056
rect 436612 269016 436618 269028
rect 491662 269016 491668 269028
rect 491720 269016 491726 269068
rect 495802 269016 495808 269068
rect 495860 269056 495866 269068
rect 576854 269056 576860 269068
rect 495860 269028 576860 269056
rect 495860 269016 495866 269028
rect 576854 269016 576860 269028
rect 576912 269016 576918 269068
rect 115750 268880 115756 268932
rect 115808 268920 115814 268932
rect 171226 268920 171232 268932
rect 115808 268892 171232 268920
rect 115808 268880 115814 268892
rect 171226 268880 171232 268892
rect 171284 268880 171290 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 415486 268920 415492 268932
rect 382424 268892 415492 268920
rect 382424 268880 382430 268892
rect 415486 268880 415492 268892
rect 415544 268880 415550 268932
rect 433702 268880 433708 268932
rect 433760 268920 433766 268932
rect 488534 268920 488540 268932
rect 433760 268892 488540 268920
rect 433760 268880 433766 268892
rect 488534 268880 488540 268892
rect 488592 268880 488598 268932
rect 498286 268880 498292 268932
rect 498344 268920 498350 268932
rect 580994 268920 581000 268932
rect 498344 268892 581000 268920
rect 498344 268880 498350 268892
rect 580994 268880 581000 268892
rect 581052 268880 581058 268932
rect 188890 268812 188896 268864
rect 188948 268852 188954 268864
rect 190454 268852 190460 268864
rect 188948 268824 190460 268852
rect 188948 268812 188954 268824
rect 190454 268812 190460 268824
rect 190512 268812 190518 268864
rect 110322 268744 110328 268796
rect 110380 268784 110386 268796
rect 167914 268784 167920 268796
rect 110380 268756 167920 268784
rect 110380 268744 110386 268756
rect 167914 268744 167920 268756
rect 167972 268744 167978 268796
rect 168282 268744 168288 268796
rect 168340 268784 168346 268796
rect 181990 268784 181996 268796
rect 168340 268756 181996 268784
rect 168340 268744 168346 268756
rect 181990 268744 181996 268756
rect 182048 268744 182054 268796
rect 200574 268744 200580 268796
rect 200632 268784 200638 268796
rect 231302 268784 231308 268796
rect 200632 268756 231308 268784
rect 200632 268744 200638 268756
rect 231302 268744 231308 268756
rect 231360 268744 231366 268796
rect 387334 268744 387340 268796
rect 387392 268784 387398 268796
rect 422294 268784 422300 268796
rect 387392 268756 422300 268784
rect 387392 268744 387398 268756
rect 422294 268744 422300 268756
rect 422352 268744 422358 268796
rect 438670 268744 438676 268796
rect 438728 268784 438734 268796
rect 495434 268784 495440 268796
rect 438728 268756 495440 268784
rect 438728 268744 438734 268756
rect 495434 268744 495440 268756
rect 495492 268744 495498 268796
rect 500770 268744 500776 268796
rect 500828 268784 500834 268796
rect 583754 268784 583760 268796
rect 500828 268756 583760 268784
rect 500828 268744 500834 268756
rect 583754 268744 583760 268756
rect 583812 268744 583818 268796
rect 104986 268608 104992 268660
rect 105044 268648 105050 268660
rect 163774 268648 163780 268660
rect 105044 268620 163780 268648
rect 105044 268608 105050 268620
rect 163774 268608 163780 268620
rect 163832 268608 163838 268660
rect 176930 268608 176936 268660
rect 176988 268648 176994 268660
rect 215110 268648 215116 268660
rect 176988 268620 215116 268648
rect 176988 268608 176994 268620
rect 215110 268608 215116 268620
rect 215168 268608 215174 268660
rect 224218 268608 224224 268660
rect 224276 268648 224282 268660
rect 243262 268648 243268 268660
rect 224276 268620 243268 268648
rect 224276 268608 224282 268620
rect 243262 268608 243268 268620
rect 243320 268608 243326 268660
rect 352558 268608 352564 268660
rect 352616 268648 352622 268660
rect 372614 268648 372620 268660
rect 352616 268620 372620 268648
rect 352616 268608 352622 268620
rect 372614 268608 372620 268620
rect 372672 268608 372678 268660
rect 393314 268608 393320 268660
rect 393372 268648 393378 268660
rect 429194 268648 429200 268660
rect 393372 268620 429200 268648
rect 393372 268608 393378 268620
rect 429194 268608 429200 268620
rect 429252 268608 429258 268660
rect 441154 268608 441160 268660
rect 441212 268648 441218 268660
rect 499574 268648 499580 268660
rect 441212 268620 499580 268648
rect 441212 268608 441218 268620
rect 499574 268608 499580 268620
rect 499632 268608 499638 268660
rect 503254 268608 503260 268660
rect 503312 268648 503318 268660
rect 587894 268648 587900 268660
rect 503312 268620 587900 268648
rect 503312 268608 503318 268620
rect 587894 268608 587900 268620
rect 587952 268608 587958 268660
rect 99282 268472 99288 268524
rect 99340 268512 99346 268524
rect 160462 268512 160468 268524
rect 99340 268484 160468 268512
rect 99340 268472 99346 268484
rect 160462 268472 160468 268484
rect 160520 268472 160526 268524
rect 180702 268472 180708 268524
rect 180760 268512 180766 268524
rect 217594 268512 217600 268524
rect 180760 268484 217600 268512
rect 180760 268472 180766 268484
rect 217594 268472 217600 268484
rect 217652 268472 217658 268524
rect 231670 268472 231676 268524
rect 231728 268512 231734 268524
rect 253198 268512 253204 268524
rect 231728 268484 253204 268512
rect 231728 268472 231734 268484
rect 253198 268472 253204 268484
rect 253256 268472 253262 268524
rect 338482 268472 338488 268524
rect 338540 268512 338546 268524
rect 352098 268512 352104 268524
rect 338540 268484 352104 268512
rect 338540 268472 338546 268484
rect 352098 268472 352104 268484
rect 352156 268472 352162 268524
rect 367462 268472 367468 268524
rect 367520 268512 367526 268524
rect 393498 268512 393504 268524
rect 367520 268484 393504 268512
rect 367520 268472 367526 268484
rect 393498 268472 393504 268484
rect 393556 268472 393562 268524
rect 397270 268472 397276 268524
rect 397328 268512 397334 268524
rect 436094 268512 436100 268524
rect 397328 268484 436100 268512
rect 397328 268472 397334 268484
rect 436094 268472 436100 268484
rect 436152 268472 436158 268524
rect 446122 268472 446128 268524
rect 446180 268512 446186 268524
rect 506474 268512 506480 268524
rect 446180 268484 506480 268512
rect 446180 268472 446186 268484
rect 506474 268472 506480 268484
rect 506532 268472 506538 268524
rect 508222 268472 508228 268524
rect 508280 268512 508286 268524
rect 594794 268512 594800 268524
rect 508280 268484 594800 268512
rect 508280 268472 508286 268484
rect 594794 268472 594800 268484
rect 594852 268472 594858 268524
rect 92382 268336 92388 268388
rect 92440 268376 92446 268388
rect 155494 268376 155500 268388
rect 92440 268348 155500 268376
rect 92440 268336 92446 268348
rect 155494 268336 155500 268348
rect 155552 268336 155558 268388
rect 161566 268336 161572 268388
rect 161624 268376 161630 268388
rect 203518 268376 203524 268388
rect 161624 268348 203524 268376
rect 161624 268336 161630 268348
rect 203518 268336 203524 268348
rect 203576 268336 203582 268388
rect 210694 268336 210700 268388
rect 210752 268376 210758 268388
rect 236638 268376 236644 268388
rect 210752 268348 236644 268376
rect 210752 268336 210758 268348
rect 236638 268336 236644 268348
rect 236696 268336 236702 268388
rect 252646 268336 252652 268388
rect 252704 268376 252710 268388
rect 268102 268376 268108 268388
rect 252704 268348 268108 268376
rect 252704 268336 252710 268348
rect 268102 268336 268108 268348
rect 268160 268336 268166 268388
rect 348786 268336 348792 268388
rect 348844 268376 348850 268388
rect 367094 268376 367100 268388
rect 348844 268348 367100 268376
rect 348844 268336 348850 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 372430 268336 372436 268388
rect 372488 268376 372494 268388
rect 400490 268376 400496 268388
rect 372488 268348 400496 268376
rect 372488 268336 372494 268348
rect 400490 268336 400496 268348
rect 400548 268336 400554 268388
rect 402238 268336 402244 268388
rect 402296 268376 402302 268388
rect 443086 268376 443092 268388
rect 402296 268348 443092 268376
rect 402296 268336 402302 268348
rect 443086 268336 443092 268348
rect 443144 268336 443150 268388
rect 461854 268336 461860 268388
rect 461912 268376 461918 268388
rect 528554 268376 528560 268388
rect 461912 268348 528560 268376
rect 461912 268336 461918 268348
rect 528554 268336 528560 268348
rect 528612 268336 528618 268388
rect 541342 268336 541348 268388
rect 541400 268376 541406 268388
rect 641714 268376 641720 268388
rect 541400 268348 641720 268376
rect 541400 268336 541406 268348
rect 641714 268336 641720 268348
rect 641772 268336 641778 268388
rect 135622 268200 135628 268252
rect 135680 268240 135686 268252
rect 140130 268240 140136 268252
rect 135680 268212 140136 268240
rect 135680 268200 135686 268212
rect 140130 268200 140136 268212
rect 140188 268200 140194 268252
rect 140682 268200 140688 268252
rect 140740 268240 140746 268252
rect 188614 268240 188620 268252
rect 140740 268212 188620 268240
rect 140740 268200 140746 268212
rect 188614 268200 188620 268212
rect 188672 268200 188678 268252
rect 416222 268200 416228 268252
rect 416280 268240 416286 268252
rect 447134 268240 447140 268252
rect 416280 268212 447140 268240
rect 416280 268200 416286 268212
rect 447134 268200 447140 268212
rect 447192 268200 447198 268252
rect 493318 268200 493324 268252
rect 493376 268240 493382 268252
rect 574094 268240 574100 268252
rect 493376 268212 574100 268240
rect 493376 268200 493382 268212
rect 574094 268200 574100 268212
rect 574152 268200 574158 268252
rect 151722 268064 151728 268116
rect 151780 268104 151786 268116
rect 196066 268104 196072 268116
rect 151780 268076 196072 268104
rect 151780 268064 151786 268076
rect 196066 268064 196072 268076
rect 196124 268064 196130 268116
rect 422294 268064 422300 268116
rect 422352 268104 422358 268116
rect 444374 268104 444380 268116
rect 422352 268076 444380 268104
rect 422352 268064 422358 268076
rect 444374 268064 444380 268076
rect 444432 268064 444438 268116
rect 448422 268064 448428 268116
rect 448480 268104 448486 268116
rect 494054 268104 494060 268116
rect 448480 268076 494060 268104
rect 448480 268064 448486 268076
rect 494054 268064 494060 268076
rect 494112 268064 494118 268116
rect 527174 268064 527180 268116
rect 527232 268104 527238 268116
rect 607398 268104 607404 268116
rect 527232 268076 607404 268104
rect 527232 268064 527238 268076
rect 607398 268064 607404 268076
rect 607456 268064 607462 268116
rect 490834 267928 490840 267980
rect 490892 267968 490898 267980
rect 570046 267968 570052 267980
rect 490892 267940 570052 267968
rect 490892 267928 490898 267940
rect 570046 267928 570052 267940
rect 570104 267928 570110 267980
rect 276474 267724 276480 267776
rect 276532 267764 276538 267776
rect 278038 267764 278044 267776
rect 276532 267736 278044 267764
rect 276532 267724 276538 267736
rect 278038 267724 278044 267736
rect 278096 267724 278102 267776
rect 119338 267656 119344 267708
rect 119396 267696 119402 267708
rect 153470 267696 153476 267708
rect 119396 267668 153476 267696
rect 119396 267656 119402 267668
rect 153470 267656 153476 267668
rect 153528 267656 153534 267708
rect 153838 267656 153844 267708
rect 153896 267696 153902 267708
rect 184474 267696 184480 267708
rect 153896 267668 184480 267696
rect 153896 267656 153902 267668
rect 184474 267656 184480 267668
rect 184532 267656 184538 267708
rect 390646 267656 390652 267708
rect 390704 267696 390710 267708
rect 408402 267696 408408 267708
rect 390704 267668 408408 267696
rect 390704 267656 390710 267668
rect 408402 267656 408408 267668
rect 408460 267656 408466 267708
rect 422938 267656 422944 267708
rect 422996 267696 423002 267708
rect 438118 267696 438124 267708
rect 422996 267668 438124 267696
rect 422996 267656 423002 267668
rect 438118 267656 438124 267668
rect 438176 267656 438182 267708
rect 445294 267656 445300 267708
rect 445352 267696 445358 267708
rect 490558 267696 490564 267708
rect 445352 267668 490564 267696
rect 445352 267656 445358 267668
rect 490558 267656 490564 267668
rect 490616 267656 490622 267708
rect 509878 267656 509884 267708
rect 509936 267696 509942 267708
rect 567838 267696 567844 267708
rect 509936 267668 567844 267696
rect 509936 267656 509942 267668
rect 567838 267656 567844 267668
rect 567896 267656 567902 267708
rect 111702 267520 111708 267572
rect 111760 267560 111766 267572
rect 168558 267560 168564 267572
rect 111760 267532 168564 267560
rect 111760 267520 111766 267532
rect 168558 267520 168564 267532
rect 168616 267520 168622 267572
rect 169018 267520 169024 267572
rect 169076 267560 169082 267572
rect 199378 267560 199384 267572
rect 169076 267532 199384 267560
rect 169076 267520 169082 267532
rect 199378 267520 199384 267532
rect 199436 267520 199442 267572
rect 215938 267520 215944 267572
rect 215996 267560 216002 267572
rect 222562 267560 222568 267572
rect 215996 267532 222568 267560
rect 215996 267520 216002 267532
rect 222562 267520 222568 267532
rect 222620 267520 222626 267572
rect 353386 267520 353392 267572
rect 353444 267560 353450 267572
rect 374454 267560 374460 267572
rect 353444 267532 374460 267560
rect 353444 267520 353450 267532
rect 374454 267520 374460 267532
rect 374512 267520 374518 267572
rect 380710 267520 380716 267572
rect 380768 267560 380774 267572
rect 398742 267560 398748 267572
rect 380768 267532 398748 267560
rect 380768 267520 380774 267532
rect 398742 267520 398748 267532
rect 398800 267520 398806 267572
rect 404722 267520 404728 267572
rect 404780 267560 404786 267572
rect 416222 267560 416228 267572
rect 404780 267532 416228 267560
rect 404780 267520 404786 267532
rect 416222 267520 416228 267532
rect 416280 267520 416286 267572
rect 421282 267520 421288 267572
rect 421340 267560 421346 267572
rect 440878 267560 440884 267572
rect 421340 267532 440884 267560
rect 421340 267520 421346 267532
rect 440878 267520 440884 267532
rect 440936 267520 440942 267572
rect 450262 267520 450268 267572
rect 450320 267560 450326 267572
rect 498838 267560 498844 267572
rect 450320 267532 498844 267560
rect 450320 267520 450326 267532
rect 498838 267520 498844 267532
rect 498896 267520 498902 267572
rect 514846 267520 514852 267572
rect 514904 267560 514910 267572
rect 578878 267560 578884 267572
rect 514904 267532 578884 267560
rect 514904 267520 514910 267532
rect 578878 267520 578884 267532
rect 578936 267520 578942 267572
rect 86218 267384 86224 267436
rect 86276 267424 86282 267436
rect 144730 267424 144736 267436
rect 86276 267396 144736 267424
rect 86276 267384 86282 267396
rect 144730 267384 144736 267396
rect 144788 267384 144794 267436
rect 145558 267384 145564 267436
rect 145616 267424 145622 267436
rect 191926 267424 191932 267436
rect 145616 267396 191932 267424
rect 145616 267384 145622 267396
rect 191926 267384 191932 267396
rect 191984 267384 191990 267436
rect 199562 267384 199568 267436
rect 199620 267424 199626 267436
rect 204346 267424 204352 267436
rect 199620 267396 204352 267424
rect 199620 267384 199626 267396
rect 204346 267384 204352 267396
rect 204404 267384 204410 267436
rect 205450 267384 205456 267436
rect 205508 267424 205514 267436
rect 218422 267424 218428 267436
rect 205508 267396 218428 267424
rect 205508 267384 205514 267396
rect 218422 267384 218428 267396
rect 218480 267384 218486 267436
rect 233878 267384 233884 267436
rect 233936 267424 233942 267436
rect 233936 267396 238754 267424
rect 233936 267384 233942 267396
rect 104802 267248 104808 267300
rect 104860 267288 104866 267300
rect 164602 267288 164608 267300
rect 104860 267260 164608 267288
rect 104860 267248 104866 267260
rect 164602 267248 164608 267260
rect 164660 267248 164666 267300
rect 186958 267248 186964 267300
rect 187016 267288 187022 267300
rect 219250 267288 219256 267300
rect 187016 267260 219256 267288
rect 187016 267248 187022 267260
rect 219250 267248 219256 267260
rect 219308 267248 219314 267300
rect 223482 267248 223488 267300
rect 223540 267288 223546 267300
rect 234154 267288 234160 267300
rect 223540 267260 234160 267288
rect 223540 267248 223546 267260
rect 234154 267248 234160 267260
rect 234212 267248 234218 267300
rect 238726 267288 238754 267396
rect 243538 267384 243544 267436
rect 243596 267424 243602 267436
rect 251542 267424 251548 267436
rect 243596 267396 251548 267424
rect 243596 267384 243602 267396
rect 251542 267384 251548 267396
rect 251600 267384 251606 267436
rect 315298 267384 315304 267436
rect 315356 267424 315362 267436
rect 319162 267424 319168 267436
rect 315356 267396 319168 267424
rect 315356 267384 315362 267396
rect 319162 267384 319168 267396
rect 319220 267384 319226 267436
rect 340966 267384 340972 267436
rect 341024 267424 341030 267436
rect 355318 267424 355324 267436
rect 341024 267396 355324 267424
rect 341024 267384 341030 267396
rect 355318 267384 355324 267396
rect 355376 267384 355382 267436
rect 368290 267384 368296 267436
rect 368348 267424 368354 267436
rect 385678 267424 385684 267436
rect 368348 267396 385684 267424
rect 368348 267384 368354 267396
rect 385678 267384 385684 267396
rect 385736 267384 385742 267436
rect 398098 267384 398104 267436
rect 398156 267424 398162 267436
rect 417418 267424 417424 267436
rect 398156 267396 417424 267424
rect 398156 267384 398162 267396
rect 417418 267384 417424 267396
rect 417476 267384 417482 267436
rect 428734 267384 428740 267436
rect 428792 267424 428798 267436
rect 447778 267424 447784 267436
rect 428792 267396 447784 267424
rect 428792 267384 428798 267396
rect 447778 267384 447784 267396
rect 447836 267384 447842 267436
rect 460198 267384 460204 267436
rect 460256 267424 460262 267436
rect 516778 267424 516784 267436
rect 460256 267396 516784 267424
rect 460256 267384 460262 267396
rect 516778 267384 516784 267396
rect 516836 267384 516842 267436
rect 519814 267384 519820 267436
rect 519872 267424 519878 267436
rect 583018 267424 583024 267436
rect 519872 267396 583024 267424
rect 519872 267384 519878 267396
rect 583018 267384 583024 267396
rect 583076 267384 583082 267436
rect 244090 267288 244096 267300
rect 238726 267260 244096 267288
rect 244090 267248 244096 267260
rect 244148 267248 244154 267300
rect 321922 267248 321928 267300
rect 321980 267288 321986 267300
rect 327718 267288 327724 267300
rect 321980 267260 327724 267288
rect 321980 267248 321986 267260
rect 327718 267248 327724 267260
rect 327776 267248 327782 267300
rect 350902 267248 350908 267300
rect 350960 267288 350966 267300
rect 362218 267288 362224 267300
rect 350960 267260 362224 267288
rect 350960 267248 350966 267260
rect 362218 267248 362224 267260
rect 362276 267248 362282 267300
rect 371602 267248 371608 267300
rect 371660 267288 371666 267300
rect 373258 267288 373264 267300
rect 371660 267260 373264 267288
rect 371660 267248 371666 267260
rect 373258 267248 373264 267260
rect 373316 267248 373322 267300
rect 373442 267248 373448 267300
rect 373500 267288 373506 267300
rect 381538 267288 381544 267300
rect 373500 267260 381544 267288
rect 373500 267248 373506 267260
rect 381538 267248 381544 267260
rect 381596 267248 381602 267300
rect 383194 267248 383200 267300
rect 383252 267288 383258 267300
rect 401686 267288 401692 267300
rect 383252 267260 401692 267288
rect 383252 267248 383258 267260
rect 401686 267248 401692 267260
rect 401744 267248 401750 267300
rect 403066 267248 403072 267300
rect 403124 267288 403130 267300
rect 422294 267288 422300 267300
rect 403124 267260 422300 267288
rect 403124 267248 403130 267260
rect 422294 267248 422300 267260
rect 422352 267248 422358 267300
rect 432874 267248 432880 267300
rect 432932 267288 432938 267300
rect 453298 267288 453304 267300
rect 432932 267260 453304 267288
rect 432932 267248 432938 267260
rect 453298 267248 453304 267260
rect 453356 267248 453362 267300
rect 462958 267288 462964 267300
rect 454972 267260 462964 267288
rect 90358 267112 90364 267164
rect 90416 267152 90422 267164
rect 151354 267152 151360 267164
rect 90416 267124 151360 267152
rect 90416 267112 90422 267124
rect 151354 267112 151360 267124
rect 151412 267112 151418 267164
rect 168098 267112 168104 267164
rect 168156 267152 168162 267164
rect 177022 267152 177028 267164
rect 168156 267124 177028 267152
rect 168156 267112 168162 267124
rect 177022 267112 177028 267124
rect 177080 267112 177086 267164
rect 177666 267112 177672 267164
rect 177724 267152 177730 267164
rect 214282 267152 214288 267164
rect 177724 267124 214288 267152
rect 177724 267112 177730 267124
rect 214282 267112 214288 267124
rect 214340 267112 214346 267164
rect 220078 267112 220084 267164
rect 220136 267152 220142 267164
rect 239122 267152 239128 267164
rect 220136 267124 239128 267152
rect 220136 267112 220142 267124
rect 239122 267112 239128 267124
rect 239180 267112 239186 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 362494 267112 362500 267164
rect 362552 267152 362558 267164
rect 369118 267152 369124 267164
rect 362552 267124 369124 267152
rect 362552 267112 362558 267124
rect 369118 267112 369124 267124
rect 369176 267112 369182 267164
rect 373258 267112 373264 267164
rect 373316 267152 373322 267164
rect 392026 267152 392032 267164
rect 373316 267124 392032 267152
rect 373316 267112 373322 267124
rect 392026 267112 392032 267124
rect 392084 267112 392090 267164
rect 394786 267112 394792 267164
rect 394844 267152 394850 267164
rect 403618 267152 403624 267164
rect 394844 267124 403624 267152
rect 394844 267112 394850 267124
rect 403618 267112 403624 267124
rect 403676 267112 403682 267164
rect 413002 267112 413008 267164
rect 413060 267152 413066 267164
rect 441614 267152 441620 267164
rect 413060 267124 441620 267152
rect 413060 267112 413066 267124
rect 441614 267112 441620 267124
rect 441672 267112 441678 267164
rect 447134 267112 447140 267164
rect 447192 267152 447198 267164
rect 448422 267152 448428 267164
rect 447192 267124 448428 267152
rect 447192 267112 447198 267124
rect 448422 267112 448428 267124
rect 448480 267112 448486 267164
rect 452746 267112 452752 267164
rect 452804 267152 452810 267164
rect 454972 267152 455000 267260
rect 462958 267248 462964 267260
rect 463016 267248 463022 267300
rect 465166 267248 465172 267300
rect 465224 267288 465230 267300
rect 523678 267288 523684 267300
rect 465224 267260 523684 267288
rect 465224 267248 465230 267260
rect 523678 267248 523684 267260
rect 523736 267248 523742 267300
rect 524782 267248 524788 267300
rect 524840 267288 524846 267300
rect 611998 267288 612004 267300
rect 524840 267260 612004 267288
rect 524840 267248 524846 267260
rect 611998 267248 612004 267260
rect 612056 267248 612062 267300
rect 452804 267124 455000 267152
rect 452804 267112 452810 267124
rect 455138 267112 455144 267164
rect 455196 267152 455202 267164
rect 515398 267152 515404 267164
rect 455196 267124 515404 267152
rect 455196 267112 455202 267124
rect 515398 267112 515404 267124
rect 515456 267112 515462 267164
rect 517238 267112 517244 267164
rect 517296 267152 517302 267164
rect 527174 267152 527180 267164
rect 517296 267124 527180 267152
rect 517296 267112 517302 267124
rect 527174 267112 527180 267124
rect 527232 267112 527238 267164
rect 529658 267112 529664 267164
rect 529716 267152 529722 267164
rect 617518 267152 617524 267164
rect 529716 267124 617524 267152
rect 529716 267112 529722 267124
rect 617518 267112 617524 267124
rect 617576 267112 617582 267164
rect 79318 266976 79324 267028
rect 79376 267016 79382 267028
rect 79376 266988 122834 267016
rect 79376 266976 79382 266988
rect 122806 266880 122834 266988
rect 140130 266976 140136 267028
rect 140188 267016 140194 267028
rect 186958 267016 186964 267028
rect 140188 266988 186964 267016
rect 140188 266976 140194 266988
rect 186958 266976 186964 266988
rect 187016 266976 187022 267028
rect 190454 266976 190460 267028
rect 190512 267016 190518 267028
rect 224218 267016 224224 267028
rect 190512 266988 224224 267016
rect 190512 266976 190518 266988
rect 224218 266976 224224 266988
rect 224276 266976 224282 267028
rect 228358 266976 228364 267028
rect 228416 267016 228422 267028
rect 228416 266988 238754 267016
rect 228416 266976 228422 266988
rect 140590 266880 140596 266892
rect 122806 266852 140596 266880
rect 140590 266840 140596 266852
rect 140648 266840 140654 266892
rect 150526 266880 150532 266892
rect 140792 266852 150532 266880
rect 137462 266704 137468 266756
rect 137520 266744 137526 266756
rect 140792 266744 140820 266852
rect 150526 266840 150532 266852
rect 150584 266840 150590 266892
rect 159450 266840 159456 266892
rect 159508 266880 159514 266892
rect 162118 266880 162124 266892
rect 159508 266852 162124 266880
rect 159508 266840 159514 266852
rect 162118 266840 162124 266852
rect 162176 266840 162182 266892
rect 178678 266840 178684 266892
rect 178736 266880 178742 266892
rect 209314 266880 209320 266892
rect 178736 266852 209320 266880
rect 178736 266840 178742 266852
rect 209314 266840 209320 266852
rect 209372 266840 209378 266892
rect 218698 266840 218704 266892
rect 218756 266880 218762 266892
rect 220906 266880 220912 266892
rect 218756 266852 220912 266880
rect 218756 266840 218762 266852
rect 220906 266840 220912 266852
rect 220964 266840 220970 266892
rect 238726 266880 238754 266988
rect 249058 266976 249064 267028
rect 249116 267016 249122 267028
rect 250714 267016 250720 267028
rect 249116 266988 250720 267016
rect 249116 266976 249122 266988
rect 250714 266976 250720 266988
rect 250772 266976 250778 267028
rect 255958 266976 255964 267028
rect 256016 267016 256022 267028
rect 258994 267016 259000 267028
rect 256016 266988 259000 267016
rect 256016 266976 256022 266988
rect 258994 266976 259000 266988
rect 259052 266976 259058 267028
rect 286318 266976 286324 267028
rect 286376 267016 286382 267028
rect 287974 267016 287980 267028
rect 286376 266988 287980 267016
rect 286376 266976 286382 266988
rect 287974 266976 287980 266988
rect 288032 266976 288038 267028
rect 312814 266976 312820 267028
rect 312872 267016 312878 267028
rect 316034 267016 316040 267028
rect 312872 266988 316040 267016
rect 312872 266976 312878 266988
rect 316034 266976 316040 266988
rect 316092 266976 316098 267028
rect 316954 266976 316960 267028
rect 317012 267016 317018 267028
rect 321554 267016 321560 267028
rect 317012 266988 321560 267016
rect 317012 266976 317018 266988
rect 321554 266976 321560 266988
rect 321612 266976 321618 267028
rect 365806 266976 365812 267028
rect 365864 267016 365870 267028
rect 373442 267016 373448 267028
rect 365864 266988 373448 267016
rect 365864 266976 365870 266988
rect 373442 266976 373448 266988
rect 373500 266976 373506 267028
rect 393130 266976 393136 267028
rect 393188 267016 393194 267028
rect 420178 267016 420184 267028
rect 393188 266988 420184 267016
rect 393188 266976 393194 266988
rect 420178 266976 420184 266988
rect 420236 266976 420242 267028
rect 457438 267016 457444 267028
rect 431926 266988 457444 267016
rect 249058 266880 249064 266892
rect 238726 266852 249064 266880
rect 249058 266840 249064 266852
rect 249116 266840 249122 266892
rect 314470 266840 314476 266892
rect 314528 266880 314534 266892
rect 318978 266880 318984 266892
rect 314528 266852 318984 266880
rect 314528 266840 314534 266852
rect 318978 266840 318984 266852
rect 319036 266840 319042 266892
rect 332686 266840 332692 266892
rect 332744 266880 332750 266892
rect 343818 266880 343824 266892
rect 332744 266852 343824 266880
rect 332744 266840 332750 266852
rect 343818 266840 343824 266852
rect 343876 266840 343882 266892
rect 378226 266840 378232 266892
rect 378284 266880 378290 266892
rect 394970 266880 394976 266892
rect 378284 266852 394976 266880
rect 378284 266840 378290 266852
rect 394970 266840 394976 266852
rect 395028 266840 395034 266892
rect 427906 266840 427912 266892
rect 427964 266880 427970 266892
rect 431926 266880 431954 266988
rect 457438 266976 457444 266988
rect 457496 266976 457502 267028
rect 470134 266976 470140 267028
rect 470192 267016 470198 267028
rect 534718 267016 534724 267028
rect 470192 266988 534724 267016
rect 470192 266976 470198 266988
rect 534718 266976 534724 266988
rect 534776 266976 534782 267028
rect 539686 266976 539692 267028
rect 539744 267016 539750 267028
rect 634078 267016 634084 267028
rect 539744 266988 634084 267016
rect 539744 266976 539750 266988
rect 634078 266976 634084 266988
rect 634136 266976 634142 267028
rect 427964 266852 431954 266880
rect 427964 266840 427970 266852
rect 442718 266840 442724 266892
rect 442776 266880 442782 266892
rect 485038 266880 485044 266892
rect 442776 266852 485044 266880
rect 442776 266840 442782 266852
rect 485038 266840 485044 266852
rect 485096 266840 485102 266892
rect 499942 266840 499948 266892
rect 500000 266880 500006 266892
rect 507854 266880 507860 266892
rect 500000 266852 507860 266880
rect 500000 266840 500006 266852
rect 507854 266840 507860 266852
rect 507912 266840 507918 266892
rect 534718 266840 534724 266892
rect 534776 266880 534782 266892
rect 589918 266880 589924 266892
rect 534776 266852 589924 266880
rect 534776 266840 534782 266852
rect 589918 266840 589924 266852
rect 589976 266840 589982 266892
rect 137520 266716 140820 266744
rect 137520 266704 137526 266716
rect 151078 266704 151084 266756
rect 151136 266744 151142 266756
rect 179506 266744 179512 266756
rect 151136 266716 179512 266744
rect 151136 266704 151142 266716
rect 179506 266704 179512 266716
rect 179564 266704 179570 266756
rect 347498 266704 347504 266756
rect 347556 266744 347562 266756
rect 351178 266744 351184 266756
rect 347556 266716 351184 266744
rect 347556 266704 347562 266716
rect 351178 266704 351184 266716
rect 351236 266704 351242 266756
rect 388162 266704 388168 266756
rect 388220 266744 388226 266756
rect 404354 266744 404360 266756
rect 388220 266716 404360 266744
rect 388220 266704 388226 266716
rect 404354 266704 404360 266716
rect 404412 266704 404418 266756
rect 408034 266704 408040 266756
rect 408092 266744 408098 266756
rect 423950 266744 423956 266756
rect 408092 266716 423956 266744
rect 408092 266704 408098 266716
rect 423950 266704 423956 266716
rect 424008 266704 424014 266756
rect 434530 266704 434536 266756
rect 434588 266744 434594 266756
rect 449158 266744 449164 266756
rect 434588 266716 449164 266744
rect 434588 266704 434594 266716
rect 449158 266704 449164 266716
rect 449216 266704 449222 266756
rect 457714 266704 457720 266756
rect 457772 266744 457778 266756
rect 476758 266744 476764 266756
rect 457772 266716 476764 266744
rect 457772 266704 457778 266716
rect 476758 266704 476764 266716
rect 476816 266704 476822 266756
rect 485038 266704 485044 266756
rect 485096 266744 485102 266756
rect 485096 266716 489914 266744
rect 485096 266704 485102 266716
rect 308674 266636 308680 266688
rect 308732 266676 308738 266688
rect 310514 266676 310520 266688
rect 308732 266648 310520 266676
rect 308732 266636 308738 266648
rect 310514 266636 310520 266648
rect 310572 266636 310578 266688
rect 313642 266636 313648 266688
rect 313700 266676 313706 266688
rect 317414 266676 317420 266688
rect 313700 266648 317420 266676
rect 313700 266636 313706 266648
rect 317414 266636 317420 266648
rect 317472 266636 317478 266688
rect 317782 266636 317788 266688
rect 317840 266676 317846 266688
rect 322934 266676 322940 266688
rect 317840 266648 322940 266676
rect 317840 266636 317846 266648
rect 322934 266636 322940 266648
rect 322992 266636 322998 266688
rect 360010 266636 360016 266688
rect 360068 266676 360074 266688
rect 366358 266676 366364 266688
rect 360068 266648 366364 266676
rect 360068 266636 360074 266648
rect 366358 266636 366364 266648
rect 366416 266636 366422 266688
rect 130378 266568 130384 266620
rect 130436 266608 130442 266620
rect 138106 266608 138112 266620
rect 130436 266580 138112 266608
rect 130436 266568 130442 266580
rect 138106 266568 138112 266580
rect 138164 266568 138170 266620
rect 149606 266568 149612 266620
rect 149664 266608 149670 266620
rect 159634 266608 159640 266620
rect 149664 266580 159640 266608
rect 149664 266568 149670 266580
rect 159634 266568 159640 266580
rect 159692 266568 159698 266620
rect 345106 266568 345112 266620
rect 345164 266608 345170 266620
rect 348418 266608 348424 266620
rect 345164 266580 348424 266608
rect 345164 266568 345170 266580
rect 348418 266568 348424 266580
rect 348476 266568 348482 266620
rect 399754 266568 399760 266620
rect 399812 266608 399818 266620
rect 407758 266608 407764 266620
rect 399812 266580 407764 266608
rect 399812 266568 399818 266580
rect 407758 266568 407764 266580
rect 407816 266568 407822 266620
rect 414658 266608 414664 266620
rect 407960 266580 414664 266608
rect 310330 266500 310336 266552
rect 310388 266540 310394 266552
rect 311894 266540 311900 266552
rect 310388 266512 311900 266540
rect 310388 266500 310394 266512
rect 311894 266500 311900 266512
rect 311952 266500 311958 266552
rect 312354 266500 312360 266552
rect 312412 266540 312418 266552
rect 314654 266540 314660 266552
rect 312412 266512 314660 266540
rect 312412 266500 312418 266512
rect 314654 266500 314660 266512
rect 314712 266500 314718 266552
rect 316126 266500 316132 266552
rect 316184 266540 316190 266552
rect 320174 266540 320180 266552
rect 316184 266512 320180 266540
rect 316184 266500 316190 266512
rect 320174 266500 320180 266512
rect 320232 266500 320238 266552
rect 327718 266500 327724 266552
rect 327776 266540 327782 266552
rect 331858 266540 331864 266552
rect 327776 266512 331864 266540
rect 327776 266500 327782 266512
rect 331858 266500 331864 266512
rect 331916 266500 331922 266552
rect 350074 266500 350080 266552
rect 350132 266540 350138 266552
rect 353938 266540 353944 266552
rect 350132 266512 353944 266540
rect 350132 266500 350138 266512
rect 353938 266500 353944 266512
rect 353996 266500 354002 266552
rect 355870 266500 355876 266552
rect 355928 266540 355934 266552
rect 360838 266540 360844 266552
rect 355928 266512 360844 266540
rect 355928 266500 355934 266512
rect 360838 266500 360844 266512
rect 360896 266500 360902 266552
rect 369946 266500 369952 266552
rect 370004 266540 370010 266552
rect 372246 266540 372252 266552
rect 370004 266512 372252 266540
rect 370004 266500 370010 266512
rect 372246 266500 372252 266512
rect 372304 266500 372310 266552
rect 374914 266500 374920 266552
rect 374972 266540 374978 266552
rect 380526 266540 380532 266552
rect 374972 266512 380532 266540
rect 374972 266500 374978 266512
rect 380526 266500 380532 266512
rect 380584 266500 380590 266552
rect 132494 266432 132500 266484
rect 132552 266472 132558 266484
rect 147214 266472 147220 266484
rect 132552 266444 147220 266472
rect 132552 266432 132558 266444
rect 147214 266432 147220 266444
rect 147272 266432 147278 266484
rect 342622 266432 342628 266484
rect 342680 266472 342686 266484
rect 345290 266472 345296 266484
rect 342680 266444 345296 266472
rect 342680 266432 342686 266444
rect 345290 266432 345296 266444
rect 345348 266432 345354 266484
rect 407206 266432 407212 266484
rect 407264 266472 407270 266484
rect 407960 266472 407988 266580
rect 414658 266568 414664 266580
rect 414716 266568 414722 266620
rect 437842 266568 437848 266620
rect 437900 266608 437906 266620
rect 447134 266608 447140 266620
rect 437900 266580 447140 266608
rect 437900 266568 437906 266580
rect 447134 266568 447140 266580
rect 447192 266568 447198 266620
rect 489886 266608 489914 266716
rect 490006 266704 490012 266756
rect 490064 266744 490070 266756
rect 509694 266744 509700 266756
rect 490064 266716 509700 266744
rect 490064 266704 490070 266716
rect 509694 266704 509700 266716
rect 509752 266704 509758 266756
rect 510706 266704 510712 266756
rect 510764 266744 510770 266756
rect 511810 266744 511816 266756
rect 510764 266716 511816 266744
rect 510764 266704 510770 266716
rect 511810 266704 511816 266716
rect 511868 266704 511874 266756
rect 512362 266704 512368 266756
rect 512420 266744 512426 266756
rect 513190 266744 513196 266756
rect 512420 266716 513196 266744
rect 512420 266704 512426 266716
rect 513190 266704 513196 266716
rect 513248 266704 513254 266756
rect 516502 266704 516508 266756
rect 516560 266744 516566 266756
rect 517422 266744 517428 266756
rect 516560 266716 517428 266744
rect 516560 266704 516566 266716
rect 517422 266704 517428 266716
rect 517480 266704 517486 266756
rect 518986 266704 518992 266756
rect 519044 266744 519050 266756
rect 520090 266744 520096 266756
rect 519044 266716 520096 266744
rect 519044 266704 519050 266716
rect 520090 266704 520096 266716
rect 520148 266704 520154 266756
rect 527266 266704 527272 266756
rect 527324 266744 527330 266756
rect 528186 266744 528192 266756
rect 527324 266716 528192 266744
rect 527324 266704 527330 266716
rect 528186 266704 528192 266716
rect 528244 266704 528250 266756
rect 528922 266704 528928 266756
rect 528980 266744 528986 266756
rect 529842 266744 529848 266756
rect 528980 266716 529848 266744
rect 528980 266704 528986 266716
rect 529842 266704 529848 266716
rect 529900 266704 529906 266756
rect 531406 266704 531412 266756
rect 531464 266744 531470 266756
rect 532510 266744 532516 266756
rect 531464 266716 532516 266744
rect 531464 266704 531470 266716
rect 532510 266704 532516 266716
rect 532568 266704 532574 266756
rect 533062 266704 533068 266756
rect 533120 266744 533126 266756
rect 533982 266744 533988 266756
rect 533120 266716 533988 266744
rect 533120 266704 533126 266716
rect 533982 266704 533988 266716
rect 534040 266704 534046 266756
rect 535546 266704 535552 266756
rect 535604 266744 535610 266756
rect 536742 266744 536748 266756
rect 535604 266716 536748 266744
rect 535604 266704 535610 266716
rect 536742 266704 536748 266716
rect 536800 266704 536806 266756
rect 542998 266704 543004 266756
rect 543056 266744 543062 266756
rect 598198 266744 598204 266756
rect 543056 266716 598204 266744
rect 543056 266704 543062 266716
rect 598198 266704 598204 266716
rect 598256 266704 598262 266756
rect 501598 266608 501604 266620
rect 489886 266580 501604 266608
rect 501598 266568 501604 266580
rect 501656 266568 501662 266620
rect 504818 266568 504824 266620
rect 504876 266608 504882 266620
rect 556798 266608 556804 266620
rect 504876 266580 556804 266608
rect 504876 266568 504882 266580
rect 556798 266568 556804 266580
rect 556856 266568 556862 266620
rect 423766 266500 423772 266552
rect 423824 266540 423830 266552
rect 425698 266540 425704 266552
rect 423824 266512 425704 266540
rect 423824 266500 423830 266512
rect 425698 266500 425704 266512
rect 425756 266500 425762 266552
rect 426250 266500 426256 266552
rect 426308 266540 426314 266552
rect 428458 266540 428464 266552
rect 426308 266512 428464 266540
rect 426308 266500 426314 266512
rect 428458 266500 428464 266512
rect 428516 266500 428522 266552
rect 447778 266500 447784 266552
rect 447836 266540 447842 266552
rect 456058 266540 456064 266552
rect 447836 266512 456064 266540
rect 447836 266500 447842 266512
rect 456058 266500 456064 266512
rect 456116 266500 456122 266552
rect 407264 266444 407988 266472
rect 407264 266432 407270 266444
rect 491662 266432 491668 266484
rect 491720 266472 491726 266484
rect 492582 266472 492588 266484
rect 491720 266444 492588 266472
rect 491720 266432 491726 266444
rect 492582 266432 492588 266444
rect 492640 266432 492646 266484
rect 494146 266432 494152 266484
rect 494204 266472 494210 266484
rect 495066 266472 495072 266484
rect 494204 266444 495072 266472
rect 494204 266432 494210 266444
rect 495066 266432 495072 266444
rect 495124 266432 495130 266484
rect 502426 266432 502432 266484
rect 502484 266472 502490 266484
rect 503438 266472 503444 266484
rect 502484 266444 503444 266472
rect 502484 266432 502490 266444
rect 503438 266432 503444 266444
rect 503496 266432 503502 266484
rect 504082 266432 504088 266484
rect 504140 266472 504146 266484
rect 505002 266472 505008 266484
rect 504140 266444 505008 266472
rect 504140 266432 504146 266444
rect 505002 266432 505008 266444
rect 505060 266432 505066 266484
rect 506566 266432 506572 266484
rect 506624 266472 506630 266484
rect 507670 266472 507676 266484
rect 506624 266444 507676 266472
rect 506624 266432 506630 266444
rect 507670 266432 507676 266444
rect 507728 266432 507734 266484
rect 507854 266432 507860 266484
rect 507912 266472 507918 266484
rect 549898 266472 549904 266484
rect 507912 266444 549904 266472
rect 507912 266432 507918 266444
rect 549898 266432 549904 266444
rect 549956 266432 549962 266484
rect 163498 266364 163504 266416
rect 163556 266404 163562 266416
rect 167086 266404 167092 266416
rect 163556 266376 167092 266404
rect 163556 266364 163562 266376
rect 167086 266364 167092 266376
rect 167144 266364 167150 266416
rect 168558 266364 168564 266416
rect 168616 266404 168622 266416
rect 169570 266404 169576 266416
rect 168616 266376 169576 266404
rect 168616 266364 168622 266376
rect 169570 266364 169576 266376
rect 169628 266364 169634 266416
rect 211154 266364 211160 266416
rect 211212 266404 211218 266416
rect 213454 266404 213460 266416
rect 211212 266376 213460 266404
rect 211212 266364 211218 266376
rect 213454 266364 213460 266376
rect 213512 266364 213518 266416
rect 214558 266364 214564 266416
rect 214616 266404 214622 266416
rect 215938 266404 215944 266416
rect 214616 266376 215944 266404
rect 214616 266364 214622 266376
rect 215938 266364 215944 266376
rect 215996 266364 216002 266416
rect 239398 266364 239404 266416
rect 239456 266404 239462 266416
rect 241606 266404 241612 266416
rect 239456 266376 241612 266404
rect 239456 266364 239462 266376
rect 241606 266364 241612 266376
rect 241664 266364 241670 266416
rect 243722 266364 243728 266416
rect 243780 266404 243786 266416
rect 246574 266404 246580 266416
rect 243780 266376 246580 266404
rect 243780 266364 243786 266376
rect 246574 266364 246580 266376
rect 246632 266364 246638 266416
rect 250438 266364 250444 266416
rect 250496 266404 250502 266416
rect 256510 266404 256516 266416
rect 250496 266376 256516 266404
rect 250496 266364 250502 266376
rect 256510 266364 256516 266376
rect 256568 266364 256574 266416
rect 300946 266364 300952 266416
rect 301004 266404 301010 266416
rect 302050 266404 302056 266416
rect 301004 266376 302056 266404
rect 301004 266364 301010 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 303706 266364 303712 266416
rect 303764 266404 303770 266416
rect 304534 266404 304540 266416
rect 303764 266376 304540 266404
rect 303764 266364 303770 266376
rect 304534 266364 304540 266376
rect 304592 266364 304598 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309134 266404 309140 266416
rect 307904 266376 309140 266404
rect 307904 266364 307910 266376
rect 309134 266364 309140 266376
rect 309192 266364 309198 266416
rect 309502 266364 309508 266416
rect 309560 266404 309566 266416
rect 310698 266404 310704 266416
rect 309560 266376 310704 266404
rect 309560 266364 309566 266376
rect 310698 266364 310704 266376
rect 310756 266364 310762 266416
rect 311158 266364 311164 266416
rect 311216 266404 311222 266416
rect 313274 266404 313280 266416
rect 311216 266376 313280 266404
rect 311216 266364 311222 266376
rect 313274 266364 313280 266376
rect 313332 266364 313338 266416
rect 320266 266364 320272 266416
rect 320324 266404 320330 266416
rect 321370 266404 321376 266416
rect 320324 266376 321376 266404
rect 320324 266364 320330 266376
rect 321370 266364 321376 266376
rect 321428 266364 321434 266416
rect 324406 266364 324412 266416
rect 324464 266404 324470 266416
rect 325326 266404 325332 266416
rect 324464 266376 325332 266404
rect 324464 266364 324470 266376
rect 325326 266364 325332 266376
rect 325384 266364 325390 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329742 266404 329748 266416
rect 328604 266376 329748 266404
rect 328604 266364 328610 266376
rect 329742 266364 329748 266376
rect 329800 266364 329806 266416
rect 336826 266364 336832 266416
rect 336884 266404 336890 266416
rect 337930 266404 337936 266416
rect 336884 266376 337936 266404
rect 336884 266364 336890 266376
rect 337930 266364 337936 266376
rect 337988 266364 337994 266416
rect 346762 266364 346768 266416
rect 346820 266404 346826 266416
rect 347682 266404 347688 266416
rect 346820 266376 347688 266404
rect 346820 266364 346826 266376
rect 347682 266364 347688 266376
rect 347740 266364 347746 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350350 266404 350356 266416
rect 349304 266376 350356 266404
rect 349304 266364 349310 266376
rect 350350 266364 350356 266376
rect 350408 266364 350414 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 359458 266404 359464 266416
rect 357584 266376 359464 266404
rect 357584 266364 357590 266376
rect 359458 266364 359464 266376
rect 359516 266364 359522 266416
rect 361666 266364 361672 266416
rect 361724 266404 361730 266416
rect 362770 266404 362776 266416
rect 361724 266376 362776 266404
rect 361724 266364 361730 266376
rect 362770 266364 362776 266376
rect 362828 266364 362834 266416
rect 369118 266364 369124 266416
rect 369176 266404 369182 266416
rect 370498 266404 370504 266416
rect 369176 266376 370504 266404
rect 369176 266364 369182 266376
rect 370498 266364 370504 266376
rect 370556 266364 370562 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375282 266404 375288 266416
rect 374144 266376 375288 266404
rect 374144 266364 374150 266376
rect 375282 266364 375288 266376
rect 375340 266364 375346 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 383010 266404 383016 266416
rect 379940 266376 383016 266404
rect 379940 266364 379946 266376
rect 383010 266364 383016 266376
rect 383068 266364 383074 266416
rect 384022 266364 384028 266416
rect 384080 266404 384086 266416
rect 384942 266404 384948 266416
rect 384080 266376 384948 266404
rect 384080 266364 384086 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387702 266404 387708 266416
rect 386564 266376 387708 266404
rect 386564 266364 386570 266376
rect 387702 266364 387708 266376
rect 387760 266364 387766 266416
rect 392302 266364 392308 266416
rect 392360 266404 392366 266416
rect 393314 266404 393320 266416
rect 392360 266376 393320 266404
rect 392360 266364 392366 266376
rect 393314 266364 393320 266376
rect 393372 266364 393378 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400030 266404 400036 266416
rect 398984 266376 400036 266404
rect 398984 266364 398990 266376
rect 400030 266364 400036 266376
rect 400088 266364 400094 266416
rect 408862 266364 408868 266416
rect 408920 266404 408926 266416
rect 409782 266404 409788 266416
rect 408920 266376 409788 266404
rect 408920 266364 408926 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412266 266404 412272 266416
rect 411404 266376 412272 266404
rect 411404 266364 411410 266376
rect 412266 266364 412272 266376
rect 412324 266364 412330 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 417970 266364 417976 266416
rect 418028 266404 418034 266416
rect 418798 266404 418804 266416
rect 418028 266376 418804 266404
rect 418028 266364 418034 266376
rect 418798 266364 418804 266376
rect 418856 266364 418862 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 427078 266404 427084 266416
rect 425480 266376 427084 266404
rect 425480 266364 425486 266376
rect 427078 266364 427084 266376
rect 427136 266364 427142 266416
rect 429562 266364 429568 266416
rect 429620 266404 429626 266416
rect 430390 266404 430396 266416
rect 429620 266376 430396 266404
rect 429620 266364 429626 266376
rect 430390 266364 430396 266376
rect 430448 266364 430454 266416
rect 432046 266364 432052 266416
rect 432104 266404 432110 266416
rect 433150 266404 433156 266416
rect 432104 266376 433156 266404
rect 432104 266364 432110 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 440326 266364 440332 266416
rect 440384 266404 440390 266416
rect 441338 266404 441344 266416
rect 440384 266376 441344 266404
rect 440384 266364 440390 266376
rect 441338 266364 441344 266376
rect 441396 266364 441402 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 444466 266364 444472 266416
rect 444524 266404 444530 266416
rect 445662 266404 445668 266416
rect 444524 266376 445668 266404
rect 444524 266364 444530 266376
rect 445662 266364 445668 266376
rect 445720 266364 445726 266416
rect 448606 266364 448612 266416
rect 448664 266404 448670 266416
rect 450538 266404 450544 266416
rect 448664 266376 450544 266404
rect 448664 266364 448670 266376
rect 450538 266364 450544 266376
rect 450596 266364 450602 266416
rect 454402 266364 454408 266416
rect 454460 266404 454466 266416
rect 455322 266404 455328 266416
rect 454460 266376 455328 266404
rect 454460 266364 454466 266376
rect 455322 266364 455328 266376
rect 455380 266364 455386 266416
rect 473446 266364 473452 266416
rect 473504 266404 473510 266416
rect 474642 266404 474648 266416
rect 473504 266376 474648 266404
rect 473504 266364 473510 266376
rect 474642 266364 474648 266376
rect 474700 266364 474706 266416
rect 475102 266364 475108 266416
rect 475160 266404 475166 266416
rect 479518 266404 479524 266416
rect 475160 266376 479524 266404
rect 475160 266364 475166 266376
rect 479518 266364 479524 266376
rect 479576 266364 479582 266416
rect 481726 266364 481732 266416
rect 481784 266404 481790 266416
rect 482830 266404 482836 266416
rect 481784 266376 482836 266404
rect 481784 266364 481790 266376
rect 482830 266364 482836 266376
rect 482888 266364 482894 266416
rect 483382 266364 483388 266416
rect 483440 266404 483446 266416
rect 484210 266404 484216 266416
rect 483440 266376 484216 266404
rect 483440 266364 483446 266376
rect 484210 266364 484216 266376
rect 484268 266364 484274 266416
rect 485866 266364 485872 266416
rect 485924 266404 485930 266416
rect 486786 266404 486792 266416
rect 485924 266376 486792 266404
rect 485924 266364 485930 266376
rect 486786 266364 486792 266376
rect 486844 266364 486850 266416
rect 487154 266296 487160 266348
rect 487212 266336 487218 266348
rect 557718 266336 557724 266348
rect 487212 266308 557724 266336
rect 487212 266296 487218 266308
rect 557718 266296 557724 266308
rect 557776 266296 557782 266348
rect 484210 266160 484216 266212
rect 484268 266200 484274 266212
rect 560662 266200 560668 266212
rect 484268 266172 560668 266200
rect 484268 266160 484274 266172
rect 560662 266160 560668 266172
rect 560720 266160 560726 266212
rect 482554 266024 482560 266076
rect 482612 266064 482618 266076
rect 487154 266064 487160 266076
rect 482612 266036 487160 266064
rect 482612 266024 482618 266036
rect 487154 266024 487160 266036
rect 487212 266024 487218 266076
rect 492490 266024 492496 266076
rect 492548 266064 492554 266076
rect 572714 266064 572720 266076
rect 492548 266036 572720 266064
rect 492548 266024 492554 266036
rect 572714 266024 572720 266036
rect 572772 266024 572778 266076
rect 513190 265888 513196 265940
rect 513248 265928 513254 265940
rect 601694 265928 601700 265940
rect 513248 265900 601700 265928
rect 513248 265888 513254 265900
rect 601694 265888 601700 265900
rect 601752 265888 601758 265940
rect 515674 265752 515680 265804
rect 515732 265792 515738 265804
rect 605834 265792 605840 265804
rect 515732 265764 605840 265792
rect 515732 265752 515738 265764
rect 605834 265752 605840 265764
rect 605892 265752 605898 265804
rect 209774 265616 209780 265668
rect 209832 265656 209838 265668
rect 210694 265656 210700 265668
rect 209832 265628 210700 265656
rect 209832 265616 209838 265628
rect 210694 265616 210700 265628
rect 210752 265616 210758 265668
rect 224954 265616 224960 265668
rect 225012 265656 225018 265668
rect 225598 265656 225604 265668
rect 225012 265628 225604 265656
rect 225012 265616 225018 265628
rect 225598 265616 225604 265628
rect 225656 265616 225662 265668
rect 280338 265616 280344 265668
rect 280396 265656 280402 265668
rect 280982 265656 280988 265668
rect 280396 265628 280988 265656
rect 280396 265616 280402 265628
rect 280982 265616 280988 265628
rect 281040 265616 281046 265668
rect 520642 265616 520648 265668
rect 520700 265656 520706 265668
rect 612734 265656 612740 265668
rect 520700 265628 612740 265656
rect 520700 265616 520706 265628
rect 612734 265616 612740 265628
rect 612792 265616 612798 265668
rect 479242 265480 479248 265532
rect 479300 265520 479306 265532
rect 553394 265520 553400 265532
rect 479300 265492 553400 265520
rect 479300 265480 479306 265492
rect 553394 265480 553400 265492
rect 553452 265480 553458 265532
rect 477586 265344 477592 265396
rect 477644 265384 477650 265396
rect 550634 265384 550640 265396
rect 477644 265356 550640 265384
rect 477644 265344 477650 265356
rect 550634 265344 550640 265356
rect 550692 265344 550698 265396
rect 469306 265208 469312 265260
rect 469364 265248 469370 265260
rect 539962 265248 539968 265260
rect 469364 265220 539968 265248
rect 469364 265208 469370 265220
rect 539962 265208 539968 265220
rect 540020 265208 540026 265260
rect 466822 265072 466828 265124
rect 466880 265112 466886 265124
rect 535730 265112 535736 265124
rect 466880 265084 535736 265112
rect 466880 265072 466886 265084
rect 535730 265072 535736 265084
rect 535788 265072 535794 265124
rect 64138 264460 64144 264512
rect 64196 264500 64202 264512
rect 668946 264500 668952 264512
rect 64196 264472 668952 264500
rect 64196 264460 64202 264472
rect 668946 264460 668952 264472
rect 669004 264460 669010 264512
rect 61378 264324 61384 264376
rect 61436 264364 61442 264376
rect 668118 264364 668124 264376
rect 61436 264336 668124 264364
rect 61436 264324 61442 264336
rect 668118 264324 668124 264336
rect 668176 264324 668182 264376
rect 55858 264188 55864 264240
rect 55916 264228 55922 264240
rect 667934 264228 667940 264240
rect 55916 264200 667940 264228
rect 55916 264188 55922 264200
rect 667934 264188 667940 264200
rect 667992 264188 667998 264240
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 563698 259468 563704 259480
rect 554372 259440 563704 259468
rect 554372 259428 554378 259440
rect 563698 259428 563704 259440
rect 563756 259428 563762 259480
rect 675846 258680 675852 258732
rect 675904 258720 675910 258732
rect 676398 258720 676404 258732
rect 675904 258692 676404 258720
rect 675904 258680 675910 258692
rect 676398 258680 676404 258692
rect 676456 258680 676462 258732
rect 35802 256776 35808 256828
rect 35860 256816 35866 256828
rect 40494 256816 40500 256828
rect 35860 256788 40500 256816
rect 35860 256776 35866 256788
rect 40494 256776 40500 256788
rect 40552 256776 40558 256828
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 560938 256748 560944 256760
rect 554004 256720 560944 256748
rect 554004 256708 554010 256720
rect 560938 256708 560944 256720
rect 560996 256708 561002 256760
rect 35802 255552 35808 255604
rect 35860 255592 35866 255604
rect 35860 255564 38654 255592
rect 35860 255552 35866 255564
rect 38626 255524 38654 255564
rect 554498 255552 554504 255604
rect 554556 255592 554562 255604
rect 558178 255592 558184 255604
rect 554556 255564 558184 255592
rect 554556 255552 554562 255564
rect 558178 255552 558184 255564
rect 558236 255552 558242 255604
rect 39574 255524 39580 255536
rect 38626 255496 39580 255524
rect 39574 255484 39580 255496
rect 39632 255484 39638 255536
rect 35618 255280 35624 255332
rect 35676 255320 35682 255332
rect 39850 255320 39856 255332
rect 35676 255292 39856 255320
rect 35676 255280 35682 255292
rect 39850 255280 39856 255292
rect 39908 255280 39914 255332
rect 35802 254056 35808 254108
rect 35860 254096 35866 254108
rect 40218 254096 40224 254108
rect 35860 254068 40224 254096
rect 35860 254056 35866 254068
rect 40218 254056 40224 254068
rect 40276 254056 40282 254108
rect 35802 252696 35808 252748
rect 35860 252736 35866 252748
rect 41322 252736 41328 252748
rect 35860 252708 41328 252736
rect 35860 252696 35866 252708
rect 41322 252696 41328 252708
rect 41380 252696 41386 252748
rect 35618 252560 35624 252612
rect 35676 252600 35682 252612
rect 41690 252600 41696 252612
rect 35676 252572 41696 252600
rect 35676 252560 35682 252572
rect 41690 252560 41696 252572
rect 41748 252560 41754 252612
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 562318 252600 562324 252612
rect 554464 252572 562324 252600
rect 554464 252560 554470 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 37918 251240 37924 251252
rect 35860 251212 37924 251240
rect 35860 251200 35866 251212
rect 37918 251200 37924 251212
rect 37976 251200 37982 251252
rect 554130 251200 554136 251252
rect 554188 251240 554194 251252
rect 556798 251240 556804 251252
rect 554188 251212 556804 251240
rect 554188 251200 554194 251212
rect 556798 251200 556804 251212
rect 556856 251200 556862 251252
rect 35802 249908 35808 249960
rect 35860 249948 35866 249960
rect 39758 249948 39764 249960
rect 35860 249920 39764 249948
rect 35860 249908 35866 249920
rect 39758 249908 39764 249920
rect 39816 249908 39822 249960
rect 674834 249704 674840 249756
rect 674892 249744 674898 249756
rect 675478 249744 675484 249756
rect 674892 249716 675484 249744
rect 674892 249704 674898 249716
rect 675478 249704 675484 249716
rect 675536 249704 675542 249756
rect 675018 247936 675024 247988
rect 675076 247936 675082 247988
rect 675036 247840 675064 247936
rect 675386 247840 675392 247852
rect 675036 247812 675392 247840
rect 675386 247800 675392 247812
rect 675444 247800 675450 247852
rect 35802 247052 35808 247104
rect 35860 247092 35866 247104
rect 41690 247092 41696 247104
rect 35860 247064 41696 247092
rect 35860 247052 35866 247064
rect 41690 247052 41696 247064
rect 41748 247052 41754 247104
rect 559558 246304 559564 246356
rect 559616 246344 559622 246356
rect 647234 246344 647240 246356
rect 559616 246316 647240 246344
rect 559616 246304 559622 246316
rect 647234 246304 647240 246316
rect 647292 246304 647298 246356
rect 671614 245964 671620 246016
rect 671672 246004 671678 246016
rect 672166 246004 672172 246016
rect 671672 245976 672172 246004
rect 671672 245964 671678 245976
rect 672166 245964 672172 245976
rect 672224 245964 672230 246016
rect 553854 245624 553860 245676
rect 553912 245664 553918 245676
rect 596818 245664 596824 245676
rect 553912 245636 596824 245664
rect 553912 245624 553918 245636
rect 596818 245624 596824 245636
rect 596876 245624 596882 245676
rect 674834 245352 674840 245404
rect 674892 245392 674898 245404
rect 675202 245392 675208 245404
rect 674892 245364 675208 245392
rect 674892 245352 674898 245364
rect 675202 245352 675208 245364
rect 675260 245352 675266 245404
rect 553486 244264 553492 244316
rect 553544 244304 553550 244316
rect 555418 244304 555424 244316
rect 553544 244276 555424 244304
rect 553544 244264 553550 244276
rect 555418 244264 555424 244276
rect 555476 244264 555482 244316
rect 37918 242700 37924 242752
rect 37976 242740 37982 242752
rect 41690 242740 41696 242752
rect 37976 242712 41696 242740
rect 37976 242700 37982 242712
rect 41690 242700 41696 242712
rect 41748 242700 41754 242752
rect 42058 242632 42064 242684
rect 42116 242672 42122 242684
rect 42702 242672 42708 242684
rect 42116 242644 42708 242672
rect 42116 242632 42122 242644
rect 42702 242632 42708 242644
rect 42760 242632 42766 242684
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553670 241476 553676 241528
rect 553728 241516 553734 241528
rect 629938 241516 629944 241528
rect 553728 241488 629944 241516
rect 553728 241476 553734 241488
rect 629938 241476 629944 241488
rect 629996 241476 630002 241528
rect 554498 240116 554504 240168
rect 554556 240156 554562 240168
rect 577498 240156 577504 240168
rect 554556 240128 577504 240156
rect 554556 240116 554562 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 672166 236988 672172 237040
rect 672224 237028 672230 237040
rect 672756 237028 672784 237082
rect 672224 237000 672784 237028
rect 672224 236988 672230 237000
rect 671246 236852 671252 236904
rect 671304 236892 671310 236904
rect 671304 236864 672888 236892
rect 671304 236852 671310 236864
rect 553762 236784 553768 236836
rect 553820 236824 553826 236836
rect 559558 236824 559564 236836
rect 553820 236796 559564 236824
rect 553820 236784 553826 236796
rect 559558 236784 559564 236796
rect 559616 236784 559622 236836
rect 672954 236768 673006 236774
rect 672954 236710 673006 236716
rect 671706 236512 671712 236564
rect 671764 236552 671770 236564
rect 671764 236524 673118 236552
rect 671764 236512 671770 236524
rect 673184 236496 673236 236502
rect 673184 236438 673236 236444
rect 672166 236172 672172 236224
rect 672224 236212 672230 236224
rect 673086 236212 673092 236224
rect 672224 236184 673092 236212
rect 672224 236172 672230 236184
rect 673086 236172 673092 236184
rect 673144 236172 673150 236224
rect 671540 236048 673330 236076
rect 671062 235900 671068 235952
rect 671120 235940 671126 235952
rect 671540 235940 671568 236048
rect 671120 235912 671568 235940
rect 671120 235900 671126 235912
rect 673408 235832 673414 235884
rect 673466 235832 673472 235884
rect 672902 235696 672908 235748
rect 672960 235736 672966 235748
rect 672960 235708 673554 235736
rect 672960 235696 672966 235708
rect 673472 235504 673670 235532
rect 673472 235124 673500 235504
rect 673196 235096 673500 235124
rect 673196 234864 673224 235096
rect 673362 234948 673368 235000
rect 673420 234988 673426 235000
rect 673764 234988 673792 235314
rect 673420 234960 673792 234988
rect 673420 234948 673426 234960
rect 673178 234812 673184 234864
rect 673236 234812 673242 234864
rect 673454 234812 673460 234864
rect 673512 234852 673518 234864
rect 673886 234852 673914 235110
rect 673512 234824 673914 234852
rect 673512 234812 673518 234824
rect 669682 234608 669688 234660
rect 669740 234648 669746 234660
rect 673978 234648 674006 234906
rect 674088 234728 674140 234734
rect 674088 234670 674140 234676
rect 669740 234620 674006 234648
rect 669740 234608 669746 234620
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 670234 234472 670240 234524
rect 670292 234512 670298 234524
rect 670292 234484 674222 234512
rect 670292 234472 670298 234484
rect 671430 234200 671436 234252
rect 671488 234240 671494 234252
rect 674082 234240 674088 234252
rect 671488 234212 674088 234240
rect 671488 234200 671494 234212
rect 674082 234200 674088 234212
rect 674140 234200 674146 234252
rect 652202 233860 652208 233912
rect 652260 233900 652266 233912
rect 670878 233900 670884 233912
rect 652260 233872 670884 233900
rect 652260 233860 652266 233872
rect 670878 233860 670884 233872
rect 670936 233860 670942 233912
rect 675846 233860 675852 233912
rect 675904 233900 675910 233912
rect 678238 233900 678244 233912
rect 675904 233872 678244 233900
rect 675904 233860 675910 233872
rect 678238 233860 678244 233872
rect 678296 233860 678302 233912
rect 672074 233248 672080 233300
rect 672132 233288 672138 233300
rect 673178 233288 673184 233300
rect 672132 233260 673184 233288
rect 672132 233248 672138 233260
rect 673178 233248 673184 233260
rect 673236 233248 673242 233300
rect 673454 233180 673460 233232
rect 673512 233220 673518 233232
rect 673960 233220 673966 233232
rect 673512 233192 673966 233220
rect 673512 233180 673518 233192
rect 673960 233180 673966 233192
rect 674018 233180 674024 233232
rect 670050 232976 670056 233028
rect 670108 233016 670114 233028
rect 672994 233016 673000 233028
rect 670108 232988 673000 233016
rect 670108 232976 670114 232988
rect 672994 232976 673000 232988
rect 673052 232976 673058 233028
rect 670878 232840 670884 232892
rect 670936 232880 670942 232892
rect 672902 232880 672908 232892
rect 670936 232852 672908 232880
rect 670936 232840 670942 232852
rect 672902 232840 672908 232852
rect 672960 232840 672966 232892
rect 663766 232716 666554 232744
rect 663058 232636 663064 232688
rect 663116 232676 663122 232688
rect 663766 232676 663794 232716
rect 663116 232648 663794 232676
rect 666526 232676 666554 232716
rect 674374 232676 674380 232688
rect 666526 232648 674380 232676
rect 663116 232636 663122 232648
rect 674374 232636 674380 232648
rect 674432 232636 674438 232688
rect 675846 232636 675852 232688
rect 675904 232676 675910 232688
rect 683206 232676 683212 232688
rect 675904 232648 683212 232676
rect 675904 232636 675910 232648
rect 683206 232636 683212 232648
rect 683264 232636 683270 232688
rect 660298 232500 660304 232552
rect 660356 232540 660362 232552
rect 674558 232540 674564 232552
rect 660356 232512 674564 232540
rect 660356 232500 660362 232512
rect 674558 232500 674564 232512
rect 674616 232500 674622 232552
rect 676030 232500 676036 232552
rect 676088 232540 676094 232552
rect 683390 232540 683396 232552
rect 676088 232512 683396 232540
rect 676088 232500 676094 232512
rect 683390 232500 683396 232512
rect 683448 232500 683454 232552
rect 156414 231548 156420 231600
rect 156472 231588 156478 231600
rect 162670 231588 162676 231600
rect 156472 231560 162676 231588
rect 156472 231548 156478 231560
rect 162670 231548 162676 231560
rect 162728 231548 162734 231600
rect 135162 231412 135168 231464
rect 135220 231452 135226 231464
rect 137646 231452 137652 231464
rect 135220 231424 137652 231452
rect 135220 231412 135226 231424
rect 137646 231412 137652 231424
rect 137704 231412 137710 231464
rect 155126 231412 155132 231464
rect 155184 231452 155190 231464
rect 156966 231452 156972 231464
rect 155184 231424 156972 231452
rect 155184 231412 155190 231424
rect 156966 231412 156972 231424
rect 157024 231412 157030 231464
rect 157242 231412 157248 231464
rect 157300 231452 157306 231464
rect 161750 231452 161756 231464
rect 157300 231424 161756 231452
rect 157300 231412 157306 231424
rect 161750 231412 161756 231424
rect 161808 231412 161814 231464
rect 662506 231412 662512 231464
rect 662564 231452 662570 231464
rect 674834 231452 674840 231464
rect 662564 231424 674840 231452
rect 662564 231412 662570 231424
rect 674834 231412 674840 231424
rect 674892 231412 674898 231464
rect 46198 231276 46204 231328
rect 46256 231316 46262 231328
rect 668394 231316 668400 231328
rect 46256 231288 668400 231316
rect 46256 231276 46262 231288
rect 668394 231276 668400 231288
rect 668452 231276 668458 231328
rect 92382 231140 92388 231192
rect 92440 231180 92446 231192
rect 170766 231180 170772 231192
rect 92440 231152 170772 231180
rect 92440 231140 92446 231152
rect 170766 231140 170772 231152
rect 170824 231140 170830 231192
rect 665082 231140 665088 231192
rect 665140 231180 665146 231192
rect 665140 231152 675326 231180
rect 665140 231140 665146 231152
rect 128262 231004 128268 231056
rect 128320 231044 128326 231056
rect 195882 231044 195888 231056
rect 128320 231016 195888 231044
rect 128320 231004 128326 231016
rect 195882 231004 195888 231016
rect 195940 231004 195946 231056
rect 673178 230936 673184 230988
rect 673236 230976 673242 230988
rect 673236 230948 675142 230976
rect 673236 230936 673242 230948
rect 118602 230868 118608 230920
rect 118660 230908 118666 230920
rect 188154 230908 188160 230920
rect 118660 230880 188160 230908
rect 118660 230868 118666 230880
rect 188154 230868 188160 230880
rect 188212 230868 188218 230920
rect 674834 230800 674840 230852
rect 674892 230840 674898 230852
rect 674892 230812 674982 230840
rect 674892 230800 674898 230812
rect 94498 230732 94504 230784
rect 94556 230772 94562 230784
rect 171410 230772 171416 230784
rect 94556 230744 171416 230772
rect 94556 230732 94562 230744
rect 171410 230732 171416 230744
rect 171468 230732 171474 230784
rect 104802 230596 104808 230648
rect 104860 230636 104866 230648
rect 179138 230636 179144 230648
rect 104860 230608 179144 230636
rect 104860 230596 104866 230608
rect 179138 230596 179144 230608
rect 179196 230596 179202 230648
rect 194410 230596 194416 230648
rect 194468 230636 194474 230648
rect 196894 230636 196900 230648
rect 194468 230608 196900 230636
rect 194468 230596 194474 230608
rect 196894 230596 196900 230608
rect 196952 230596 196958 230648
rect 665266 230596 665272 230648
rect 665324 230636 665330 230648
rect 665324 230608 674820 230636
rect 665324 230596 665330 230608
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 137646 230460 137652 230512
rect 137704 230500 137710 230512
rect 201034 230500 201040 230512
rect 137704 230472 201040 230500
rect 137704 230460 137710 230472
rect 201034 230460 201040 230472
rect 201092 230460 201098 230512
rect 42426 230392 42432 230444
rect 42484 230432 42490 230444
rect 43254 230432 43260 230444
rect 42484 230404 43260 230432
rect 42484 230392 42490 230404
rect 43254 230392 43260 230404
rect 43312 230392 43318 230444
rect 133782 230392 133788 230444
rect 133840 230432 133846 230444
rect 137462 230432 137468 230444
rect 133840 230404 137468 230432
rect 133840 230392 133846 230404
rect 137462 230392 137468 230404
rect 137520 230392 137526 230444
rect 213086 230392 213092 230444
rect 213144 230432 213150 230444
rect 261570 230432 261576 230444
rect 213144 230404 261576 230432
rect 213144 230392 213150 230404
rect 261570 230392 261576 230404
rect 261628 230392 261634 230444
rect 311986 230392 311992 230444
rect 312044 230432 312050 230444
rect 313090 230432 313096 230444
rect 312044 230404 313096 230432
rect 312044 230392 312050 230404
rect 313090 230392 313096 230404
rect 313148 230392 313154 230444
rect 374638 230392 374644 230444
rect 374696 230432 374702 230444
rect 376202 230432 376208 230444
rect 374696 230404 376208 230432
rect 374696 230392 374702 230404
rect 376202 230392 376208 230404
rect 376260 230392 376266 230444
rect 439516 230432 439544 230540
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 451550 230392 451556 230444
rect 451608 230432 451614 230444
rect 453298 230432 453304 230444
rect 451608 230404 453304 230432
rect 451608 230392 451614 230404
rect 453298 230392 453304 230404
rect 453356 230392 453362 230444
rect 476114 230392 476120 230444
rect 476172 230432 476178 230444
rect 478598 230432 478604 230444
rect 476172 230404 478604 230432
rect 476172 230392 476178 230404
rect 478598 230392 478604 230404
rect 478656 230392 478662 230444
rect 539594 230432 539600 230444
rect 532528 230404 539600 230432
rect 387426 230324 387432 230376
rect 387484 230364 387490 230376
rect 388438 230364 388444 230376
rect 387484 230336 388444 230364
rect 387484 230324 387490 230336
rect 388438 230324 388444 230336
rect 388496 230324 388502 230376
rect 398098 230324 398104 230376
rect 398156 230364 398162 230376
rect 399386 230364 399392 230376
rect 398156 230336 399392 230364
rect 398156 230324 398162 230336
rect 399386 230324 399392 230336
rect 399444 230324 399450 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 470870 230324 470876 230376
rect 470928 230364 470934 230376
rect 471882 230364 471888 230376
rect 470928 230336 471888 230364
rect 470928 230324 470934 230336
rect 471882 230324 471888 230336
rect 471940 230324 471946 230376
rect 493410 230324 493416 230376
rect 493468 230364 493474 230376
rect 496354 230364 496360 230376
rect 493468 230336 496360 230364
rect 493468 230324 493474 230336
rect 496354 230324 496360 230336
rect 496412 230324 496418 230376
rect 497274 230324 497280 230376
rect 497332 230364 497338 230376
rect 498102 230364 498108 230376
rect 497332 230336 498108 230364
rect 497332 230324 497338 230336
rect 498102 230324 498108 230336
rect 498160 230324 498166 230376
rect 510798 230324 510804 230376
rect 510856 230364 510862 230376
rect 511902 230364 511908 230376
rect 510856 230336 511908 230364
rect 510856 230324 510862 230336
rect 511902 230324 511908 230336
rect 511960 230324 511966 230376
rect 521102 230324 521108 230376
rect 521160 230364 521166 230376
rect 526438 230364 526444 230376
rect 521160 230336 526444 230364
rect 521160 230324 521166 230336
rect 526438 230324 526444 230336
rect 526496 230324 526502 230376
rect 530118 230324 530124 230376
rect 530176 230364 530182 230376
rect 531130 230364 531136 230376
rect 530176 230336 531136 230364
rect 530176 230324 530182 230336
rect 531130 230324 531136 230336
rect 531188 230324 531194 230376
rect 126882 230256 126888 230308
rect 126940 230296 126946 230308
rect 194410 230296 194416 230308
rect 126940 230268 194416 230296
rect 126940 230256 126946 230268
rect 194410 230256 194416 230268
rect 194468 230256 194474 230308
rect 194870 230256 194876 230308
rect 194928 230296 194934 230308
rect 195422 230296 195428 230308
rect 194928 230268 195428 230296
rect 194928 230256 194934 230268
rect 195422 230256 195428 230268
rect 195480 230256 195486 230308
rect 195606 230256 195612 230308
rect 195664 230296 195670 230308
rect 204898 230296 204904 230308
rect 195664 230268 204904 230296
rect 195664 230256 195670 230268
rect 204898 230256 204904 230268
rect 204956 230256 204962 230308
rect 206554 230256 206560 230308
rect 206612 230296 206618 230308
rect 256418 230296 256424 230308
rect 206612 230268 256424 230296
rect 206612 230256 206618 230268
rect 256418 230256 256424 230268
rect 256476 230256 256482 230308
rect 256602 230256 256608 230308
rect 256660 230296 256666 230308
rect 297634 230296 297640 230308
rect 256660 230268 297640 230296
rect 256660 230256 256666 230268
rect 297634 230256 297640 230268
rect 297692 230256 297698 230308
rect 297818 230256 297824 230308
rect 297876 230296 297882 230308
rect 323394 230296 323400 230308
rect 297876 230268 323400 230296
rect 297876 230256 297882 230268
rect 323394 230256 323400 230268
rect 323452 230256 323458 230308
rect 452838 230188 452844 230240
rect 452896 230228 452902 230240
rect 454310 230228 454316 230240
rect 452896 230200 454316 230228
rect 452896 230188 452902 230200
rect 454310 230188 454316 230200
rect 454368 230188 454374 230240
rect 468294 230188 468300 230240
rect 468352 230228 468358 230240
rect 469122 230228 469128 230240
rect 468352 230200 469128 230228
rect 468352 230188 468358 230200
rect 469122 230188 469128 230200
rect 469180 230188 469186 230240
rect 487614 230188 487620 230240
rect 487672 230228 487678 230240
rect 488442 230228 488448 230240
rect 487672 230200 488448 230228
rect 487672 230188 487678 230200
rect 488442 230188 488448 230200
rect 488500 230188 488506 230240
rect 495158 230228 495164 230240
rect 489886 230200 495164 230228
rect 95234 230120 95240 230172
rect 95292 230160 95298 230172
rect 157610 230160 157616 230172
rect 95292 230132 157616 230160
rect 95292 230120 95298 230132
rect 157610 230120 157616 230132
rect 157668 230120 157674 230172
rect 157794 230120 157800 230172
rect 157852 230160 157858 230172
rect 158530 230160 158536 230172
rect 157852 230132 158536 230160
rect 157852 230120 157858 230132
rect 158530 230120 158536 230132
rect 158588 230120 158594 230172
rect 162486 230120 162492 230172
rect 162544 230160 162550 230172
rect 185578 230160 185584 230172
rect 162544 230132 185584 230160
rect 162544 230120 162550 230132
rect 185578 230120 185584 230132
rect 185636 230120 185642 230172
rect 186038 230120 186044 230172
rect 186096 230160 186102 230172
rect 235810 230160 235816 230172
rect 186096 230132 235816 230160
rect 186096 230120 186102 230132
rect 235810 230120 235816 230132
rect 235868 230120 235874 230172
rect 240318 230120 240324 230172
rect 240376 230160 240382 230172
rect 282178 230160 282184 230172
rect 240376 230132 282184 230160
rect 240376 230120 240382 230132
rect 282178 230120 282184 230132
rect 282236 230120 282242 230172
rect 282638 230120 282644 230172
rect 282696 230160 282702 230172
rect 307938 230160 307944 230172
rect 282696 230132 307944 230160
rect 282696 230120 282702 230132
rect 307938 230120 307944 230132
rect 307996 230120 308002 230172
rect 308122 230120 308128 230172
rect 308180 230160 308186 230172
rect 334986 230160 334992 230172
rect 308180 230132 334992 230160
rect 308180 230120 308186 230132
rect 334986 230120 334992 230132
rect 335044 230120 335050 230172
rect 335170 230120 335176 230172
rect 335228 230160 335234 230172
rect 350442 230160 350448 230172
rect 335228 230132 350448 230160
rect 335228 230120 335234 230132
rect 350442 230120 350448 230132
rect 350500 230120 350506 230172
rect 444466 230120 444472 230172
rect 444524 230160 444530 230172
rect 447686 230160 447692 230172
rect 444524 230132 447692 230160
rect 444524 230120 444530 230132
rect 447686 230120 447692 230132
rect 447744 230120 447750 230172
rect 454126 230052 454132 230104
rect 454184 230092 454190 230104
rect 455322 230092 455328 230104
rect 454184 230064 455328 230092
rect 454184 230052 454190 230064
rect 455322 230052 455328 230064
rect 455380 230052 455386 230104
rect 82078 229984 82084 230036
rect 82136 230024 82142 230036
rect 82136 229996 84194 230024
rect 82136 229984 82142 229996
rect 84166 229888 84194 229996
rect 86218 229984 86224 230036
rect 86276 230024 86282 230036
rect 137278 230024 137284 230036
rect 86276 229996 137284 230024
rect 86276 229984 86282 229996
rect 137278 229984 137284 229996
rect 137336 229984 137342 230036
rect 137462 229984 137468 230036
rect 137520 230024 137526 230036
rect 156782 230024 156788 230036
rect 137520 229996 156788 230024
rect 137520 229984 137526 229996
rect 156782 229984 156788 229996
rect 156840 229984 156846 230036
rect 157426 229984 157432 230036
rect 157484 230024 157490 230036
rect 195054 230024 195060 230036
rect 157484 229996 195060 230024
rect 157484 229984 157490 229996
rect 195054 229984 195060 229996
rect 195112 229984 195118 230036
rect 195422 229984 195428 230036
rect 195480 230024 195486 230036
rect 215202 230024 215208 230036
rect 195480 229996 215208 230024
rect 195480 229984 195486 229996
rect 215202 229984 215208 229996
rect 215260 229984 215266 230036
rect 230474 229984 230480 230036
rect 230532 230024 230538 230036
rect 277026 230024 277032 230036
rect 230532 229996 277032 230024
rect 230532 229984 230538 229996
rect 277026 229984 277032 229996
rect 277084 229984 277090 230036
rect 277210 229984 277216 230036
rect 277268 230024 277274 230036
rect 302786 230024 302792 230036
rect 277268 229996 302792 230024
rect 277268 229984 277274 229996
rect 302786 229984 302792 229996
rect 302844 229984 302850 230036
rect 303246 229984 303252 230036
rect 303304 230024 303310 230036
rect 329834 230024 329840 230036
rect 303304 229996 329840 230024
rect 303304 229984 303310 229996
rect 329834 229984 329840 229996
rect 329892 229984 329898 230036
rect 330938 229984 330944 230036
rect 330996 230024 331002 230036
rect 355594 230024 355600 230036
rect 330996 229996 355600 230024
rect 330996 229984 331002 229996
rect 355594 229984 355600 229996
rect 355652 229984 355658 230036
rect 484394 229984 484400 230036
rect 484452 230024 484458 230036
rect 489886 230024 489914 230200
rect 495158 230188 495164 230200
rect 495216 230188 495222 230240
rect 511442 230188 511448 230240
rect 511500 230228 511506 230240
rect 517514 230228 517520 230240
rect 511500 230200 517520 230228
rect 511500 230188 511506 230200
rect 517514 230188 517520 230200
rect 517572 230188 517578 230240
rect 530762 230188 530768 230240
rect 530820 230228 530826 230240
rect 532528 230228 532556 230404
rect 539594 230392 539600 230404
rect 539652 230392 539658 230444
rect 674676 230308 674728 230314
rect 533522 230256 533528 230308
rect 533580 230296 533586 230308
rect 538306 230296 538312 230308
rect 533580 230268 538312 230296
rect 533580 230256 533586 230268
rect 538306 230256 538312 230268
rect 538364 230256 538370 230308
rect 674676 230250 674728 230256
rect 530820 230200 532556 230228
rect 530820 230188 530826 230200
rect 673454 230188 673460 230240
rect 673512 230228 673518 230240
rect 673512 230200 674590 230228
rect 673512 230188 673518 230200
rect 532694 230120 532700 230172
rect 532752 230160 532758 230172
rect 547138 230160 547144 230172
rect 532752 230132 547144 230160
rect 532752 230120 532758 230132
rect 547138 230120 547144 230132
rect 547196 230120 547202 230172
rect 491478 230052 491484 230104
rect 491536 230092 491542 230104
rect 492490 230092 492496 230104
rect 491536 230064 492496 230092
rect 491536 230052 491542 230064
rect 492490 230052 492496 230064
rect 492548 230052 492554 230104
rect 560938 230052 560944 230104
rect 560996 230092 561002 230104
rect 568114 230092 568120 230104
rect 560996 230064 568120 230092
rect 560996 230052 561002 230064
rect 568114 230052 568120 230064
rect 568172 230052 568178 230104
rect 484452 229996 489914 230024
rect 484452 229984 484458 229996
rect 517238 229984 517244 230036
rect 517296 230024 517302 230036
rect 524598 230024 524604 230036
rect 517296 229996 524604 230024
rect 517296 229984 517302 229996
rect 524598 229984 524604 229996
rect 524656 229984 524662 230036
rect 528830 229984 528836 230036
rect 528888 230024 528894 230036
rect 533522 230024 533528 230036
rect 528888 229996 533528 230024
rect 528888 229984 528894 229996
rect 533522 229984 533528 229996
rect 533580 229984 533586 230036
rect 534626 229984 534632 230036
rect 534684 230024 534690 230036
rect 549254 230024 549260 230036
rect 534684 229996 549260 230024
rect 534684 229984 534690 229996
rect 549254 229984 549260 229996
rect 549312 229984 549318 230036
rect 674452 229968 674504 229974
rect 453482 229916 453488 229968
rect 453540 229956 453546 229968
rect 455782 229956 455788 229968
rect 453540 229928 455788 229956
rect 453540 229916 453546 229928
rect 455782 229916 455788 229928
rect 455840 229916 455846 229968
rect 674452 229910 674504 229916
rect 151446 229888 151452 229900
rect 84166 229860 151452 229888
rect 151446 229848 151452 229860
rect 151504 229848 151510 229900
rect 151630 229848 151636 229900
rect 151688 229888 151694 229900
rect 157242 229888 157248 229900
rect 151688 229860 157248 229888
rect 151688 229848 151694 229860
rect 157242 229848 157248 229860
rect 157300 229848 157306 229900
rect 162302 229848 162308 229900
rect 162360 229888 162366 229900
rect 166258 229888 166264 229900
rect 162360 229860 166264 229888
rect 162360 229848 162366 229860
rect 166258 229848 166264 229860
rect 166316 229848 166322 229900
rect 225506 229888 225512 229900
rect 171106 229860 225512 229888
rect 68278 229712 68284 229764
rect 68336 229752 68342 229764
rect 144454 229752 144460 229764
rect 68336 229724 144460 229752
rect 68336 229712 68342 229724
rect 144454 229712 144460 229724
rect 144512 229712 144518 229764
rect 144822 229712 144828 229764
rect 144880 229752 144886 229764
rect 146294 229752 146300 229764
rect 144880 229724 146300 229752
rect 144880 229712 144886 229724
rect 146294 229712 146300 229724
rect 146352 229712 146358 229764
rect 156782 229752 156788 229764
rect 146956 229724 156788 229752
rect 137278 229576 137284 229628
rect 137336 229616 137342 229628
rect 146956 229616 146984 229724
rect 156782 229712 156788 229724
rect 156840 229712 156846 229764
rect 162118 229752 162124 229764
rect 157812 229724 162124 229752
rect 137336 229588 146984 229616
rect 137336 229576 137342 229588
rect 148134 229576 148140 229628
rect 148192 229616 148198 229628
rect 150802 229616 150808 229628
rect 148192 229588 150808 229616
rect 148192 229576 148198 229588
rect 150802 229576 150808 229588
rect 150860 229576 150866 229628
rect 150986 229576 150992 229628
rect 151044 229616 151050 229628
rect 153378 229616 153384 229628
rect 151044 229588 153384 229616
rect 151044 229576 151050 229588
rect 153378 229576 153384 229588
rect 153436 229576 153442 229628
rect 154390 229576 154396 229628
rect 154448 229616 154454 229628
rect 157812 229616 157840 229724
rect 162118 229712 162124 229724
rect 162176 229712 162182 229764
rect 163958 229712 163964 229764
rect 164016 229752 164022 229764
rect 171106 229752 171134 229860
rect 225506 229848 225512 229860
rect 225564 229848 225570 229900
rect 225690 229848 225696 229900
rect 225748 229888 225754 229900
rect 271874 229888 271880 229900
rect 225748 229860 271880 229888
rect 225748 229848 225754 229860
rect 271874 229848 271880 229860
rect 271932 229848 271938 229900
rect 275646 229848 275652 229900
rect 275704 229888 275710 229900
rect 311986 229888 311992 229900
rect 275704 229860 311992 229888
rect 275704 229848 275710 229860
rect 311986 229848 311992 229860
rect 312044 229848 312050 229900
rect 312630 229848 312636 229900
rect 312688 229888 312694 229900
rect 340138 229888 340144 229900
rect 312688 229860 340144 229888
rect 312688 229848 312694 229860
rect 340138 229848 340144 229860
rect 340196 229848 340202 229900
rect 345658 229848 345664 229900
rect 345716 229888 345722 229900
rect 360746 229888 360752 229900
rect 345716 229860 360752 229888
rect 345716 229848 345722 229860
rect 360746 229848 360752 229860
rect 360804 229848 360810 229900
rect 361206 229848 361212 229900
rect 361264 229888 361270 229900
rect 378778 229888 378784 229900
rect 361264 229860 378784 229888
rect 361264 229848 361270 229860
rect 378778 229848 378784 229860
rect 378836 229848 378842 229900
rect 410886 229848 410892 229900
rect 410944 229888 410950 229900
rect 417418 229888 417424 229900
rect 410944 229860 417424 229888
rect 410944 229848 410950 229860
rect 417418 229848 417424 229860
rect 417476 229848 417482 229900
rect 449618 229848 449624 229900
rect 449676 229888 449682 229900
rect 450538 229888 450544 229900
rect 449676 229860 450544 229888
rect 449676 229848 449682 229860
rect 450538 229848 450544 229860
rect 450596 229848 450602 229900
rect 467006 229848 467012 229900
rect 467064 229888 467070 229900
rect 473998 229888 474004 229900
rect 467064 229860 474004 229888
rect 467064 229848 467070 229860
rect 473998 229848 474004 229860
rect 474056 229848 474062 229900
rect 476666 229848 476672 229900
rect 476724 229888 476730 229900
rect 481634 229888 481640 229900
rect 476724 229860 481640 229888
rect 476724 229848 476730 229860
rect 481634 229848 481640 229860
rect 481692 229848 481698 229900
rect 481818 229848 481824 229900
rect 481876 229888 481882 229900
rect 493686 229888 493692 229900
rect 481876 229860 493692 229888
rect 481876 229848 481882 229860
rect 493686 229848 493692 229860
rect 493744 229848 493750 229900
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 506382 229888 506388 229900
rect 496044 229860 506388 229888
rect 496044 229848 496050 229860
rect 506382 229848 506388 229860
rect 506440 229848 506446 229900
rect 507578 229848 507584 229900
rect 507636 229888 507642 229900
rect 516778 229888 516784 229900
rect 507636 229860 516784 229888
rect 507636 229848 507642 229860
rect 516778 229848 516784 229860
rect 516836 229848 516842 229900
rect 519170 229848 519176 229900
rect 519228 229888 519234 229900
rect 528554 229888 528560 229900
rect 519228 229860 528560 229888
rect 519228 229848 519234 229860
rect 528554 229848 528560 229860
rect 528612 229848 528618 229900
rect 536558 229848 536564 229900
rect 536616 229888 536622 229900
rect 559558 229888 559564 229900
rect 536616 229860 559564 229888
rect 536616 229848 536622 229860
rect 559558 229848 559564 229860
rect 559616 229848 559622 229900
rect 668578 229848 668584 229900
rect 668636 229888 668642 229900
rect 672718 229888 672724 229900
rect 668636 229860 672724 229888
rect 668636 229848 668642 229860
rect 672718 229848 672724 229860
rect 672776 229848 672782 229900
rect 674334 229832 674386 229838
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 674334 229774 674386 229780
rect 164016 229724 171134 229752
rect 164016 229712 164022 229724
rect 173894 229712 173900 229764
rect 173952 229752 173958 229764
rect 175918 229752 175924 229764
rect 173952 229724 175924 229752
rect 173952 229712 173958 229724
rect 175918 229712 175924 229724
rect 175976 229712 175982 229764
rect 176378 229712 176384 229764
rect 176436 229752 176442 229764
rect 185394 229752 185400 229764
rect 176436 229724 185400 229752
rect 176436 229712 176442 229724
rect 185394 229712 185400 229724
rect 185452 229712 185458 229764
rect 185578 229712 185584 229764
rect 185636 229752 185642 229764
rect 194870 229752 194876 229764
rect 185636 229724 194876 229752
rect 185636 229712 185642 229724
rect 194870 229712 194876 229724
rect 194928 229712 194934 229764
rect 195054 229712 195060 229764
rect 195112 229752 195118 229764
rect 202322 229752 202328 229764
rect 195112 229724 202328 229752
rect 195112 229712 195118 229724
rect 202322 229712 202328 229724
rect 202380 229712 202386 229764
rect 204898 229712 204904 229764
rect 204956 229752 204962 229764
rect 246114 229752 246120 229764
rect 204956 229724 246120 229752
rect 204956 229712 204962 229724
rect 246114 229712 246120 229724
rect 246172 229712 246178 229764
rect 246482 229712 246488 229764
rect 246540 229752 246546 229764
rect 287330 229752 287336 229764
rect 246540 229724 287336 229752
rect 246540 229712 246546 229724
rect 287330 229712 287336 229724
rect 287388 229712 287394 229764
rect 287698 229712 287704 229764
rect 287756 229752 287762 229764
rect 318242 229752 318248 229764
rect 287756 229724 318248 229752
rect 287756 229712 287762 229724
rect 318242 229712 318248 229724
rect 318300 229712 318306 229764
rect 345290 229752 345296 229764
rect 325666 229724 345296 229752
rect 154448 229588 157840 229616
rect 154448 229576 154454 229588
rect 157978 229576 157984 229628
rect 158036 229616 158042 229628
rect 160738 229616 160744 229628
rect 158036 229588 160744 229616
rect 158036 229576 158042 229588
rect 160738 229576 160744 229588
rect 160796 229576 160802 229628
rect 160922 229576 160928 229628
rect 160980 229616 160986 229628
rect 220354 229616 220360 229628
rect 160980 229588 220360 229616
rect 160980 229576 160986 229588
rect 220354 229576 220360 229588
rect 220412 229576 220418 229628
rect 251266 229616 251272 229628
rect 229066 229588 251272 229616
rect 147048 229520 147812 229548
rect 102134 229440 102140 229492
rect 102192 229480 102198 229492
rect 145650 229480 145656 229492
rect 102192 229452 145656 229480
rect 102192 229440 102198 229452
rect 145650 229440 145656 229452
rect 145708 229440 145714 229492
rect 146018 229372 146024 229424
rect 146076 229412 146082 229424
rect 147048 229412 147076 229520
rect 147784 229480 147812 229520
rect 210050 229480 210056 229492
rect 147784 229452 210056 229480
rect 210050 229440 210056 229452
rect 210108 229440 210114 229492
rect 220078 229440 220084 229492
rect 220136 229480 220142 229492
rect 229066 229480 229094 229588
rect 251266 229576 251272 229588
rect 251324 229576 251330 229628
rect 251726 229576 251732 229628
rect 251784 229616 251790 229628
rect 292482 229616 292488 229628
rect 251784 229588 292488 229616
rect 251784 229576 251790 229588
rect 292482 229576 292488 229588
rect 292540 229576 292546 229628
rect 318058 229576 318064 229628
rect 318116 229616 318122 229628
rect 325666 229616 325694 229724
rect 345290 229712 345296 229724
rect 345348 229712 345354 229764
rect 351730 229712 351736 229764
rect 351788 229752 351794 229764
rect 371050 229752 371056 229764
rect 351788 229724 371056 229752
rect 351788 229712 351794 229724
rect 371050 229712 371056 229724
rect 371108 229712 371114 229764
rect 377674 229712 377680 229764
rect 377732 229752 377738 229764
rect 389082 229752 389088 229764
rect 377732 229724 389088 229752
rect 377732 229712 377738 229724
rect 389082 229712 389088 229724
rect 389140 229712 389146 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 457346 229712 457352 229764
rect 457404 229752 457410 229764
rect 463878 229752 463884 229764
rect 457404 229724 463884 229752
rect 457404 229712 457410 229724
rect 463878 229712 463884 229724
rect 463936 229712 463942 229764
rect 465442 229712 465448 229764
rect 465500 229752 465506 229764
rect 467466 229752 467472 229764
rect 465500 229724 467472 229752
rect 465500 229712 465506 229724
rect 467466 229712 467472 229724
rect 467524 229712 467530 229764
rect 469582 229712 469588 229764
rect 469640 229752 469646 229764
rect 476758 229752 476764 229764
rect 469640 229724 476764 229752
rect 469640 229712 469646 229724
rect 476758 229712 476764 229724
rect 476816 229712 476822 229764
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 489914 229752 489920 229764
rect 479300 229724 489920 229752
rect 479300 229712 479306 229724
rect 489914 229712 489920 229724
rect 489972 229712 489978 229764
rect 492122 229712 492128 229764
rect 492180 229752 492186 229764
rect 507118 229752 507124 229764
rect 492180 229724 507124 229752
rect 492180 229712 492186 229724
rect 507118 229712 507124 229724
rect 507176 229712 507182 229764
rect 523034 229712 523040 229764
rect 523092 229752 523098 229764
rect 534810 229752 534816 229764
rect 523092 229724 534816 229752
rect 523092 229712 523098 229724
rect 534810 229712 534816 229724
rect 534868 229712 534874 229764
rect 538490 229712 538496 229764
rect 538548 229752 538554 229764
rect 566826 229752 566832 229764
rect 538548 229724 566832 229752
rect 538548 229712 538554 229724
rect 566826 229712 566832 229724
rect 566884 229712 566890 229764
rect 662322 229712 662328 229764
rect 662380 229752 662386 229764
rect 673178 229752 673184 229764
rect 662380 229724 673184 229752
rect 662380 229712 662386 229724
rect 673178 229712 673184 229724
rect 673236 229712 673242 229764
rect 509510 229644 509516 229696
rect 509568 229684 509574 229696
rect 515490 229684 515496 229696
rect 509568 229656 515496 229684
rect 509568 229644 509574 229656
rect 515490 229644 515496 229656
rect 515548 229644 515554 229696
rect 318116 229588 325694 229616
rect 318116 229576 318122 229588
rect 388622 229576 388628 229628
rect 388680 229616 388686 229628
rect 398742 229616 398748 229628
rect 388680 229588 398748 229616
rect 388680 229576 388686 229588
rect 398742 229576 398748 229588
rect 398800 229576 398806 229628
rect 526898 229576 526904 229628
rect 526956 229616 526962 229628
rect 536098 229616 536104 229628
rect 526956 229588 536104 229616
rect 526956 229576 526962 229588
rect 536098 229576 536104 229588
rect 536156 229576 536162 229628
rect 672810 229576 672816 229628
rect 672868 229616 672874 229628
rect 672868 229588 674268 229616
rect 672868 229576 672874 229588
rect 448974 229508 448980 229560
rect 449032 229548 449038 229560
rect 451918 229548 451924 229560
rect 449032 229520 451924 229548
rect 449032 229508 449038 229520
rect 451918 229508 451924 229520
rect 451976 229508 451982 229560
rect 220136 229452 229094 229480
rect 220136 229440 220142 229452
rect 660942 229440 660948 229492
rect 661000 229480 661006 229492
rect 662506 229480 662512 229492
rect 661000 229452 662512 229480
rect 661000 229440 661006 229452
rect 662506 229440 662512 229452
rect 662564 229440 662570 229492
rect 146076 229384 147076 229412
rect 146076 229372 146082 229384
rect 446398 229372 446404 229424
rect 446456 229412 446462 229424
rect 448974 229412 448980 229424
rect 446456 229384 448980 229412
rect 446456 229372 446462 229384
rect 448974 229372 448980 229384
rect 449032 229372 449038 229424
rect 505646 229372 505652 229424
rect 505704 229412 505710 229424
rect 510614 229412 510620 229424
rect 505704 229384 510620 229412
rect 505704 229372 505710 229384
rect 510614 229372 510620 229384
rect 510672 229372 510678 229424
rect 673270 229372 673276 229424
rect 673328 229412 673334 229424
rect 673328 229384 674130 229412
rect 673328 229372 673334 229384
rect 110322 229304 110328 229356
rect 110380 229344 110386 229356
rect 145834 229344 145840 229356
rect 110380 229316 145840 229344
rect 110380 229304 110386 229316
rect 145834 229304 145840 229316
rect 145892 229304 145898 229356
rect 151446 229304 151452 229356
rect 151504 229344 151510 229356
rect 155954 229344 155960 229356
rect 151504 229316 155960 229344
rect 151504 229304 151510 229316
rect 155954 229304 155960 229316
rect 156012 229304 156018 229356
rect 157794 229344 157800 229356
rect 156156 229316 157800 229344
rect 123478 229168 123484 229220
rect 123536 229208 123542 229220
rect 148134 229208 148140 229220
rect 123536 229180 148140 229208
rect 123536 229168 123542 229180
rect 148134 229168 148140 229180
rect 148192 229168 148198 229220
rect 148318 229168 148324 229220
rect 148376 229208 148382 229220
rect 154022 229208 154028 229220
rect 148376 229180 154028 229208
rect 148376 229168 148382 229180
rect 154022 229168 154028 229180
rect 154080 229168 154086 229220
rect 154206 229168 154212 229220
rect 154264 229208 154270 229220
rect 156156 229208 156184 229316
rect 157794 229304 157800 229316
rect 157852 229304 157858 229356
rect 157978 229304 157984 229356
rect 158036 229344 158042 229356
rect 163682 229344 163688 229356
rect 158036 229316 163688 229344
rect 158036 229304 158042 229316
rect 163682 229304 163688 229316
rect 163740 229304 163746 229356
rect 166810 229304 166816 229356
rect 166868 229344 166874 229356
rect 169110 229344 169116 229356
rect 166868 229316 169116 229344
rect 166868 229304 166874 229316
rect 169110 229304 169116 229316
rect 169168 229304 169174 229356
rect 170950 229304 170956 229356
rect 171008 229344 171014 229356
rect 230658 229344 230664 229356
rect 171008 229316 230664 229344
rect 171008 229304 171014 229316
rect 230658 229304 230664 229316
rect 230716 229304 230722 229356
rect 413830 229304 413836 229356
rect 413888 229344 413894 229356
rect 419994 229344 420000 229356
rect 413888 229316 420000 229344
rect 413888 229304 413894 229316
rect 419994 229304 420000 229316
rect 420052 229304 420058 229356
rect 443822 229304 443828 229356
rect 443880 229344 443886 229356
rect 444834 229344 444840 229356
rect 443880 229316 444840 229344
rect 443880 229304 443886 229316
rect 444834 229304 444840 229316
rect 444892 229304 444898 229356
rect 472158 229304 472164 229356
rect 472216 229344 472222 229356
rect 472986 229344 472992 229356
rect 472216 229316 472992 229344
rect 472216 229304 472222 229316
rect 472986 229304 472992 229316
rect 473044 229304 473050 229356
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451734 229276 451740 229288
rect 450320 229248 451740 229276
rect 450320 229236 450326 229248
rect 451734 229236 451740 229248
rect 451792 229236 451798 229288
rect 495342 229236 495348 229288
rect 495400 229276 495406 229288
rect 500218 229276 500224 229288
rect 495400 229248 500224 229276
rect 495400 229236 495406 229248
rect 500218 229236 500224 229248
rect 500276 229236 500282 229288
rect 513374 229236 513380 229288
rect 513432 229276 513438 229288
rect 519078 229276 519084 229288
rect 513432 229248 519084 229276
rect 513432 229236 513438 229248
rect 519078 229236 519084 229248
rect 519136 229236 519142 229288
rect 154264 229180 156184 229208
rect 154264 229168 154270 229180
rect 162118 229168 162124 229220
rect 162176 229208 162182 229220
rect 173894 229208 173900 229220
rect 162176 229180 173900 229208
rect 162176 229168 162182 229180
rect 173894 229168 173900 229180
rect 173952 229168 173958 229220
rect 174096 229180 174860 229208
rect 106182 229032 106188 229084
rect 106240 229072 106246 229084
rect 174096 229072 174124 229180
rect 106240 229044 174124 229072
rect 174832 229072 174860 229180
rect 175918 229168 175924 229220
rect 175976 229208 175982 229220
rect 180426 229208 180432 229220
rect 175976 229180 180432 229208
rect 175976 229168 175982 229180
rect 180426 229168 180432 229180
rect 180484 229168 180490 229220
rect 183370 229168 183376 229220
rect 183428 229208 183434 229220
rect 240962 229208 240968 229220
rect 183428 229180 240968 229208
rect 183428 229168 183434 229180
rect 240962 229168 240968 229180
rect 241020 229168 241026 229220
rect 423490 229100 423496 229152
rect 423548 229140 423554 229152
rect 427722 229140 427728 229152
rect 423548 229112 427728 229140
rect 423548 229100 423554 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 450906 229100 450912 229152
rect 450964 229140 450970 229152
rect 452746 229140 452752 229152
rect 450964 229112 452752 229140
rect 450964 229100 450970 229112
rect 452746 229100 452752 229112
rect 452804 229100 452810 229152
rect 503714 229100 503720 229152
rect 503772 229140 503778 229152
rect 509878 229140 509884 229152
rect 503772 229112 509884 229140
rect 503772 229100 503778 229112
rect 509878 229100 509884 229112
rect 509936 229100 509942 229152
rect 515306 229100 515312 229152
rect 515364 229140 515370 229152
rect 520918 229140 520924 229152
rect 515364 229112 520924 229140
rect 515364 229100 515370 229112
rect 520918 229100 520924 229112
rect 520976 229100 520982 229152
rect 524966 229100 524972 229152
rect 525024 229140 525030 229152
rect 529934 229140 529940 229152
rect 525024 229112 529940 229140
rect 525024 229100 525030 229112
rect 529934 229100 529940 229112
rect 529992 229100 529998 229152
rect 673564 229112 674038 229140
rect 179782 229072 179788 229084
rect 174832 229044 179788 229072
rect 106240 229032 106246 229044
rect 179782 229032 179788 229044
rect 179840 229032 179846 229084
rect 180058 229032 180064 229084
rect 180116 229072 180122 229084
rect 185578 229072 185584 229084
rect 180116 229044 185584 229072
rect 180116 229032 180122 229044
rect 185578 229032 185584 229044
rect 185636 229032 185642 229084
rect 189718 229032 189724 229084
rect 189776 229072 189782 229084
rect 189776 229044 190454 229072
rect 189776 229032 189782 229044
rect 100662 228896 100668 228948
rect 100720 228936 100726 228948
rect 174630 228936 174636 228948
rect 100720 228908 174636 228936
rect 100720 228896 100726 228908
rect 174630 228896 174636 228908
rect 174688 228896 174694 228948
rect 184842 228936 184848 228948
rect 175936 228908 184848 228936
rect 93578 228760 93584 228812
rect 93636 228800 93642 228812
rect 159358 228800 159364 228812
rect 93636 228772 159364 228800
rect 93636 228760 93642 228772
rect 159358 228760 159364 228772
rect 159416 228760 159422 228812
rect 162670 228760 162676 228812
rect 162728 228800 162734 228812
rect 175936 228800 175964 228908
rect 184842 228896 184848 228908
rect 184900 228896 184906 228948
rect 185210 228896 185216 228948
rect 185268 228936 185274 228948
rect 190086 228936 190092 228948
rect 185268 228908 190092 228936
rect 185268 228896 185274 228908
rect 190086 228896 190092 228908
rect 190144 228896 190150 228948
rect 190426 228936 190454 229044
rect 192478 229032 192484 229084
rect 192536 229072 192542 229084
rect 200390 229072 200396 229084
rect 192536 229044 200396 229072
rect 192536 229032 192542 229044
rect 200390 229032 200396 229044
rect 200448 229032 200454 229084
rect 201402 229032 201408 229084
rect 201460 229072 201466 229084
rect 252554 229072 252560 229084
rect 201460 229044 252560 229072
rect 201460 229032 201466 229044
rect 252554 229032 252560 229044
rect 252612 229032 252618 229084
rect 257522 229032 257528 229084
rect 257580 229072 257586 229084
rect 296346 229072 296352 229084
rect 257580 229044 296352 229072
rect 257580 229032 257586 229044
rect 296346 229032 296352 229044
rect 296404 229032 296410 229084
rect 305546 229032 305552 229084
rect 305604 229072 305610 229084
rect 315666 229072 315672 229084
rect 305604 229044 315672 229072
rect 305604 229032 305610 229044
rect 315666 229032 315672 229044
rect 315724 229032 315730 229084
rect 326890 229032 326896 229084
rect 326948 229072 326954 229084
rect 351086 229072 351092 229084
rect 326948 229044 351092 229072
rect 326948 229032 326954 229044
rect 351086 229032 351092 229044
rect 351144 229032 351150 229084
rect 195238 228936 195244 228948
rect 190426 228908 195244 228936
rect 195238 228896 195244 228908
rect 195296 228896 195302 228948
rect 195422 228896 195428 228948
rect 195480 228936 195486 228948
rect 246758 228936 246764 228948
rect 195480 228908 246764 228936
rect 195480 228896 195486 228908
rect 246758 228896 246764 228908
rect 246816 228896 246822 228948
rect 253842 228936 253848 228948
rect 246960 228908 253848 228936
rect 162728 228772 175964 228800
rect 162728 228760 162734 228772
rect 176102 228760 176108 228812
rect 176160 228800 176166 228812
rect 231302 228800 231308 228812
rect 176160 228772 231308 228800
rect 176160 228760 176166 228772
rect 231302 228760 231308 228772
rect 231360 228760 231366 228812
rect 246298 228760 246304 228812
rect 246356 228800 246362 228812
rect 246960 228800 246988 228908
rect 253842 228896 253848 228908
rect 253900 228896 253906 228948
rect 255222 228896 255228 228948
rect 255280 228936 255286 228948
rect 295702 228936 295708 228948
rect 255280 228908 295708 228936
rect 255280 228896 255286 228908
rect 295702 228896 295708 228908
rect 295760 228896 295766 228948
rect 302142 228896 302148 228948
rect 302200 228936 302206 228948
rect 331214 228936 331220 228948
rect 302200 228908 331220 228936
rect 302200 228896 302206 228908
rect 331214 228896 331220 228908
rect 331272 228896 331278 228948
rect 506382 228896 506388 228948
rect 506440 228936 506446 228948
rect 512730 228936 512736 228948
rect 506440 228908 512736 228936
rect 506440 228896 506446 228908
rect 512730 228896 512736 228908
rect 512788 228896 512794 228948
rect 526438 228896 526444 228948
rect 526496 228936 526502 228948
rect 544286 228936 544292 228948
rect 526496 228908 544292 228936
rect 526496 228896 526502 228908
rect 544286 228896 544292 228908
rect 544344 228896 544350 228948
rect 246356 228772 246988 228800
rect 246356 228760 246362 228772
rect 248230 228760 248236 228812
rect 248288 228800 248294 228812
rect 291838 228800 291844 228812
rect 248288 228772 291844 228800
rect 248288 228760 248294 228772
rect 291838 228760 291844 228772
rect 291896 228760 291902 228812
rect 300210 228800 300216 228812
rect 292132 228772 300216 228800
rect 67542 228624 67548 228676
rect 67600 228664 67606 228676
rect 146202 228664 146208 228676
rect 67600 228636 146208 228664
rect 67600 228624 67606 228636
rect 146202 228624 146208 228636
rect 146260 228624 146266 228676
rect 162302 228664 162308 228676
rect 146956 228636 162308 228664
rect 61378 228488 61384 228540
rect 61436 228528 61442 228540
rect 61436 228500 137232 228528
rect 61436 228488 61442 228500
rect 57238 228352 57244 228404
rect 57296 228392 57302 228404
rect 136818 228392 136824 228404
rect 57296 228364 136824 228392
rect 57296 228352 57302 228364
rect 136818 228352 136824 228364
rect 136876 228352 136882 228404
rect 137204 228392 137232 228500
rect 137370 228488 137376 228540
rect 137428 228528 137434 228540
rect 146956 228528 146984 228636
rect 162302 228624 162308 228636
rect 162360 228624 162366 228676
rect 162486 228624 162492 228676
rect 162544 228664 162550 228676
rect 166810 228664 166816 228676
rect 162544 228636 166816 228664
rect 162544 228624 162550 228636
rect 166810 228624 166816 228636
rect 166868 228624 166874 228676
rect 166948 228624 166954 228676
rect 167006 228664 167012 228676
rect 185394 228664 185400 228676
rect 167006 228636 185400 228664
rect 167006 228624 167012 228636
rect 185394 228624 185400 228636
rect 185452 228624 185458 228676
rect 185578 228624 185584 228676
rect 185636 228664 185642 228676
rect 226150 228664 226156 228676
rect 185636 228636 226156 228664
rect 185636 228624 185642 228636
rect 226150 228624 226156 228636
rect 226208 228624 226214 228676
rect 226334 228624 226340 228676
rect 226392 228664 226398 228676
rect 272518 228664 272524 228676
rect 226392 228636 272524 228664
rect 226392 228624 226398 228636
rect 272518 228624 272524 228636
rect 272576 228624 272582 228676
rect 291654 228624 291660 228676
rect 291712 228664 291718 228676
rect 292132 228664 292160 228772
rect 300210 228760 300216 228772
rect 300268 228760 300274 228812
rect 300670 228760 300676 228812
rect 300728 228800 300734 228812
rect 330478 228800 330484 228812
rect 300728 228772 330484 228800
rect 300728 228760 300734 228772
rect 330478 228760 330484 228772
rect 330536 228760 330542 228812
rect 376018 228760 376024 228812
rect 376076 228800 376082 228812
rect 387794 228800 387800 228812
rect 376076 228772 387800 228800
rect 376076 228760 376082 228772
rect 387794 228760 387800 228772
rect 387852 228760 387858 228812
rect 478874 228760 478880 228812
rect 478932 228800 478938 228812
rect 490374 228800 490380 228812
rect 478932 228772 490380 228800
rect 478932 228760 478938 228772
rect 490374 228760 490380 228772
rect 490432 228760 490438 228812
rect 499850 228760 499856 228812
rect 499908 228800 499914 228812
rect 518158 228800 518164 228812
rect 499908 228772 518164 228800
rect 499908 228760 499914 228772
rect 518158 228760 518164 228772
rect 518216 228760 518222 228812
rect 518526 228760 518532 228812
rect 518584 228800 518590 228812
rect 541618 228800 541624 228812
rect 518584 228772 541624 228800
rect 518584 228760 518590 228772
rect 541618 228760 541624 228772
rect 541676 228760 541682 228812
rect 291712 228636 292160 228664
rect 291712 228624 291718 228636
rect 296622 228624 296628 228676
rect 296680 228664 296686 228676
rect 329190 228664 329196 228676
rect 296680 228636 329196 228664
rect 296680 228624 296686 228636
rect 329190 228624 329196 228636
rect 329248 228624 329254 228676
rect 336458 228624 336464 228676
rect 336516 228664 336522 228676
rect 358814 228664 358820 228676
rect 336516 228636 358820 228664
rect 336516 228624 336522 228636
rect 358814 228624 358820 228636
rect 358872 228624 358878 228676
rect 359918 228624 359924 228676
rect 359976 228664 359982 228676
rect 376846 228664 376852 228676
rect 359976 228636 376852 228664
rect 359976 228624 359982 228636
rect 376846 228624 376852 228636
rect 376904 228624 376910 228676
rect 485682 228624 485688 228676
rect 485740 228664 485746 228676
rect 498286 228664 498292 228676
rect 485740 228636 498292 228664
rect 485740 228624 485746 228636
rect 498286 228624 498292 228636
rect 498344 228624 498350 228676
rect 498562 228624 498568 228676
rect 498620 228664 498626 228676
rect 515766 228664 515772 228676
rect 498620 228636 515772 228664
rect 498620 228624 498626 228636
rect 515766 228624 515772 228636
rect 515824 228624 515830 228676
rect 517882 228624 517888 228676
rect 517940 228664 517946 228676
rect 539410 228664 539416 228676
rect 517940 228636 539416 228664
rect 517940 228624 517946 228636
rect 539410 228624 539416 228636
rect 539468 228624 539474 228676
rect 539594 228624 539600 228676
rect 539652 228664 539658 228676
rect 557166 228664 557172 228676
rect 539652 228636 557172 228664
rect 539652 228624 539658 228636
rect 557166 228624 557172 228636
rect 557224 228624 557230 228676
rect 137428 228500 146984 228528
rect 137428 228488 137434 228500
rect 147122 228488 147128 228540
rect 147180 228528 147186 228540
rect 200390 228528 200396 228540
rect 147180 228500 200396 228528
rect 147180 228488 147186 228500
rect 200390 228488 200396 228500
rect 200448 228488 200454 228540
rect 204898 228488 204904 228540
rect 204956 228528 204962 228540
rect 220998 228528 221004 228540
rect 204956 228500 221004 228528
rect 204956 228488 204962 228500
rect 220998 228488 221004 228500
rect 221056 228488 221062 228540
rect 264790 228528 264796 228540
rect 222672 228500 264796 228528
rect 137204 228364 137416 228392
rect 112990 228216 112996 228268
rect 113048 228256 113054 228268
rect 137186 228256 137192 228268
rect 113048 228228 137192 228256
rect 113048 228216 113054 228228
rect 137186 228216 137192 228228
rect 137244 228216 137250 228268
rect 137388 228256 137416 228364
rect 139302 228352 139308 228404
rect 139360 228392 139366 228404
rect 139360 228364 152504 228392
rect 139360 228352 139366 228364
rect 143074 228256 143080 228268
rect 137388 228228 143080 228256
rect 143074 228216 143080 228228
rect 143132 228216 143138 228268
rect 143442 228216 143448 228268
rect 143500 228256 143506 228268
rect 146018 228256 146024 228268
rect 143500 228228 146024 228256
rect 143500 228216 143506 228228
rect 146018 228216 146024 228228
rect 146076 228216 146082 228268
rect 146202 228216 146208 228268
rect 146260 228256 146266 228268
rect 148870 228256 148876 228268
rect 146260 228228 148876 228256
rect 146260 228216 146266 228228
rect 148870 228216 148876 228228
rect 148928 228216 148934 228268
rect 152476 228256 152504 228364
rect 153010 228352 153016 228404
rect 153068 228392 153074 228404
rect 215846 228392 215852 228404
rect 153068 228364 215852 228392
rect 153068 228352 153074 228364
rect 215846 228352 215852 228364
rect 215904 228352 215910 228404
rect 216490 228352 216496 228404
rect 216548 228392 216554 228404
rect 222672 228392 222700 228500
rect 264790 228488 264796 228500
rect 264848 228488 264854 228540
rect 272518 228488 272524 228540
rect 272576 228528 272582 228540
rect 309870 228528 309876 228540
rect 272576 228500 309876 228528
rect 272576 228488 272582 228500
rect 309870 228488 309876 228500
rect 309928 228488 309934 228540
rect 313918 228488 313924 228540
rect 313976 228528 313982 228540
rect 320818 228528 320824 228540
rect 313976 228500 320824 228528
rect 313976 228488 313982 228500
rect 320818 228488 320824 228500
rect 320876 228488 320882 228540
rect 325418 228488 325424 228540
rect 325476 228528 325482 228540
rect 349154 228528 349160 228540
rect 325476 228500 349160 228528
rect 325476 228488 325482 228500
rect 349154 228488 349160 228500
rect 349212 228488 349218 228540
rect 350442 228488 350448 228540
rect 350500 228528 350506 228540
rect 369118 228528 369124 228540
rect 350500 228500 369124 228528
rect 350500 228488 350506 228500
rect 369118 228488 369124 228500
rect 369176 228488 369182 228540
rect 371050 228488 371056 228540
rect 371108 228528 371114 228540
rect 385218 228528 385224 228540
rect 371108 228500 385224 228528
rect 371108 228488 371114 228500
rect 385218 228488 385224 228500
rect 385276 228488 385282 228540
rect 386046 228488 386052 228540
rect 386104 228528 386110 228540
rect 397454 228528 397460 228540
rect 386104 228500 397460 228528
rect 386104 228488 386110 228500
rect 397454 228488 397460 228500
rect 397512 228488 397518 228540
rect 407758 228528 407764 228540
rect 400232 228500 407764 228528
rect 216548 228364 222700 228392
rect 216548 228352 216554 228364
rect 224678 228352 224684 228404
rect 224736 228392 224742 228404
rect 273806 228392 273812 228404
rect 224736 228364 273812 228392
rect 224736 228352 224742 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 285490 228352 285496 228404
rect 285548 228392 285554 228404
rect 318886 228392 318892 228404
rect 285548 228364 318892 228392
rect 285548 228352 285554 228364
rect 318886 228352 318892 228364
rect 318944 228352 318950 228404
rect 330478 228352 330484 228404
rect 330536 228392 330542 228404
rect 354950 228392 354956 228404
rect 330536 228364 354956 228392
rect 330536 228352 330542 228364
rect 354950 228352 354956 228364
rect 355008 228352 355014 228404
rect 355318 228352 355324 228404
rect 355376 228392 355382 228404
rect 372982 228392 372988 228404
rect 355376 228364 372988 228392
rect 355376 228352 355382 228364
rect 372982 228352 372988 228364
rect 373040 228352 373046 228404
rect 373442 228352 373448 228404
rect 373500 228392 373506 228404
rect 387150 228392 387156 228404
rect 373500 228364 387156 228392
rect 373500 228352 373506 228364
rect 387150 228352 387156 228364
rect 387208 228352 387214 228404
rect 390002 228352 390008 228404
rect 390060 228392 390066 228404
rect 400030 228392 400036 228404
rect 390060 228364 400036 228392
rect 390060 228352 390066 228364
rect 400030 228352 400036 228364
rect 400088 228352 400094 228404
rect 205542 228256 205548 228268
rect 152476 228228 205548 228256
rect 205542 228216 205548 228228
rect 205600 228216 205606 228268
rect 205910 228216 205916 228268
rect 205968 228256 205974 228268
rect 257062 228256 257068 228268
rect 205968 228228 257068 228256
rect 205968 228216 205974 228228
rect 257062 228216 257068 228228
rect 257120 228216 257126 228268
rect 268930 228216 268936 228268
rect 268988 228256 268994 228268
rect 306006 228256 306012 228268
rect 268988 228228 306012 228256
rect 268988 228216 268994 228228
rect 306006 228216 306012 228228
rect 306064 228216 306070 228268
rect 400232 228256 400260 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 409782 228488 409788 228540
rect 409840 228528 409846 228540
rect 415486 228528 415492 228540
rect 409840 228500 415492 228528
rect 409840 228488 409846 228500
rect 415486 228488 415492 228500
rect 415544 228488 415550 228540
rect 485038 228488 485044 228540
rect 485096 228528 485102 228540
rect 498654 228528 498660 228540
rect 485096 228500 498660 228528
rect 485096 228488 485102 228500
rect 498654 228488 498660 228500
rect 498712 228488 498718 228540
rect 502426 228488 502432 228540
rect 502484 228528 502490 228540
rect 521102 228528 521108 228540
rect 502484 228500 521108 228528
rect 502484 228488 502490 228500
rect 521102 228488 521108 228500
rect 521160 228488 521166 228540
rect 527542 228488 527548 228540
rect 527600 228528 527606 228540
rect 553210 228528 553216 228540
rect 527600 228500 553216 228528
rect 527600 228488 527606 228500
rect 553210 228488 553216 228500
rect 553268 228488 553274 228540
rect 556798 228488 556804 228540
rect 556856 228528 556862 228540
rect 570598 228528 570604 228540
rect 556856 228500 570604 228528
rect 556856 228488 556862 228500
rect 570598 228488 570604 228500
rect 570656 228488 570662 228540
rect 673564 228404 673592 229112
rect 402790 228352 402796 228404
rect 402848 228392 402854 228404
rect 411622 228392 411628 228404
rect 402848 228364 411628 228392
rect 402848 228352 402854 228364
rect 411622 228352 411628 228364
rect 411680 228352 411686 228404
rect 474458 228352 474464 228404
rect 474516 228392 474522 228404
rect 484486 228392 484492 228404
rect 474516 228364 484492 228392
rect 474516 228352 474522 228364
rect 484486 228352 484492 228364
rect 484544 228352 484550 228404
rect 490190 228352 490196 228404
rect 490248 228392 490254 228404
rect 505186 228392 505192 228404
rect 490248 228364 505192 228392
rect 490248 228352 490254 228364
rect 505186 228352 505192 228364
rect 505244 228352 505250 228404
rect 512086 228352 512092 228404
rect 512144 228392 512150 228404
rect 532970 228392 532976 228404
rect 512144 228364 532976 228392
rect 512144 228352 512150 228364
rect 532970 228352 532976 228364
rect 533028 228352 533034 228404
rect 537202 228352 537208 228404
rect 537260 228392 537266 228404
rect 565630 228392 565636 228404
rect 537260 228364 565636 228392
rect 537260 228352 537266 228364
rect 565630 228352 565636 228364
rect 565688 228352 565694 228404
rect 673546 228352 673552 228404
rect 673604 228352 673610 228404
rect 400140 228228 400260 228256
rect 400140 228132 400168 228228
rect 539410 228216 539416 228268
rect 539468 228256 539474 228268
rect 540790 228256 540796 228268
rect 539468 228228 540796 228256
rect 539468 228216 539474 228228
rect 540790 228216 540796 228228
rect 540848 228216 540854 228268
rect 119982 228080 119988 228132
rect 120040 228120 120046 228132
rect 185210 228120 185216 228132
rect 120040 228092 185216 228120
rect 120040 228080 120046 228092
rect 185210 228080 185216 228092
rect 185268 228080 185274 228132
rect 185394 228080 185400 228132
rect 185452 228120 185458 228132
rect 185452 228092 194180 228120
rect 185452 228080 185458 228092
rect 126698 227944 126704 227996
rect 126756 227984 126762 227996
rect 194152 227984 194180 228092
rect 195238 228080 195244 228132
rect 195296 228120 195302 228132
rect 239030 228120 239036 228132
rect 195296 228092 239036 228120
rect 195296 228080 195302 228092
rect 239030 228080 239036 228092
rect 239088 228080 239094 228132
rect 400122 228080 400128 228132
rect 400180 228080 400186 228132
rect 415026 228012 415032 228064
rect 415084 228052 415090 228064
rect 421926 228052 421932 228064
rect 415084 228024 421932 228052
rect 415084 228012 415090 228024
rect 421926 228012 421932 228024
rect 421984 228012 421990 228064
rect 126756 227956 192892 227984
rect 194152 227956 200114 227984
rect 126756 227944 126762 227956
rect 88242 227808 88248 227860
rect 88300 227848 88306 227860
rect 95234 227848 95240 227860
rect 88300 227820 95240 227848
rect 88300 227808 88306 227820
rect 95234 227808 95240 227820
rect 95292 227808 95298 227860
rect 133506 227808 133512 227860
rect 133564 227848 133570 227860
rect 136634 227848 136640 227860
rect 133564 227820 136640 227848
rect 133564 227808 133570 227820
rect 136634 227808 136640 227820
rect 136692 227808 136698 227860
rect 136818 227808 136824 227860
rect 136876 227848 136882 227860
rect 141142 227848 141148 227860
rect 136876 227820 141148 227848
rect 136876 227808 136882 227820
rect 141142 227808 141148 227820
rect 141200 227808 141206 227860
rect 141510 227808 141516 227860
rect 141568 227848 141574 227860
rect 192478 227848 192484 227860
rect 141568 227820 192484 227848
rect 141568 227808 141574 227820
rect 192478 227808 192484 227820
rect 192536 227808 192542 227860
rect 192864 227848 192892 227956
rect 195054 227848 195060 227860
rect 192864 227820 195060 227848
rect 195054 227808 195060 227820
rect 195112 227808 195118 227860
rect 200086 227848 200114 227956
rect 200390 227944 200396 227996
rect 200448 227984 200454 227996
rect 210694 227984 210700 227996
rect 200448 227956 210700 227984
rect 200448 227944 200454 227956
rect 210694 227944 210700 227956
rect 210752 227944 210758 227996
rect 238386 227984 238392 227996
rect 219406 227956 238392 227984
rect 204898 227848 204904 227860
rect 200086 227820 204904 227848
rect 204898 227808 204904 227820
rect 204956 227808 204962 227860
rect 205450 227808 205456 227860
rect 205508 227848 205514 227860
rect 205910 227848 205916 227860
rect 205508 227820 205916 227848
rect 205508 227808 205514 227820
rect 205910 227808 205916 227820
rect 205968 227808 205974 227860
rect 210326 227808 210332 227860
rect 210384 227848 210390 227860
rect 219406 227848 219434 227956
rect 238386 227944 238392 227956
rect 238444 227944 238450 227996
rect 238662 227944 238668 227996
rect 238720 227984 238726 227996
rect 282822 227984 282828 227996
rect 238720 227956 282828 227984
rect 238720 227944 238726 227956
rect 282822 227944 282828 227956
rect 282880 227944 282886 227996
rect 416682 227876 416688 227928
rect 416740 227916 416746 227928
rect 420638 227916 420644 227928
rect 416740 227888 420644 227916
rect 416740 227876 416746 227888
rect 420638 227876 420644 227888
rect 420696 227876 420702 227928
rect 447042 227876 447048 227928
rect 447100 227916 447106 227928
rect 450538 227916 450544 227928
rect 447100 227888 450544 227916
rect 447100 227876 447106 227888
rect 450538 227876 450544 227888
rect 450596 227876 450602 227928
rect 210384 227820 219434 227848
rect 210384 227808 210390 227820
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 420638 227740 420644 227792
rect 420696 227780 420702 227792
rect 423858 227780 423864 227792
rect 420696 227752 423864 227780
rect 420696 227740 420702 227752
rect 423858 227740 423864 227752
rect 423916 227740 423922 227792
rect 471514 227740 471520 227792
rect 471572 227780 471578 227792
rect 479518 227780 479524 227792
rect 471572 227752 479524 227780
rect 471572 227740 471578 227752
rect 479518 227740 479524 227752
rect 479576 227740 479582 227792
rect 64782 227672 64788 227724
rect 64840 227712 64846 227724
rect 110322 227712 110328 227724
rect 64840 227684 110328 227712
rect 64840 227672 64846 227684
rect 110322 227672 110328 227684
rect 110380 227672 110386 227724
rect 110506 227672 110512 227724
rect 110564 227712 110570 227724
rect 182358 227712 182364 227724
rect 110564 227684 182364 227712
rect 110564 227672 110570 227684
rect 182358 227672 182364 227684
rect 182416 227672 182422 227724
rect 185210 227712 185216 227724
rect 182560 227684 185216 227712
rect 60642 227536 60648 227588
rect 60700 227576 60706 227588
rect 102134 227576 102140 227588
rect 60700 227548 102140 227576
rect 60700 227536 60706 227548
rect 102134 227536 102140 227548
rect 102192 227536 102198 227588
rect 103422 227536 103428 227588
rect 103480 227576 103486 227588
rect 175182 227576 175188 227588
rect 103480 227548 175188 227576
rect 103480 227536 103486 227548
rect 175182 227536 175188 227548
rect 175240 227536 175246 227588
rect 181530 227536 181536 227588
rect 181588 227576 181594 227588
rect 182560 227576 182588 227684
rect 185210 227672 185216 227684
rect 185268 227672 185274 227724
rect 185394 227672 185400 227724
rect 185452 227712 185458 227724
rect 192662 227712 192668 227724
rect 185452 227684 192668 227712
rect 185452 227672 185458 227684
rect 192662 227672 192668 227684
rect 192720 227672 192726 227724
rect 195238 227672 195244 227724
rect 195296 227712 195302 227724
rect 214742 227712 214748 227724
rect 195296 227684 214748 227712
rect 195296 227672 195302 227684
rect 214742 227672 214748 227684
rect 214800 227672 214806 227724
rect 214926 227672 214932 227724
rect 214984 227712 214990 227724
rect 262214 227712 262220 227724
rect 214984 227684 262220 227712
rect 214984 227672 214990 227684
rect 262214 227672 262220 227684
rect 262272 227672 262278 227724
rect 277026 227672 277032 227724
rect 277084 227712 277090 227724
rect 311802 227712 311808 227724
rect 277084 227684 311808 227712
rect 277084 227672 277090 227684
rect 311802 227672 311808 227684
rect 311860 227672 311866 227724
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 181588 227548 182588 227576
rect 181588 227536 181594 227548
rect 184106 227536 184112 227588
rect 184164 227576 184170 227588
rect 187510 227576 187516 227588
rect 184164 227548 187516 227576
rect 184164 227536 184170 227548
rect 187510 227536 187516 227548
rect 187568 227536 187574 227588
rect 189902 227536 189908 227588
rect 189960 227576 189966 227588
rect 205082 227576 205088 227588
rect 189960 227548 205088 227576
rect 189960 227536 189966 227548
rect 205082 227536 205088 227548
rect 205140 227536 205146 227588
rect 205266 227536 205272 227588
rect 205324 227576 205330 227588
rect 251910 227576 251916 227588
rect 205324 227548 251916 227576
rect 205324 227536 205330 227548
rect 251910 227536 251916 227548
rect 251968 227536 251974 227588
rect 259270 227536 259276 227588
rect 259328 227576 259334 227588
rect 298278 227576 298284 227588
rect 259328 227548 298284 227576
rect 259328 227536 259334 227548
rect 298278 227536 298284 227548
rect 298336 227536 298342 227588
rect 301498 227536 301504 227588
rect 301556 227576 301562 227588
rect 308582 227576 308588 227588
rect 301556 227548 308588 227576
rect 301556 227536 301562 227548
rect 308582 227536 308588 227548
rect 308640 227536 308646 227588
rect 524598 227536 524604 227588
rect 524656 227576 524662 227588
rect 539962 227576 539968 227588
rect 524656 227548 539968 227576
rect 524656 227536 524662 227548
rect 539962 227536 539968 227548
rect 540020 227536 540026 227588
rect 175918 227508 175924 227520
rect 175476 227480 175924 227508
rect 96430 227400 96436 227452
rect 96488 227440 96494 227452
rect 170766 227440 170772 227452
rect 96488 227412 170772 227440
rect 96488 227400 96494 227412
rect 170766 227400 170772 227412
rect 170824 227400 170830 227452
rect 171088 227400 171094 227452
rect 171146 227440 171152 227452
rect 175476 227440 175504 227480
rect 175918 227468 175924 227480
rect 175976 227468 175982 227520
rect 185578 227440 185584 227452
rect 171146 227412 175504 227440
rect 176304 227412 185584 227440
rect 171146 227400 171152 227412
rect 176304 227372 176332 227412
rect 185578 227400 185584 227412
rect 185636 227400 185642 227452
rect 185762 227400 185768 227452
rect 185820 227440 185826 227452
rect 223574 227440 223580 227452
rect 185820 227412 223580 227440
rect 185820 227400 185826 227412
rect 223574 227400 223580 227412
rect 223632 227400 223638 227452
rect 224218 227400 224224 227452
rect 224276 227440 224282 227452
rect 241606 227440 241612 227452
rect 224276 227412 241612 227440
rect 224276 227400 224282 227412
rect 241606 227400 241612 227412
rect 241664 227400 241670 227452
rect 257890 227400 257896 227452
rect 257948 227440 257954 227452
rect 299566 227440 299572 227452
rect 257948 227412 299572 227440
rect 257948 227400 257954 227412
rect 299566 227400 299572 227412
rect 299624 227400 299630 227452
rect 304902 227400 304908 227452
rect 304960 227440 304966 227452
rect 333698 227440 333704 227452
rect 304960 227412 333704 227440
rect 304960 227400 304966 227412
rect 333698 227400 333704 227412
rect 333756 227400 333762 227452
rect 333882 227400 333888 227452
rect 333940 227440 333946 227452
rect 356238 227440 356244 227452
rect 333940 227412 356244 227440
rect 333940 227400 333946 227412
rect 356238 227400 356244 227412
rect 356296 227400 356302 227452
rect 357066 227400 357072 227452
rect 357124 227440 357130 227452
rect 374270 227440 374276 227452
rect 357124 227412 374276 227440
rect 357124 227400 357130 227412
rect 374270 227400 374276 227412
rect 374328 227400 374334 227452
rect 514018 227400 514024 227452
rect 514076 227440 514082 227452
rect 535730 227440 535736 227452
rect 514076 227412 535736 227440
rect 514076 227400 514082 227412
rect 535730 227400 535736 227412
rect 535788 227400 535794 227452
rect 538306 227400 538312 227452
rect 538364 227440 538370 227452
rect 556062 227440 556068 227452
rect 538364 227412 556068 227440
rect 538364 227400 538370 227412
rect 556062 227400 556068 227412
rect 556120 227400 556126 227452
rect 176120 227344 176332 227372
rect 89622 227264 89628 227316
rect 89680 227304 89686 227316
rect 157288 227304 157294 227316
rect 89680 227276 157294 227304
rect 89680 227264 89686 227276
rect 157288 227264 157294 227276
rect 157346 227264 157352 227316
rect 157518 227264 157524 227316
rect 157576 227304 157582 227316
rect 176120 227304 176148 227344
rect 157576 227276 176148 227304
rect 157576 227264 157582 227276
rect 176746 227264 176752 227316
rect 176804 227304 176810 227316
rect 222470 227304 222476 227316
rect 176804 227276 222476 227304
rect 176804 227264 176810 227276
rect 222470 227264 222476 227276
rect 222528 227264 222534 227316
rect 233878 227304 233884 227316
rect 222672 227276 233884 227304
rect 63310 227128 63316 227180
rect 63368 227168 63374 227180
rect 144822 227168 144828 227180
rect 63368 227140 144828 227168
rect 63368 227128 63374 227140
rect 144822 227128 144828 227140
rect 144880 227128 144886 227180
rect 150066 227128 150072 227180
rect 150124 227168 150130 227180
rect 213270 227168 213276 227180
rect 150124 227140 213276 227168
rect 150124 227128 150130 227140
rect 213270 227128 213276 227140
rect 213328 227128 213334 227180
rect 214374 227128 214380 227180
rect 214432 227168 214438 227180
rect 222672 227168 222700 227276
rect 233878 227264 233884 227276
rect 233936 227264 233942 227316
rect 235810 227264 235816 227316
rect 235868 227304 235874 227316
rect 280246 227304 280252 227316
rect 235868 227276 280252 227304
rect 235868 227264 235874 227276
rect 280246 227264 280252 227276
rect 280304 227264 280310 227316
rect 306190 227264 306196 227316
rect 306248 227304 306254 227316
rect 336918 227304 336924 227316
rect 306248 227276 336924 227304
rect 306248 227264 306254 227276
rect 336918 227264 336924 227276
rect 336976 227264 336982 227316
rect 340690 227264 340696 227316
rect 340748 227304 340754 227316
rect 361390 227304 361396 227316
rect 340748 227276 361396 227304
rect 340748 227264 340754 227276
rect 361390 227264 361396 227276
rect 361448 227264 361454 227316
rect 382090 227264 382096 227316
rect 382148 227304 382154 227316
rect 392946 227304 392952 227316
rect 382148 227276 392952 227304
rect 382148 227264 382154 227276
rect 392946 227264 392952 227276
rect 393004 227264 393010 227316
rect 402606 227304 402612 227316
rect 393286 227276 402612 227304
rect 214432 227140 222700 227168
rect 214432 227128 214438 227140
rect 224034 227128 224040 227180
rect 224092 227168 224098 227180
rect 262858 227168 262864 227180
rect 224092 227140 262864 227168
rect 224092 227128 224098 227140
rect 262858 227128 262864 227140
rect 262916 227128 262922 227180
rect 263502 227128 263508 227180
rect 263560 227168 263566 227180
rect 277210 227168 277216 227180
rect 263560 227140 277216 227168
rect 263560 227128 263566 227140
rect 277210 227128 277216 227140
rect 277268 227128 277274 227180
rect 281350 227128 281356 227180
rect 281408 227168 281414 227180
rect 317598 227168 317604 227180
rect 281408 227140 317604 227168
rect 281408 227128 281414 227140
rect 317598 227128 317604 227140
rect 317656 227128 317662 227180
rect 322842 227128 322848 227180
rect 322900 227168 322906 227180
rect 349798 227168 349804 227180
rect 322900 227140 349804 227168
rect 322900 227128 322906 227140
rect 349798 227128 349804 227140
rect 349856 227128 349862 227180
rect 355870 227128 355876 227180
rect 355928 227168 355934 227180
rect 375558 227168 375564 227180
rect 355928 227140 375564 227168
rect 355928 227128 355934 227140
rect 375558 227128 375564 227140
rect 375616 227128 375622 227180
rect 376662 227128 376668 227180
rect 376720 227168 376726 227180
rect 389726 227168 389732 227180
rect 376720 227140 389732 227168
rect 376720 227128 376726 227140
rect 389726 227128 389732 227140
rect 389784 227128 389790 227180
rect 393130 227128 393136 227180
rect 393188 227168 393194 227180
rect 393286 227168 393314 227276
rect 402606 227264 402612 227276
rect 402664 227264 402670 227316
rect 494698 227264 494704 227316
rect 494756 227304 494762 227316
rect 494756 227276 504404 227304
rect 494756 227264 494762 227276
rect 393188 227140 393314 227168
rect 393188 227128 393194 227140
rect 402238 227128 402244 227180
rect 402296 227168 402302 227180
rect 408402 227168 408408 227180
rect 402296 227140 408408 227168
rect 402296 227128 402302 227140
rect 408402 227128 408408 227140
rect 408460 227128 408466 227180
rect 478598 227128 478604 227180
rect 478656 227168 478662 227180
rect 486786 227168 486792 227180
rect 478656 227140 486792 227168
rect 478656 227128 478662 227140
rect 486786 227128 486792 227140
rect 486844 227128 486850 227180
rect 489546 227128 489552 227180
rect 489604 227168 489610 227180
rect 504174 227168 504180 227180
rect 489604 227140 504180 227168
rect 489604 227128 489610 227140
rect 504174 227128 504180 227140
rect 504232 227128 504238 227180
rect 56502 226992 56508 227044
rect 56560 227032 56566 227044
rect 142430 227032 142436 227044
rect 56560 227004 142436 227032
rect 56560 226992 56566 227004
rect 142430 226992 142436 227004
rect 142488 226992 142494 227044
rect 143258 226992 143264 227044
rect 143316 227032 143322 227044
rect 204070 227032 204076 227044
rect 143316 227004 204076 227032
rect 143316 226992 143322 227004
rect 204070 226992 204076 227004
rect 204128 226992 204134 227044
rect 204916 227004 214696 227032
rect 117222 226856 117228 226908
rect 117280 226896 117286 226908
rect 184106 226896 184112 226908
rect 117280 226868 184112 226896
rect 117280 226856 117286 226868
rect 184106 226856 184112 226868
rect 184164 226856 184170 226908
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 204916 226896 204944 227004
rect 185636 226868 204944 226896
rect 185636 226856 185642 226868
rect 205082 226856 205088 226908
rect 205140 226896 205146 226908
rect 214374 226896 214380 226908
rect 205140 226868 214380 226896
rect 205140 226856 205146 226868
rect 214374 226856 214380 226868
rect 214432 226856 214438 226908
rect 214668 226896 214696 227004
rect 215110 226992 215116 227044
rect 215168 227032 215174 227044
rect 224218 227032 224224 227044
rect 215168 227004 224224 227032
rect 215168 226992 215174 227004
rect 224218 226992 224224 227004
rect 224276 226992 224282 227044
rect 271230 227032 271236 227044
rect 228928 227004 271236 227032
rect 218422 226896 218428 226908
rect 214668 226868 218428 226896
rect 218422 226856 218428 226868
rect 218480 226856 218486 226908
rect 222470 226856 222476 226908
rect 222528 226896 222534 226908
rect 228726 226896 228732 226908
rect 222528 226868 228732 226896
rect 222528 226856 222534 226868
rect 228726 226856 228732 226868
rect 228784 226856 228790 226908
rect 122742 226720 122748 226772
rect 122800 226760 122806 226772
rect 185394 226760 185400 226772
rect 122800 226732 185400 226760
rect 122800 226720 122806 226732
rect 185394 226720 185400 226732
rect 185452 226720 185458 226772
rect 186130 226720 186136 226772
rect 186188 226760 186194 226772
rect 195238 226760 195244 226772
rect 186188 226732 195244 226760
rect 186188 226720 186194 226732
rect 195238 226720 195244 226732
rect 195296 226720 195302 226772
rect 200022 226720 200028 226772
rect 200080 226760 200086 226772
rect 205266 226760 205272 226772
rect 200080 226732 205272 226760
rect 200080 226720 200086 226732
rect 205266 226720 205272 226732
rect 205324 226720 205330 226772
rect 222930 226760 222936 226772
rect 209746 226732 222936 226760
rect 129550 226584 129556 226636
rect 129608 226624 129614 226636
rect 197354 226624 197360 226636
rect 129608 226596 197360 226624
rect 129608 226584 129614 226596
rect 197354 226584 197360 226596
rect 197412 226584 197418 226636
rect 204070 226584 204076 226636
rect 204128 226624 204134 226636
rect 208118 226624 208124 226636
rect 204128 226596 208124 226624
rect 204128 226584 204134 226596
rect 208118 226584 208124 226596
rect 208176 226584 208182 226636
rect 136542 226448 136548 226500
rect 136600 226488 136606 226500
rect 141602 226488 141608 226500
rect 136600 226460 141608 226488
rect 136600 226448 136606 226460
rect 141602 226448 141608 226460
rect 141660 226448 141666 226500
rect 142246 226448 142252 226500
rect 142304 226488 142310 226500
rect 202966 226488 202972 226500
rect 142304 226460 202972 226488
rect 142304 226448 142310 226460
rect 202966 226448 202972 226460
rect 203024 226448 203030 226500
rect 203518 226448 203524 226500
rect 203576 226488 203582 226500
rect 209746 226488 209774 226732
rect 222930 226720 222936 226732
rect 222988 226720 222994 226772
rect 223114 226720 223120 226772
rect 223172 226760 223178 226772
rect 228928 226760 228956 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 301498 227032 301504 227044
rect 271840 227004 301504 227032
rect 271840 226992 271846 227004
rect 301498 226992 301504 227004
rect 301556 226992 301562 227044
rect 310422 226992 310428 227044
rect 310480 227032 310486 227044
rect 338206 227032 338212 227044
rect 310480 227004 338212 227032
rect 310480 226992 310486 227004
rect 338206 226992 338212 227004
rect 338264 226992 338270 227044
rect 338666 226992 338672 227044
rect 338724 227032 338730 227044
rect 360102 227032 360108 227044
rect 338724 227004 360108 227032
rect 338724 226992 338730 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 362770 226992 362776 227044
rect 362828 227032 362834 227044
rect 379422 227032 379428 227044
rect 362828 227004 379428 227032
rect 362828 226992 362834 227004
rect 379422 226992 379428 227004
rect 379480 226992 379486 227044
rect 391842 226992 391848 227044
rect 391900 227032 391906 227044
rect 403526 227032 403532 227044
rect 391900 227004 403532 227032
rect 391900 226992 391906 227004
rect 403526 226992 403532 227004
rect 403584 226992 403590 227044
rect 412542 226992 412548 227044
rect 412600 227032 412606 227044
rect 419350 227032 419356 227044
rect 412600 227004 419356 227032
rect 412600 226992 412606 227004
rect 419350 226992 419356 227004
rect 419408 226992 419414 227044
rect 486970 226992 486976 227044
rect 487028 227032 487034 227044
rect 500954 227032 500960 227044
rect 487028 227004 500960 227032
rect 487028 226992 487034 227004
rect 500954 226992 500960 227004
rect 501012 226992 501018 227044
rect 267366 226896 267372 226908
rect 223172 226732 228956 226760
rect 229066 226868 267372 226896
rect 223172 226720 223178 226732
rect 212166 226584 212172 226636
rect 212224 226624 212230 226636
rect 214926 226624 214932 226636
rect 212224 226596 214932 226624
rect 212224 226584 212230 226596
rect 214926 226584 214932 226596
rect 214984 226584 214990 226636
rect 219342 226584 219348 226636
rect 219400 226624 219406 226636
rect 229066 226624 229094 226868
rect 267366 226856 267372 226868
rect 267424 226856 267430 226908
rect 293770 226856 293776 226908
rect 293828 226896 293834 226908
rect 324958 226896 324964 226908
rect 293828 226868 324964 226896
rect 293828 226856 293834 226868
rect 324958 226856 324964 226868
rect 325016 226856 325022 226908
rect 504376 226896 504404 227276
rect 510614 227264 510620 227316
rect 510672 227304 510678 227316
rect 524414 227304 524420 227316
rect 510672 227276 524420 227304
rect 510672 227264 510678 227276
rect 524414 227264 524420 227276
rect 524472 227264 524478 227316
rect 526254 227264 526260 227316
rect 526312 227304 526318 227316
rect 551554 227304 551560 227316
rect 526312 227276 551560 227304
rect 526312 227264 526318 227276
rect 551554 227264 551560 227276
rect 551612 227264 551618 227316
rect 506198 227128 506204 227180
rect 506256 227168 506262 227180
rect 525978 227168 525984 227180
rect 506256 227140 525984 227168
rect 506256 227128 506262 227140
rect 525978 227128 525984 227140
rect 526036 227128 526042 227180
rect 533338 227128 533344 227180
rect 533396 227168 533402 227180
rect 560938 227168 560944 227180
rect 533396 227140 560944 227168
rect 533396 227128 533402 227140
rect 560938 227128 560944 227140
rect 560996 227128 561002 227180
rect 505002 226992 505008 227044
rect 505060 227032 505066 227044
rect 523034 227032 523040 227044
rect 505060 227004 523040 227032
rect 505060 226992 505066 227004
rect 523034 226992 523040 227004
rect 523092 226992 523098 227044
rect 523678 226992 523684 227044
rect 523736 227032 523742 227044
rect 548702 227032 548708 227044
rect 523736 227004 548708 227032
rect 523736 226992 523742 227004
rect 548702 226992 548708 227004
rect 548760 226992 548766 227044
rect 555418 226992 555424 227044
rect 555476 227032 555482 227044
rect 633710 227032 633716 227044
rect 555476 227004 633716 227032
rect 555476 226992 555482 227004
rect 633710 226992 633716 227004
rect 633768 226992 633774 227044
rect 510982 226896 510988 226908
rect 504376 226868 510988 226896
rect 510982 226856 510988 226868
rect 511040 226856 511046 226908
rect 672442 226856 672448 226908
rect 672500 226896 672506 226908
rect 673086 226896 673092 226908
rect 672500 226868 673092 226896
rect 672500 226856 672506 226868
rect 673086 226856 673092 226868
rect 673144 226856 673150 226908
rect 231026 226720 231032 226772
rect 231084 226760 231090 226772
rect 243262 226760 243268 226772
rect 231084 226732 243268 226760
rect 231084 226720 231090 226732
rect 243262 226720 243268 226732
rect 243320 226720 243326 226772
rect 249610 226720 249616 226772
rect 249668 226760 249674 226772
rect 290550 226760 290556 226772
rect 249668 226732 290556 226760
rect 249668 226720 249674 226732
rect 290550 226720 290556 226732
rect 290608 226720 290614 226772
rect 243446 226652 243452 226704
rect 243504 226692 243510 226704
rect 248690 226692 248696 226704
rect 243504 226664 248696 226692
rect 243504 226652 243510 226664
rect 248690 226652 248696 226664
rect 248748 226652 248754 226704
rect 219400 226596 229094 226624
rect 219400 226584 219406 226596
rect 264146 226516 264152 226568
rect 264204 226556 264210 226568
rect 269298 226556 269304 226568
rect 264204 226528 269304 226556
rect 264204 226516 264210 226528
rect 269298 226516 269304 226528
rect 269356 226516 269362 226568
rect 673270 226556 673276 226568
rect 672842 226528 673276 226556
rect 673270 226516 673276 226528
rect 673328 226516 673334 226568
rect 203576 226460 209774 226488
rect 203576 226448 203582 226460
rect 213822 226448 213828 226500
rect 213880 226488 213886 226500
rect 224034 226488 224040 226500
rect 213880 226460 224040 226488
rect 213880 226448 213886 226460
rect 224034 226448 224040 226460
rect 224092 226448 224098 226500
rect 351086 226448 351092 226500
rect 351144 226488 351150 226500
rect 353018 226488 353024 226500
rect 351144 226460 353024 226488
rect 351144 226448 351150 226460
rect 353018 226448 353024 226460
rect 353076 226448 353082 226500
rect 403986 226448 403992 226500
rect 404044 226488 404050 226500
rect 412266 226488 412272 226500
rect 404044 226460 412272 226488
rect 404044 226448 404050 226460
rect 412266 226448 412272 226460
rect 412324 226448 412330 226500
rect 474734 226448 474740 226500
rect 474792 226488 474798 226500
rect 482738 226488 482744 226500
rect 474792 226460 482744 226488
rect 474792 226448 474798 226460
rect 482738 226448 482744 226460
rect 482796 226448 482802 226500
rect 672724 226432 672776 226438
rect 141786 226380 141792 226432
rect 141844 226420 141850 226432
rect 142108 226420 142114 226432
rect 141844 226392 142114 226420
rect 141844 226380 141850 226392
rect 142108 226380 142114 226392
rect 142166 226380 142172 226432
rect 271138 226380 271144 226432
rect 271196 226420 271202 226432
rect 279602 226420 279608 226432
rect 271196 226392 279608 226420
rect 271196 226380 271202 226392
rect 279602 226380 279608 226392
rect 279660 226380 279666 226432
rect 672724 226374 672776 226380
rect 350258 226312 350264 226364
rect 350316 226352 350322 226364
rect 351730 226352 351736 226364
rect 350316 226324 351736 226352
rect 350316 226312 350322 226324
rect 351730 226312 351736 226324
rect 351788 226312 351794 226364
rect 388530 226312 388536 226364
rect 388588 226352 388594 226364
rect 391658 226352 391664 226364
rect 388588 226324 391664 226352
rect 388588 226312 388594 226324
rect 391658 226312 391664 226324
rect 391716 226312 391722 226364
rect 407758 226312 407764 226364
rect 407816 226352 407822 226364
rect 408678 226352 408684 226364
rect 407816 226324 408684 226352
rect 407816 226312 407822 226324
rect 408678 226312 408684 226324
rect 408736 226312 408742 226364
rect 481634 226312 481640 226364
rect 481692 226352 481698 226364
rect 487798 226352 487804 226364
rect 481692 226324 487804 226352
rect 481692 226312 481698 226324
rect 487798 226312 487804 226324
rect 487856 226312 487862 226364
rect 663518 226312 663524 226364
rect 663576 226352 663582 226364
rect 665266 226352 665272 226364
rect 663576 226324 665272 226352
rect 663576 226312 663582 226324
rect 665266 226312 665272 226324
rect 665324 226312 665330 226364
rect 122558 226244 122564 226296
rect 122616 226284 122622 226296
rect 193950 226284 193956 226296
rect 122616 226256 193956 226284
rect 122616 226244 122622 226256
rect 193950 226244 193956 226256
rect 194008 226244 194014 226296
rect 194134 226244 194140 226296
rect 194192 226284 194198 226296
rect 244182 226284 244188 226296
rect 194192 226256 244188 226284
rect 194192 226244 194198 226256
rect 244182 226244 244188 226256
rect 244240 226244 244246 226296
rect 266998 226244 267004 226296
rect 267056 226284 267062 226296
rect 274450 226284 274456 226296
rect 267056 226256 274456 226284
rect 267056 226244 267062 226256
rect 274450 226244 274456 226256
rect 274508 226244 274514 226296
rect 286318 226244 286324 226296
rect 286376 226284 286382 226296
rect 289906 226284 289912 226296
rect 286376 226256 289912 226284
rect 286376 226244 286382 226256
rect 289906 226244 289912 226256
rect 289964 226244 289970 226296
rect 291010 226244 291016 226296
rect 291068 226284 291074 226296
rect 322106 226284 322112 226296
rect 291068 226256 322112 226284
rect 291068 226244 291074 226256
rect 322106 226244 322112 226256
rect 322164 226244 322170 226296
rect 458634 226244 458640 226296
rect 458692 226284 458698 226296
rect 462958 226284 462964 226296
rect 458692 226256 462964 226284
rect 458692 226244 458698 226256
rect 462958 226244 462964 226256
rect 463016 226244 463022 226296
rect 672604 226160 672656 226166
rect 127618 226108 127624 226160
rect 127676 226148 127682 226160
rect 142108 226148 142114 226160
rect 127676 226120 142114 226148
rect 127676 226108 127682 226120
rect 142108 226108 142114 226120
rect 142166 226108 142172 226160
rect 142246 226108 142252 226160
rect 142304 226148 142310 226160
rect 209406 226148 209412 226160
rect 142304 226120 209412 226148
rect 142304 226108 142310 226120
rect 209406 226108 209412 226120
rect 209464 226108 209470 226160
rect 209682 226108 209688 226160
rect 209740 226148 209746 226160
rect 259638 226148 259644 226160
rect 209740 226120 259644 226148
rect 209740 226108 209746 226120
rect 259638 226108 259644 226120
rect 259696 226108 259702 226160
rect 261846 226108 261852 226160
rect 261904 226148 261910 226160
rect 300854 226148 300860 226160
rect 261904 226120 300860 226148
rect 261904 226108 261910 226120
rect 300854 226108 300860 226120
rect 300912 226108 300918 226160
rect 309042 226108 309048 226160
rect 309100 226148 309106 226160
rect 336274 226148 336280 226160
rect 309100 226120 336280 226148
rect 309100 226108 309106 226120
rect 336274 226108 336280 226120
rect 336332 226108 336338 226160
rect 528554 226108 528560 226160
rect 528612 226148 528618 226160
rect 542630 226148 542636 226160
rect 528612 226120 542636 226148
rect 528612 226108 528618 226120
rect 542630 226108 542636 226120
rect 542688 226108 542694 226160
rect 672604 226102 672656 226108
rect 66162 225972 66168 226024
rect 66220 226012 66226 226024
rect 142614 226012 142620 226024
rect 66220 225984 142620 226012
rect 66220 225972 66226 225984
rect 142614 225972 142620 225984
rect 142672 225972 142678 226024
rect 142798 225972 142804 226024
rect 142856 226012 142862 226024
rect 147582 226012 147588 226024
rect 142856 225984 147588 226012
rect 142856 225972 142862 225984
rect 147582 225972 147588 225984
rect 147640 225972 147646 226024
rect 147766 225972 147772 226024
rect 147824 226012 147830 226024
rect 147824 225984 157104 226012
rect 147824 225972 147830 225984
rect 83458 225836 83464 225888
rect 83516 225876 83522 225888
rect 156414 225876 156420 225888
rect 83516 225848 156420 225876
rect 83516 225836 83522 225848
rect 156414 225836 156420 225848
rect 156472 225836 156478 225888
rect 157076 225808 157104 225984
rect 157334 225972 157340 226024
rect 157392 226012 157398 226024
rect 217134 226012 217140 226024
rect 157392 225984 217140 226012
rect 157392 225972 157398 225984
rect 217134 225972 217140 225984
rect 217192 225972 217198 226024
rect 222010 225972 222016 226024
rect 222068 226012 222074 226024
rect 269942 226012 269948 226024
rect 222068 225984 269948 226012
rect 222068 225972 222074 225984
rect 269942 225972 269948 225984
rect 270000 225972 270006 226024
rect 278406 225972 278412 226024
rect 278464 226012 278470 226024
rect 313274 226012 313280 226024
rect 278464 225984 313280 226012
rect 278464 225972 278470 225984
rect 313274 225972 313280 225984
rect 313332 225972 313338 226024
rect 329742 225972 329748 226024
rect 329800 226012 329806 226024
rect 353662 226012 353668 226024
rect 329800 225984 353668 226012
rect 329800 225972 329806 225984
rect 353662 225972 353668 225984
rect 353720 225972 353726 226024
rect 354582 225972 354588 226024
rect 354640 226012 354646 226024
rect 372338 226012 372344 226024
rect 354640 225984 372344 226012
rect 354640 225972 354646 225984
rect 372338 225972 372344 225984
rect 372396 225972 372402 226024
rect 498102 225972 498108 226024
rect 498160 226012 498166 226024
rect 514294 226012 514300 226024
rect 498160 225984 514300 226012
rect 498160 225972 498166 225984
rect 514294 225972 514300 225984
rect 514352 225972 514358 226024
rect 516594 225972 516600 226024
rect 516652 226012 516658 226024
rect 538674 226012 538680 226024
rect 516652 225984 538680 226012
rect 516652 225972 516658 225984
rect 538674 225972 538680 225984
rect 538732 225972 538738 226024
rect 672494 225956 672546 225962
rect 672494 225898 672546 225904
rect 183646 225836 183652 225888
rect 183704 225876 183710 225888
rect 183704 225848 190454 225876
rect 183704 225836 183710 225848
rect 157076 225780 164234 225808
rect 76558 225700 76564 225752
rect 76616 225740 76622 225752
rect 164206 225740 164234 225780
rect 184290 225740 184296 225752
rect 76616 225712 147904 225740
rect 164206 225712 184296 225740
rect 76616 225700 76622 225712
rect 147876 225672 147904 225712
rect 184290 225700 184296 225712
rect 184348 225700 184354 225752
rect 190426 225740 190454 225848
rect 197998 225836 198004 225888
rect 198056 225876 198062 225888
rect 198056 225848 204944 225876
rect 198056 225836 198062 225848
rect 204714 225740 204720 225752
rect 190426 225712 204720 225740
rect 204714 225700 204720 225712
rect 204772 225700 204778 225752
rect 204916 225740 204944 225848
rect 205082 225836 205088 225888
rect 205140 225876 205146 225888
rect 236454 225876 236460 225888
rect 205140 225848 236460 225876
rect 205140 225836 205146 225848
rect 236454 225836 236460 225848
rect 236512 225836 236518 225888
rect 237282 225836 237288 225888
rect 237340 225876 237346 225888
rect 240318 225876 240324 225888
rect 237340 225848 240324 225876
rect 237340 225836 237346 225848
rect 240318 225836 240324 225848
rect 240376 225836 240382 225888
rect 252462 225836 252468 225888
rect 252520 225876 252526 225888
rect 293126 225876 293132 225888
rect 252520 225848 293132 225876
rect 252520 225836 252526 225848
rect 293126 225836 293132 225848
rect 293184 225836 293190 225888
rect 296438 225836 296444 225888
rect 296496 225876 296502 225888
rect 327534 225876 327540 225888
rect 296496 225848 327540 225876
rect 296496 225836 296502 225848
rect 327534 225836 327540 225848
rect 327592 225836 327598 225888
rect 332226 225836 332232 225888
rect 332284 225876 332290 225888
rect 357526 225876 357532 225888
rect 332284 225848 357532 225876
rect 332284 225836 332290 225848
rect 357526 225836 357532 225848
rect 357584 225836 357590 225888
rect 373810 225836 373816 225888
rect 373868 225876 373874 225888
rect 377674 225876 377680 225888
rect 373868 225848 377680 225876
rect 373868 225836 373874 225848
rect 377674 225836 377680 225848
rect 377732 225836 377738 225888
rect 377858 225836 377864 225888
rect 377916 225876 377922 225888
rect 390370 225876 390376 225888
rect 377916 225848 390376 225876
rect 377916 225836 377922 225848
rect 390370 225836 390376 225848
rect 390428 225836 390434 225888
rect 394326 225836 394332 225888
rect 394384 225876 394390 225888
rect 403250 225876 403256 225888
rect 394384 225848 403256 225876
rect 394384 225836 394390 225848
rect 403250 225836 403256 225848
rect 403308 225836 403314 225888
rect 483750 225836 483756 225888
rect 483808 225876 483814 225888
rect 497274 225876 497280 225888
rect 483808 225848 497280 225876
rect 483808 225836 483814 225848
rect 497274 225836 497280 225848
rect 497332 225836 497338 225888
rect 501138 225836 501144 225888
rect 501196 225876 501202 225888
rect 519262 225876 519268 225888
rect 501196 225848 519268 225876
rect 501196 225836 501202 225848
rect 519262 225836 519268 225848
rect 519320 225836 519326 225888
rect 521746 225836 521752 225888
rect 521804 225876 521810 225888
rect 545758 225876 545764 225888
rect 521804 225848 545764 225876
rect 521804 225836 521810 225848
rect 545758 225836 545764 225848
rect 545816 225836 545822 225888
rect 558178 225836 558184 225888
rect 558236 225876 558242 225888
rect 571334 225876 571340 225888
rect 558236 225848 571340 225876
rect 558236 225836 558242 225848
rect 571334 225836 571340 225848
rect 571392 225836 571398 225888
rect 672380 225752 672432 225758
rect 249334 225740 249340 225752
rect 204916 225712 249340 225740
rect 249334 225700 249340 225712
rect 249392 225700 249398 225752
rect 255038 225700 255044 225752
rect 255096 225740 255102 225752
rect 296990 225740 296996 225752
rect 255096 225712 296996 225740
rect 255096 225700 255102 225712
rect 296990 225700 296996 225712
rect 297048 225700 297054 225752
rect 315666 225700 315672 225752
rect 315724 225740 315730 225752
rect 344646 225740 344652 225752
rect 315724 225712 344652 225740
rect 315724 225700 315730 225712
rect 344646 225700 344652 225712
rect 344704 225700 344710 225752
rect 352926 225700 352932 225752
rect 352984 225740 352990 225752
rect 371602 225740 371608 225752
rect 352984 225712 371608 225740
rect 352984 225700 352990 225712
rect 371602 225700 371608 225712
rect 371660 225700 371666 225752
rect 371786 225700 371792 225752
rect 371844 225740 371850 225752
rect 382734 225740 382740 225752
rect 371844 225712 382740 225740
rect 371844 225700 371850 225712
rect 382734 225700 382740 225712
rect 382792 225700 382798 225752
rect 382918 225700 382924 225752
rect 382976 225740 382982 225752
rect 396166 225740 396172 225752
rect 382976 225712 396172 225740
rect 382976 225700 382982 225712
rect 396166 225700 396172 225712
rect 396224 225700 396230 225752
rect 488902 225700 488908 225752
rect 488960 225740 488966 225752
rect 503622 225740 503628 225752
rect 488960 225712 503628 225740
rect 488960 225700 488966 225712
rect 503622 225700 503628 225712
rect 503680 225700 503686 225752
rect 508866 225700 508872 225752
rect 508924 225740 508930 225752
rect 529198 225740 529204 225752
rect 508924 225712 529204 225740
rect 508924 225700 508930 225712
rect 529198 225700 529204 225712
rect 529256 225700 529262 225752
rect 535914 225700 535920 225752
rect 535972 225740 535978 225752
rect 563974 225740 563980 225752
rect 535972 225712 563980 225740
rect 535972 225700 535978 225712
rect 563974 225700 563980 225712
rect 564032 225700 564038 225752
rect 672380 225694 672432 225700
rect 156598 225672 156604 225684
rect 147876 225644 156604 225672
rect 156598 225632 156604 225644
rect 156656 225632 156662 225684
rect 671890 225632 671896 225684
rect 671948 225672 671954 225684
rect 671948 225644 672290 225672
rect 671948 225632 671954 225644
rect 72418 225564 72424 225616
rect 72476 225604 72482 225616
rect 142108 225604 142114 225616
rect 72476 225576 142114 225604
rect 72476 225564 72482 225576
rect 142108 225564 142114 225576
rect 142166 225564 142172 225616
rect 142246 225564 142252 225616
rect 142304 225604 142310 225616
rect 147674 225604 147680 225616
rect 142304 225576 147680 225604
rect 142304 225564 142310 225576
rect 147674 225564 147680 225576
rect 147732 225564 147738 225616
rect 157334 225564 157340 225616
rect 157392 225604 157398 225616
rect 214558 225604 214564 225616
rect 157392 225576 214564 225604
rect 157392 225564 157398 225576
rect 214558 225564 214564 225576
rect 214616 225564 214622 225616
rect 215202 225564 215208 225616
rect 215260 225604 215266 225616
rect 266078 225604 266084 225616
rect 215260 225576 266084 225604
rect 215260 225564 215266 225576
rect 266078 225564 266084 225576
rect 266136 225564 266142 225616
rect 270034 225564 270040 225616
rect 270092 225604 270098 225616
rect 282638 225604 282644 225616
rect 270092 225576 282644 225604
rect 270092 225564 270098 225576
rect 282638 225564 282644 225576
rect 282696 225564 282702 225616
rect 284110 225564 284116 225616
rect 284168 225604 284174 225616
rect 320174 225604 320180 225616
rect 284168 225576 320180 225604
rect 284168 225564 284174 225576
rect 320174 225564 320180 225576
rect 320232 225564 320238 225616
rect 321370 225564 321376 225616
rect 321428 225604 321434 225616
rect 346578 225604 346584 225616
rect 321428 225576 346584 225604
rect 321428 225564 321434 225576
rect 346578 225564 346584 225576
rect 346636 225564 346642 225616
rect 347038 225564 347044 225616
rect 347096 225604 347102 225616
rect 367830 225604 367836 225616
rect 347096 225576 367836 225604
rect 347096 225564 347102 225576
rect 367830 225564 367836 225576
rect 367888 225564 367894 225616
rect 372522 225564 372528 225616
rect 372580 225604 372586 225616
rect 387426 225604 387432 225616
rect 372580 225576 387432 225604
rect 372580 225564 372586 225576
rect 387426 225564 387432 225576
rect 387484 225564 387490 225616
rect 390186 225564 390192 225616
rect 390244 225604 390250 225616
rect 401962 225604 401968 225616
rect 390244 225576 401968 225604
rect 390244 225564 390250 225576
rect 401962 225564 401968 225576
rect 402020 225564 402026 225616
rect 410978 225564 410984 225616
rect 411036 225604 411042 225616
rect 416130 225604 416136 225616
rect 411036 225576 416136 225604
rect 411036 225564 411042 225576
rect 416130 225564 416136 225576
rect 416188 225564 416194 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 488810 225604 488816 225616
rect 477368 225576 488816 225604
rect 477368 225564 477374 225576
rect 488810 225564 488816 225576
rect 488868 225564 488874 225616
rect 494054 225564 494060 225616
rect 494112 225604 494118 225616
rect 509510 225604 509516 225616
rect 494112 225576 509516 225604
rect 494112 225564 494118 225576
rect 509510 225564 509516 225576
rect 509568 225564 509574 225616
rect 510154 225564 510160 225616
rect 510212 225604 510218 225616
rect 530946 225604 530952 225616
rect 510212 225576 530952 225604
rect 510212 225564 510218 225576
rect 530946 225564 530952 225576
rect 531004 225564 531010 225616
rect 531406 225564 531412 225616
rect 531464 225604 531470 225616
rect 558270 225604 558276 225616
rect 531464 225576 558276 225604
rect 531464 225564 531470 225576
rect 558270 225564 558276 225576
rect 558328 225564 558334 225616
rect 110138 225428 110144 225480
rect 110196 225468 110202 225480
rect 127618 225468 127624 225480
rect 110196 225440 127624 225468
rect 110196 225428 110202 225440
rect 127618 225428 127624 225440
rect 127676 225428 127682 225480
rect 196158 225468 196164 225480
rect 127820 225440 196164 225468
rect 125226 225292 125232 225344
rect 125284 225332 125290 225344
rect 127820 225332 127848 225440
rect 196158 225428 196164 225440
rect 196216 225428 196222 225480
rect 196342 225428 196348 225480
rect 196400 225468 196406 225480
rect 196400 225440 200114 225468
rect 196400 225428 196406 225440
rect 125284 225304 127848 225332
rect 125284 225292 125290 225304
rect 129366 225292 129372 225344
rect 129424 225332 129430 225344
rect 199102 225332 199108 225344
rect 129424 225304 199108 225332
rect 129424 225292 129430 225304
rect 199102 225292 199108 225304
rect 199160 225292 199166 225344
rect 200086 225332 200114 225440
rect 204714 225428 204720 225480
rect 204772 225468 204778 225480
rect 212534 225468 212540 225480
rect 204772 225440 212540 225468
rect 204772 225428 204778 225440
rect 212534 225428 212540 225440
rect 212592 225428 212598 225480
rect 257706 225468 257712 225480
rect 219406 225440 257712 225468
rect 205082 225332 205088 225344
rect 200086 225304 205088 225332
rect 205082 225292 205088 225304
rect 205140 225292 205146 225344
rect 208118 225292 208124 225344
rect 208176 225332 208182 225344
rect 219406 225332 219434 225440
rect 257706 225428 257712 225440
rect 257764 225428 257770 225480
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 672156 225344 672208 225350
rect 208176 225304 219434 225332
rect 208176 225292 208182 225304
rect 241146 225292 241152 225344
rect 241204 225332 241210 225344
rect 286686 225332 286692 225344
rect 241204 225304 286692 225332
rect 241204 225292 241210 225304
rect 286686 225292 286692 225304
rect 286744 225292 286750 225344
rect 563026 225304 572714 225332
rect 135070 225156 135076 225208
rect 135128 225196 135134 225208
rect 204254 225196 204260 225208
rect 135128 225168 204260 225196
rect 135128 225156 135134 225168
rect 204254 225156 204260 225168
rect 204312 225156 204318 225208
rect 242710 225156 242716 225208
rect 242768 225196 242774 225208
rect 285030 225196 285036 225208
rect 242768 225168 285036 225196
rect 242768 225156 242774 225168
rect 285030 225156 285036 225168
rect 285088 225156 285094 225208
rect 557626 225088 557632 225140
rect 557684 225128 557690 225140
rect 561950 225128 561956 225140
rect 557684 225100 561956 225128
rect 557684 225088 557690 225100
rect 561950 225088 561956 225100
rect 562008 225088 562014 225140
rect 132402 225020 132408 225072
rect 132460 225060 132466 225072
rect 201678 225060 201684 225072
rect 132460 225032 201684 225060
rect 132460 225020 132466 225032
rect 201678 225020 201684 225032
rect 201736 225020 201742 225072
rect 202690 225020 202696 225072
rect 202748 225060 202754 225072
rect 254486 225060 254492 225072
rect 202748 225032 254492 225060
rect 202748 225020 202754 225032
rect 254486 225020 254492 225032
rect 254544 225020 254550 225072
rect 297266 225020 297272 225072
rect 297324 225060 297330 225072
rect 305362 225060 305368 225072
rect 297324 225032 305368 225060
rect 297324 225020 297330 225032
rect 305362 225020 305368 225032
rect 305420 225020 305426 225072
rect 327718 224952 327724 225004
rect 327776 224992 327782 225004
rect 332042 224992 332048 225004
rect 327776 224964 332048 224992
rect 327776 224952 327782 224964
rect 332042 224952 332048 224964
rect 332100 224952 332106 225004
rect 369118 224952 369124 225004
rect 369176 224992 369182 225004
rect 373626 224992 373632 225004
rect 369176 224964 373632 224992
rect 369176 224952 369182 224964
rect 373626 224952 373632 224964
rect 373684 224952 373690 225004
rect 404170 224952 404176 225004
rect 404228 224992 404234 225004
rect 410610 224992 410616 225004
rect 404228 224964 410616 224992
rect 404228 224952 404234 224964
rect 410610 224952 410616 224964
rect 410668 224952 410674 225004
rect 416498 224952 416504 225004
rect 416556 224992 416562 225004
rect 422202 224992 422208 225004
rect 416556 224964 422208 224992
rect 416556 224952 416562 224964
rect 422202 224952 422208 224964
rect 422260 224952 422266 225004
rect 493686 224952 493692 225004
rect 493744 224992 493750 225004
rect 494698 224992 494704 225004
rect 493744 224964 494704 224992
rect 493744 224952 493750 224964
rect 494698 224952 494704 224964
rect 494756 224952 494762 225004
rect 495158 224952 495164 225004
rect 495216 224992 495222 225004
rect 563026 224992 563054 225304
rect 567010 225020 567016 225072
rect 567068 225060 567074 225072
rect 569126 225060 569132 225072
rect 567068 225032 569132 225060
rect 567068 225020 567074 225032
rect 569126 225020 569132 225032
rect 569184 225020 569190 225072
rect 572686 225060 572714 225304
rect 672156 225286 672208 225292
rect 672034 225276 672086 225282
rect 672034 225218 672086 225224
rect 572686 225032 576854 225060
rect 495216 224964 563054 224992
rect 495216 224952 495222 224964
rect 563698 224952 563704 225004
rect 563756 224992 563762 225004
rect 576826 224992 576854 225032
rect 666462 225020 666468 225072
rect 666520 225060 666526 225072
rect 666520 225032 671968 225060
rect 666520 225020 666526 225032
rect 630858 224992 630864 225004
rect 563756 224964 566780 224992
rect 576826 224964 630864 224992
rect 563756 224952 563762 224964
rect 96246 224884 96252 224936
rect 96304 224924 96310 224936
rect 172974 224924 172980 224936
rect 96304 224896 172980 224924
rect 96304 224884 96310 224896
rect 172974 224884 172980 224896
rect 173032 224884 173038 224936
rect 178494 224924 178500 224936
rect 176626 224896 178500 224924
rect 102042 224748 102048 224800
rect 102100 224788 102106 224800
rect 176626 224788 176654 224896
rect 178494 224884 178500 224896
rect 178552 224884 178558 224936
rect 178678 224884 178684 224936
rect 178736 224924 178742 224936
rect 185578 224924 185584 224936
rect 178736 224896 185584 224924
rect 178736 224884 178742 224896
rect 185578 224884 185584 224896
rect 185636 224884 185642 224936
rect 185762 224884 185768 224936
rect 185820 224924 185826 224936
rect 195238 224924 195244 224936
rect 185820 224896 195244 224924
rect 185820 224884 185826 224896
rect 195238 224884 195244 224896
rect 195296 224884 195302 224936
rect 195422 224884 195428 224936
rect 195480 224924 195486 224936
rect 242894 224924 242900 224936
rect 195480 224896 242900 224924
rect 195480 224884 195486 224896
rect 242894 224884 242900 224896
rect 242952 224884 242958 224936
rect 274266 224884 274272 224936
rect 274324 224924 274330 224936
rect 312446 224924 312452 224936
rect 274324 224896 312452 224924
rect 274324 224884 274330 224896
rect 312446 224884 312452 224896
rect 312504 224884 312510 224936
rect 460566 224884 460572 224936
rect 460624 224924 460630 224936
rect 463142 224924 463148 224936
rect 460624 224896 463148 224924
rect 460624 224884 460630 224896
rect 463142 224884 463148 224896
rect 463200 224884 463206 224936
rect 566752 224924 566780 224964
rect 630858 224952 630864 224964
rect 630916 224952 630922 225004
rect 568850 224924 568856 224936
rect 566752 224896 568856 224924
rect 568850 224884 568856 224896
rect 568908 224884 568914 224936
rect 572438 224924 572444 224936
rect 569052 224896 572444 224924
rect 102100 224760 176654 224788
rect 102100 224748 102106 224760
rect 178034 224748 178040 224800
rect 178092 224788 178098 224800
rect 204530 224788 204536 224800
rect 178092 224760 204536 224788
rect 178092 224748 178098 224760
rect 204530 224748 204536 224760
rect 204588 224748 204594 224800
rect 204714 224748 204720 224800
rect 204772 224788 204778 224800
rect 237742 224788 237748 224800
rect 204772 224760 237748 224788
rect 204772 224748 204778 224760
rect 237742 224748 237748 224760
rect 237800 224748 237806 224800
rect 245286 224748 245292 224800
rect 245344 224788 245350 224800
rect 287974 224788 287980 224800
rect 245344 224760 287980 224788
rect 245344 224748 245350 224760
rect 287974 224748 287980 224760
rect 288032 224748 288038 224800
rect 319990 224748 319996 224800
rect 320048 224788 320054 224800
rect 345934 224788 345940 224800
rect 320048 224760 345940 224788
rect 320048 224748 320054 224760
rect 345934 224748 345940 224760
rect 345992 224748 345998 224800
rect 462498 224748 462504 224800
rect 462556 224788 462562 224800
rect 469306 224788 469312 224800
rect 462556 224760 469312 224788
rect 462556 224748 462562 224760
rect 469306 224748 469312 224760
rect 469364 224748 469370 224800
rect 506934 224748 506940 224800
rect 506992 224788 506998 224800
rect 526714 224788 526720 224800
rect 506992 224760 526720 224788
rect 506992 224748 506998 224760
rect 526714 224748 526720 224760
rect 526772 224748 526778 224800
rect 529934 224748 529940 224800
rect 529992 224788 529998 224800
rect 548058 224788 548064 224800
rect 529992 224760 548064 224788
rect 529992 224748 529998 224760
rect 548058 224748 548064 224760
rect 548116 224748 548122 224800
rect 548242 224748 548248 224800
rect 548300 224788 548306 224800
rect 548300 224760 549162 224788
rect 548300 224748 548306 224760
rect 85482 224612 85488 224664
rect 85540 224652 85546 224664
rect 165614 224652 165620 224664
rect 85540 224624 165620 224652
rect 85540 224612 85546 224624
rect 165614 224612 165620 224624
rect 165672 224612 165678 224664
rect 174906 224612 174912 224664
rect 174964 224652 174970 224664
rect 178678 224652 178684 224664
rect 174964 224624 178684 224652
rect 174964 224612 174970 224624
rect 178678 224612 178684 224624
rect 178736 224612 178742 224664
rect 179322 224612 179328 224664
rect 179380 224652 179386 224664
rect 185394 224652 185400 224664
rect 179380 224624 185400 224652
rect 179380 224612 179386 224624
rect 185394 224612 185400 224624
rect 185452 224612 185458 224664
rect 185578 224612 185584 224664
rect 185636 224652 185642 224664
rect 235166 224652 235172 224664
rect 185636 224624 235172 224652
rect 185636 224612 185642 224624
rect 235166 224612 235172 224624
rect 235224 224612 235230 224664
rect 251082 224612 251088 224664
rect 251140 224652 251146 224664
rect 294414 224652 294420 224664
rect 251140 224624 294420 224652
rect 251140 224612 251146 224624
rect 294414 224612 294420 224624
rect 294472 224612 294478 224664
rect 299290 224612 299296 224664
rect 299348 224652 299354 224664
rect 331766 224652 331772 224664
rect 299348 224624 331772 224652
rect 299348 224612 299354 224624
rect 331766 224612 331772 224624
rect 331824 224612 331830 224664
rect 335170 224612 335176 224664
rect 335228 224652 335234 224664
rect 356882 224652 356888 224664
rect 335228 224624 356888 224652
rect 335228 224612 335234 224624
rect 356882 224612 356888 224624
rect 356940 224612 356946 224664
rect 363598 224612 363604 224664
rect 363656 224652 363662 224664
rect 368474 224652 368480 224664
rect 363656 224624 368480 224652
rect 363656 224612 363662 224624
rect 368474 224612 368480 224624
rect 368532 224612 368538 224664
rect 520458 224612 520464 224664
rect 520516 224652 520522 224664
rect 544102 224652 544108 224664
rect 520516 224624 544108 224652
rect 520516 224612 520522 224624
rect 544102 224612 544108 224624
rect 544160 224612 544166 224664
rect 544286 224612 544292 224664
rect 544344 224652 544350 224664
rect 545022 224652 545028 224664
rect 544344 224624 545028 224652
rect 544344 224612 544350 224624
rect 545022 224612 545028 224624
rect 545080 224652 545086 224664
rect 549134 224652 549162 224760
rect 549254 224748 549260 224800
rect 549312 224788 549318 224800
rect 557626 224788 557632 224800
rect 549312 224760 557632 224788
rect 549312 224748 549318 224760
rect 557626 224748 557632 224760
rect 557684 224748 557690 224800
rect 557810 224748 557816 224800
rect 557868 224788 557874 224800
rect 562134 224788 562140 224800
rect 557868 224760 562140 224788
rect 557868 224748 557874 224760
rect 562134 224748 562140 224760
rect 562192 224748 562198 224800
rect 562318 224748 562324 224800
rect 562376 224788 562382 224800
rect 567010 224788 567016 224800
rect 562376 224760 567016 224788
rect 562376 224748 562382 224760
rect 567010 224748 567016 224760
rect 567068 224748 567074 224800
rect 567194 224748 567200 224800
rect 567252 224788 567258 224800
rect 569052 224788 569080 224896
rect 572438 224884 572444 224896
rect 572496 224884 572502 224936
rect 671820 224800 671872 224806
rect 567252 224760 569080 224788
rect 567252 224748 567258 224760
rect 569218 224748 569224 224800
rect 569276 224788 569282 224800
rect 571334 224788 571340 224800
rect 569276 224760 571340 224788
rect 569276 224748 569282 224760
rect 571334 224748 571340 224760
rect 571392 224748 571398 224800
rect 571702 224748 571708 224800
rect 571760 224788 571766 224800
rect 616046 224788 616052 224800
rect 571760 224760 616052 224788
rect 571760 224748 571766 224760
rect 616046 224748 616052 224760
rect 616104 224748 616110 224800
rect 671820 224742 671872 224748
rect 550634 224652 550640 224664
rect 545080 224624 548656 224652
rect 549134 224624 550640 224652
rect 545080 224612 545086 224624
rect 79962 224476 79968 224528
rect 80020 224516 80026 224528
rect 160462 224516 160468 224528
rect 80020 224488 160468 224516
rect 80020 224476 80026 224488
rect 160462 224476 160468 224488
rect 160520 224476 160526 224528
rect 161658 224476 161664 224528
rect 161716 224516 161722 224528
rect 224862 224516 224868 224528
rect 161716 224488 224868 224516
rect 161716 224476 161722 224488
rect 224862 224476 224868 224488
rect 224920 224476 224926 224528
rect 228726 224476 228732 224528
rect 228784 224516 228790 224528
rect 274910 224516 274916 224528
rect 228784 224488 274916 224516
rect 228784 224476 228790 224488
rect 274910 224476 274916 224488
rect 274968 224476 274974 224528
rect 275094 224476 275100 224528
rect 275152 224516 275158 224528
rect 311158 224516 311164 224528
rect 275152 224488 311164 224516
rect 275152 224476 275158 224488
rect 311158 224476 311164 224488
rect 311216 224476 311222 224528
rect 311526 224476 311532 224528
rect 311584 224516 311590 224528
rect 338850 224516 338856 224528
rect 311584 224488 338856 224516
rect 311584 224476 311590 224488
rect 338850 224476 338856 224488
rect 338908 224476 338914 224528
rect 346210 224476 346216 224528
rect 346268 224516 346274 224528
rect 366542 224516 366548 224528
rect 346268 224488 366548 224516
rect 346268 224476 346274 224488
rect 366542 224476 366548 224488
rect 366600 224476 366606 224528
rect 387702 224476 387708 224528
rect 387760 224516 387766 224528
rect 397822 224516 397828 224528
rect 387760 224488 397828 224516
rect 387760 224476 387766 224488
rect 397822 224476 397828 224488
rect 397880 224476 397886 224528
rect 456058 224476 456064 224528
rect 456116 224516 456122 224528
rect 459738 224516 459744 224528
rect 456116 224488 459744 224516
rect 456116 224476 456122 224488
rect 459738 224476 459744 224488
rect 459796 224476 459802 224528
rect 491294 224476 491300 224528
rect 491352 224516 491358 224528
rect 506014 224516 506020 224528
rect 491352 224488 506020 224516
rect 491352 224476 491358 224488
rect 506014 224476 506020 224488
rect 506072 224476 506078 224528
rect 515950 224476 515956 224528
rect 516008 224516 516014 224528
rect 538858 224516 538864 224528
rect 516008 224488 538864 224516
rect 516008 224476 516014 224488
rect 538858 224476 538864 224488
rect 538916 224476 538922 224528
rect 539962 224476 539968 224528
rect 540020 224516 540026 224528
rect 542446 224516 542452 224528
rect 540020 224488 542452 224516
rect 540020 224476 540026 224488
rect 542446 224476 542452 224488
rect 542504 224476 542510 224528
rect 542814 224476 542820 224528
rect 542872 224516 542878 224528
rect 548628 224516 548656 224624
rect 550634 224612 550640 224624
rect 550692 224612 550698 224664
rect 550772 224612 550778 224664
rect 550830 224652 550836 224664
rect 625246 224652 625252 224664
rect 550830 224624 625252 224652
rect 550830 224612 550836 224624
rect 625246 224612 625252 224624
rect 625304 224612 625310 224664
rect 666830 224612 666836 224664
rect 666888 224652 666894 224664
rect 666888 224624 671738 224652
rect 666888 224612 666894 224624
rect 623774 224516 623780 224528
rect 542872 224488 548564 224516
rect 548628 224488 623780 224516
rect 542872 224476 542878 224488
rect 73706 224340 73712 224392
rect 73764 224380 73770 224392
rect 88978 224380 88984 224392
rect 73764 224352 88984 224380
rect 73764 224340 73770 224352
rect 88978 224340 88984 224352
rect 89036 224340 89042 224392
rect 89438 224340 89444 224392
rect 89496 224380 89502 224392
rect 167822 224380 167828 224392
rect 89496 224352 167828 224380
rect 89496 224340 89502 224352
rect 167822 224340 167828 224352
rect 167880 224340 167886 224392
rect 168282 224340 168288 224392
rect 168340 224380 168346 224392
rect 230014 224380 230020 224392
rect 168340 224352 230020 224380
rect 168340 224340 168346 224352
rect 230014 224340 230020 224352
rect 230072 224340 230078 224392
rect 233142 224340 233148 224392
rect 233200 224380 233206 224392
rect 277670 224380 277676 224392
rect 233200 224352 277676 224380
rect 233200 224340 233206 224352
rect 277670 224340 277676 224352
rect 277728 224340 277734 224392
rect 286686 224340 286692 224392
rect 286744 224380 286750 224392
rect 319530 224380 319536 224392
rect 286744 224352 319536 224380
rect 286744 224340 286750 224352
rect 319530 224340 319536 224352
rect 319588 224340 319594 224392
rect 319806 224340 319812 224392
rect 319864 224380 319870 224392
rect 347222 224380 347228 224392
rect 319864 224352 347228 224380
rect 319864 224340 319870 224352
rect 347222 224340 347228 224352
rect 347280 224340 347286 224392
rect 361206 224340 361212 224392
rect 361264 224380 361270 224392
rect 377490 224380 377496 224392
rect 361264 224352 377496 224380
rect 361264 224340 361270 224352
rect 377490 224340 377496 224352
rect 377548 224340 377554 224392
rect 379238 224340 379244 224392
rect 379296 224380 379302 224392
rect 393590 224380 393596 224392
rect 379296 224352 393596 224380
rect 379296 224340 379302 224352
rect 393590 224340 393596 224352
rect 393648 224340 393654 224392
rect 480530 224340 480536 224392
rect 480588 224380 480594 224392
rect 492766 224380 492772 224392
rect 480588 224352 492772 224380
rect 480588 224340 480594 224352
rect 492766 224340 492772 224352
rect 492824 224340 492830 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516778 224380 516784 224392
rect 499264 224352 516784 224380
rect 499264 224340 499270 224352
rect 516778 224340 516784 224352
rect 516836 224340 516842 224392
rect 525610 224340 525616 224392
rect 525668 224380 525674 224392
rect 548242 224380 548248 224392
rect 525668 224352 548248 224380
rect 525668 224340 525674 224352
rect 548242 224340 548248 224352
rect 548300 224340 548306 224392
rect 548536 224380 548564 224488
rect 623774 224476 623780 224488
rect 623832 224476 623838 224528
rect 667750 224408 667756 224460
rect 667808 224448 667814 224460
rect 667808 224420 671622 224448
rect 667808 224408 667814 224420
rect 548536 224352 553394 224380
rect 426434 224272 426440 224324
rect 426492 224312 426498 224324
rect 426986 224312 426992 224324
rect 426492 224284 426992 224312
rect 426492 224272 426498 224284
rect 426986 224272 426992 224284
rect 427044 224272 427050 224324
rect 553366 224312 553394 224352
rect 557994 224340 558000 224392
rect 558052 224380 558058 224392
rect 625430 224380 625436 224392
rect 558052 224352 625436 224380
rect 558052 224340 558058 224352
rect 625430 224340 625436 224352
rect 625488 224340 625494 224392
rect 553366 224284 557764 224312
rect 151630 224244 151636 224256
rect 84166 224216 151636 224244
rect 68922 224068 68928 224120
rect 68980 224108 68986 224120
rect 84166 224108 84194 224216
rect 151630 224204 151636 224216
rect 151688 224204 151694 224256
rect 151768 224204 151774 224256
rect 151826 224244 151832 224256
rect 155310 224244 155316 224256
rect 151826 224216 155316 224244
rect 151826 224204 151832 224216
rect 155310 224204 155316 224216
rect 155368 224204 155374 224256
rect 157242 224204 157248 224256
rect 157300 224244 157306 224256
rect 160922 224244 160928 224256
rect 157300 224216 160928 224244
rect 157300 224204 157306 224216
rect 160922 224204 160928 224216
rect 160980 224204 160986 224256
rect 165154 224204 165160 224256
rect 165212 224244 165218 224256
rect 227438 224244 227444 224256
rect 165212 224216 227444 224244
rect 165212 224204 165218 224216
rect 227438 224204 227444 224216
rect 227496 224204 227502 224256
rect 231670 224204 231676 224256
rect 231728 224244 231734 224256
rect 278958 224244 278964 224256
rect 231728 224216 278964 224244
rect 231728 224204 231734 224216
rect 278958 224204 278964 224216
rect 279016 224204 279022 224256
rect 290826 224204 290832 224256
rect 290884 224244 290890 224256
rect 323670 224244 323676 224256
rect 290884 224216 323676 224244
rect 290884 224204 290890 224216
rect 323670 224204 323676 224216
rect 323728 224204 323734 224256
rect 323946 224204 323952 224256
rect 324004 224244 324010 224256
rect 334986 224244 334992 224256
rect 324004 224216 334992 224244
rect 324004 224204 324010 224216
rect 334986 224204 334992 224216
rect 335044 224204 335050 224256
rect 339402 224204 339408 224256
rect 339460 224244 339466 224256
rect 339460 224216 354674 224244
rect 339460 224204 339466 224216
rect 68980 224080 84194 224108
rect 68980 224068 68986 224080
rect 88978 224068 88984 224120
rect 89036 224108 89042 224120
rect 142108 224108 142114 224120
rect 89036 224080 142114 224108
rect 89036 224068 89042 224080
rect 142108 224068 142114 224080
rect 142166 224068 142172 224120
rect 142246 224068 142252 224120
rect 142304 224108 142310 224120
rect 194594 224108 194600 224120
rect 142304 224080 194600 224108
rect 142304 224068 142310 224080
rect 194594 224068 194600 224080
rect 194652 224068 194658 224120
rect 195238 224068 195244 224120
rect 195296 224108 195302 224120
rect 204622 224108 204628 224120
rect 195296 224080 204628 224108
rect 195296 224068 195302 224080
rect 204622 224068 204628 224080
rect 204680 224068 204686 224120
rect 255774 224108 255780 224120
rect 204916 224080 255780 224108
rect 204916 224040 204944 224080
rect 255774 224068 255780 224080
rect 255832 224068 255838 224120
rect 266170 224068 266176 224120
rect 266228 224108 266234 224120
rect 303430 224108 303436 224120
rect 266228 224080 303436 224108
rect 266228 224068 266234 224080
rect 303430 224068 303436 224080
rect 303488 224068 303494 224120
rect 354646 224108 354674 224216
rect 358078 224204 358084 224256
rect 358136 224244 358142 224256
rect 363322 224244 363328 224256
rect 358136 224216 363328 224244
rect 358136 224204 358142 224216
rect 363322 224204 363328 224216
rect 363380 224204 363386 224256
rect 366726 224204 366732 224256
rect 366784 224244 366790 224256
rect 381630 224244 381636 224256
rect 366784 224216 381636 224244
rect 366784 224204 366790 224216
rect 381630 224204 381636 224216
rect 381688 224204 381694 224256
rect 394510 224204 394516 224256
rect 394568 224244 394574 224256
rect 404538 224244 404544 224256
rect 394568 224216 404544 224244
rect 394568 224204 394574 224216
rect 404538 224204 404544 224216
rect 404596 224204 404602 224256
rect 405550 224204 405556 224256
rect 405608 224244 405614 224256
rect 414198 224244 414204 224256
rect 405608 224216 414204 224244
rect 405608 224204 405614 224216
rect 414198 224204 414204 224216
rect 414256 224204 414262 224256
rect 427906 224204 427912 224256
rect 427964 224244 427970 224256
rect 428734 224244 428740 224256
rect 427964 224216 428740 224244
rect 427964 224204 427970 224216
rect 428734 224204 428740 224216
rect 428792 224204 428798 224256
rect 447502 224204 447508 224256
rect 447560 224244 447566 224256
rect 448054 224244 448060 224256
rect 447560 224216 448060 224244
rect 447560 224204 447566 224216
rect 448054 224204 448060 224216
rect 448112 224204 448118 224256
rect 470226 224204 470232 224256
rect 470284 224244 470290 224256
rect 480438 224244 480444 224256
rect 470284 224216 480444 224244
rect 470284 224204 470290 224216
rect 480438 224204 480444 224216
rect 480496 224204 480502 224256
rect 486602 224204 486608 224256
rect 486660 224244 486666 224256
rect 500034 224244 500040 224256
rect 486660 224216 500040 224244
rect 486660 224204 486666 224216
rect 500034 224204 500040 224216
rect 500092 224204 500098 224256
rect 504450 224204 504456 224256
rect 504508 224244 504514 224256
rect 523494 224244 523500 224256
rect 504508 224216 523500 224244
rect 504508 224204 504514 224216
rect 523494 224204 523500 224216
rect 523552 224204 523558 224256
rect 535270 224204 535276 224256
rect 535328 224244 535334 224256
rect 535328 224216 543734 224244
rect 535328 224204 535334 224216
rect 543706 224176 543734 224216
rect 557534 224176 557540 224188
rect 543706 224148 557540 224176
rect 557534 224136 557540 224148
rect 557592 224136 557598 224188
rect 557736 224176 557764 224284
rect 571702 224176 571708 224188
rect 557736 224148 571708 224176
rect 571702 224136 571708 224148
rect 571760 224136 571766 224188
rect 572438 224136 572444 224188
rect 572496 224176 572502 224188
rect 628742 224176 628748 224188
rect 572496 224148 628748 224176
rect 572496 224136 572502 224148
rect 628742 224136 628748 224148
rect 628800 224136 628806 224188
rect 671482 224120 671534 224126
rect 362310 224108 362316 224120
rect 354646 224080 362316 224108
rect 362310 224068 362316 224080
rect 362368 224068 362374 224120
rect 377398 224068 377404 224120
rect 377456 224108 377462 224120
rect 385862 224108 385868 224120
rect 377456 224080 385868 224108
rect 377456 224068 377462 224080
rect 385862 224068 385868 224080
rect 385920 224068 385926 224120
rect 519078 224068 519084 224120
rect 519136 224108 519142 224120
rect 534994 224108 535000 224120
rect 519136 224080 535000 224108
rect 519136 224068 519142 224080
rect 534994 224068 535000 224080
rect 535052 224108 535058 224120
rect 535052 224080 538214 224108
rect 535052 224068 535058 224080
rect 204824 224012 204944 224040
rect 538186 224040 538214 224080
rect 671482 224062 671534 224068
rect 542998 224040 543004 224052
rect 538186 224012 543004 224040
rect 105906 223932 105912 223984
rect 105964 223972 105970 223984
rect 181070 223972 181076 223984
rect 105964 223944 181076 223972
rect 105964 223932 105970 223944
rect 181070 223932 181076 223944
rect 181128 223932 181134 223984
rect 201218 223932 201224 223984
rect 201276 223972 201282 223984
rect 204824 223972 204852 224012
rect 542998 224000 543004 224012
rect 543056 224000 543062 224052
rect 543182 224000 543188 224052
rect 543240 224040 543246 224052
rect 622670 224040 622676 224052
rect 543240 224012 622676 224040
rect 543240 224000 543246 224012
rect 622670 224000 622676 224012
rect 622728 224000 622734 224052
rect 670712 224012 671398 224040
rect 201276 223944 204852 223972
rect 201276 223932 201282 223944
rect 205082 223932 205088 223984
rect 205140 223972 205146 223984
rect 250622 223972 250628 223984
rect 205140 223944 250628 223972
rect 205140 223932 205146 223944
rect 250622 223932 250628 223944
rect 250680 223932 250686 223984
rect 667750 223932 667756 223984
rect 667808 223972 667814 223984
rect 670712 223972 670740 224012
rect 667808 223944 670740 223972
rect 667808 223932 667814 223944
rect 279418 223864 279424 223916
rect 279476 223904 279482 223916
rect 284754 223904 284760 223916
rect 279476 223876 284760 223904
rect 279476 223864 279482 223876
rect 284754 223864 284760 223876
rect 284812 223864 284818 223916
rect 524414 223864 524420 223916
rect 524472 223904 524478 223916
rect 525058 223904 525064 223916
rect 524472 223876 525064 223904
rect 524472 223864 524478 223876
rect 525058 223864 525064 223876
rect 525116 223904 525122 223916
rect 619634 223904 619640 223916
rect 525116 223876 619640 223904
rect 525116 223864 525122 223876
rect 619634 223864 619640 223876
rect 619692 223864 619698 223916
rect 108666 223796 108672 223848
rect 108724 223836 108730 223848
rect 183830 223836 183836 223848
rect 108724 223808 183836 223836
rect 108724 223796 108730 223808
rect 183830 223796 183836 223808
rect 183888 223796 183894 223848
rect 185946 223836 185952 223848
rect 184032 223808 185952 223836
rect 112806 223660 112812 223712
rect 112864 223700 112870 223712
rect 184032 223700 184060 223808
rect 185946 223796 185952 223808
rect 186004 223796 186010 223848
rect 186958 223796 186964 223848
rect 187016 223836 187022 223848
rect 217778 223836 217784 223848
rect 187016 223808 217784 223836
rect 187016 223796 187022 223808
rect 217778 223796 217784 223808
rect 217836 223796 217842 223848
rect 224586 223796 224592 223848
rect 224644 223836 224650 223848
rect 270586 223836 270592 223848
rect 224644 223808 270592 223836
rect 224644 223796 224650 223808
rect 270586 223796 270592 223808
rect 270644 223796 270650 223848
rect 667014 223796 667020 223848
rect 667072 223836 667078 223848
rect 667072 223808 671278 223836
rect 667072 223796 667078 223808
rect 509510 223728 509516 223780
rect 509568 223768 509574 223780
rect 510154 223768 510160 223780
rect 509568 223740 510160 223768
rect 509568 223728 509574 223740
rect 510154 223728 510160 223740
rect 510212 223768 510218 223780
rect 542814 223768 542820 223780
rect 510212 223740 542820 223768
rect 510212 223728 510218 223740
rect 542814 223728 542820 223740
rect 542872 223728 542878 223780
rect 542998 223728 543004 223780
rect 543056 223768 543062 223780
rect 621566 223768 621572 223780
rect 543056 223740 621572 223768
rect 543056 223728 543062 223740
rect 621566 223728 621572 223740
rect 621624 223728 621630 223780
rect 112864 223672 184060 223700
rect 112864 223660 112870 223672
rect 184842 223660 184848 223712
rect 184900 223700 184906 223712
rect 195422 223700 195428 223712
rect 184900 223672 195428 223700
rect 184900 223660 184906 223672
rect 195422 223660 195428 223672
rect 195480 223660 195486 223712
rect 195882 223660 195888 223712
rect 195940 223700 195946 223712
rect 205082 223700 205088 223712
rect 195940 223672 205088 223700
rect 195940 223660 195946 223672
rect 205082 223660 205088 223672
rect 205140 223660 205146 223712
rect 238018 223660 238024 223712
rect 238076 223700 238082 223712
rect 266722 223700 266728 223712
rect 238076 223672 266728 223700
rect 238076 223660 238082 223672
rect 266722 223660 266728 223672
rect 266780 223660 266786 223712
rect 505186 223592 505192 223644
rect 505244 223632 505250 223644
rect 614942 223632 614948 223644
rect 505244 223604 614948 223632
rect 505244 223592 505250 223604
rect 614942 223592 614948 223604
rect 615000 223592 615006 223644
rect 669590 223592 669596 223644
rect 669648 223632 669654 223644
rect 669648 223604 671186 223632
rect 669648 223592 669654 223604
rect 81342 223524 81348 223576
rect 81400 223564 81406 223576
rect 153194 223564 153200 223576
rect 81400 223536 153200 223564
rect 81400 223524 81406 223536
rect 153194 223524 153200 223536
rect 153252 223524 153258 223576
rect 154942 223564 154948 223576
rect 153396 223536 154948 223564
rect 75822 223388 75828 223440
rect 75880 223428 75886 223440
rect 153396 223428 153424 223536
rect 154942 223524 154948 223536
rect 155000 223524 155006 223576
rect 155770 223524 155776 223576
rect 155828 223564 155834 223576
rect 159818 223564 159824 223576
rect 155828 223536 159824 223564
rect 155828 223524 155834 223536
rect 159818 223524 159824 223536
rect 159876 223524 159882 223576
rect 165614 223524 165620 223576
rect 165672 223564 165678 223576
rect 171962 223564 171968 223576
rect 165672 223536 171968 223564
rect 165672 223524 165678 223536
rect 171962 223524 171968 223536
rect 172020 223524 172026 223576
rect 175274 223524 175280 223576
rect 175332 223564 175338 223576
rect 176562 223564 176568 223576
rect 175332 223536 176568 223564
rect 175332 223524 175338 223536
rect 176562 223524 176568 223536
rect 176620 223524 176626 223576
rect 186590 223564 186596 223576
rect 183756 223536 186596 223564
rect 75880 223400 153424 223428
rect 75880 223388 75886 223400
rect 154206 223388 154212 223440
rect 154264 223428 154270 223440
rect 156782 223428 156788 223440
rect 154264 223400 156788 223428
rect 154264 223388 154270 223400
rect 156782 223388 156788 223400
rect 156840 223388 156846 223440
rect 158714 223388 158720 223440
rect 158772 223428 158778 223440
rect 181714 223428 181720 223440
rect 158772 223400 181720 223428
rect 158772 223388 158778 223400
rect 181714 223388 181720 223400
rect 181772 223388 181778 223440
rect 69566 223252 69572 223304
rect 69624 223292 69630 223304
rect 142108 223292 142114 223304
rect 69624 223264 142114 223292
rect 69624 223252 69630 223264
rect 142108 223252 142114 223264
rect 142166 223252 142172 223304
rect 146662 223292 146668 223304
rect 142264 223264 146668 223292
rect 66898 223116 66904 223168
rect 66956 223156 66962 223168
rect 142264 223156 142292 223264
rect 146662 223252 146668 223264
rect 146720 223252 146726 223304
rect 146938 223252 146944 223304
rect 146996 223292 147002 223304
rect 152090 223292 152096 223304
rect 146996 223264 152096 223292
rect 146996 223252 147002 223264
rect 152090 223252 152096 223264
rect 152148 223252 152154 223304
rect 153194 223252 153200 223304
rect 153252 223292 153258 223304
rect 155770 223292 155776 223304
rect 153252 223264 155776 223292
rect 153252 223252 153258 223264
rect 155770 223252 155776 223264
rect 155828 223252 155834 223304
rect 156414 223252 156420 223304
rect 156472 223292 156478 223304
rect 161934 223292 161940 223304
rect 156472 223264 161940 223292
rect 156472 223252 156478 223264
rect 161934 223252 161940 223264
rect 161992 223252 161998 223304
rect 162486 223252 162492 223304
rect 162544 223292 162550 223304
rect 183756 223292 183784 223536
rect 186590 223524 186596 223536
rect 186648 223524 186654 223576
rect 187326 223524 187332 223576
rect 187384 223564 187390 223576
rect 242250 223564 242256 223576
rect 187384 223536 242256 223564
rect 187384 223524 187390 223536
rect 242250 223524 242256 223536
rect 242308 223524 242314 223576
rect 250898 223524 250904 223576
rect 250956 223564 250962 223576
rect 291194 223564 291200 223576
rect 250956 223536 291200 223564
rect 250956 223524 250962 223536
rect 291194 223524 291200 223536
rect 291252 223524 291258 223576
rect 297910 223524 297916 223576
rect 297968 223564 297974 223576
rect 303246 223564 303252 223576
rect 297968 223536 303252 223564
rect 297968 223524 297974 223536
rect 303246 223524 303252 223536
rect 303304 223524 303310 223576
rect 307662 223524 307668 223576
rect 307720 223564 307726 223576
rect 335630 223564 335636 223576
rect 307720 223536 335636 223564
rect 307720 223524 307726 223536
rect 335630 223524 335636 223536
rect 335688 223524 335694 223576
rect 406746 223524 406752 223576
rect 406804 223564 406810 223576
rect 414842 223564 414848 223576
rect 406804 223536 414848 223564
rect 406804 223524 406810 223536
rect 414842 223524 414848 223536
rect 414900 223524 414906 223576
rect 454862 223524 454868 223576
rect 454920 223564 454926 223576
rect 460474 223564 460480 223576
rect 454920 223536 460480 223564
rect 454920 223524 454926 223536
rect 460474 223524 460480 223536
rect 460532 223524 460538 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 342070 223496 342076 223508
rect 335832 223468 342076 223496
rect 184658 223388 184664 223440
rect 184716 223428 184722 223440
rect 239674 223428 239680 223440
rect 184716 223400 239680 223428
rect 184716 223388 184722 223400
rect 239674 223388 239680 223400
rect 239732 223388 239738 223440
rect 244090 223388 244096 223440
rect 244148 223428 244154 223440
rect 286042 223428 286048 223440
rect 244148 223400 286048 223428
rect 244148 223388 244154 223400
rect 286042 223388 286048 223400
rect 286100 223388 286106 223440
rect 304718 223388 304724 223440
rect 304776 223428 304782 223440
rect 308122 223428 308128 223440
rect 304776 223400 308128 223428
rect 304776 223388 304782 223400
rect 308122 223388 308128 223400
rect 308180 223388 308186 223440
rect 312906 223388 312912 223440
rect 312964 223428 312970 223440
rect 312964 223400 335354 223428
rect 312964 223388 312970 223400
rect 335326 223360 335354 223400
rect 335832 223360 335860 223468
rect 342070 223456 342076 223468
rect 342128 223456 342134 223508
rect 670712 223468 671048 223496
rect 342806 223388 342812 223440
rect 342864 223428 342870 223440
rect 347866 223428 347872 223440
rect 342864 223400 347872 223428
rect 342864 223388 342870 223400
rect 347866 223388 347872 223400
rect 347924 223388 347930 223440
rect 517514 223388 517520 223440
rect 517572 223428 517578 223440
rect 531498 223428 531504 223440
rect 517572 223400 531504 223428
rect 517572 223388 517578 223400
rect 531498 223388 531504 223400
rect 531556 223388 531562 223440
rect 534810 223388 534816 223440
rect 534868 223428 534874 223440
rect 547414 223428 547420 223440
rect 534868 223400 547420 223428
rect 534868 223388 534874 223400
rect 547414 223388 547420 223400
rect 547472 223388 547478 223440
rect 669268 223388 669274 223440
rect 669326 223428 669332 223440
rect 670712 223428 670740 223468
rect 669326 223400 670740 223428
rect 669326 223388 669332 223400
rect 335326 223332 335860 223360
rect 335998 223320 336004 223372
rect 336056 223360 336062 223372
rect 342254 223360 342260 223372
rect 336056 223332 342260 223360
rect 336056 223320 336062 223332
rect 342254 223320 342260 223332
rect 342312 223320 342318 223372
rect 162544 223264 183784 223292
rect 162544 223252 162550 223264
rect 185394 223252 185400 223304
rect 185452 223292 185458 223304
rect 185452 223264 185808 223292
rect 185452 223252 185458 223264
rect 66956 223128 142292 223156
rect 66956 223116 66962 223128
rect 142430 223116 142436 223168
rect 142488 223156 142494 223168
rect 143994 223156 144000 223168
rect 142488 223128 144000 223156
rect 142488 223116 142494 223128
rect 143994 223116 144000 223128
rect 144052 223116 144058 223168
rect 146570 223116 146576 223168
rect 146628 223156 146634 223168
rect 171594 223156 171600 223168
rect 146628 223128 171600 223156
rect 146628 223116 146634 223128
rect 171594 223116 171600 223128
rect 171652 223116 171658 223168
rect 171778 223116 171784 223168
rect 171836 223156 171842 223168
rect 185578 223156 185584 223168
rect 171836 223128 185584 223156
rect 171836 223116 171842 223128
rect 185578 223116 185584 223128
rect 185636 223116 185642 223168
rect 185780 223156 185808 223264
rect 188890 223252 188896 223304
rect 188948 223292 188954 223304
rect 245102 223292 245108 223304
rect 188948 223264 245108 223292
rect 188948 223252 188954 223264
rect 245102 223252 245108 223264
rect 245160 223252 245166 223304
rect 246850 223252 246856 223304
rect 246908 223292 246914 223304
rect 288618 223292 288624 223304
rect 246908 223264 288624 223292
rect 246908 223252 246914 223264
rect 288618 223252 288624 223264
rect 288676 223252 288682 223304
rect 289722 223252 289728 223304
rect 289780 223292 289786 223304
rect 297726 223292 297732 223304
rect 289780 223264 297732 223292
rect 289780 223252 289786 223264
rect 297726 223252 297732 223264
rect 297784 223252 297790 223304
rect 299106 223252 299112 223304
rect 299164 223292 299170 223304
rect 328546 223292 328552 223304
rect 299164 223264 328552 223292
rect 299164 223252 299170 223264
rect 328546 223252 328552 223264
rect 328604 223252 328610 223304
rect 347222 223252 347228 223304
rect 347280 223292 347286 223304
rect 357894 223292 357900 223304
rect 347280 223264 357900 223292
rect 347280 223252 347286 223264
rect 357894 223252 357900 223264
rect 357952 223252 357958 223304
rect 483106 223252 483112 223304
rect 483164 223292 483170 223304
rect 496078 223292 496084 223304
rect 483164 223264 496084 223292
rect 483164 223252 483170 223264
rect 496078 223252 496084 223264
rect 496136 223252 496142 223304
rect 503346 223252 503352 223304
rect 503404 223292 503410 223304
rect 503404 223264 514064 223292
rect 503404 223252 503410 223264
rect 192018 223156 192024 223168
rect 185780 223128 192024 223156
rect 192018 223116 192024 223128
rect 192076 223116 192082 223168
rect 194318 223116 194324 223168
rect 194376 223156 194382 223168
rect 199746 223156 199752 223168
rect 194376 223128 199752 223156
rect 194376 223116 194382 223128
rect 199746 223116 199752 223128
rect 199804 223116 199810 223168
rect 204254 223116 204260 223168
rect 204312 223156 204318 223168
rect 211982 223156 211988 223168
rect 204312 223128 211988 223156
rect 204312 223116 204318 223128
rect 211982 223116 211988 223128
rect 212040 223116 212046 223168
rect 215386 223116 215392 223168
rect 215444 223156 215450 223168
rect 216214 223156 216220 223168
rect 215444 223128 216220 223156
rect 215444 223116 215450 223128
rect 216214 223116 216220 223128
rect 216272 223116 216278 223168
rect 241330 223116 241336 223168
rect 241388 223156 241394 223168
rect 283466 223156 283472 223168
rect 241388 223128 283472 223156
rect 241388 223116 241394 223128
rect 283466 223116 283472 223128
rect 283524 223116 283530 223168
rect 288250 223116 288256 223168
rect 288308 223156 288314 223168
rect 321094 223156 321100 223168
rect 288308 223128 321100 223156
rect 288308 223116 288314 223128
rect 321094 223116 321100 223128
rect 321152 223116 321158 223168
rect 344646 223116 344652 223168
rect 344704 223156 344710 223168
rect 364610 223156 364616 223168
rect 344704 223128 364616 223156
rect 344704 223116 344710 223128
rect 364610 223116 364616 223128
rect 364668 223116 364674 223168
rect 365530 223116 365536 223168
rect 365588 223156 365594 223168
rect 379606 223156 379612 223168
rect 365588 223128 379612 223156
rect 365588 223116 365594 223128
rect 379606 223116 379612 223128
rect 379664 223116 379670 223168
rect 380066 223116 380072 223168
rect 380124 223156 380130 223168
rect 386506 223156 386512 223168
rect 380124 223128 386512 223156
rect 380124 223116 380130 223128
rect 386506 223116 386512 223128
rect 386564 223116 386570 223168
rect 488626 223116 488632 223168
rect 488684 223156 488690 223168
rect 502702 223156 502708 223168
rect 488684 223128 502708 223156
rect 488684 223116 488690 223128
rect 502702 223116 502708 223128
rect 502760 223116 502766 223168
rect 508222 223116 508228 223168
rect 508280 223156 508286 223168
rect 514036 223156 514064 223264
rect 514662 223252 514668 223304
rect 514720 223292 514726 223304
rect 535454 223292 535460 223304
rect 514720 223264 535460 223292
rect 514720 223252 514726 223264
rect 535454 223252 535460 223264
rect 535512 223252 535518 223304
rect 561950 223252 561956 223304
rect 562008 223292 562014 223304
rect 567838 223292 567844 223304
rect 562008 223264 567844 223292
rect 562008 223252 562014 223264
rect 567838 223252 567844 223264
rect 567896 223252 567902 223304
rect 586974 223252 586980 223304
rect 587032 223292 587038 223304
rect 593966 223292 593972 223304
rect 587032 223264 593972 223292
rect 587032 223252 587038 223264
rect 593966 223252 593972 223264
rect 594024 223252 594030 223304
rect 521746 223156 521752 223168
rect 508280 223128 509234 223156
rect 514036 223128 521752 223156
rect 508280 223116 508286 223128
rect 71406 222980 71412 223032
rect 71464 223020 71470 223032
rect 146938 223020 146944 223032
rect 71464 222992 146944 223020
rect 71464 222980 71470 222992
rect 146938 222980 146944 222992
rect 146996 222980 147002 223032
rect 147122 222980 147128 223032
rect 147180 223020 147186 223032
rect 162118 223020 162124 223032
rect 147180 222992 162124 223020
rect 147180 222980 147186 222992
rect 162118 222980 162124 222992
rect 162176 222980 162182 223032
rect 162302 222980 162308 223032
rect 162360 223020 162366 223032
rect 219710 223020 219716 223032
rect 162360 222992 219716 223020
rect 162360 222980 162366 222992
rect 219710 222980 219716 222992
rect 219768 222980 219774 223032
rect 230198 222980 230204 223032
rect 230256 223020 230262 223032
rect 275462 223020 275468 223032
rect 230256 222992 275468 223020
rect 230256 222980 230262 222992
rect 275462 222980 275468 222992
rect 275520 222980 275526 223032
rect 278590 222980 278596 223032
rect 278648 223020 278654 223032
rect 315022 223020 315028 223032
rect 278648 222992 315028 223020
rect 278648 222980 278654 222992
rect 315022 222980 315028 222992
rect 315080 222980 315086 223032
rect 316678 222980 316684 223032
rect 316736 223020 316742 223032
rect 327258 223020 327264 223032
rect 316736 222992 327264 223020
rect 316736 222980 316742 222992
rect 327258 222980 327264 222992
rect 327316 222980 327322 223032
rect 328086 222980 328092 223032
rect 328144 223020 328150 223032
rect 351454 223020 351460 223032
rect 328144 222992 351460 223020
rect 328144 222980 328150 222992
rect 351454 222980 351460 222992
rect 351512 222980 351518 223032
rect 353938 222980 353944 223032
rect 353996 223020 354002 223032
rect 365898 223020 365904 223032
rect 353996 222992 365904 223020
rect 353996 222980 354002 222992
rect 365898 222980 365904 222992
rect 365956 222980 365962 223032
rect 366910 222980 366916 223032
rect 366968 223020 366974 223032
rect 383838 223020 383844 223032
rect 366968 222992 383844 223020
rect 366968 222980 366974 222992
rect 383838 222980 383844 222992
rect 383896 222980 383902 223032
rect 384206 222980 384212 223032
rect 384264 223020 384270 223032
rect 393958 223020 393964 223032
rect 384264 222992 393964 223020
rect 384264 222980 384270 222992
rect 393958 222980 393964 222992
rect 394016 222980 394022 223032
rect 493042 222980 493048 223032
rect 493100 223020 493106 223032
rect 508590 223020 508596 223032
rect 493100 222992 508596 223020
rect 493100 222980 493106 222992
rect 508590 222980 508596 222992
rect 508648 222980 508654 223032
rect 509206 223020 509234 223128
rect 521746 223116 521752 223128
rect 521804 223116 521810 223168
rect 532050 223116 532056 223168
rect 532108 223156 532114 223168
rect 559006 223156 559012 223168
rect 532108 223128 559012 223156
rect 532108 223116 532114 223128
rect 559006 223116 559012 223128
rect 559064 223116 559070 223168
rect 562318 223116 562324 223168
rect 562376 223156 562382 223168
rect 587158 223156 587164 223168
rect 562376 223128 587164 223156
rect 562376 223116 562382 223128
rect 587158 223116 587164 223128
rect 587216 223116 587222 223168
rect 667750 223116 667756 223168
rect 667808 223156 667814 223168
rect 667808 223128 670956 223156
rect 667808 223116 667814 223128
rect 527818 223020 527824 223032
rect 509206 222992 527824 223020
rect 527818 222980 527824 222992
rect 527876 222980 527882 223032
rect 529474 222980 529480 223032
rect 529532 223020 529538 223032
rect 555694 223020 555700 223032
rect 529532 222992 555700 223020
rect 529532 222980 529538 222992
rect 555694 222980 555700 222992
rect 555752 222980 555758 223032
rect 557534 222980 557540 223032
rect 557592 223020 557598 223032
rect 559834 223020 559840 223032
rect 557592 222992 559840 223020
rect 557592 222980 557598 222992
rect 559834 222980 559840 222992
rect 559892 223020 559898 223032
rect 627086 223020 627092 223032
rect 559892 222992 627092 223020
rect 559892 222980 559898 222992
rect 627086 222980 627092 222992
rect 627144 222980 627150 223032
rect 62758 222844 62764 222896
rect 62816 222884 62822 222896
rect 141970 222884 141976 222896
rect 62816 222856 141976 222884
rect 62816 222844 62822 222856
rect 141970 222844 141976 222856
rect 142028 222844 142034 222896
rect 142154 222844 142160 222896
rect 142212 222884 142218 222896
rect 156598 222884 156604 222896
rect 142212 222856 156604 222884
rect 142212 222844 142218 222856
rect 156598 222844 156604 222856
rect 156656 222844 156662 222896
rect 156782 222844 156788 222896
rect 156840 222884 156846 222896
rect 215386 222884 215392 222896
rect 156840 222856 215392 222884
rect 156840 222844 156846 222856
rect 215386 222844 215392 222856
rect 215444 222844 215450 222896
rect 215938 222844 215944 222896
rect 215996 222884 216002 222896
rect 233326 222884 233332 222896
rect 215996 222856 233332 222884
rect 215996 222844 216002 222856
rect 233326 222844 233332 222856
rect 233384 222844 233390 222896
rect 234522 222844 234528 222896
rect 234580 222884 234586 222896
rect 281534 222884 281540 222896
rect 234580 222856 281540 222884
rect 234580 222844 234586 222856
rect 281534 222844 281540 222856
rect 281592 222844 281598 222896
rect 282454 222844 282460 222896
rect 282512 222884 282518 222896
rect 316310 222884 316316 222896
rect 282512 222856 316316 222884
rect 282512 222844 282518 222856
rect 316310 222844 316316 222856
rect 316368 222844 316374 222896
rect 324130 222844 324136 222896
rect 324188 222884 324194 222896
rect 348510 222884 348516 222896
rect 324188 222856 348516 222884
rect 324188 222844 324194 222856
rect 348510 222844 348516 222856
rect 348568 222844 348574 222896
rect 349062 222844 349068 222896
rect 349120 222884 349126 222896
rect 367186 222884 367192 222896
rect 349120 222856 367192 222884
rect 349120 222844 349126 222856
rect 367186 222844 367192 222856
rect 367244 222844 367250 222896
rect 368382 222844 368388 222896
rect 368440 222884 368446 222896
rect 382366 222884 382372 222896
rect 368440 222856 382372 222884
rect 368440 222844 368446 222856
rect 382366 222844 382372 222856
rect 382424 222844 382430 222896
rect 383470 222844 383476 222896
rect 383528 222884 383534 222896
rect 394878 222884 394884 222896
rect 383528 222856 394884 222884
rect 383528 222844 383534 222856
rect 394878 222844 394884 222856
rect 394936 222844 394942 222896
rect 395798 222844 395804 222896
rect 395856 222884 395862 222896
rect 406470 222884 406476 222896
rect 395856 222856 406476 222884
rect 395856 222844 395862 222856
rect 406470 222844 406476 222856
rect 406528 222844 406534 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 479886 222844 479892 222896
rect 479944 222884 479950 222896
rect 491938 222884 491944 222896
rect 479944 222856 491944 222884
rect 479944 222844 479950 222856
rect 491938 222844 491944 222856
rect 491996 222844 492002 222896
rect 500770 222844 500776 222896
rect 500828 222884 500834 222896
rect 517514 222884 517520 222896
rect 500828 222856 517520 222884
rect 500828 222844 500834 222856
rect 517514 222844 517520 222856
rect 517572 222844 517578 222896
rect 519814 222844 519820 222896
rect 519872 222884 519878 222896
rect 543366 222884 543372 222896
rect 519872 222856 543372 222884
rect 519872 222844 519878 222856
rect 543366 222844 543372 222856
rect 543424 222844 543430 222896
rect 554038 222844 554044 222896
rect 554096 222884 554102 222896
rect 632698 222884 632704 222896
rect 554096 222856 632704 222884
rect 554096 222844 554102 222856
rect 632698 222844 632704 222856
rect 632756 222844 632762 222896
rect 651282 222844 651288 222896
rect 651340 222884 651346 222896
rect 666462 222884 666468 222896
rect 651340 222856 666468 222884
rect 651340 222844 651346 222856
rect 666462 222844 666468 222856
rect 666520 222844 666526 222896
rect 78582 222708 78588 222760
rect 78640 222748 78646 222760
rect 155126 222748 155132 222760
rect 78640 222720 155132 222748
rect 78640 222708 78646 222720
rect 155126 222708 155132 222720
rect 155184 222708 155190 222760
rect 155678 222708 155684 222760
rect 155736 222748 155742 222760
rect 161934 222748 161940 222760
rect 155736 222720 161940 222748
rect 155736 222708 155742 222720
rect 161934 222708 161940 222720
rect 161992 222708 161998 222760
rect 162118 222708 162124 222760
rect 162176 222748 162182 222760
rect 171778 222748 171784 222760
rect 162176 222720 171784 222748
rect 162176 222708 162182 222720
rect 171778 222708 171784 222720
rect 171836 222708 171842 222760
rect 171962 222708 171968 222760
rect 172020 222748 172026 222760
rect 185394 222748 185400 222760
rect 172020 222720 185400 222748
rect 172020 222708 172026 222720
rect 185394 222708 185400 222720
rect 185452 222708 185458 222760
rect 185578 222708 185584 222760
rect 185636 222748 185642 222760
rect 204254 222748 204260 222760
rect 185636 222720 204260 222748
rect 185636 222708 185642 222720
rect 204254 222708 204260 222720
rect 204312 222708 204318 222760
rect 204438 222708 204444 222760
rect 204496 222748 204502 222760
rect 247402 222748 247408 222760
rect 204496 222720 247408 222748
rect 204496 222708 204502 222720
rect 247402 222708 247408 222720
rect 247460 222708 247466 222760
rect 264790 222708 264796 222760
rect 264848 222748 264854 222760
rect 304350 222748 304356 222760
rect 264848 222720 304356 222748
rect 264848 222708 264854 222720
rect 304350 222708 304356 222720
rect 304408 222708 304414 222760
rect 543826 222708 543832 222760
rect 543884 222748 543890 222760
rect 552382 222748 552388 222760
rect 543884 222720 552388 222748
rect 543884 222708 543890 222720
rect 552382 222708 552388 222720
rect 552440 222748 552446 222760
rect 625614 222748 625620 222760
rect 552440 222720 625620 222748
rect 552440 222708 552446 222720
rect 625614 222708 625620 222720
rect 625672 222708 625678 222760
rect 99282 222572 99288 222624
rect 99340 222612 99346 222624
rect 99340 222584 166994 222612
rect 99340 222572 99346 222584
rect 87966 222436 87972 222488
rect 88024 222476 88030 222488
rect 164970 222476 164976 222488
rect 88024 222448 164976 222476
rect 88024 222436 88030 222448
rect 164970 222436 164976 222448
rect 165028 222436 165034 222488
rect 166966 222476 166994 222584
rect 171594 222572 171600 222624
rect 171652 222612 171658 222624
rect 175274 222612 175280 222624
rect 171652 222584 175280 222612
rect 171652 222572 171658 222584
rect 175274 222572 175280 222584
rect 175332 222572 175338 222624
rect 197170 222572 197176 222624
rect 197228 222612 197234 222624
rect 249978 222612 249984 222624
rect 197228 222584 249984 222612
rect 197228 222572 197234 222584
rect 249978 222572 249984 222584
rect 250036 222572 250042 222624
rect 529842 222572 529848 222624
rect 529900 222612 529906 222624
rect 619910 222612 619916 222624
rect 529900 222584 619916 222612
rect 529900 222572 529906 222584
rect 619910 222572 619916 222584
rect 619968 222572 619974 222624
rect 176010 222504 176016 222556
rect 176068 222544 176074 222556
rect 176068 222516 190454 222544
rect 176068 222504 176074 222516
rect 175642 222476 175648 222488
rect 166966 222448 175648 222476
rect 175642 222436 175648 222448
rect 175700 222436 175706 222488
rect 190426 222476 190454 222516
rect 207474 222476 207480 222488
rect 190426 222448 207480 222476
rect 207474 222436 207480 222448
rect 207532 222436 207538 222488
rect 207658 222436 207664 222488
rect 207716 222476 207722 222488
rect 258350 222476 258356 222488
rect 207716 222448 258356 222476
rect 207716 222436 207722 222448
rect 258350 222436 258356 222448
rect 258408 222436 258414 222488
rect 562318 222476 562324 222488
rect 485746 222448 562324 222476
rect 175826 222368 175832 222420
rect 175884 222408 175890 222420
rect 175884 222380 185716 222408
rect 175884 222368 175890 222380
rect 85298 222300 85304 222352
rect 85356 222340 85362 222352
rect 156414 222340 156420 222352
rect 85356 222312 156420 222340
rect 85356 222300 85362 222312
rect 156414 222300 156420 222312
rect 156472 222300 156478 222352
rect 185688 222340 185716 222380
rect 194318 222340 194324 222352
rect 185688 222312 194324 222340
rect 194318 222300 194324 222312
rect 194376 222300 194382 222352
rect 194502 222300 194508 222352
rect 194560 222340 194566 222352
rect 204438 222340 204444 222352
rect 194560 222312 204444 222340
rect 194560 222300 194566 222312
rect 204438 222300 204444 222312
rect 204496 222300 204502 222352
rect 211798 222300 211804 222352
rect 211856 222340 211862 222352
rect 228082 222340 228088 222352
rect 211856 222312 228088 222340
rect 211856 222300 211862 222312
rect 228082 222300 228088 222312
rect 228140 222300 228146 222352
rect 287882 222300 287888 222352
rect 287940 222340 287946 222352
rect 295058 222340 295064 222352
rect 287940 222312 295064 222340
rect 287940 222300 287946 222312
rect 295058 222300 295064 222312
rect 295116 222300 295122 222352
rect 484486 222300 484492 222352
rect 484544 222340 484550 222352
rect 485746 222340 485774 222448
rect 562318 222436 562324 222448
rect 562376 222436 562382 222488
rect 567838 222436 567844 222488
rect 567896 222476 567902 222488
rect 627914 222476 627920 222488
rect 567896 222448 627920 222476
rect 567896 222436 567902 222448
rect 627914 222436 627920 222448
rect 627972 222436 627978 222488
rect 484544 222312 485774 222340
rect 484544 222300 484550 222312
rect 489914 222300 489920 222352
rect 489972 222340 489978 222352
rect 491110 222340 491116 222352
rect 489972 222312 491116 222340
rect 489972 222300 489978 222312
rect 491110 222300 491116 222312
rect 491168 222340 491174 222352
rect 629846 222340 629852 222352
rect 491168 222312 629852 222340
rect 491168 222300 491174 222312
rect 629846 222300 629852 222312
rect 629904 222300 629910 222352
rect 156598 222232 156604 222284
rect 156656 222272 156662 222284
rect 156656 222244 185624 222272
rect 156656 222232 156662 222244
rect 185596 222204 185624 222244
rect 191006 222204 191012 222216
rect 185596 222176 191012 222204
rect 191006 222164 191012 222176
rect 191064 222164 191070 222216
rect 482738 222164 482744 222216
rect 482796 222204 482802 222216
rect 586974 222204 586980 222216
rect 482796 222176 586980 222204
rect 482796 222164 482802 222176
rect 586974 222164 586980 222176
rect 587032 222164 587038 222216
rect 587158 222164 587164 222216
rect 587216 222204 587222 222216
rect 631502 222204 631508 222216
rect 587216 222176 631508 222204
rect 587216 222164 587222 222176
rect 631502 222164 631508 222176
rect 631560 222164 631566 222216
rect 97902 222096 97908 222148
rect 97960 222136 97966 222148
rect 104342 222136 104348 222148
rect 97960 222108 104348 222136
rect 97960 222096 97966 222108
rect 104342 222096 104348 222108
rect 104400 222096 104406 222148
rect 106366 222096 106372 222148
rect 106424 222136 106430 222148
rect 157426 222136 157432 222148
rect 106424 222108 157432 222136
rect 106424 222096 106430 222108
rect 157426 222096 157432 222108
rect 157484 222096 157490 222148
rect 172698 222136 172704 222148
rect 158088 222108 172704 222136
rect 158088 222068 158116 222108
rect 172698 222096 172704 222108
rect 172756 222096 172762 222148
rect 174078 222096 174084 222148
rect 174136 222136 174142 222148
rect 174136 222108 180932 222136
rect 174136 222096 174142 222108
rect 157904 222040 158116 222068
rect 94682 221960 94688 222012
rect 94740 222000 94746 222012
rect 157610 222000 157616 222012
rect 94740 221972 157616 222000
rect 94740 221960 94746 221972
rect 157610 221960 157616 221972
rect 157668 221960 157674 222012
rect 157904 222000 157932 222040
rect 157812 221972 157932 222000
rect 104342 221824 104348 221876
rect 104400 221864 104406 221876
rect 157812 221864 157840 221972
rect 158346 221960 158352 222012
rect 158404 222000 158410 222012
rect 166810 222000 166816 222012
rect 158404 221972 166816 222000
rect 158404 221960 158410 221972
rect 166810 221960 166816 221972
rect 166868 221960 166874 222012
rect 166994 221960 167000 222012
rect 167052 222000 167058 222012
rect 169754 222000 169760 222012
rect 167052 221972 169760 222000
rect 167052 221960 167058 221972
rect 169754 221960 169760 221972
rect 169812 221960 169818 222012
rect 171778 221960 171784 222012
rect 171836 222000 171842 222012
rect 180904 222000 180932 222108
rect 181254 222096 181260 222148
rect 181312 222136 181318 222148
rect 182634 222136 182640 222148
rect 181312 222108 182640 222136
rect 181312 222096 181318 222108
rect 182634 222096 182640 222108
rect 182692 222096 182698 222148
rect 191466 222096 191472 222148
rect 191524 222136 191530 222148
rect 247586 222136 247592 222148
rect 191524 222108 247592 222136
rect 191524 222096 191530 222108
rect 247586 222096 247592 222108
rect 247644 222096 247650 222148
rect 258074 222096 258080 222148
rect 258132 222136 258138 222148
rect 263686 222136 263692 222148
rect 258132 222108 263692 222136
rect 258132 222096 258138 222108
rect 263686 222096 263692 222108
rect 263744 222096 263750 222148
rect 270218 222096 270224 222148
rect 270276 222136 270282 222148
rect 306374 222136 306380 222148
rect 270276 222108 306380 222136
rect 270276 222096 270282 222108
rect 306374 222096 306380 222108
rect 306432 222096 306438 222148
rect 310698 222096 310704 222148
rect 310756 222136 310762 222148
rect 312630 222136 312636 222148
rect 310756 222108 312636 222136
rect 310756 222096 310762 222108
rect 312630 222096 312636 222108
rect 312688 222096 312694 222148
rect 331398 222096 331404 222148
rect 331456 222136 331462 222148
rect 353754 222136 353760 222148
rect 331456 222108 353760 222136
rect 331456 222096 331462 222108
rect 353754 222096 353760 222108
rect 353812 222096 353818 222148
rect 424962 222096 424968 222148
rect 425020 222136 425026 222148
rect 429286 222136 429292 222148
rect 425020 222108 429292 222136
rect 425020 222096 425026 222108
rect 429286 222096 429292 222108
rect 429344 222096 429350 222148
rect 452562 222096 452568 222148
rect 452620 222136 452626 222148
rect 455598 222136 455604 222148
rect 452620 222108 455604 222136
rect 452620 222096 452626 222108
rect 455598 222096 455604 222108
rect 455656 222096 455662 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 495158 222028 495164 222080
rect 495216 222068 495222 222080
rect 497734 222068 497740 222080
rect 495216 222040 497740 222068
rect 495216 222028 495222 222040
rect 497734 222028 497740 222040
rect 497792 222028 497798 222080
rect 515490 222028 515496 222080
rect 515548 222068 515554 222080
rect 529842 222068 529848 222080
rect 515548 222040 529848 222068
rect 515548 222028 515554 222040
rect 529842 222028 529848 222040
rect 529900 222028 529906 222080
rect 533982 222028 533988 222080
rect 534040 222068 534046 222080
rect 559374 222068 559380 222080
rect 534040 222040 559380 222068
rect 534040 222028 534046 222040
rect 559374 222028 559380 222040
rect 559432 222028 559438 222080
rect 559558 222028 559564 222080
rect 559616 222068 559622 222080
rect 564802 222068 564808 222080
rect 559616 222040 564808 222068
rect 559616 222028 559622 222040
rect 564802 222028 564808 222040
rect 564860 222028 564866 222080
rect 231854 222000 231860 222012
rect 171836 221972 180794 222000
rect 180904 221972 231860 222000
rect 171836 221960 171842 221972
rect 104400 221836 157840 221864
rect 104400 221824 104406 221836
rect 158162 221824 158168 221876
rect 158220 221864 158226 221876
rect 176562 221864 176568 221876
rect 158220 221836 176568 221864
rect 158220 221824 158226 221836
rect 176562 221824 176568 221836
rect 176620 221824 176626 221876
rect 180766 221864 180794 221972
rect 231854 221960 231860 221972
rect 231912 221960 231918 222012
rect 233694 221960 233700 222012
rect 233752 222000 233758 222012
rect 277946 222000 277952 222012
rect 233752 221972 277952 222000
rect 233752 221960 233758 221972
rect 277946 221960 277952 221972
rect 278004 221960 278010 222012
rect 280062 221960 280068 222012
rect 280120 222000 280126 222012
rect 313734 222000 313740 222012
rect 280120 221972 313740 222000
rect 280120 221960 280126 221972
rect 313734 221960 313740 221972
rect 313792 221960 313798 222012
rect 318242 221960 318248 222012
rect 318300 222000 318306 222012
rect 343818 222000 343824 222012
rect 318300 221972 343824 222000
rect 318300 221960 318306 221972
rect 343818 221960 343824 221972
rect 343876 221960 343882 222012
rect 367646 221960 367652 222012
rect 367704 222000 367710 222012
rect 380250 222000 380256 222012
rect 367704 221972 380256 222000
rect 367704 221960 367710 221972
rect 380250 221960 380256 221972
rect 380308 221960 380314 222012
rect 600590 222000 600596 222012
rect 582346 221972 600596 222000
rect 536098 221892 536104 221944
rect 536156 221932 536162 221944
rect 543688 221932 543694 221944
rect 536156 221904 543694 221932
rect 536156 221892 536162 221904
rect 543688 221892 543694 221904
rect 543746 221892 543752 221944
rect 547138 221892 547144 221944
rect 547196 221932 547202 221944
rect 556982 221932 556988 221944
rect 547196 221904 556988 221932
rect 547196 221892 547202 221904
rect 556982 221892 556988 221904
rect 557040 221892 557046 221944
rect 562318 221932 562324 221944
rect 557506 221904 562324 221932
rect 181254 221864 181260 221876
rect 180766 221836 181260 221864
rect 181254 221824 181260 221836
rect 181312 221824 181318 221876
rect 181622 221824 181628 221876
rect 181680 221864 181686 221876
rect 240134 221864 240140 221876
rect 181680 221836 240140 221864
rect 181680 221824 181686 221836
rect 240134 221824 240140 221836
rect 240192 221824 240198 221876
rect 263318 221824 263324 221876
rect 263376 221864 263382 221876
rect 301222 221864 301228 221876
rect 263376 221836 301228 221864
rect 263376 221824 263382 221836
rect 301222 221824 301228 221836
rect 301280 221824 301286 221876
rect 301958 221824 301964 221876
rect 302016 221864 302022 221876
rect 310882 221864 310888 221876
rect 302016 221836 310888 221864
rect 302016 221824 302022 221836
rect 310882 221824 310888 221836
rect 310940 221824 310946 221876
rect 313182 221824 313188 221876
rect 313240 221864 313246 221876
rect 340414 221864 340420 221876
rect 313240 221836 340420 221864
rect 313240 221824 313246 221836
rect 340414 221824 340420 221836
rect 340472 221824 340478 221876
rect 351270 221824 351276 221876
rect 351328 221864 351334 221876
rect 369302 221864 369308 221876
rect 351328 221836 369308 221864
rect 351328 221824 351334 221836
rect 369302 221824 369308 221836
rect 369360 221824 369366 221876
rect 509878 221824 509884 221876
rect 509936 221864 509942 221876
rect 522574 221864 522580 221876
rect 509936 221836 522580 221864
rect 509936 221824 509942 221836
rect 522574 221824 522580 221836
rect 522632 221824 522638 221876
rect 546954 221864 546960 221876
rect 544166 221836 546960 221864
rect 544166 221796 544194 221836
rect 546954 221824 546960 221836
rect 547012 221824 547018 221876
rect 557350 221824 557356 221876
rect 557408 221864 557414 221876
rect 557506 221864 557534 221904
rect 562318 221892 562324 221904
rect 562376 221892 562382 221944
rect 582346 221864 582374 221972
rect 600590 221960 600596 221972
rect 600648 221960 600654 222012
rect 600958 221960 600964 222012
rect 601016 222000 601022 222012
rect 606662 222000 606668 222012
rect 601016 221972 606668 222000
rect 601016 221960 601022 221972
rect 606662 221960 606668 221972
rect 606720 221960 606726 222012
rect 557408 221836 557534 221864
rect 562520 221836 582374 221864
rect 557408 221824 557414 221836
rect 543844 221768 544194 221796
rect 80514 221688 80520 221740
rect 80572 221728 80578 221740
rect 86218 221728 86224 221740
rect 80572 221700 86224 221728
rect 80572 221688 80578 221700
rect 86218 221688 86224 221700
rect 86276 221688 86282 221740
rect 91278 221688 91284 221740
rect 91336 221728 91342 221740
rect 167178 221728 167184 221740
rect 91336 221700 167184 221728
rect 91336 221688 91342 221700
rect 167178 221688 167184 221700
rect 167236 221688 167242 221740
rect 167454 221688 167460 221740
rect 167512 221728 167518 221740
rect 171410 221728 171416 221740
rect 167512 221700 171416 221728
rect 167512 221688 167518 221700
rect 171410 221688 171416 221700
rect 171468 221688 171474 221740
rect 171594 221688 171600 221740
rect 171652 221728 171658 221740
rect 232222 221728 232228 221740
rect 171652 221700 232228 221728
rect 171652 221688 171658 221700
rect 232222 221688 232228 221700
rect 232280 221688 232286 221740
rect 239306 221688 239312 221740
rect 239364 221728 239370 221740
rect 283650 221728 283656 221740
rect 239364 221700 283656 221728
rect 239364 221688 239370 221700
rect 283650 221688 283656 221700
rect 283708 221688 283714 221740
rect 303246 221688 303252 221740
rect 303304 221728 303310 221740
rect 332778 221728 332784 221740
rect 303304 221700 332784 221728
rect 303304 221688 303310 221700
rect 332778 221688 332784 221700
rect 332836 221688 332842 221740
rect 357158 221688 357164 221740
rect 357216 221728 357222 221740
rect 374638 221728 374644 221740
rect 357216 221700 374644 221728
rect 357216 221688 357222 221700
rect 374638 221688 374644 221700
rect 374696 221688 374702 221740
rect 391014 221688 391020 221740
rect 391072 221728 391078 221740
rect 400398 221728 400404 221740
rect 391072 221700 400404 221728
rect 391072 221688 391078 221700
rect 400398 221688 400404 221700
rect 400456 221688 400462 221740
rect 475930 221688 475936 221740
rect 475988 221728 475994 221740
rect 486142 221728 486148 221740
rect 475988 221700 486148 221728
rect 475988 221688 475994 221700
rect 486142 221688 486148 221700
rect 486200 221688 486206 221740
rect 496262 221688 496268 221740
rect 496320 221728 496326 221740
rect 513558 221728 513564 221740
rect 496320 221700 513564 221728
rect 496320 221688 496326 221700
rect 513558 221688 513564 221700
rect 513616 221688 513622 221740
rect 524230 221688 524236 221740
rect 524288 221728 524294 221740
rect 543844 221728 543872 221768
rect 524288 221700 543872 221728
rect 524288 221688 524294 221700
rect 544286 221688 544292 221740
rect 544344 221728 544350 221740
rect 562520 221728 562548 221836
rect 596818 221824 596824 221876
rect 596876 221864 596882 221876
rect 633434 221864 633440 221876
rect 596876 221836 633440 221864
rect 596876 221824 596882 221836
rect 633434 221824 633440 221836
rect 633492 221824 633498 221876
rect 544344 221700 562548 221728
rect 544344 221688 544350 221700
rect 562686 221688 562692 221740
rect 562744 221728 562750 221740
rect 608594 221728 608600 221740
rect 562744 221700 608600 221728
rect 562744 221688 562750 221700
rect 608594 221688 608600 221700
rect 608652 221688 608658 221740
rect 73890 221552 73896 221604
rect 73948 221592 73954 221604
rect 82078 221592 82084 221604
rect 73948 221564 82084 221592
rect 73948 221552 73954 221564
rect 82078 221552 82084 221564
rect 82136 221552 82142 221604
rect 86310 221552 86316 221604
rect 86368 221592 86374 221604
rect 160830 221592 160836 221604
rect 86368 221564 160836 221592
rect 86368 221552 86374 221564
rect 160830 221552 160836 221564
rect 160888 221552 160894 221604
rect 162118 221552 162124 221604
rect 162176 221592 162182 221604
rect 202506 221592 202512 221604
rect 162176 221564 202512 221592
rect 162176 221552 162182 221564
rect 202506 221552 202512 221564
rect 202564 221552 202570 221604
rect 205726 221592 205732 221604
rect 202892 221564 205732 221592
rect 59354 221416 59360 221468
rect 59412 221456 59418 221468
rect 140774 221456 140780 221468
rect 59412 221428 140780 221456
rect 59412 221416 59418 221428
rect 140774 221416 140780 221428
rect 140832 221416 140838 221468
rect 140958 221416 140964 221468
rect 141016 221456 141022 221468
rect 202892 221456 202920 221564
rect 205726 221552 205732 221564
rect 205784 221552 205790 221604
rect 208394 221552 208400 221604
rect 208452 221592 208458 221604
rect 260834 221592 260840 221604
rect 208452 221564 260840 221592
rect 208452 221552 208458 221564
rect 260834 221552 260840 221564
rect 260892 221552 260898 221604
rect 261018 221552 261024 221604
rect 261076 221592 261082 221604
rect 301774 221592 301780 221604
rect 261076 221564 301780 221592
rect 261076 221552 261082 221564
rect 301774 221552 301780 221564
rect 301832 221552 301838 221604
rect 308858 221552 308864 221604
rect 308916 221592 308922 221604
rect 339678 221592 339684 221604
rect 308916 221564 339684 221592
rect 308916 221552 308922 221564
rect 339678 221552 339684 221564
rect 339736 221552 339742 221604
rect 341334 221552 341340 221604
rect 341392 221592 341398 221604
rect 361758 221592 361764 221604
rect 341392 221564 361764 221592
rect 341392 221552 341398 221564
rect 361758 221552 361764 221564
rect 361816 221552 361822 221604
rect 369486 221552 369492 221604
rect 369544 221592 369550 221604
rect 384022 221592 384028 221604
rect 369544 221564 384028 221592
rect 369544 221552 369550 221564
rect 384022 221552 384028 221564
rect 384080 221552 384086 221604
rect 384390 221552 384396 221604
rect 384448 221592 384454 221604
rect 395154 221592 395160 221604
rect 384448 221564 395160 221592
rect 384448 221552 384454 221564
rect 395154 221552 395160 221564
rect 395212 221552 395218 221604
rect 400582 221552 400588 221604
rect 400640 221592 400646 221604
rect 405826 221592 405832 221604
rect 400640 221564 405832 221592
rect 400640 221552 400646 221564
rect 405826 221552 405832 221564
rect 405884 221552 405890 221604
rect 480806 221552 480812 221604
rect 480864 221592 480870 221604
rect 492950 221592 492956 221604
rect 480864 221564 492956 221592
rect 480864 221552 480870 221564
rect 492950 221552 492956 221564
rect 493008 221552 493014 221604
rect 497458 221552 497464 221604
rect 497516 221592 497522 221604
rect 515122 221592 515128 221604
rect 497516 221564 515128 221592
rect 497516 221552 497522 221564
rect 515122 221552 515128 221564
rect 515180 221552 515186 221604
rect 522850 221552 522856 221604
rect 522908 221592 522914 221604
rect 522908 221564 533476 221592
rect 522908 221552 522914 221564
rect 226518 221456 226524 221468
rect 141016 221428 202920 221456
rect 203352 221428 226524 221456
rect 141016 221416 141022 221428
rect 104526 221280 104532 221332
rect 104584 221320 104590 221332
rect 106366 221320 106372 221332
rect 104584 221292 106372 221320
rect 104584 221280 104590 221292
rect 106366 221280 106372 221292
rect 106424 221280 106430 221332
rect 111150 221280 111156 221332
rect 111208 221320 111214 221332
rect 171778 221320 171784 221332
rect 111208 221292 171784 221320
rect 111208 221280 111214 221292
rect 171778 221280 171784 221292
rect 171836 221280 171842 221332
rect 171962 221280 171968 221332
rect 172020 221320 172026 221332
rect 203352 221320 203380 221428
rect 226518 221416 226524 221428
rect 226576 221416 226582 221468
rect 227898 221416 227904 221468
rect 227956 221456 227962 221468
rect 276106 221456 276112 221468
rect 227956 221428 276112 221456
rect 227956 221416 227962 221428
rect 276106 221416 276112 221428
rect 276164 221416 276170 221468
rect 292482 221416 292488 221468
rect 292540 221456 292546 221468
rect 326246 221456 326252 221468
rect 292540 221428 326252 221456
rect 292540 221416 292546 221428
rect 326246 221416 326252 221428
rect 326304 221416 326310 221468
rect 342162 221416 342168 221468
rect 342220 221456 342226 221468
rect 364794 221456 364800 221468
rect 342220 221428 364800 221456
rect 342220 221416 342226 221428
rect 364794 221416 364800 221428
rect 364852 221416 364858 221468
rect 375282 221416 375288 221468
rect 375340 221456 375346 221468
rect 390738 221456 390744 221468
rect 375340 221428 390744 221456
rect 375340 221416 375346 221428
rect 390738 221416 390744 221428
rect 390796 221416 390802 221468
rect 396810 221416 396816 221468
rect 396868 221456 396874 221468
rect 407298 221456 407304 221468
rect 396868 221428 407304 221456
rect 396868 221416 396874 221428
rect 407298 221416 407304 221428
rect 407356 221416 407362 221468
rect 408402 221416 408408 221468
rect 408460 221456 408466 221468
rect 416866 221456 416872 221468
rect 408460 221428 416872 221456
rect 408460 221416 408466 221428
rect 416866 221416 416872 221428
rect 416924 221416 416930 221468
rect 468938 221416 468944 221468
rect 468996 221456 469002 221468
rect 476206 221456 476212 221468
rect 468996 221428 476212 221456
rect 468996 221416 469002 221428
rect 476206 221416 476212 221428
rect 476264 221416 476270 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 533448 221456 533476 221564
rect 533614 221552 533620 221604
rect 533672 221592 533678 221604
rect 601786 221592 601792 221604
rect 533672 221564 601792 221592
rect 533672 221552 533678 221564
rect 601786 221552 601792 221564
rect 601844 221552 601850 221604
rect 546586 221456 546592 221468
rect 483808 221428 533384 221456
rect 533448 221428 546592 221456
rect 483808 221416 483814 221428
rect 172020 221292 203380 221320
rect 172020 221280 172026 221292
rect 204162 221280 204168 221332
rect 204220 221320 204226 221332
rect 252738 221320 252744 221332
rect 204220 221292 252744 221320
rect 204220 221280 204226 221292
rect 252738 221280 252744 221292
rect 252796 221280 252802 221332
rect 266814 221280 266820 221332
rect 266872 221320 266878 221332
rect 303798 221320 303804 221332
rect 266872 221292 303804 221320
rect 266872 221280 266878 221292
rect 303798 221280 303804 221292
rect 303856 221280 303862 221332
rect 525978 221280 525984 221332
rect 526036 221320 526042 221332
rect 533154 221320 533160 221332
rect 526036 221292 533160 221320
rect 526036 221280 526042 221292
rect 533154 221280 533160 221292
rect 533212 221280 533218 221332
rect 533356 221320 533384 221428
rect 546586 221416 546592 221428
rect 546644 221416 546650 221468
rect 546954 221416 546960 221468
rect 547012 221456 547018 221468
rect 549070 221456 549076 221468
rect 547012 221428 549076 221456
rect 547012 221416 547018 221428
rect 549070 221416 549076 221428
rect 549128 221416 549134 221468
rect 549254 221416 549260 221468
rect 549312 221456 549318 221468
rect 600958 221456 600964 221468
rect 549312 221428 600964 221456
rect 549312 221416 549318 221428
rect 600958 221416 600964 221428
rect 601016 221416 601022 221468
rect 538306 221320 538312 221332
rect 533356 221292 538312 221320
rect 538306 221280 538312 221292
rect 538364 221280 538370 221332
rect 538490 221212 538496 221264
rect 538548 221252 538554 221264
rect 604822 221252 604828 221264
rect 538548 221224 604828 221252
rect 538548 221212 538554 221224
rect 604822 221212 604828 221224
rect 604880 221212 604886 221264
rect 138474 221144 138480 221196
rect 138532 221184 138538 221196
rect 162118 221184 162124 221196
rect 138532 221156 162124 221184
rect 138532 221144 138538 221156
rect 162118 221144 162124 221156
rect 162176 221144 162182 221196
rect 162302 221144 162308 221196
rect 162360 221184 162366 221196
rect 221274 221184 221280 221196
rect 162360 221156 221280 221184
rect 162360 221144 162366 221156
rect 221274 221144 221280 221156
rect 221332 221144 221338 221196
rect 222746 221144 222752 221196
rect 222804 221184 222810 221196
rect 268286 221184 268292 221196
rect 222804 221156 268292 221184
rect 222804 221144 222810 221156
rect 268286 221144 268292 221156
rect 268344 221144 268350 221196
rect 523494 221076 523500 221128
rect 523552 221116 523558 221128
rect 601970 221116 601976 221128
rect 523552 221088 601976 221116
rect 523552 221076 523558 221088
rect 601970 221076 601976 221088
rect 602028 221076 602034 221128
rect 124398 221008 124404 221060
rect 124456 221048 124462 221060
rect 193398 221048 193404 221060
rect 124456 221020 193404 221048
rect 124456 221008 124462 221020
rect 193398 221008 193404 221020
rect 193456 221008 193462 221060
rect 202506 221008 202512 221060
rect 202564 221048 202570 221060
rect 206370 221048 206376 221060
rect 202564 221020 206376 221048
rect 202564 221008 202570 221020
rect 206370 221008 206376 221020
rect 206428 221008 206434 221060
rect 219802 221008 219808 221060
rect 219860 221048 219866 221060
rect 263042 221048 263048 221060
rect 219860 221020 263048 221048
rect 219860 221008 219866 221020
rect 263042 221008 263048 221020
rect 263100 221008 263106 221060
rect 521102 220940 521108 220992
rect 521160 220980 521166 220992
rect 600406 220980 600412 220992
rect 521160 220952 600412 220980
rect 521160 220940 521166 220952
rect 600406 220940 600412 220952
rect 600464 220940 600470 220992
rect 600590 220940 600596 220992
rect 600648 220980 600654 220992
rect 604638 220980 604644 220992
rect 600648 220952 604644 220980
rect 600648 220940 600654 220952
rect 604638 220940 604644 220952
rect 604696 220940 604702 220992
rect 82998 220872 83004 220924
rect 83056 220912 83062 220924
rect 142108 220912 142114 220924
rect 83056 220884 142114 220912
rect 83056 220872 83062 220884
rect 142108 220872 142114 220884
rect 142166 220872 142172 220924
rect 142246 220872 142252 220924
rect 142304 220912 142310 220924
rect 148318 220912 148324 220924
rect 142304 220884 148324 220912
rect 142304 220872 142310 220884
rect 148318 220872 148324 220884
rect 148376 220872 148382 220924
rect 148502 220872 148508 220924
rect 148560 220912 148566 220924
rect 151170 220912 151176 220924
rect 148560 220884 151176 220912
rect 148560 220872 148566 220884
rect 151170 220872 151176 220884
rect 151228 220872 151234 220924
rect 158346 220872 158352 220924
rect 158404 220912 158410 220924
rect 160646 220912 160652 220924
rect 158404 220884 160652 220912
rect 158404 220872 158410 220884
rect 160646 220872 160652 220884
rect 160704 220872 160710 220924
rect 160830 220872 160836 220924
rect 160888 220912 160894 220924
rect 164326 220912 164332 220924
rect 160888 220884 164332 220912
rect 160888 220872 160894 220884
rect 164326 220872 164332 220884
rect 164384 220872 164390 220924
rect 164510 220872 164516 220924
rect 164568 220912 164574 220924
rect 222286 220912 222292 220924
rect 164568 220884 222292 220912
rect 164568 220872 164574 220884
rect 222286 220872 222292 220884
rect 222344 220872 222350 220924
rect 282638 220872 282644 220924
rect 282696 220912 282702 220924
rect 287698 220912 287704 220924
rect 282696 220884 287704 220912
rect 282696 220872 282702 220884
rect 287698 220872 287704 220884
rect 287756 220872 287762 220924
rect 456702 220872 456708 220924
rect 456760 220912 456766 220924
rect 456760 220884 460934 220912
rect 456760 220872 456766 220884
rect 253842 220804 253848 220856
rect 253900 220844 253906 220856
rect 258626 220844 258632 220856
rect 253900 220816 258632 220844
rect 253900 220804 253906 220816
rect 258626 220804 258632 220816
rect 258684 220804 258690 220856
rect 418338 220804 418344 220856
rect 418396 220844 418402 220856
rect 424042 220844 424048 220856
rect 418396 220816 424048 220844
rect 418396 220804 418402 220816
rect 424042 220804 424048 220816
rect 424100 220804 424106 220856
rect 460906 220844 460934 220884
rect 466086 220872 466092 220924
rect 466144 220912 466150 220924
rect 471422 220912 471428 220924
rect 466144 220884 471428 220912
rect 466144 220872 466150 220884
rect 471422 220872 471428 220884
rect 471480 220872 471486 220924
rect 462130 220844 462136 220856
rect 460906 220816 462136 220844
rect 462130 220804 462136 220816
rect 462188 220804 462194 220856
rect 517514 220804 517520 220856
rect 517572 220844 517578 220856
rect 518526 220844 518532 220856
rect 517572 220816 518532 220844
rect 517572 220804 517578 220816
rect 518526 220804 518532 220816
rect 518584 220844 518590 220856
rect 600682 220844 600688 220856
rect 518584 220816 600688 220844
rect 518584 220804 518590 220816
rect 600682 220804 600688 220816
rect 600740 220804 600746 220856
rect 114278 220736 114284 220788
rect 114336 220776 114342 220788
rect 146754 220776 146760 220788
rect 114336 220748 146760 220776
rect 114336 220736 114342 220748
rect 146754 220736 146760 220748
rect 146812 220736 146818 220788
rect 146938 220736 146944 220788
rect 146996 220776 147002 220788
rect 180748 220776 180754 220788
rect 146996 220748 180754 220776
rect 146996 220736 147002 220748
rect 180748 220736 180754 220748
rect 180806 220736 180812 220788
rect 181254 220736 181260 220788
rect 181312 220776 181318 220788
rect 190270 220776 190276 220788
rect 181312 220748 190276 220776
rect 181312 220736 181318 220748
rect 190270 220736 190276 220748
rect 190328 220736 190334 220788
rect 190408 220736 190414 220788
rect 190466 220776 190472 220788
rect 236638 220776 236644 220788
rect 190466 220748 236644 220776
rect 190466 220736 190472 220748
rect 236638 220736 236644 220748
rect 236696 220736 236702 220788
rect 242618 220736 242624 220788
rect 242676 220776 242682 220788
rect 246482 220776 246488 220788
rect 242676 220748 246488 220776
rect 242676 220736 242682 220748
rect 246482 220736 246488 220748
rect 246540 220736 246546 220788
rect 260190 220736 260196 220788
rect 260248 220776 260254 220788
rect 298554 220776 298560 220788
rect 260248 220748 298560 220776
rect 260248 220736 260254 220748
rect 298554 220736 298560 220748
rect 298612 220736 298618 220788
rect 321554 220736 321560 220788
rect 321612 220776 321618 220788
rect 324498 220776 324504 220788
rect 321612 220748 324504 220776
rect 321612 220736 321618 220748
rect 324498 220736 324504 220748
rect 324556 220736 324562 220788
rect 385218 220736 385224 220788
rect 385276 220776 385282 220788
rect 388714 220776 388720 220788
rect 385276 220748 388720 220776
rect 385276 220736 385282 220748
rect 388714 220736 388720 220748
rect 388772 220736 388778 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418154 220776 418160 220788
rect 414256 220748 418160 220776
rect 414256 220736 414262 220748
rect 418154 220736 418160 220748
rect 418212 220736 418218 220788
rect 455322 220736 455328 220788
rect 455380 220776 455386 220788
rect 458818 220776 458824 220788
rect 455380 220748 458824 220776
rect 455380 220736 455386 220748
rect 458818 220736 458824 220748
rect 458876 220736 458882 220788
rect 465718 220736 465724 220788
rect 465776 220776 465782 220788
rect 469582 220776 469588 220788
rect 465776 220748 469588 220776
rect 465776 220736 465782 220748
rect 469582 220736 469588 220748
rect 469640 220736 469646 220788
rect 473998 220736 474004 220788
rect 474056 220776 474062 220788
rect 475378 220776 475384 220788
rect 474056 220748 475384 220776
rect 474056 220736 474062 220748
rect 475378 220736 475384 220748
rect 475436 220736 475442 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 511810 220736 511816 220788
rect 511868 220776 511874 220788
rect 511868 220748 512040 220776
rect 511868 220736 511874 220748
rect 512012 220708 512040 220748
rect 538490 220708 538496 220720
rect 512012 220680 518894 220708
rect 101214 220600 101220 220652
rect 101272 220640 101278 220652
rect 175458 220640 175464 220652
rect 101272 220612 175464 220640
rect 101272 220600 101278 220612
rect 175458 220600 175464 220612
rect 175516 220600 175522 220652
rect 177390 220600 177396 220652
rect 177448 220640 177454 220652
rect 180794 220640 180800 220652
rect 177448 220612 180800 220640
rect 177448 220600 177454 220612
rect 180794 220600 180800 220612
rect 180852 220600 180858 220652
rect 181070 220600 181076 220652
rect 181128 220640 181134 220652
rect 224218 220640 224224 220652
rect 181128 220612 224224 220640
rect 181128 220600 181134 220612
rect 224218 220600 224224 220612
rect 224276 220600 224282 220652
rect 253566 220600 253572 220652
rect 253624 220640 253630 220652
rect 293310 220640 293316 220652
rect 253624 220612 293316 220640
rect 253624 220600 253630 220612
rect 293310 220600 293316 220612
rect 293368 220600 293374 220652
rect 302418 220600 302424 220652
rect 302476 220640 302482 220652
rect 334066 220640 334072 220652
rect 302476 220612 334072 220640
rect 302476 220600 302482 220612
rect 334066 220600 334072 220612
rect 334124 220600 334130 220652
rect 357894 220600 357900 220652
rect 357952 220640 357958 220652
rect 374454 220640 374460 220652
rect 357952 220612 374460 220640
rect 357952 220600 357958 220612
rect 374454 220600 374460 220612
rect 374512 220600 374518 220652
rect 500218 220600 500224 220652
rect 500276 220640 500282 220652
rect 511810 220640 511816 220652
rect 500276 220612 511816 220640
rect 500276 220600 500282 220612
rect 511810 220600 511816 220612
rect 511868 220600 511874 220652
rect 69750 220464 69756 220516
rect 69808 220504 69814 220516
rect 136910 220504 136916 220516
rect 69808 220476 136916 220504
rect 69808 220464 69814 220476
rect 136910 220464 136916 220476
rect 136968 220464 136974 220516
rect 137094 220464 137100 220516
rect 137152 220504 137158 220516
rect 146938 220504 146944 220516
rect 137152 220476 146944 220504
rect 137152 220464 137158 220476
rect 146938 220464 146944 220476
rect 146996 220464 147002 220516
rect 147582 220464 147588 220516
rect 147640 220504 147646 220516
rect 150710 220504 150716 220516
rect 147640 220476 150716 220504
rect 147640 220464 147646 220476
rect 150710 220464 150716 220476
rect 150768 220464 150774 220516
rect 150894 220464 150900 220516
rect 150952 220504 150958 220516
rect 150952 220476 151814 220504
rect 150952 220464 150958 220476
rect 73062 220328 73068 220380
rect 73120 220368 73126 220380
rect 142108 220368 142114 220380
rect 73120 220340 142114 220368
rect 73120 220328 73126 220340
rect 142108 220328 142114 220340
rect 142166 220328 142172 220380
rect 142246 220328 142252 220380
rect 142304 220368 142310 220380
rect 144638 220368 144644 220380
rect 142304 220340 144644 220368
rect 142304 220328 142310 220340
rect 144638 220328 144644 220340
rect 144696 220328 144702 220380
rect 146754 220328 146760 220380
rect 146812 220368 146818 220380
rect 151630 220368 151636 220380
rect 146812 220340 151636 220368
rect 146812 220328 146818 220340
rect 151630 220328 151636 220340
rect 151688 220328 151694 220380
rect 151786 220368 151814 220476
rect 151906 220464 151912 220516
rect 151964 220504 151970 220516
rect 211338 220504 211344 220516
rect 151964 220476 211344 220504
rect 151964 220464 151970 220476
rect 211338 220464 211344 220476
rect 211396 220464 211402 220516
rect 214098 220504 214104 220516
rect 211908 220476 214104 220504
rect 211908 220368 211936 220476
rect 214098 220464 214104 220476
rect 214156 220464 214162 220516
rect 214282 220464 214288 220516
rect 214340 220504 214346 220516
rect 218698 220504 218704 220516
rect 214340 220476 218704 220504
rect 214340 220464 214346 220476
rect 218698 220464 218704 220476
rect 218756 220464 218762 220516
rect 223666 220464 223672 220516
rect 223724 220504 223730 220516
rect 265158 220504 265164 220516
rect 223724 220476 265164 220504
rect 223724 220464 223730 220476
rect 265158 220464 265164 220476
rect 265216 220464 265222 220516
rect 267642 220464 267648 220516
rect 267700 220504 267706 220516
rect 306834 220504 306840 220516
rect 267700 220476 306840 220504
rect 267700 220464 267706 220476
rect 306834 220464 306840 220476
rect 306892 220464 306898 220516
rect 338022 220464 338028 220516
rect 338080 220504 338086 220516
rect 358998 220504 359004 220516
rect 338080 220476 359004 220504
rect 338080 220464 338086 220476
rect 358998 220464 359004 220476
rect 359056 220464 359062 220516
rect 469122 220464 469128 220516
rect 469180 220504 469186 220516
rect 474550 220504 474556 220516
rect 469180 220476 474556 220504
rect 469180 220464 469186 220476
rect 474550 220464 474556 220476
rect 474608 220464 474614 220516
rect 488442 220464 488448 220516
rect 488500 220504 488506 220516
rect 501874 220504 501880 220516
rect 488500 220476 501880 220504
rect 488500 220464 488506 220476
rect 501874 220464 501880 220476
rect 501932 220464 501938 220516
rect 518866 220504 518894 220680
rect 538186 220680 538496 220708
rect 520918 220600 520924 220652
rect 520976 220640 520982 220652
rect 537478 220640 537484 220652
rect 520976 220612 537484 220640
rect 520976 220600 520982 220612
rect 537478 220600 537484 220612
rect 537536 220600 537542 220652
rect 531682 220504 531688 220516
rect 518866 220476 531688 220504
rect 531682 220464 531688 220476
rect 531740 220464 531746 220516
rect 535730 220464 535736 220516
rect 535788 220504 535794 220516
rect 538186 220504 538214 220680
rect 538490 220668 538496 220680
rect 538548 220668 538554 220720
rect 538858 220668 538864 220720
rect 538916 220708 538922 220720
rect 544286 220708 544292 220720
rect 538916 220680 544292 220708
rect 538916 220668 538922 220680
rect 544286 220668 544292 220680
rect 544344 220668 544350 220720
rect 550634 220600 550640 220652
rect 550692 220640 550698 220652
rect 554222 220640 554228 220652
rect 550692 220612 554228 220640
rect 550692 220600 550698 220612
rect 554222 220600 554228 220612
rect 554280 220600 554286 220652
rect 555694 220600 555700 220652
rect 555752 220640 555758 220652
rect 608870 220640 608876 220652
rect 555752 220612 608876 220640
rect 555752 220600 555758 220612
rect 608870 220600 608876 220612
rect 608928 220600 608934 220652
rect 556522 220504 556528 220516
rect 535788 220476 538214 220504
rect 543706 220476 556528 220504
rect 535788 220464 535794 220476
rect 151786 220340 211936 220368
rect 213638 220328 213644 220380
rect 213696 220368 213702 220380
rect 213696 220340 224264 220368
rect 213696 220328 213702 220340
rect 79686 220192 79692 220244
rect 79744 220232 79750 220244
rect 151722 220232 151728 220244
rect 79744 220204 151728 220232
rect 79744 220192 79750 220204
rect 151722 220192 151728 220204
rect 151780 220192 151786 220244
rect 151906 220192 151912 220244
rect 151964 220232 151970 220244
rect 154022 220232 154028 220244
rect 151964 220204 154028 220232
rect 151964 220192 151970 220204
rect 154022 220192 154028 220204
rect 154080 220192 154086 220244
rect 156322 220192 156328 220244
rect 156380 220232 156386 220244
rect 158898 220232 158904 220244
rect 156380 220204 158904 220232
rect 156380 220192 156386 220204
rect 158898 220192 158904 220204
rect 158956 220192 158962 220244
rect 164142 220192 164148 220244
rect 164200 220232 164206 220244
rect 223850 220232 223856 220244
rect 164200 220204 223856 220232
rect 164200 220192 164206 220204
rect 223850 220192 223856 220204
rect 223908 220192 223914 220244
rect 224236 220232 224264 220340
rect 224402 220328 224408 220380
rect 224460 220368 224466 220380
rect 267918 220368 267924 220380
rect 224460 220340 267924 220368
rect 224460 220328 224466 220340
rect 267918 220328 267924 220340
rect 267976 220328 267982 220380
rect 273438 220328 273444 220380
rect 273496 220368 273502 220380
rect 309226 220368 309232 220380
rect 273496 220340 309232 220368
rect 273496 220328 273502 220340
rect 309226 220328 309232 220340
rect 309284 220328 309290 220380
rect 314838 220328 314844 220380
rect 314896 220368 314902 220380
rect 341058 220368 341064 220380
rect 314896 220340 341064 220368
rect 314896 220328 314902 220340
rect 341058 220328 341064 220340
rect 341116 220328 341122 220380
rect 342990 220328 342996 220380
rect 343048 220368 343054 220380
rect 363414 220368 363420 220380
rect 343048 220340 363420 220368
rect 343048 220328 343054 220340
rect 363414 220328 363420 220340
rect 363472 220328 363478 220380
rect 472986 220328 472992 220380
rect 473044 220368 473050 220380
rect 481174 220368 481180 220380
rect 473044 220340 481180 220368
rect 473044 220328 473050 220340
rect 481174 220328 481180 220340
rect 481232 220328 481238 220380
rect 496446 220328 496452 220380
rect 496504 220368 496510 220380
rect 509326 220368 509332 220380
rect 496504 220340 509332 220368
rect 496504 220328 496510 220340
rect 509326 220328 509332 220340
rect 509384 220328 509390 220380
rect 516962 220328 516968 220380
rect 517020 220368 517026 220380
rect 527542 220368 527548 220380
rect 517020 220340 527548 220368
rect 517020 220328 517026 220340
rect 527542 220328 527548 220340
rect 527600 220328 527606 220380
rect 531130 220328 531136 220380
rect 531188 220368 531194 220380
rect 543706 220368 543734 220476
rect 556522 220464 556528 220476
rect 556580 220464 556586 220516
rect 558270 220464 558276 220516
rect 558328 220504 558334 220516
rect 561766 220504 561772 220516
rect 558328 220476 561772 220504
rect 558328 220464 558334 220476
rect 561766 220464 561772 220476
rect 561824 220464 561830 220516
rect 561950 220464 561956 220516
rect 562008 220504 562014 220516
rect 562008 220476 563054 220504
rect 562008 220464 562014 220476
rect 554038 220368 554044 220380
rect 531188 220340 543734 220368
rect 548536 220340 554044 220368
rect 531188 220328 531194 220340
rect 234154 220232 234160 220244
rect 224236 220204 234160 220232
rect 234154 220192 234160 220204
rect 234212 220192 234218 220244
rect 237006 220192 237012 220244
rect 237064 220232 237070 220244
rect 280430 220232 280436 220244
rect 237064 220204 280436 220232
rect 237064 220192 237070 220204
rect 280430 220192 280436 220204
rect 280488 220192 280494 220244
rect 283374 220192 283380 220244
rect 283432 220232 283438 220244
rect 316310 220232 316316 220244
rect 283432 220204 316316 220232
rect 283432 220192 283438 220204
rect 316310 220192 316316 220204
rect 316368 220192 316374 220244
rect 316494 220192 316500 220244
rect 316552 220232 316558 220244
rect 342622 220232 342628 220244
rect 316552 220204 342628 220232
rect 316552 220192 316558 220204
rect 342622 220192 342628 220204
rect 342680 220192 342686 220244
rect 348786 220192 348792 220244
rect 348844 220232 348850 220244
rect 369946 220232 369952 220244
rect 348844 220204 369952 220232
rect 348844 220192 348850 220204
rect 369946 220192 369952 220204
rect 370004 220192 370010 220244
rect 370498 220192 370504 220244
rect 370556 220232 370562 220244
rect 381078 220232 381084 220244
rect 370556 220204 381084 220232
rect 370556 220192 370562 220204
rect 381078 220192 381084 220204
rect 381136 220192 381142 220244
rect 388714 220192 388720 220244
rect 388772 220232 388778 220244
rect 400950 220232 400956 220244
rect 388772 220204 400956 220232
rect 388772 220192 388778 220204
rect 400950 220192 400956 220204
rect 401008 220192 401014 220244
rect 430114 220192 430120 220244
rect 430172 220232 430178 220244
rect 432046 220232 432052 220244
rect 430172 220204 432052 220232
rect 430172 220192 430178 220204
rect 432046 220192 432052 220204
rect 432104 220192 432110 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 473170 220192 473176 220244
rect 473228 220232 473234 220244
rect 482002 220232 482008 220244
rect 473228 220204 482008 220232
rect 473228 220192 473234 220204
rect 482002 220192 482008 220204
rect 482060 220192 482066 220244
rect 482922 220192 482928 220244
rect 482980 220232 482986 220244
rect 495250 220232 495256 220244
rect 482980 220204 495256 220232
rect 482980 220192 482986 220204
rect 495250 220192 495256 220204
rect 495308 220192 495314 220244
rect 501322 220192 501328 220244
rect 501380 220232 501386 220244
rect 520182 220232 520188 220244
rect 501380 220204 520188 220232
rect 501380 220192 501386 220204
rect 520182 220192 520188 220204
rect 520240 220192 520246 220244
rect 528370 220192 528376 220244
rect 528428 220232 528434 220244
rect 548536 220232 548564 220340
rect 554038 220328 554044 220340
rect 554096 220328 554102 220380
rect 554222 220328 554228 220380
rect 554280 220368 554286 220380
rect 562318 220368 562324 220380
rect 554280 220340 562324 220368
rect 554280 220328 554286 220340
rect 562318 220328 562324 220340
rect 562376 220328 562382 220380
rect 563026 220368 563054 220476
rect 563146 220464 563152 220516
rect 563204 220504 563210 220516
rect 609422 220504 609428 220516
rect 563204 220476 609428 220504
rect 563204 220464 563210 220476
rect 609422 220464 609428 220476
rect 609480 220464 609486 220516
rect 566458 220368 566464 220380
rect 563026 220340 566464 220368
rect 566458 220328 566464 220340
rect 566516 220328 566522 220380
rect 566826 220328 566832 220380
rect 566884 220368 566890 220380
rect 567286 220368 567292 220380
rect 566884 220340 567292 220368
rect 566884 220328 566890 220340
rect 567286 220328 567292 220340
rect 567344 220328 567350 220380
rect 568574 220328 568580 220380
rect 568632 220368 568638 220380
rect 569770 220368 569776 220380
rect 568632 220340 569776 220368
rect 568632 220328 568638 220340
rect 569770 220328 569776 220340
rect 569828 220328 569834 220380
rect 572668 220328 572674 220380
rect 572726 220368 572732 220380
rect 610526 220368 610532 220380
rect 572726 220340 610532 220368
rect 572726 220328 572732 220340
rect 610526 220328 610532 220340
rect 610584 220328 610590 220380
rect 569954 220260 569960 220312
rect 570012 220300 570018 220312
rect 570012 220272 572484 220300
rect 570012 220260 570018 220272
rect 528428 220204 548564 220232
rect 528428 220192 528434 220204
rect 548702 220192 548708 220244
rect 548760 220232 548766 220244
rect 548760 220204 562364 220232
rect 548760 220192 548766 220204
rect 154390 220124 154396 220176
rect 154448 220164 154454 220176
rect 156138 220164 156144 220176
rect 154448 220136 156144 220164
rect 154448 220124 154454 220136
rect 156138 220124 156144 220136
rect 156196 220124 156202 220176
rect 562336 220164 562364 220204
rect 572070 220164 572076 220176
rect 562336 220136 572076 220164
rect 572070 220124 572076 220136
rect 572128 220124 572134 220176
rect 572456 220164 572484 220272
rect 611446 220232 611452 220244
rect 572686 220204 611452 220232
rect 572686 220164 572714 220204
rect 611446 220192 611452 220204
rect 611504 220192 611510 220244
rect 648614 220192 648620 220244
rect 648672 220232 648678 220244
rect 652754 220232 652760 220244
rect 648672 220204 652760 220232
rect 648672 220192 648678 220204
rect 652754 220192 652760 220204
rect 652812 220192 652818 220244
rect 572456 220136 572714 220164
rect 76374 220056 76380 220108
rect 76432 220096 76438 220108
rect 152182 220096 152188 220108
rect 76432 220068 152188 220096
rect 76432 220056 76438 220068
rect 152182 220056 152188 220068
rect 152240 220056 152246 220108
rect 152366 220056 152372 220108
rect 152424 220096 152430 220108
rect 153838 220096 153844 220108
rect 152424 220068 153844 220096
rect 152424 220056 152430 220068
rect 153838 220056 153844 220068
rect 153896 220056 153902 220108
rect 157518 220056 157524 220108
rect 157576 220096 157582 220108
rect 214282 220096 214288 220108
rect 157576 220068 214288 220096
rect 157576 220056 157582 220068
rect 214282 220056 214288 220068
rect 214340 220056 214346 220108
rect 244274 220096 244280 220108
rect 214576 220068 244280 220096
rect 107838 219920 107844 219972
rect 107896 219960 107902 219972
rect 114278 219960 114284 219972
rect 107896 219932 114284 219960
rect 107896 219920 107902 219932
rect 114278 219920 114284 219932
rect 114336 219920 114342 219972
rect 114462 219920 114468 219972
rect 114520 219960 114526 219972
rect 114520 219932 126744 219960
rect 114520 219920 114526 219932
rect 121086 219784 121092 219836
rect 121144 219824 121150 219836
rect 126716 219824 126744 219932
rect 127618 219920 127624 219972
rect 127676 219960 127682 219972
rect 190270 219960 190276 219972
rect 127676 219932 190276 219960
rect 127676 219920 127682 219932
rect 190270 219920 190276 219932
rect 190328 219920 190334 219972
rect 190408 219920 190414 219972
rect 190466 219960 190472 219972
rect 213638 219960 213644 219972
rect 190466 219932 213644 219960
rect 190466 219920 190472 219932
rect 213638 219920 213644 219932
rect 213696 219920 213702 219972
rect 137094 219824 137100 219836
rect 121144 219796 122834 219824
rect 126716 219796 137100 219824
rect 121144 219784 121150 219796
rect 122806 219688 122834 219796
rect 137094 219784 137100 219796
rect 137152 219784 137158 219836
rect 197630 219824 197636 219836
rect 137296 219796 197636 219824
rect 127618 219688 127624 219700
rect 122806 219660 127624 219688
rect 127618 219648 127624 219660
rect 127676 219648 127682 219700
rect 131022 219648 131028 219700
rect 131080 219688 131086 219700
rect 137296 219688 137324 219796
rect 197630 219784 197636 219796
rect 197688 219784 197694 219836
rect 197814 219784 197820 219836
rect 197872 219824 197878 219836
rect 214576 219824 214604 220068
rect 244274 220056 244280 220068
rect 244332 220056 244338 220108
rect 244458 220056 244464 220108
rect 244516 220096 244522 220108
rect 288526 220096 288532 220108
rect 244516 220068 288532 220096
rect 244516 220056 244522 220068
rect 288526 220056 288532 220068
rect 288584 220056 288590 220108
rect 288710 220056 288716 220108
rect 288768 220096 288774 220108
rect 322382 220096 322388 220108
rect 288768 220068 322388 220096
rect 288768 220056 288774 220068
rect 322382 220056 322388 220068
rect 322440 220056 322446 220108
rect 325602 220056 325608 220108
rect 325660 220096 325666 220108
rect 352098 220096 352104 220108
rect 325660 220068 352104 220096
rect 325660 220056 325666 220068
rect 352098 220056 352104 220068
rect 352156 220056 352162 220108
rect 358814 220056 358820 220108
rect 358872 220096 358878 220108
rect 378318 220096 378324 220108
rect 358872 220068 378324 220096
rect 358872 220056 358878 220068
rect 378318 220056 378324 220068
rect 378376 220056 378382 220108
rect 379422 220056 379428 220108
rect 379480 220096 379486 220108
rect 392118 220096 392124 220108
rect 379480 220068 392124 220096
rect 379480 220056 379486 220068
rect 392118 220056 392124 220068
rect 392176 220056 392182 220108
rect 395982 220056 395988 220108
rect 396040 220096 396046 220108
rect 404722 220096 404728 220108
rect 396040 220068 404728 220096
rect 396040 220056 396046 220068
rect 404722 220056 404728 220068
rect 404780 220056 404786 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426802 220096 426808 220108
rect 421708 220068 426808 220096
rect 421708 220056 421714 220068
rect 426802 220056 426808 220068
rect 426860 220056 426866 220108
rect 431954 220056 431960 220108
rect 432012 220096 432018 220108
rect 434806 220096 434812 220108
rect 432012 220068 434812 220096
rect 432012 220056 432018 220068
rect 434806 220056 434812 220068
rect 434864 220056 434870 220108
rect 478322 220056 478328 220108
rect 478380 220096 478386 220108
rect 489454 220096 489460 220108
rect 478380 220068 489460 220096
rect 478380 220056 478386 220068
rect 489454 220056 489460 220068
rect 489512 220056 489518 220108
rect 492490 220056 492496 220108
rect 492548 220096 492554 220108
rect 506842 220096 506848 220108
rect 492548 220068 506848 220096
rect 492548 220056 492554 220068
rect 506842 220056 506848 220068
rect 506900 220056 506906 220108
rect 513098 220056 513104 220108
rect 513156 220096 513162 220108
rect 534166 220096 534172 220108
rect 513156 220068 534172 220096
rect 513156 220056 513162 220068
rect 534166 220056 534172 220068
rect 534224 220056 534230 220108
rect 538122 220056 538128 220108
rect 538180 220096 538186 220108
rect 561950 220096 561956 220108
rect 538180 220068 561956 220096
rect 538180 220056 538186 220068
rect 561950 220056 561956 220068
rect 562008 220056 562014 220108
rect 562318 219988 562324 220040
rect 562376 220028 562382 220040
rect 607306 220028 607312 220040
rect 562376 220000 607312 220028
rect 562376 219988 562382 220000
rect 607306 219988 607312 220000
rect 607364 219988 607370 220040
rect 214742 219920 214748 219972
rect 214800 219960 214806 219972
rect 254762 219960 254768 219972
rect 214800 219932 254768 219960
rect 214800 219920 214806 219932
rect 254762 219920 254768 219932
rect 254820 219920 254826 219972
rect 294966 219920 294972 219972
rect 295024 219960 295030 219972
rect 325878 219960 325884 219972
rect 295024 219932 325884 219960
rect 295024 219920 295030 219932
rect 325878 219920 325884 219932
rect 325936 219920 325942 219972
rect 548702 219892 548708 219904
rect 528526 219864 548708 219892
rect 259914 219824 259920 219836
rect 197872 219796 214604 219824
rect 214760 219796 259920 219824
rect 197872 219784 197878 219796
rect 142108 219688 142114 219700
rect 131080 219660 137324 219688
rect 137388 219660 142114 219688
rect 131080 219648 131086 219660
rect 123478 219552 123484 219564
rect 120092 219524 123484 219552
rect 70578 219376 70584 219428
rect 70636 219416 70642 219428
rect 70636 219388 103514 219416
rect 70636 219376 70642 219388
rect 93762 219240 93768 219292
rect 93820 219280 93826 219292
rect 94406 219280 94412 219292
rect 93820 219252 94412 219280
rect 93820 219240 93826 219252
rect 94406 219240 94412 219252
rect 94464 219240 94470 219292
rect 103486 219280 103514 219388
rect 109494 219376 109500 219428
rect 109552 219416 109558 219428
rect 110414 219416 110420 219428
rect 109552 219388 110420 219416
rect 109552 219376 109558 219388
rect 110414 219376 110420 219388
rect 110472 219376 110478 219428
rect 117774 219376 117780 219428
rect 117832 219416 117838 219428
rect 118694 219416 118700 219428
rect 117832 219388 118700 219416
rect 117832 219376 117838 219388
rect 118694 219376 118700 219388
rect 118752 219376 118758 219428
rect 120092 219280 120120 219524
rect 123478 219512 123484 219524
rect 123536 219512 123542 219564
rect 131684 219524 133920 219552
rect 120258 219376 120264 219428
rect 120316 219416 120322 219428
rect 120316 219388 122834 219416
rect 120316 219376 120322 219388
rect 103486 219252 120120 219280
rect 122806 219280 122834 219388
rect 123570 219376 123576 219428
rect 123628 219416 123634 219428
rect 129826 219416 129832 219428
rect 123628 219388 129832 219416
rect 123628 219376 123634 219388
rect 129826 219376 129832 219388
rect 129884 219376 129890 219428
rect 130194 219376 130200 219428
rect 130252 219416 130258 219428
rect 131684 219416 131712 219524
rect 130252 219388 131712 219416
rect 130252 219376 130258 219388
rect 131850 219376 131856 219428
rect 131908 219416 131914 219428
rect 132402 219416 132408 219428
rect 131908 219388 132408 219416
rect 131908 219376 131914 219388
rect 132402 219376 132408 219388
rect 132460 219376 132466 219428
rect 133892 219416 133920 219524
rect 136910 219512 136916 219564
rect 136968 219552 136974 219564
rect 137388 219552 137416 219660
rect 142108 219648 142114 219660
rect 142166 219648 142172 219700
rect 203150 219688 203156 219700
rect 142264 219660 203156 219688
rect 136968 219524 137416 219552
rect 136968 219512 136974 219524
rect 137646 219512 137652 219564
rect 137704 219552 137710 219564
rect 142264 219552 142292 219660
rect 203150 219648 203156 219660
rect 203208 219648 203214 219700
rect 208578 219688 208584 219700
rect 203720 219660 208584 219688
rect 137704 219524 142292 219552
rect 137704 219512 137710 219524
rect 144270 219512 144276 219564
rect 144328 219552 144334 219564
rect 203720 219552 203748 219660
rect 208578 219648 208584 219660
rect 208636 219648 208642 219700
rect 210510 219648 210516 219700
rect 210568 219688 210574 219700
rect 214760 219688 214788 219796
rect 259914 219784 259920 219796
rect 259972 219784 259978 219836
rect 527542 219716 527548 219768
rect 527600 219756 527606 219768
rect 528526 219756 528554 219864
rect 548702 219852 548708 219864
rect 548760 219852 548766 219904
rect 548886 219852 548892 219904
rect 548944 219892 548950 219904
rect 598566 219892 598572 219904
rect 548944 219864 598572 219892
rect 548944 219852 548950 219864
rect 598566 219852 598572 219864
rect 598624 219852 598630 219904
rect 606018 219892 606024 219904
rect 598768 219864 606024 219892
rect 527600 219728 528554 219756
rect 527600 219716 527606 219728
rect 540790 219716 540796 219768
rect 540848 219756 540854 219768
rect 598768 219756 598796 219864
rect 606018 219852 606024 219864
rect 606076 219852 606082 219904
rect 620094 219756 620100 219768
rect 540848 219728 598796 219756
rect 600976 219728 620100 219756
rect 540848 219716 540854 219728
rect 210568 219660 214788 219688
rect 210568 219648 210574 219660
rect 217134 219648 217140 219700
rect 217192 219688 217198 219700
rect 223666 219688 223672 219700
rect 217192 219660 223672 219688
rect 217192 219648 217198 219660
rect 223666 219648 223672 219660
rect 223724 219648 223730 219700
rect 224402 219688 224408 219700
rect 223868 219660 224408 219688
rect 144328 219524 203748 219552
rect 144328 219512 144334 219524
rect 203886 219512 203892 219564
rect 203944 219552 203950 219564
rect 214742 219552 214748 219564
rect 203944 219524 214748 219552
rect 203944 219512 203950 219524
rect 214742 219512 214748 219524
rect 214800 219512 214806 219564
rect 220446 219512 220452 219564
rect 220504 219552 220510 219564
rect 223868 219552 223896 219660
rect 224402 219648 224408 219660
rect 224460 219648 224466 219700
rect 227070 219648 227076 219700
rect 227128 219688 227134 219700
rect 272702 219688 272708 219700
rect 227128 219660 272708 219688
rect 227128 219648 227134 219660
rect 272702 219648 272708 219660
rect 272760 219648 272766 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 503622 219580 503628 219632
rect 503680 219620 503686 219632
rect 591850 219620 591856 219632
rect 503680 219592 591856 219620
rect 503680 219580 503686 219592
rect 591850 219580 591856 219592
rect 591908 219580 591914 219632
rect 591988 219580 591994 219632
rect 592046 219620 592052 219632
rect 600976 219620 601004 219728
rect 620094 219716 620100 219728
rect 620152 219716 620158 219768
rect 592046 219592 601004 219620
rect 592046 219580 592052 219592
rect 220504 219524 223896 219552
rect 220504 219512 220510 219524
rect 224218 219512 224224 219564
rect 224276 219552 224282 219564
rect 229278 219552 229284 219564
rect 224276 219524 229284 219552
rect 224276 219512 224282 219524
rect 229278 219512 229284 219524
rect 229336 219512 229342 219564
rect 332686 219512 332692 219564
rect 332744 219552 332750 219564
rect 337194 219552 337200 219564
rect 332744 219524 337200 219552
rect 332744 219512 332750 219524
rect 337194 219512 337200 219524
rect 337252 219512 337258 219564
rect 135824 219456 136772 219484
rect 135824 219416 135852 219456
rect 133892 219388 135852 219416
rect 136744 219416 136772 219456
rect 142448 219456 143442 219484
rect 142448 219416 142476 219456
rect 136744 219388 142476 219416
rect 143414 219416 143442 219456
rect 240152 219456 241514 219484
rect 146754 219416 146760 219428
rect 143414 219388 146760 219416
rect 146754 219376 146760 219388
rect 146812 219376 146818 219428
rect 146938 219376 146944 219428
rect 146996 219416 147002 219428
rect 152366 219416 152372 219428
rect 146996 219388 152372 219416
rect 146996 219376 147002 219388
rect 152366 219376 152372 219388
rect 152424 219376 152430 219428
rect 152550 219376 152556 219428
rect 152608 219416 152614 219428
rect 156230 219416 156236 219428
rect 152608 219388 156236 219416
rect 152608 219376 152614 219388
rect 156230 219376 156236 219388
rect 156288 219376 156294 219428
rect 156414 219376 156420 219428
rect 156472 219416 156478 219428
rect 158990 219416 158996 219428
rect 156472 219388 158996 219416
rect 156472 219376 156478 219388
rect 158990 219376 158996 219388
rect 159048 219376 159054 219428
rect 159174 219376 159180 219428
rect 159232 219416 159238 219428
rect 160002 219416 160008 219428
rect 159232 219388 160008 219416
rect 159232 219376 159238 219388
rect 160002 219376 160008 219388
rect 160060 219376 160066 219428
rect 162394 219416 162400 219428
rect 162044 219388 162400 219416
rect 162044 219280 162072 219388
rect 162394 219376 162400 219388
rect 162452 219376 162458 219428
rect 163314 219376 163320 219428
rect 163372 219416 163378 219428
rect 163958 219416 163964 219428
rect 163372 219388 163964 219416
rect 163372 219376 163378 219388
rect 163958 219376 163964 219388
rect 164016 219376 164022 219428
rect 178034 219416 178040 219428
rect 166966 219388 178040 219416
rect 166966 219280 166994 219388
rect 178034 219376 178040 219388
rect 178092 219376 178098 219428
rect 178218 219376 178224 219428
rect 178276 219416 178282 219428
rect 178276 219388 180380 219416
rect 178276 219376 178282 219388
rect 122806 219252 162072 219280
rect 162228 219252 166994 219280
rect 64598 219104 64604 219156
rect 64656 219144 64662 219156
rect 66898 219144 66904 219156
rect 64656 219116 66904 219144
rect 64656 219104 64662 219116
rect 66898 219104 66904 219116
rect 66956 219104 66962 219156
rect 83826 219104 83832 219156
rect 83884 219144 83890 219156
rect 157978 219144 157984 219156
rect 83884 219116 157984 219144
rect 83884 219104 83890 219116
rect 157978 219104 157984 219116
rect 158036 219104 158042 219156
rect 62298 218968 62304 219020
rect 62356 219008 62362 219020
rect 72418 219008 72424 219020
rect 62356 218980 72424 219008
rect 62356 218968 62362 218980
rect 72418 218968 72424 218980
rect 72476 218968 72482 219020
rect 77202 218968 77208 219020
rect 77260 219008 77266 219020
rect 146938 219008 146944 219020
rect 77260 218980 146944 219008
rect 77260 218968 77266 218980
rect 146938 218968 146944 218980
rect 146996 218968 147002 219020
rect 147122 218968 147128 219020
rect 147180 219008 147186 219020
rect 156414 219008 156420 219020
rect 147180 218980 156420 219008
rect 147180 218968 147186 218980
rect 156414 218968 156420 218980
rect 156472 218968 156478 219020
rect 162228 219008 162256 219252
rect 169110 219240 169116 219292
rect 169168 219280 169174 219292
rect 169570 219280 169576 219292
rect 169168 219252 169576 219280
rect 169168 219240 169174 219252
rect 169570 219240 169576 219252
rect 169628 219240 169634 219292
rect 169938 219240 169944 219292
rect 169996 219280 170002 219292
rect 170950 219280 170956 219292
rect 169996 219252 170956 219280
rect 169996 219240 170002 219252
rect 170950 219240 170956 219252
rect 171008 219240 171014 219292
rect 171410 219240 171416 219292
rect 171468 219280 171474 219292
rect 172238 219280 172244 219292
rect 171468 219252 172244 219280
rect 171468 219240 171474 219252
rect 172238 219240 172244 219252
rect 172296 219240 172302 219292
rect 172422 219240 172428 219292
rect 172480 219280 172486 219292
rect 173158 219280 173164 219292
rect 172480 219252 173164 219280
rect 172480 219240 172486 219252
rect 173158 219240 173164 219252
rect 173216 219240 173222 219292
rect 175734 219240 175740 219292
rect 175792 219280 175798 219292
rect 180352 219280 180380 219388
rect 180702 219376 180708 219428
rect 180760 219416 180766 219428
rect 185854 219416 185860 219428
rect 180760 219388 185860 219416
rect 180760 219376 180766 219388
rect 185854 219376 185860 219388
rect 185912 219376 185918 219428
rect 186498 219376 186504 219428
rect 186556 219416 186562 219428
rect 224402 219416 224408 219428
rect 186556 219388 224408 219416
rect 186556 219376 186562 219388
rect 224402 219376 224408 219388
rect 224460 219376 224466 219428
rect 229554 219376 229560 219428
rect 229612 219416 229618 219428
rect 230474 219416 230480 219428
rect 229612 219388 230480 219416
rect 229612 219376 229618 219388
rect 230474 219376 230480 219388
rect 230532 219376 230538 219428
rect 237834 219376 237840 219428
rect 237892 219416 237898 219428
rect 239306 219416 239312 219428
rect 237892 219388 239312 219416
rect 237892 219376 237898 219388
rect 239306 219376 239312 219388
rect 239364 219376 239370 219428
rect 239490 219376 239496 219428
rect 239548 219416 239554 219428
rect 240152 219416 240180 219456
rect 239548 219388 240180 219416
rect 241486 219416 241514 219456
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 241790 219416 241796 219428
rect 241486 219388 241796 219416
rect 239548 219376 239554 219388
rect 241790 219376 241796 219388
rect 241848 219376 241854 219428
rect 241974 219376 241980 219428
rect 242032 219416 242038 219428
rect 242894 219416 242900 219428
rect 242032 219388 242900 219416
rect 242032 219376 242038 219388
rect 242894 219376 242900 219388
rect 242952 219376 242958 219428
rect 244918 219376 244924 219428
rect 244976 219416 244982 219428
rect 272334 219416 272340 219428
rect 244976 219388 272340 219416
rect 244976 219376 244982 219388
rect 272334 219376 272340 219388
rect 272392 219376 272398 219428
rect 272702 219376 272708 219428
rect 272760 219416 272766 219428
rect 272760 219388 277394 219416
rect 272760 219376 272766 219388
rect 215938 219280 215944 219292
rect 175792 219252 180288 219280
rect 180352 219252 215944 219280
rect 175792 219240 175798 219252
rect 162394 219104 162400 219156
rect 162452 219144 162458 219156
rect 165614 219144 165620 219156
rect 162452 219116 165620 219144
rect 162452 219104 162458 219116
rect 165614 219104 165620 219116
rect 165672 219104 165678 219156
rect 165798 219104 165804 219156
rect 165856 219144 165862 219156
rect 180058 219144 180064 219156
rect 165856 219116 180064 219144
rect 165856 219104 165862 219116
rect 180058 219104 180064 219116
rect 180116 219104 180122 219156
rect 180260 219144 180288 219252
rect 215938 219240 215944 219252
rect 215996 219240 216002 219292
rect 219618 219240 219624 219292
rect 219676 219280 219682 219292
rect 264146 219280 264152 219292
rect 219676 219252 264152 219280
rect 219676 219240 219682 219252
rect 264146 219240 264152 219252
rect 264204 219240 264210 219292
rect 277366 219280 277394 219388
rect 285858 219376 285864 219428
rect 285916 219416 285922 219428
rect 285916 219388 306374 219416
rect 285916 219376 285922 219388
rect 301958 219280 301964 219292
rect 277366 219252 301964 219280
rect 301958 219240 301964 219252
rect 302016 219240 302022 219292
rect 306346 219280 306374 219388
rect 308214 219376 308220 219428
rect 308272 219416 308278 219428
rect 309134 219416 309140 219428
rect 308272 219388 309140 219416
rect 308272 219376 308278 219388
rect 309134 219376 309140 219388
rect 309192 219376 309198 219428
rect 333698 219376 333704 219428
rect 333756 219416 333762 219428
rect 347222 219416 347228 219428
rect 333756 219388 347228 219416
rect 333756 219376 333762 219388
rect 347222 219376 347228 219388
rect 347280 219376 347286 219428
rect 349614 219376 349620 219428
rect 349672 219416 349678 219428
rect 350534 219416 350540 219428
rect 349672 219388 350540 219416
rect 349672 219376 349678 219388
rect 350534 219376 350540 219388
rect 350592 219376 350598 219428
rect 352098 219376 352104 219428
rect 352156 219416 352162 219428
rect 355318 219416 355324 219428
rect 352156 219388 355324 219416
rect 352156 219376 352162 219388
rect 355318 219376 355324 219388
rect 355376 219376 355382 219428
rect 362034 219376 362040 219428
rect 362092 219416 362098 219428
rect 367646 219416 367652 219428
rect 362092 219388 367652 219416
rect 362092 219376 362098 219388
rect 367646 219376 367652 219388
rect 367704 219376 367710 219428
rect 380250 219376 380256 219428
rect 380308 219416 380314 219428
rect 384206 219416 384212 219428
rect 380308 219388 384212 219416
rect 380308 219376 380314 219388
rect 384206 219376 384212 219388
rect 384264 219376 384270 219428
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 501138 219444 501144 219496
rect 501196 219484 501202 219496
rect 596174 219484 596180 219496
rect 501196 219456 596180 219484
rect 501196 219444 501202 219456
rect 596174 219444 596180 219456
rect 596232 219444 596238 219496
rect 597738 219484 597744 219496
rect 596376 219456 597744 219484
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 572530 219348 572536 219360
rect 563026 219320 572536 219348
rect 313918 219280 313924 219292
rect 306346 219252 313924 219280
rect 313918 219240 313924 219252
rect 313976 219240 313982 219292
rect 320634 219240 320640 219292
rect 320692 219280 320698 219292
rect 342806 219280 342812 219292
rect 320692 219252 342812 219280
rect 320692 219240 320698 219252
rect 342806 219240 342812 219252
rect 342864 219240 342870 219292
rect 419166 219240 419172 219292
rect 419224 219280 419230 219292
rect 422662 219280 422668 219292
rect 419224 219252 422668 219280
rect 419224 219240 419230 219252
rect 422662 219240 422668 219252
rect 422720 219240 422726 219292
rect 548242 219240 548248 219292
rect 548300 219280 548306 219292
rect 548300 219252 553394 219280
rect 548300 219240 548306 219252
rect 189902 219144 189908 219156
rect 180260 219116 189908 219144
rect 189902 219104 189908 219116
rect 189960 219104 189966 219156
rect 190638 219104 190644 219156
rect 190696 219144 190702 219156
rect 197814 219144 197820 219156
rect 190696 219116 197820 219144
rect 190696 219104 190702 219116
rect 197814 219104 197820 219116
rect 197872 219104 197878 219156
rect 208854 219104 208860 219156
rect 208912 219144 208918 219156
rect 209682 219144 209688 219156
rect 208912 219116 209688 219144
rect 208912 219104 208918 219116
rect 209682 219104 209688 219116
rect 209740 219104 209746 219156
rect 218790 219104 218796 219156
rect 218848 219144 218854 219156
rect 219342 219144 219348 219156
rect 218848 219116 219348 219144
rect 218848 219104 218854 219116
rect 219342 219104 219348 219116
rect 219400 219104 219406 219156
rect 224218 219104 224224 219156
rect 224276 219144 224282 219156
rect 253198 219144 253204 219156
rect 224276 219116 253204 219144
rect 224276 219104 224282 219116
rect 253198 219104 253204 219116
rect 253256 219104 253262 219156
rect 265986 219104 265992 219156
rect 266044 219144 266050 219156
rect 266044 219116 291884 219144
rect 266044 219104 266050 219116
rect 156616 218980 162256 219008
rect 59814 218832 59820 218884
rect 59872 218872 59878 218884
rect 139946 218872 139952 218884
rect 59872 218844 139952 218872
rect 59872 218832 59878 218844
rect 139946 218832 139952 218844
rect 140004 218832 140010 218884
rect 140130 218832 140136 218884
rect 140188 218872 140194 218884
rect 156616 218872 156644 218980
rect 162670 218968 162676 219020
rect 162728 219008 162734 219020
rect 203518 219008 203524 219020
rect 162728 218980 203524 219008
rect 162728 218968 162734 218980
rect 203518 218968 203524 218980
rect 203576 218968 203582 219020
rect 206462 218968 206468 219020
rect 206520 219008 206526 219020
rect 253842 219008 253848 219020
rect 206520 218980 253848 219008
rect 206520 218968 206526 218980
rect 253842 218968 253848 218980
rect 253900 218968 253906 219020
rect 259086 218968 259092 219020
rect 259144 219008 259150 219020
rect 291654 219008 291660 219020
rect 259144 218980 291660 219008
rect 259144 218968 259150 218980
rect 291654 218968 291660 218980
rect 291712 218968 291718 219020
rect 291856 219008 291884 219116
rect 295794 219104 295800 219156
rect 295852 219144 295858 219156
rect 296714 219144 296720 219156
rect 295852 219116 296720 219144
rect 295852 219104 295858 219116
rect 296714 219104 296720 219116
rect 296772 219104 296778 219156
rect 314010 219104 314016 219156
rect 314068 219144 314074 219156
rect 335998 219144 336004 219156
rect 314068 219116 336004 219144
rect 314068 219104 314074 219116
rect 335998 219104 336004 219116
rect 336056 219104 336062 219156
rect 343818 219104 343824 219156
rect 343876 219144 343882 219156
rect 353938 219144 353944 219156
rect 343876 219116 353944 219144
rect 343876 219104 343882 219116
rect 353938 219104 353944 219116
rect 353996 219104 354002 219156
rect 542538 219104 542544 219156
rect 542596 219144 542602 219156
rect 542998 219144 543004 219156
rect 542596 219116 543004 219144
rect 542596 219104 542602 219116
rect 542998 219104 543004 219116
rect 543056 219144 543062 219156
rect 548794 219144 548800 219156
rect 543056 219116 548800 219144
rect 543056 219104 543062 219116
rect 548794 219104 548800 219116
rect 548852 219104 548858 219156
rect 553366 219144 553394 219252
rect 557350 219240 557356 219292
rect 557408 219280 557414 219292
rect 560662 219280 560668 219292
rect 557408 219252 560668 219280
rect 557408 219240 557414 219252
rect 560662 219240 560668 219252
rect 560720 219240 560726 219292
rect 563026 219280 563054 219320
rect 572530 219308 572536 219320
rect 572588 219308 572594 219360
rect 572668 219308 572674 219360
rect 572726 219348 572732 219360
rect 591666 219348 591672 219360
rect 572726 219320 591672 219348
rect 572726 219308 572732 219320
rect 591666 219308 591672 219320
rect 591724 219308 591730 219360
rect 591850 219308 591856 219360
rect 591908 219348 591914 219360
rect 596376 219348 596404 219456
rect 597738 219444 597744 219456
rect 597796 219444 597802 219496
rect 598566 219444 598572 219496
rect 598624 219484 598630 219496
rect 607490 219484 607496 219496
rect 598624 219456 607496 219484
rect 598624 219444 598630 219456
rect 607490 219444 607496 219456
rect 607548 219444 607554 219496
rect 591908 219320 596404 219348
rect 591908 219308 591914 219320
rect 561140 219252 563054 219280
rect 561140 219144 561168 219252
rect 553366 219116 561168 219144
rect 561232 219116 576854 219144
rect 297266 219008 297272 219020
rect 291856 218980 297272 219008
rect 297266 218968 297272 218980
rect 297324 218968 297330 219020
rect 307386 218968 307392 219020
rect 307444 219008 307450 219020
rect 332686 219008 332692 219020
rect 307444 218980 332692 219008
rect 307444 218968 307450 218980
rect 332686 218968 332692 218980
rect 332744 218968 332750 219020
rect 337194 218968 337200 219020
rect 337252 219008 337258 219020
rect 345658 219008 345664 219020
rect 337252 218980 345664 219008
rect 337252 218968 337258 218980
rect 345658 218968 345664 218980
rect 345716 218968 345722 219020
rect 347222 218968 347228 219020
rect 347280 219008 347286 219020
rect 363598 219008 363604 219020
rect 347280 218980 363604 219008
rect 347280 218968 347286 218980
rect 363598 218968 363604 218980
rect 363656 218968 363662 219020
rect 368658 218968 368664 219020
rect 368716 219008 368722 219020
rect 377398 219008 377404 219020
rect 368716 218980 377404 219008
rect 368716 218968 368722 218980
rect 377398 218968 377404 218980
rect 377456 218968 377462 219020
rect 377600 218980 383654 219008
rect 140188 218844 156644 218872
rect 140188 218832 140194 218844
rect 156782 218832 156788 218884
rect 156840 218872 156846 218884
rect 158714 218872 158720 218884
rect 156840 218844 158720 218872
rect 156840 218832 156846 218844
rect 158714 218832 158720 218844
rect 158772 218832 158778 218884
rect 158990 218832 158996 218884
rect 159048 218872 159054 218884
rect 171410 218872 171416 218884
rect 159048 218844 171416 218872
rect 159048 218832 159054 218844
rect 171410 218832 171416 218844
rect 171468 218832 171474 218884
rect 171778 218832 171784 218884
rect 171836 218872 171842 218884
rect 179506 218872 179512 218884
rect 171836 218844 179512 218872
rect 171836 218832 171842 218844
rect 179506 218832 179512 218844
rect 179564 218832 179570 218884
rect 182358 218832 182364 218884
rect 182416 218872 182422 218884
rect 189718 218872 189724 218884
rect 182416 218844 189724 218872
rect 182416 218832 182422 218844
rect 189718 218832 189724 218844
rect 189776 218832 189782 218884
rect 192846 218832 192852 218884
rect 192904 218872 192910 218884
rect 192904 218844 195468 218872
rect 192904 218832 192910 218844
rect 58986 218696 58992 218748
rect 59044 218736 59050 218748
rect 145006 218736 145012 218748
rect 59044 218708 145012 218736
rect 59044 218696 59050 218708
rect 145006 218696 145012 218708
rect 145064 218696 145070 218748
rect 146754 218696 146760 218748
rect 146812 218736 146818 218748
rect 183738 218736 183744 218748
rect 146812 218708 183744 218736
rect 146812 218696 146818 218708
rect 183738 218696 183744 218708
rect 183796 218696 183802 218748
rect 192110 218696 192116 218748
rect 192168 218736 192174 218748
rect 195238 218736 195244 218748
rect 192168 218708 195244 218736
rect 192168 218696 192174 218708
rect 195238 218696 195244 218708
rect 195296 218696 195302 218748
rect 195440 218736 195468 218844
rect 198918 218832 198924 218884
rect 198976 218872 198982 218884
rect 200022 218872 200028 218884
rect 198976 218844 200028 218872
rect 198976 218832 198982 218844
rect 200022 218832 200028 218844
rect 200080 218832 200086 218884
rect 200206 218832 200212 218884
rect 200264 218872 200270 218884
rect 241606 218872 241612 218884
rect 200264 218844 241612 218872
rect 200264 218832 200270 218844
rect 241606 218832 241612 218844
rect 241664 218832 241670 218884
rect 241790 218832 241796 218884
rect 241848 218872 241854 218884
rect 244918 218872 244924 218884
rect 241848 218844 244924 218872
rect 241848 218832 241854 218844
rect 244918 218832 244924 218844
rect 244976 218832 244982 218884
rect 249426 218832 249432 218884
rect 249484 218872 249490 218884
rect 251726 218872 251732 218884
rect 249484 218844 251732 218872
rect 249484 218832 249490 218844
rect 251726 218832 251732 218844
rect 251784 218832 251790 218884
rect 252738 218832 252744 218884
rect 252796 218872 252802 218884
rect 287882 218872 287888 218884
rect 252796 218844 287888 218872
rect 252796 218832 252802 218844
rect 287882 218832 287888 218844
rect 287940 218832 287946 218884
rect 291654 218832 291660 218884
rect 291712 218872 291718 218884
rect 291712 218844 296714 218872
rect 291712 218832 291718 218844
rect 243446 218736 243452 218748
rect 195440 218708 243452 218736
rect 243446 218696 243452 218708
rect 243504 218696 243510 218748
rect 251726 218696 251732 218748
rect 251784 218736 251790 218748
rect 286318 218736 286324 218748
rect 251784 218708 286324 218736
rect 251784 218696 251790 218708
rect 286318 218696 286324 218708
rect 286376 218696 286382 218748
rect 296686 218736 296714 218844
rect 300486 218832 300492 218884
rect 300544 218872 300550 218884
rect 327718 218872 327724 218884
rect 300544 218844 327724 218872
rect 300544 218832 300550 218844
rect 327718 218832 327724 218844
rect 327776 218832 327782 218884
rect 340506 218832 340512 218884
rect 340564 218872 340570 218884
rect 358078 218872 358084 218884
rect 340564 218844 358084 218872
rect 340564 218832 340570 218844
rect 358078 218832 358084 218844
rect 358136 218832 358142 218884
rect 363690 218832 363696 218884
rect 363748 218872 363754 218884
rect 370498 218872 370504 218884
rect 363748 218844 370504 218872
rect 363748 218832 363754 218844
rect 370498 218832 370504 218844
rect 370556 218832 370562 218884
rect 376938 218832 376944 218884
rect 376996 218872 377002 218884
rect 377600 218872 377628 218980
rect 376996 218844 377628 218872
rect 376996 218832 377002 218844
rect 382734 218832 382740 218884
rect 382792 218872 382798 218884
rect 383470 218872 383476 218884
rect 382792 218844 383476 218872
rect 382792 218832 382798 218844
rect 383470 218832 383476 218844
rect 383528 218832 383534 218884
rect 383626 218872 383654 218980
rect 386874 218968 386880 219020
rect 386932 219008 386938 219020
rect 398098 219008 398104 219020
rect 386932 218980 398104 219008
rect 386932 218968 386938 218980
rect 398098 218968 398104 218980
rect 398156 218968 398162 219020
rect 537478 218968 537484 219020
rect 537536 219008 537542 219020
rect 543182 219008 543188 219020
rect 537536 218980 543188 219008
rect 537536 218968 537542 218980
rect 543182 218968 543188 218980
rect 543240 218968 543246 219020
rect 561232 219008 561260 219116
rect 548444 218980 561260 219008
rect 388530 218872 388536 218884
rect 383626 218844 388536 218872
rect 388530 218832 388536 218844
rect 388588 218832 388594 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412542 218872 412548 218884
rect 411772 218844 412548 218872
rect 411772 218832 411778 218844
rect 412542 218832 412548 218844
rect 412600 218832 412606 218884
rect 512730 218832 512736 218884
rect 512788 218872 512794 218884
rect 548242 218872 548248 218884
rect 512788 218844 528554 218872
rect 512788 218832 512794 218844
rect 321554 218736 321560 218748
rect 296686 218708 321560 218736
rect 321554 218696 321560 218708
rect 321612 218696 321618 218748
rect 327258 218696 327264 218748
rect 327316 218736 327322 218748
rect 351086 218736 351092 218748
rect 327316 218708 351092 218736
rect 327316 218696 327322 218708
rect 351086 218696 351092 218708
rect 351144 218696 351150 218748
rect 353754 218696 353760 218748
rect 353812 218736 353818 218748
rect 369118 218736 369124 218748
rect 353812 218708 369124 218736
rect 353812 218696 353818 218708
rect 369118 218696 369124 218708
rect 369176 218696 369182 218748
rect 370314 218696 370320 218748
rect 370372 218736 370378 218748
rect 380066 218736 380072 218748
rect 370372 218708 380072 218736
rect 370372 218696 370378 218708
rect 380066 218696 380072 218708
rect 380124 218696 380130 218748
rect 383562 218696 383568 218748
rect 383620 218736 383626 218748
rect 396258 218736 396264 218748
rect 383620 218708 396264 218736
rect 383620 218696 383626 218708
rect 396258 218696 396264 218708
rect 396316 218696 396322 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 429930 218696 429936 218748
rect 429988 218736 429994 218748
rect 432690 218736 432696 218748
rect 429988 218708 432696 218736
rect 429988 218696 429994 218708
rect 432690 218696 432696 218708
rect 432748 218696 432754 218748
rect 482738 218696 482744 218748
rect 482796 218736 482802 218748
rect 485314 218736 485320 218748
rect 482796 218708 485320 218736
rect 482796 218696 482802 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 513834 218696 513840 218748
rect 513892 218736 513898 218748
rect 513892 218708 514248 218736
rect 513892 218696 513898 218708
rect 113634 218560 113640 218612
rect 113692 218600 113698 218612
rect 162210 218600 162216 218612
rect 113692 218572 162216 218600
rect 113692 218560 113698 218572
rect 162210 218560 162216 218572
rect 162268 218560 162274 218612
rect 162486 218560 162492 218612
rect 162544 218600 162550 218612
rect 171778 218600 171784 218612
rect 162544 218572 171784 218600
rect 162544 218560 162550 218572
rect 171778 218560 171784 218572
rect 171836 218560 171842 218612
rect 171962 218560 171968 218612
rect 172020 218600 172026 218612
rect 176010 218600 176016 218612
rect 172020 218572 176016 218600
rect 172020 218560 172026 218572
rect 176010 218560 176016 218572
rect 176068 218560 176074 218612
rect 179874 218560 179880 218612
rect 179932 218600 179938 218612
rect 210326 218600 210332 218612
rect 179932 218572 210332 218600
rect 179932 218560 179938 218572
rect 210326 218560 210332 218572
rect 210384 218560 210390 218612
rect 220078 218600 220084 218612
rect 214576 218572 220084 218600
rect 142430 218464 142436 218476
rect 103486 218436 142436 218464
rect 100386 218288 100392 218340
rect 100444 218328 100450 218340
rect 103486 218328 103514 218436
rect 142430 218424 142436 218436
rect 142488 218424 142494 218476
rect 142614 218424 142620 218476
rect 142672 218464 142678 218476
rect 143258 218464 143264 218476
rect 142672 218436 143264 218464
rect 142672 218424 142678 218436
rect 143258 218424 143264 218436
rect 143316 218424 143322 218476
rect 145098 218424 145104 218476
rect 145156 218464 145162 218476
rect 145926 218464 145932 218476
rect 145156 218436 145932 218464
rect 145156 218424 145162 218436
rect 145926 218424 145932 218436
rect 145984 218424 145990 218476
rect 148410 218424 148416 218476
rect 148468 218464 148474 218476
rect 148870 218464 148876 218476
rect 148468 218436 148876 218464
rect 148468 218424 148474 218436
rect 148870 218424 148876 218436
rect 148928 218424 148934 218476
rect 149238 218424 149244 218476
rect 149296 218464 149302 218476
rect 150066 218464 150072 218476
rect 149296 218436 150072 218464
rect 149296 218424 149302 218436
rect 150066 218424 150072 218436
rect 150124 218424 150130 218476
rect 153378 218424 153384 218476
rect 153436 218464 153442 218476
rect 186958 218464 186964 218476
rect 153436 218436 186964 218464
rect 153436 218424 153442 218436
rect 186958 218424 186964 218436
rect 187016 218424 187022 218476
rect 188706 218424 188712 218476
rect 188764 218464 188770 218476
rect 193766 218464 193772 218476
rect 188764 218436 193772 218464
rect 188764 218424 188770 218436
rect 193766 218424 193772 218436
rect 193824 218424 193830 218476
rect 195606 218424 195612 218476
rect 195664 218464 195670 218476
rect 197998 218464 198004 218476
rect 195664 218436 198004 218464
rect 195664 218424 195670 218436
rect 197998 218424 198004 218436
rect 198056 218424 198062 218476
rect 198274 218424 198280 218476
rect 198332 218464 198338 218476
rect 214576 218464 214604 218572
rect 220078 218560 220084 218572
rect 220136 218560 220142 218612
rect 225966 218560 225972 218612
rect 226024 218600 226030 218612
rect 266998 218600 267004 218612
rect 226024 218572 267004 218600
rect 226024 218560 226030 218572
rect 266998 218560 267004 218572
rect 267056 218560 267062 218612
rect 272334 218560 272340 218612
rect 272392 218600 272398 218612
rect 279418 218600 279424 218612
rect 272392 218572 279424 218600
rect 272392 218560 272398 218572
rect 279418 218560 279424 218572
rect 279476 218560 279482 218612
rect 305546 218600 305552 218612
rect 287026 218572 305552 218600
rect 224218 218464 224224 218476
rect 198332 218436 214604 218464
rect 214668 218436 224224 218464
rect 198332 218424 198338 218436
rect 100444 218300 103514 218328
rect 100444 218288 100450 218300
rect 116118 218288 116124 218340
rect 116176 218328 116182 218340
rect 117222 218328 117228 218340
rect 116176 218300 117228 218328
rect 116176 218288 116182 218300
rect 117222 218288 117228 218300
rect 117280 218288 117286 218340
rect 119430 218288 119436 218340
rect 119488 218328 119494 218340
rect 119982 218328 119988 218340
rect 119488 218300 119988 218328
rect 119488 218288 119494 218300
rect 119982 218288 119988 218300
rect 120040 218288 120046 218340
rect 121914 218288 121920 218340
rect 121972 218328 121978 218340
rect 122558 218328 122564 218340
rect 121972 218300 122564 218328
rect 121972 218288 121978 218300
rect 122558 218288 122564 218300
rect 122616 218288 122622 218340
rect 126054 218288 126060 218340
rect 126112 218328 126118 218340
rect 126698 218328 126704 218340
rect 126112 218300 126704 218328
rect 126112 218288 126118 218300
rect 126698 218288 126704 218300
rect 126756 218288 126762 218340
rect 127710 218288 127716 218340
rect 127768 218328 127774 218340
rect 128262 218328 128268 218340
rect 127768 218300 128268 218328
rect 127768 218288 127774 218300
rect 128262 218288 128268 218300
rect 128320 218288 128326 218340
rect 128538 218288 128544 218340
rect 128596 218328 128602 218340
rect 129366 218328 129372 218340
rect 128596 218300 129372 218328
rect 128596 218288 128602 218300
rect 129366 218288 129372 218300
rect 129424 218288 129430 218340
rect 129826 218288 129832 218340
rect 129884 218328 129890 218340
rect 132494 218328 132500 218340
rect 129884 218300 132500 218328
rect 129884 218288 129890 218300
rect 132494 218288 132500 218300
rect 132552 218288 132558 218340
rect 132678 218288 132684 218340
rect 132736 218328 132742 218340
rect 133506 218328 133512 218340
rect 132736 218300 133512 218328
rect 132736 218288 132742 218300
rect 133506 218288 133512 218300
rect 133564 218288 133570 218340
rect 135990 218288 135996 218340
rect 136048 218328 136054 218340
rect 136542 218328 136548 218340
rect 136048 218300 136548 218328
rect 136048 218288 136054 218300
rect 136542 218288 136548 218300
rect 136600 218288 136606 218340
rect 136910 218288 136916 218340
rect 136968 218328 136974 218340
rect 139946 218328 139952 218340
rect 136968 218300 139952 218328
rect 136968 218288 136974 218300
rect 139946 218288 139952 218300
rect 140004 218288 140010 218340
rect 140130 218288 140136 218340
rect 140188 218328 140194 218340
rect 170582 218328 170588 218340
rect 140188 218300 170588 218328
rect 140188 218288 140194 218300
rect 170582 218288 170588 218300
rect 170640 218288 170646 218340
rect 170766 218288 170772 218340
rect 170824 218328 170830 218340
rect 176562 218328 176568 218340
rect 170824 218300 176568 218328
rect 170824 218288 170830 218300
rect 176562 218288 176568 218300
rect 176620 218288 176626 218340
rect 179046 218288 179052 218340
rect 179104 218328 179110 218340
rect 196250 218328 196256 218340
rect 179104 218300 196256 218328
rect 179104 218288 179110 218300
rect 196250 218288 196256 218300
rect 196308 218288 196314 218340
rect 198090 218288 198096 218340
rect 198148 218328 198154 218340
rect 204162 218328 204168 218340
rect 198148 218300 204168 218328
rect 198148 218288 198154 218300
rect 204162 218288 204168 218300
rect 204220 218288 204226 218340
rect 204714 218288 204720 218340
rect 204772 218328 204778 218340
rect 207658 218328 207664 218340
rect 204772 218300 207664 218328
rect 204772 218288 204778 218300
rect 207658 218288 207664 218300
rect 207716 218288 207722 218340
rect 209682 218288 209688 218340
rect 209740 218328 209746 218340
rect 212810 218328 212816 218340
rect 209740 218300 212816 218328
rect 209740 218288 209746 218300
rect 212810 218288 212816 218300
rect 212868 218288 212874 218340
rect 212994 218288 213000 218340
rect 213052 218328 213058 218340
rect 214668 218328 214696 218436
rect 224218 218424 224224 218436
rect 224276 218424 224282 218476
rect 224402 218424 224408 218476
rect 224460 218464 224466 218476
rect 231026 218464 231032 218476
rect 224460 218436 231032 218464
rect 224460 218424 224466 218436
rect 231026 218424 231032 218436
rect 231084 218424 231090 218476
rect 238018 218464 238024 218476
rect 232700 218436 238024 218464
rect 213052 218300 214696 218328
rect 213052 218288 213058 218300
rect 216306 218288 216312 218340
rect 216364 218328 216370 218340
rect 232700 218328 232728 218436
rect 238018 218424 238024 218436
rect 238076 218424 238082 218476
rect 271138 218464 271144 218476
rect 238726 218436 271144 218464
rect 216364 218300 232728 218328
rect 216364 218288 216370 218300
rect 232866 218288 232872 218340
rect 232924 218328 232930 218340
rect 238726 218328 238754 218436
rect 271138 218424 271144 218436
rect 271196 218424 271202 218476
rect 279234 218424 279240 218476
rect 279292 218464 279298 218476
rect 287026 218464 287054 218572
rect 305546 218560 305552 218572
rect 305604 218560 305610 218612
rect 398466 218560 398472 218612
rect 398524 218600 398530 218612
rect 407758 218600 407764 218612
rect 398524 218572 407764 218600
rect 398524 218560 398530 218572
rect 407758 218560 407764 218572
rect 407816 218560 407822 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 475562 218560 475568 218612
rect 475620 218600 475626 218612
rect 482830 218600 482836 218612
rect 475620 218572 482836 218600
rect 475620 218560 475626 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 502702 218560 502708 218612
rect 502760 218600 502766 218612
rect 514018 218600 514024 218612
rect 502760 218572 514024 218600
rect 502760 218560 502766 218572
rect 514018 218560 514024 218572
rect 514076 218560 514082 218612
rect 514220 218600 514248 218708
rect 517698 218696 517704 218748
rect 517756 218736 517762 218748
rect 518158 218736 518164 218748
rect 517756 218708 518164 218736
rect 517756 218696 517762 218708
rect 518158 218696 518164 218708
rect 518216 218736 518222 218748
rect 519998 218736 520004 218748
rect 518216 218708 520004 218736
rect 518216 218696 518222 218708
rect 519998 218696 520004 218708
rect 520056 218696 520062 218748
rect 528526 218736 528554 218844
rect 542924 218844 548248 218872
rect 542924 218736 542952 218844
rect 548242 218832 548248 218844
rect 548300 218832 548306 218884
rect 548444 218736 548472 218980
rect 561674 218968 561680 219020
rect 561732 219008 561738 219020
rect 563008 219008 563014 219020
rect 561732 218980 563014 219008
rect 561732 218968 561738 218980
rect 563008 218968 563014 218980
rect 563066 218968 563072 219020
rect 563146 218968 563152 219020
rect 563204 219008 563210 219020
rect 567654 219008 567660 219020
rect 563204 218980 567660 219008
rect 563204 218968 563210 218980
rect 567654 218968 567660 218980
rect 567712 218968 567718 219020
rect 567838 218968 567844 219020
rect 567896 219008 567902 219020
rect 574554 219008 574560 219020
rect 567896 218980 574560 219008
rect 567896 218968 567902 218980
rect 574554 218968 574560 218980
rect 574612 218968 574618 219020
rect 576826 219008 576854 219116
rect 586974 219104 586980 219156
rect 587032 219144 587038 219156
rect 594794 219144 594800 219156
rect 587032 219116 594800 219144
rect 587032 219104 587038 219116
rect 594794 219104 594800 219116
rect 594852 219104 594858 219156
rect 587158 219008 587164 219020
rect 576826 218980 587164 219008
rect 587158 218968 587164 218980
rect 587216 218968 587222 219020
rect 548794 218832 548800 218884
rect 548852 218872 548858 218884
rect 560478 218872 560484 218884
rect 548852 218844 560484 218872
rect 548852 218832 548858 218844
rect 560478 218832 560484 218844
rect 560536 218832 560542 218884
rect 560662 218832 560668 218884
rect 560720 218872 560726 218884
rect 614114 218872 614120 218884
rect 560720 218844 614120 218872
rect 560720 218832 560726 218844
rect 614114 218832 614120 218844
rect 614172 218832 614178 218884
rect 528526 218708 542952 218736
rect 543016 218708 548472 218736
rect 543016 218600 543044 218708
rect 548610 218696 548616 218748
rect 548668 218736 548674 218748
rect 567838 218736 567844 218748
rect 548668 218708 567844 218736
rect 548668 218696 548674 218708
rect 567838 218696 567844 218708
rect 567896 218696 567902 218748
rect 568298 218696 568304 218748
rect 568356 218736 568362 218748
rect 571702 218736 571708 218748
rect 568356 218708 571708 218736
rect 568356 218696 568362 218708
rect 571702 218696 571708 218708
rect 571760 218696 571766 218748
rect 571886 218696 571892 218748
rect 571944 218736 571950 218748
rect 603074 218736 603080 218748
rect 571944 218708 603080 218736
rect 571944 218696 571950 218708
rect 603074 218696 603080 218708
rect 603132 218696 603138 218748
rect 514220 218572 543044 218600
rect 543182 218560 543188 218612
rect 543240 218600 543246 218612
rect 598842 218600 598848 218612
rect 543240 218572 598848 218600
rect 543240 218560 543246 218572
rect 598842 218560 598848 218572
rect 598900 218560 598906 218612
rect 604454 218600 604460 218612
rect 600792 218572 604460 218600
rect 279292 218436 287054 218464
rect 279292 218424 279298 218436
rect 294138 218424 294144 218476
rect 294196 218464 294202 218476
rect 316678 218464 316684 218476
rect 294196 218436 316684 218464
rect 294196 218424 294202 218436
rect 316678 218424 316684 218436
rect 316736 218424 316742 218476
rect 426618 218424 426624 218476
rect 426676 218464 426682 218476
rect 429562 218464 429568 218476
rect 426676 218436 429568 218464
rect 426676 218424 426682 218436
rect 429562 218424 429568 218436
rect 429620 218424 429626 218476
rect 500034 218424 500040 218476
rect 500092 218464 500098 218476
rect 600792 218464 600820 218572
rect 604454 218560 604460 218572
rect 604512 218560 604518 218612
rect 601234 218464 601240 218476
rect 500092 218436 600820 218464
rect 600884 218436 601240 218464
rect 500092 218424 500098 218436
rect 458174 218356 458180 218408
rect 458232 218396 458238 218408
rect 458232 218368 460934 218396
rect 458232 218356 458238 218368
rect 232924 218300 238754 218328
rect 232924 218288 232930 218300
rect 241606 218288 241612 218340
rect 241664 218328 241670 218340
rect 246298 218328 246304 218340
rect 241664 218300 246304 218328
rect 241664 218288 241670 218300
rect 246298 218288 246304 218300
rect 246356 218288 246362 218340
rect 253198 218288 253204 218340
rect 253256 218328 253262 218340
rect 258074 218328 258080 218340
rect 253256 218300 258080 218328
rect 253256 218288 253262 218300
rect 258074 218288 258080 218300
rect 258132 218288 258138 218340
rect 425790 218288 425796 218340
rect 425848 218328 425854 218340
rect 428458 218328 428464 218340
rect 425848 218300 428464 218328
rect 425848 218288 425854 218300
rect 428458 218288 428464 218300
rect 428516 218288 428522 218340
rect 450722 218288 450728 218340
rect 450780 218328 450786 218340
rect 453850 218328 453856 218340
rect 450780 218300 453856 218328
rect 450780 218288 450786 218300
rect 453850 218288 453856 218300
rect 453908 218288 453914 218340
rect 460906 218328 460934 218368
rect 461302 218328 461308 218340
rect 460906 218300 461308 218328
rect 461302 218288 461308 218300
rect 461360 218288 461366 218340
rect 496998 218288 497004 218340
rect 497056 218328 497062 218340
rect 586974 218328 586980 218340
rect 497056 218300 586980 218328
rect 497056 218288 497062 218300
rect 586974 218288 586980 218300
rect 587032 218288 587038 218340
rect 587158 218288 587164 218340
rect 587216 218328 587222 218340
rect 600884 218328 600912 218436
rect 601234 218424 601240 218436
rect 601292 218424 601298 218476
rect 670234 218424 670240 218476
rect 670292 218424 670298 218476
rect 587216 218300 600912 218328
rect 587216 218288 587222 218300
rect 601050 218288 601056 218340
rect 601108 218328 601114 218340
rect 607122 218328 607128 218340
rect 601108 218300 607128 218328
rect 601108 218288 601114 218300
rect 607122 218288 607128 218300
rect 607180 218288 607186 218340
rect 107010 218220 107016 218272
rect 107068 218260 107074 218272
rect 107068 218232 113174 218260
rect 107068 218220 107074 218232
rect 55674 218152 55680 218204
rect 55732 218192 55738 218204
rect 56502 218192 56508 218204
rect 55732 218164 56508 218192
rect 55732 218152 55738 218164
rect 56502 218152 56508 218164
rect 56560 218152 56566 218204
rect 57422 218152 57428 218204
rect 57480 218192 57486 218204
rect 61378 218192 61384 218204
rect 57480 218164 61384 218192
rect 57480 218152 57486 218164
rect 61378 218152 61384 218164
rect 61436 218152 61442 218204
rect 66438 218152 66444 218204
rect 66496 218192 66502 218204
rect 67542 218192 67548 218204
rect 66496 218164 67548 218192
rect 66496 218152 66502 218164
rect 67542 218152 67548 218164
rect 67600 218152 67606 218204
rect 68094 218152 68100 218204
rect 68152 218192 68158 218204
rect 69566 218192 69572 218204
rect 68152 218164 69572 218192
rect 68152 218152 68158 218164
rect 69566 218152 69572 218164
rect 69624 218152 69630 218204
rect 75546 218152 75552 218204
rect 75604 218192 75610 218204
rect 76558 218192 76564 218204
rect 75604 218164 76564 218192
rect 75604 218152 75610 218164
rect 76558 218152 76564 218164
rect 76616 218152 76622 218204
rect 97074 218152 97080 218204
rect 97132 218192 97138 218204
rect 113146 218192 113174 218232
rect 152366 218192 152372 218204
rect 97132 218164 100892 218192
rect 113146 218164 152372 218192
rect 97132 218152 97138 218164
rect 56502 218016 56508 218068
rect 56560 218056 56566 218068
rect 57238 218056 57244 218068
rect 56560 218028 57244 218056
rect 56560 218016 56566 218028
rect 57238 218016 57244 218028
rect 57296 218016 57302 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 59354 218056 59360 218068
rect 58216 218028 59360 218056
rect 58216 218016 58222 218028
rect 59354 218016 59360 218028
rect 59412 218016 59418 218068
rect 61470 218016 61476 218068
rect 61528 218056 61534 218068
rect 62758 218056 62764 218068
rect 61528 218028 62764 218056
rect 61528 218016 61534 218028
rect 62758 218016 62764 218028
rect 62816 218016 62822 218068
rect 63954 218016 63960 218068
rect 64012 218056 64018 218068
rect 64782 218056 64788 218068
rect 64012 218028 64788 218056
rect 64012 218016 64018 218028
rect 64782 218016 64788 218028
rect 64840 218016 64846 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 67266 218016 67272 218068
rect 67324 218056 67330 218068
rect 68278 218056 68284 218068
rect 67324 218028 68284 218056
rect 67324 218016 67330 218028
rect 68278 218016 68284 218028
rect 68336 218016 68342 218068
rect 72234 218016 72240 218068
rect 72292 218056 72298 218068
rect 73706 218056 73712 218068
rect 72292 218028 73712 218056
rect 72292 218016 72298 218028
rect 73706 218016 73712 218028
rect 73764 218016 73770 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 83458 218056 83464 218068
rect 82228 218028 83464 218056
rect 82228 218016 82234 218028
rect 83458 218016 83464 218028
rect 83516 218016 83522 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85298 218056 85304 218068
rect 84712 218028 85304 218056
rect 84712 218016 84718 218028
rect 85298 218016 85304 218028
rect 85356 218016 85362 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 92934 218016 92940 218068
rect 92992 218056 92998 218068
rect 93578 218056 93584 218068
rect 92992 218028 93584 218056
rect 92992 218016 92998 218028
rect 93578 218016 93584 218028
rect 93636 218016 93642 218068
rect 95418 218016 95424 218068
rect 95476 218056 95482 218068
rect 96246 218056 96252 218068
rect 95476 218028 96252 218056
rect 95476 218016 95482 218028
rect 96246 218016 96252 218028
rect 96304 218016 96310 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 100864 217988 100892 218164
rect 152366 218152 152372 218164
rect 152424 218152 152430 218204
rect 160002 218152 160008 218204
rect 160060 218192 160066 218204
rect 162670 218192 162676 218204
rect 160060 218164 162676 218192
rect 160060 218152 160066 218164
rect 162670 218152 162676 218164
rect 162728 218152 162734 218204
rect 166626 218152 166632 218204
rect 166684 218192 166690 218204
rect 166684 218164 200114 218192
rect 166684 218152 166690 218164
rect 102870 218084 102876 218136
rect 102928 218124 102934 218136
rect 103422 218124 103428 218136
rect 102928 218096 103428 218124
rect 102928 218084 102934 218096
rect 103422 218084 103428 218096
rect 103480 218084 103486 218136
rect 103698 218084 103704 218136
rect 103756 218124 103762 218136
rect 104802 218124 104808 218136
rect 103756 218096 104808 218124
rect 103756 218084 103762 218096
rect 104802 218084 104808 218096
rect 104860 218084 104866 218136
rect 105354 218084 105360 218136
rect 105412 218124 105418 218136
rect 105998 218124 106004 218136
rect 105412 218096 106004 218124
rect 105412 218084 105418 218096
rect 105998 218084 106004 218096
rect 106056 218084 106062 218136
rect 111978 218084 111984 218136
rect 112036 218124 112042 218136
rect 112806 218124 112812 218136
rect 112036 218096 112812 218124
rect 112036 218084 112042 218096
rect 112806 218084 112812 218096
rect 112864 218084 112870 218136
rect 152550 218084 152556 218136
rect 152608 218124 152614 218136
rect 153102 218124 153108 218136
rect 152608 218096 153108 218124
rect 152608 218084 152614 218096
rect 153102 218084 153108 218096
rect 153160 218084 153166 218136
rect 155034 218084 155040 218136
rect 155092 218124 155098 218136
rect 155678 218124 155684 218136
rect 155092 218096 155684 218124
rect 155092 218084 155098 218096
rect 155678 218084 155684 218096
rect 155736 218084 155742 218136
rect 156690 218084 156696 218136
rect 156748 218124 156754 218136
rect 157242 218124 157248 218136
rect 156748 218096 157248 218124
rect 156748 218084 156754 218096
rect 157242 218084 157248 218096
rect 157300 218084 157306 218136
rect 170582 218016 170588 218068
rect 170640 218056 170646 218068
rect 171962 218056 171968 218068
rect 170640 218028 171968 218056
rect 170640 218016 170646 218028
rect 171962 218016 171968 218028
rect 172020 218016 172026 218068
rect 173250 218016 173256 218068
rect 173308 218056 173314 218068
rect 178034 218056 178040 218068
rect 173308 218028 178040 218056
rect 173308 218016 173314 218028
rect 178034 218016 178040 218028
rect 178092 218016 178098 218068
rect 178218 218016 178224 218068
rect 178276 218056 178282 218068
rect 179322 218056 179328 218068
rect 178276 218028 179328 218056
rect 178276 218016 178282 218028
rect 179322 218016 179328 218028
rect 179380 218016 179386 218068
rect 179506 218016 179512 218068
rect 179564 218056 179570 218068
rect 181346 218056 181352 218068
rect 179564 218028 181352 218056
rect 179564 218016 179570 218028
rect 181346 218016 181352 218028
rect 181404 218016 181410 218068
rect 184014 218016 184020 218068
rect 184072 218056 184078 218068
rect 184658 218056 184664 218068
rect 184072 218028 184664 218056
rect 184072 218016 184078 218028
rect 184658 218016 184664 218028
rect 184716 218016 184722 218068
rect 185670 218016 185676 218068
rect 185728 218056 185734 218068
rect 186130 218056 186136 218068
rect 185728 218028 186136 218056
rect 185728 218016 185734 218028
rect 186130 218016 186136 218028
rect 186188 218016 186194 218068
rect 188154 218016 188160 218068
rect 188212 218056 188218 218068
rect 188890 218056 188896 218068
rect 188212 218028 188896 218056
rect 188212 218016 188218 218028
rect 188890 218016 188896 218028
rect 188948 218016 188954 218068
rect 189810 218016 189816 218068
rect 189868 218056 189874 218068
rect 192110 218056 192116 218068
rect 189868 218028 192116 218056
rect 189868 218016 189874 218028
rect 192110 218016 192116 218028
rect 192168 218016 192174 218068
rect 192294 218016 192300 218068
rect 192352 218056 192358 218068
rect 193030 218056 193036 218068
rect 192352 218028 193036 218056
rect 192352 218016 192358 218028
rect 193030 218016 193036 218028
rect 193088 218016 193094 218068
rect 193950 218016 193956 218068
rect 194008 218056 194014 218068
rect 194502 218056 194508 218068
rect 194008 218028 194508 218056
rect 194008 218016 194014 218028
rect 194502 218016 194508 218028
rect 194560 218016 194566 218068
rect 194778 218016 194784 218068
rect 194836 218056 194842 218068
rect 195882 218056 195888 218068
rect 194836 218028 195888 218056
rect 194836 218016 194842 218028
rect 195882 218016 195888 218028
rect 195940 218016 195946 218068
rect 196434 218016 196440 218068
rect 196492 218056 196498 218068
rect 198274 218056 198280 218068
rect 196492 218028 198280 218056
rect 196492 218016 196498 218028
rect 198274 218016 198280 218028
rect 198332 218016 198338 218068
rect 200086 218056 200114 218164
rect 200574 218152 200580 218204
rect 200632 218192 200638 218204
rect 201494 218192 201500 218204
rect 200632 218164 201500 218192
rect 200632 218152 200638 218164
rect 201494 218152 201500 218164
rect 201552 218152 201558 218204
rect 202230 218152 202236 218204
rect 202288 218192 202294 218204
rect 202690 218192 202696 218204
rect 202288 218164 202696 218192
rect 202288 218152 202294 218164
rect 202690 218152 202696 218164
rect 202748 218152 202754 218204
rect 203058 218152 203064 218204
rect 203116 218192 203122 218204
rect 206278 218192 206284 218204
rect 203116 218164 206284 218192
rect 203116 218152 203122 218164
rect 206278 218152 206284 218164
rect 206336 218152 206342 218204
rect 207198 218152 207204 218204
rect 207256 218192 207262 218204
rect 208118 218192 208124 218204
rect 207256 218164 208124 218192
rect 207256 218152 207262 218164
rect 208118 218152 208124 218164
rect 208176 218152 208182 218204
rect 211338 218152 211344 218204
rect 211396 218192 211402 218204
rect 211396 218164 216720 218192
rect 211396 218152 211402 218164
rect 211798 218056 211804 218068
rect 200086 218028 211804 218056
rect 211798 218016 211804 218028
rect 211856 218016 211862 218068
rect 214650 218016 214656 218068
rect 214708 218056 214714 218068
rect 215202 218056 215208 218068
rect 214708 218028 215208 218056
rect 214708 218016 214714 218028
rect 215202 218016 215208 218028
rect 215260 218016 215266 218068
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216490 218056 216496 218068
rect 215536 218028 216496 218056
rect 215536 218016 215542 218028
rect 216490 218016 216496 218028
rect 216548 218016 216554 218068
rect 216692 218056 216720 218164
rect 217962 218152 217968 218204
rect 218020 218192 218026 218204
rect 222746 218192 222752 218204
rect 218020 218164 222752 218192
rect 218020 218152 218026 218164
rect 222746 218152 222752 218164
rect 222804 218152 222810 218204
rect 222930 218152 222936 218204
rect 222988 218192 222994 218204
rect 225598 218192 225604 218204
rect 222988 218164 225604 218192
rect 222988 218152 222994 218164
rect 225598 218152 225604 218164
rect 225656 218152 225662 218204
rect 246114 218152 246120 218204
rect 246172 218192 246178 218204
rect 251726 218192 251732 218204
rect 246172 218164 251732 218192
rect 246172 218152 246178 218164
rect 251726 218152 251732 218164
rect 251784 218152 251790 218204
rect 328914 218152 328920 218204
rect 328972 218192 328978 218204
rect 330478 218192 330484 218204
rect 328972 218164 330484 218192
rect 328972 218152 328978 218164
rect 330478 218152 330484 218164
rect 330536 218152 330542 218204
rect 365346 218152 365352 218204
rect 365404 218192 365410 218204
rect 371786 218192 371792 218204
rect 365404 218164 371792 218192
rect 365404 218152 365410 218164
rect 371786 218152 371792 218164
rect 371844 218152 371850 218204
rect 374454 218152 374460 218204
rect 374512 218192 374518 218204
rect 376018 218192 376024 218204
rect 374512 218164 376024 218192
rect 374512 218152 374518 218164
rect 376018 218152 376024 218164
rect 376076 218152 376082 218204
rect 381906 218152 381912 218204
rect 381964 218192 381970 218204
rect 382918 218192 382924 218204
rect 381964 218164 382924 218192
rect 381964 218152 381970 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 401778 218152 401784 218204
rect 401836 218192 401842 218204
rect 402790 218192 402796 218204
rect 401836 218164 402796 218192
rect 401836 218152 401842 218164
rect 402790 218152 402796 218164
rect 402848 218152 402854 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 428274 218152 428280 218204
rect 428332 218192 428338 218204
rect 430114 218192 430120 218204
rect 428332 218164 430120 218192
rect 428332 218152 428338 218164
rect 430114 218152 430120 218164
rect 430172 218152 430178 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 434714 218192 434720 218204
rect 433300 218164 434720 218192
rect 433300 218152 433306 218164
rect 434714 218152 434720 218164
rect 434772 218152 434778 218204
rect 434898 218152 434904 218204
rect 434956 218192 434962 218204
rect 436830 218192 436836 218204
rect 434956 218164 436836 218192
rect 434956 218152 434962 218164
rect 436830 218152 436836 218164
rect 436888 218152 436894 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 491938 218152 491944 218204
rect 491996 218192 492002 218204
rect 500954 218192 500960 218204
rect 491996 218164 500960 218192
rect 491996 218152 492002 218164
rect 500954 218152 500960 218164
rect 501012 218152 501018 218204
rect 507118 218152 507124 218204
rect 507176 218192 507182 218204
rect 507670 218192 507676 218204
rect 507176 218164 507676 218192
rect 507176 218152 507182 218164
rect 507670 218152 507676 218164
rect 507728 218192 507734 218204
rect 513834 218192 513840 218204
rect 507728 218164 513840 218192
rect 507728 218152 507734 218164
rect 513834 218152 513840 218164
rect 513892 218152 513898 218204
rect 514018 218152 514024 218204
rect 514076 218192 514082 218204
rect 560294 218192 560300 218204
rect 514076 218164 560300 218192
rect 514076 218152 514082 218164
rect 560294 218152 560300 218164
rect 560352 218152 560358 218204
rect 560478 218152 560484 218204
rect 560536 218192 560542 218204
rect 563008 218192 563014 218204
rect 560536 218164 563014 218192
rect 560536 218152 560542 218164
rect 563008 218152 563014 218164
rect 563066 218152 563072 218204
rect 572668 218152 572674 218204
rect 572726 218192 572732 218204
rect 613562 218192 613568 218204
rect 572726 218164 613568 218192
rect 572726 218152 572732 218164
rect 613562 218152 613568 218164
rect 613620 218152 613626 218204
rect 563348 218096 572346 218124
rect 219802 218056 219808 218068
rect 216692 218028 219808 218056
rect 219802 218016 219808 218028
rect 219860 218016 219866 218068
rect 221274 218016 221280 218068
rect 221332 218056 221338 218068
rect 221826 218056 221832 218068
rect 221332 218028 221832 218056
rect 221332 218016 221338 218028
rect 221826 218016 221832 218028
rect 221884 218016 221890 218068
rect 223758 218016 223764 218068
rect 223816 218056 223822 218068
rect 224586 218056 224592 218068
rect 223816 218028 224592 218056
rect 223816 218016 223822 218028
rect 224586 218016 224592 218028
rect 224644 218016 224650 218068
rect 225414 218016 225420 218068
rect 225472 218056 225478 218068
rect 226150 218056 226156 218068
rect 225472 218028 226156 218056
rect 225472 218016 225478 218028
rect 226150 218016 226156 218028
rect 226208 218016 226214 218068
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233142 218056 233148 218068
rect 232096 218028 233148 218056
rect 232096 218016 232102 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235810 218056 235816 218068
rect 235408 218028 235816 218056
rect 235408 218016 235414 218028
rect 235810 218016 235816 218028
rect 235868 218016 235874 218068
rect 236178 218016 236184 218068
rect 236236 218056 236242 218068
rect 237282 218056 237288 218068
rect 236236 218028 237288 218056
rect 236236 218016 236242 218028
rect 237282 218016 237288 218028
rect 237340 218016 237346 218068
rect 240318 218016 240324 218068
rect 240376 218056 240382 218068
rect 241330 218056 241336 218068
rect 240376 218028 241336 218056
rect 240376 218016 240382 218028
rect 241330 218016 241336 218028
rect 241388 218016 241394 218068
rect 243630 218016 243636 218068
rect 243688 218056 243694 218068
rect 244090 218056 244096 218068
rect 243688 218028 244096 218056
rect 243688 218016 243694 218028
rect 244090 218016 244096 218028
rect 244148 218016 244154 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248230 218056 248236 218068
rect 247828 218028 248236 218056
rect 247828 218016 247834 218028
rect 248230 218016 248236 218028
rect 248288 218016 248294 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249610 218056 249616 218068
rect 248656 218028 249616 218056
rect 248656 218016 248662 218028
rect 249610 218016 249616 218028
rect 249668 218016 249674 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 250898 218056 250904 218068
rect 250312 218028 250904 218056
rect 250312 218016 250318 218028
rect 250898 218016 250904 218028
rect 250956 218016 250962 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 254394 218016 254400 218068
rect 254452 218056 254458 218068
rect 255038 218056 255044 218068
rect 254452 218028 255044 218056
rect 254452 218016 254458 218028
rect 255038 218016 255044 218028
rect 255096 218016 255102 218068
rect 256050 218016 256056 218068
rect 256108 218056 256114 218068
rect 256510 218056 256516 218068
rect 256108 218028 256516 218056
rect 256108 218016 256114 218028
rect 256510 218016 256516 218028
rect 256568 218016 256574 218068
rect 256878 218016 256884 218068
rect 256936 218056 256942 218068
rect 257522 218056 257528 218068
rect 256936 218028 257528 218056
rect 256936 218016 256942 218028
rect 257522 218016 257528 218028
rect 257580 218016 257586 218068
rect 258534 218016 258540 218068
rect 258592 218056 258598 218068
rect 259270 218056 259276 218068
rect 258592 218028 259276 218056
rect 258592 218016 258598 218028
rect 259270 218016 259276 218028
rect 259328 218016 259334 218068
rect 262674 218016 262680 218068
rect 262732 218056 262738 218068
rect 263594 218056 263600 218068
rect 262732 218028 263600 218056
rect 262732 218016 262738 218028
rect 263594 218016 263600 218028
rect 263652 218016 263658 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266170 218056 266176 218068
rect 265216 218028 266176 218056
rect 265216 218016 265222 218028
rect 266170 218016 266176 218028
rect 266228 218016 266234 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 268930 218056 268936 218068
rect 268528 218028 268936 218056
rect 268528 218016 268534 218028
rect 268930 218016 268936 218028
rect 268988 218016 268994 218068
rect 269298 218016 269304 218068
rect 269356 218056 269362 218068
rect 270034 218056 270040 218068
rect 269356 218028 270040 218056
rect 269356 218016 269362 218028
rect 270034 218016 270040 218028
rect 270092 218016 270098 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 272518 218056 272524 218068
rect 271012 218028 272524 218056
rect 271012 218016 271018 218028
rect 272518 218016 272524 218028
rect 272576 218016 272582 218068
rect 276750 218016 276756 218068
rect 276808 218056 276814 218068
rect 277210 218056 277216 218068
rect 276808 218028 277216 218056
rect 276808 218016 276814 218028
rect 277210 218016 277216 218028
rect 277268 218016 277274 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278590 218056 278596 218068
rect 277636 218028 278596 218056
rect 277636 218016 277642 218028
rect 278590 218016 278596 218028
rect 278648 218016 278654 218068
rect 280890 218016 280896 218068
rect 280948 218056 280954 218068
rect 281442 218056 281448 218068
rect 280948 218028 281448 218056
rect 280948 218016 280954 218028
rect 281442 218016 281448 218028
rect 281500 218016 281506 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282454 218056 282460 218068
rect 281776 218028 282460 218056
rect 281776 218016 281782 218028
rect 282454 218016 282460 218028
rect 282512 218016 282518 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288710 218056 288716 218068
rect 287572 218028 288716 218056
rect 287572 218016 287578 218028
rect 288710 218016 288716 218028
rect 288768 218016 288774 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289722 218056 289728 218068
rect 289228 218028 289728 218056
rect 289228 218016 289234 218028
rect 289722 218016 289728 218028
rect 289780 218016 289786 218068
rect 289998 218016 290004 218068
rect 290056 218056 290062 218068
rect 291102 218056 291108 218068
rect 290056 218028 291108 218056
rect 290056 218016 290062 218028
rect 291102 218016 291108 218028
rect 291160 218016 291166 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 297450 218016 297456 218068
rect 297508 218056 297514 218068
rect 297910 218056 297916 218068
rect 297508 218028 297916 218056
rect 297508 218016 297514 218028
rect 297910 218016 297916 218028
rect 297968 218016 297974 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299106 218056 299112 218068
rect 298336 218028 299112 218056
rect 298336 218016 298342 218028
rect 299106 218016 299112 218028
rect 299164 218016 299170 218068
rect 299934 218016 299940 218068
rect 299992 218056 299998 218068
rect 300670 218056 300676 218068
rect 299992 218028 300676 218056
rect 299992 218016 299998 218028
rect 300670 218016 300676 218028
rect 300728 218016 300734 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 304074 218016 304080 218068
rect 304132 218056 304138 218068
rect 304718 218056 304724 218068
rect 304132 218028 304724 218056
rect 304132 218016 304138 218028
rect 304718 218016 304724 218028
rect 304776 218016 304782 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306190 218056 306196 218068
rect 305788 218028 306196 218056
rect 305788 218016 305794 218028
rect 306190 218016 306196 218028
rect 306248 218016 306254 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 309870 218016 309876 218068
rect 309928 218056 309934 218068
rect 310422 218056 310428 218068
rect 309928 218028 310428 218056
rect 309928 218016 309934 218028
rect 310422 218016 310428 218028
rect 310480 218016 310486 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 312906 218056 312912 218068
rect 312412 218028 312912 218056
rect 312412 218016 312418 218028
rect 312906 218016 312912 218028
rect 312964 218016 312970 218068
rect 317322 218016 317328 218068
rect 317380 218056 317386 218068
rect 317966 218056 317972 218068
rect 317380 218028 317972 218056
rect 317380 218016 317386 218028
rect 317966 218016 317972 218028
rect 318024 218016 318030 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 319806 218056 319812 218068
rect 319036 218028 319812 218056
rect 319036 218016 319042 218028
rect 319806 218016 319812 218028
rect 319864 218016 319870 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 323118 218016 323124 218068
rect 323176 218056 323182 218068
rect 324130 218056 324136 218068
rect 323176 218028 324136 218056
rect 323176 218016 323182 218028
rect 324130 218016 324136 218028
rect 324188 218016 324194 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325418 218056 325424 218068
rect 324832 218028 325424 218056
rect 324832 218016 324838 218028
rect 325418 218016 325424 218028
rect 325476 218016 325482 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 330570 218016 330576 218068
rect 330628 218056 330634 218068
rect 331030 218056 331036 218068
rect 330628 218028 331036 218056
rect 330628 218016 330634 218028
rect 331030 218016 331036 218028
rect 331088 218016 331094 218068
rect 333054 218016 333060 218068
rect 333112 218056 333118 218068
rect 333882 218056 333888 218068
rect 333112 218028 333888 218056
rect 333112 218016 333118 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335170 218056 335176 218068
rect 334768 218028 335176 218056
rect 334768 218016 334774 218028
rect 335170 218016 335176 218028
rect 335228 218016 335234 218068
rect 335538 218016 335544 218068
rect 335596 218056 335602 218068
rect 338666 218056 338672 218068
rect 335596 218028 338672 218056
rect 335596 218016 335602 218028
rect 338666 218016 338672 218028
rect 338724 218016 338730 218068
rect 338850 218016 338856 218068
rect 338908 218056 338914 218068
rect 339402 218056 339408 218068
rect 338908 218028 339408 218056
rect 338908 218016 338914 218028
rect 339402 218016 339408 218028
rect 339460 218016 339466 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 345474 218016 345480 218068
rect 345532 218056 345538 218068
rect 347038 218056 347044 218068
rect 345532 218028 347044 218056
rect 345532 218016 345538 218028
rect 347038 218016 347044 218028
rect 347096 218016 347102 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 355410 218016 355416 218068
rect 355468 218056 355474 218068
rect 355870 218056 355876 218068
rect 355468 218028 355876 218056
rect 355468 218016 355474 218028
rect 355870 218016 355876 218028
rect 355928 218016 355934 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 356974 218056 356980 218068
rect 356296 218028 356980 218056
rect 356296 218016 356302 218028
rect 356974 218016 356980 218028
rect 357032 218016 357038 218068
rect 359550 218016 359556 218068
rect 359608 218056 359614 218068
rect 360102 218056 360108 218068
rect 359608 218028 360108 218056
rect 359608 218016 359614 218028
rect 360102 218016 360108 218028
rect 360160 218016 360166 218068
rect 360378 218016 360384 218068
rect 360436 218056 360442 218068
rect 361022 218056 361028 218068
rect 360436 218028 361028 218056
rect 360436 218016 360442 218028
rect 361022 218016 361028 218028
rect 361080 218016 361086 218068
rect 364518 218016 364524 218068
rect 364576 218056 364582 218068
rect 365530 218056 365536 218068
rect 364576 218028 365536 218056
rect 364576 218016 364582 218028
rect 365530 218016 365536 218028
rect 365588 218016 365594 218068
rect 366174 218016 366180 218068
rect 366232 218056 366238 218068
rect 366726 218056 366732 218068
rect 366232 218028 366732 218056
rect 366232 218016 366238 218028
rect 366726 218016 366732 218028
rect 366784 218016 366790 218068
rect 367830 218016 367836 218068
rect 367888 218056 367894 218068
rect 368382 218056 368388 218068
rect 367888 218028 368388 218056
rect 367888 218016 367894 218028
rect 368382 218016 368388 218028
rect 368440 218016 368446 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373442 218056 373448 218068
rect 372856 218028 373448 218056
rect 372856 218016 372862 218028
rect 373442 218016 373448 218028
rect 373500 218016 373506 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376662 218056 376668 218068
rect 376168 218028 376668 218056
rect 376168 218016 376174 218028
rect 376662 218016 376668 218028
rect 376720 218016 376726 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379238 218056 379244 218068
rect 378652 218028 379244 218056
rect 378652 218016 378658 218028
rect 379238 218016 379244 218028
rect 379296 218016 379302 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 382090 218056 382096 218068
rect 381136 218028 382096 218056
rect 381136 218016 381142 218028
rect 382090 218016 382096 218028
rect 382148 218016 382154 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390002 218056 390008 218068
rect 389416 218028 390008 218056
rect 389416 218016 389422 218028
rect 390002 218016 390008 218028
rect 390060 218016 390066 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393130 218056 393136 218068
rect 392728 218028 393136 218056
rect 392728 218016 392734 218028
rect 393130 218016 393136 218028
rect 393188 218016 393194 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394510 218056 394516 218068
rect 393556 218028 394516 218056
rect 393556 218016 393562 218028
rect 394510 218016 394516 218028
rect 394568 218016 394574 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395798 218056 395804 218068
rect 395212 218028 395804 218056
rect 395212 218016 395218 218028
rect 395798 218016 395804 218028
rect 395856 218016 395862 218068
rect 397638 218016 397644 218068
rect 397696 218056 397702 218068
rect 400582 218056 400588 218068
rect 397696 218028 400588 218056
rect 397696 218016 397702 218028
rect 400582 218016 400588 218028
rect 400640 218016 400646 218068
rect 400950 218016 400956 218068
rect 401008 218056 401014 218068
rect 402238 218056 402244 218068
rect 401008 218028 402244 218056
rect 401008 218016 401014 218028
rect 402238 218016 402244 218028
rect 402296 218016 402302 218068
rect 403434 218016 403440 218068
rect 403492 218056 403498 218068
rect 403986 218056 403992 218068
rect 403492 218028 403992 218056
rect 403492 218016 403498 218028
rect 403986 218016 403992 218028
rect 404044 218016 404050 218068
rect 405090 218016 405096 218068
rect 405148 218056 405154 218068
rect 405550 218056 405556 218068
rect 405148 218028 405556 218056
rect 405148 218016 405154 218028
rect 405550 218016 405556 218028
rect 405608 218016 405614 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 427906 218056 427912 218068
rect 427504 218028 427912 218056
rect 427504 218016 427510 218028
rect 427906 218016 427912 218028
rect 427964 218016 427970 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430574 218056 430580 218068
rect 429160 218028 430580 218056
rect 429160 218016 429166 218028
rect 430574 218016 430580 218028
rect 430632 218016 430638 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 435726 218016 435732 218068
rect 435784 218056 435790 218068
rect 436278 218056 436284 218068
rect 435784 218028 436284 218056
rect 435784 218016 435790 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436462 218016 436468 218068
rect 436520 218056 436526 218068
rect 437474 218056 437480 218068
rect 436520 218028 437480 218056
rect 436520 218016 436526 218028
rect 437474 218016 437480 218028
rect 437532 218016 437538 218068
rect 438210 218016 438216 218068
rect 438268 218056 438274 218068
rect 438854 218056 438860 218068
rect 438268 218028 438860 218056
rect 438268 218016 438274 218028
rect 438854 218016 438860 218028
rect 438912 218016 438918 218068
rect 439866 218016 439872 218068
rect 439924 218056 439930 218068
rect 440326 218056 440332 218068
rect 439924 218028 440332 218056
rect 439924 218016 439930 218028
rect 440326 218016 440332 218028
rect 440384 218016 440390 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 455598 218016 455604 218068
rect 455656 218056 455662 218068
rect 457162 218056 457168 218068
rect 455656 218028 457168 218056
rect 455656 218016 455662 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 471422 218016 471428 218068
rect 471480 218056 471486 218068
rect 472894 218056 472900 218068
rect 471480 218028 472900 218056
rect 471480 218016 471486 218028
rect 472894 218016 472900 218028
rect 472952 218016 472958 218068
rect 490374 218016 490380 218068
rect 490432 218056 490438 218068
rect 563348 218056 563376 218096
rect 490432 218028 563100 218056
rect 490432 218016 490438 218028
rect 563072 217988 563100 218028
rect 563210 218028 563376 218056
rect 572318 218056 572346 218096
rect 601050 218056 601056 218068
rect 572318 218028 601056 218056
rect 563210 217988 563238 218028
rect 601050 218016 601056 218028
rect 601108 218016 601114 218068
rect 601234 218016 601240 218068
rect 601292 218056 601298 218068
rect 601292 218028 610664 218056
rect 601292 218016 601298 218028
rect 100864 217960 157334 217988
rect 563072 217960 563238 217988
rect 157306 217920 157334 217960
rect 563514 217948 563520 218000
rect 563572 217988 563578 218000
rect 572162 217988 572168 218000
rect 563572 217960 572168 217988
rect 563572 217948 563578 217960
rect 572162 217948 572168 217960
rect 572220 217948 572226 218000
rect 610636 217988 610664 218028
rect 615678 217988 615684 218000
rect 610636 217960 615684 217988
rect 615678 217948 615684 217960
rect 615736 217948 615742 218000
rect 174262 217920 174268 217932
rect 157306 217892 174268 217920
rect 174262 217880 174268 217892
rect 174320 217880 174326 217932
rect 523034 217812 523040 217864
rect 523092 217852 523098 217864
rect 524230 217852 524236 217864
rect 523092 217824 524236 217852
rect 523092 217812 523098 217824
rect 524230 217812 524236 217824
rect 524288 217812 524294 217864
rect 535454 217812 535460 217864
rect 535512 217852 535518 217864
rect 536650 217852 536656 217864
rect 535512 217824 536656 217852
rect 535512 217812 535518 217824
rect 536650 217812 536656 217824
rect 536708 217812 536714 217864
rect 603994 217852 604000 217864
rect 536852 217824 604000 217852
rect 533430 217676 533436 217728
rect 533488 217716 533494 217728
rect 536852 217716 536880 217824
rect 603994 217812 604000 217824
rect 604052 217812 604058 217864
rect 670252 217784 670280 218424
rect 670418 218288 670424 218340
rect 670476 218328 670482 218340
rect 670476 218300 670648 218328
rect 670476 218288 670482 218300
rect 670620 218068 670648 218300
rect 670602 218016 670608 218068
rect 670660 218016 670666 218068
rect 675846 217948 675852 218000
rect 675904 217988 675910 218000
rect 676766 217988 676772 218000
rect 675904 217960 676772 217988
rect 675904 217948 675910 217960
rect 676766 217948 676772 217960
rect 676824 217948 676830 218000
rect 670418 217784 670424 217796
rect 670252 217756 670424 217784
rect 670418 217744 670424 217756
rect 670476 217744 670482 217796
rect 603442 217716 603448 217728
rect 533488 217688 536880 217716
rect 536944 217688 603448 217716
rect 533488 217676 533494 217688
rect 116946 217540 116952 217592
rect 117004 217580 117010 217592
rect 189166 217580 189172 217592
rect 117004 217552 189172 217580
rect 117004 217540 117010 217552
rect 189166 217540 189172 217552
rect 189224 217540 189230 217592
rect 530946 217540 530952 217592
rect 531004 217580 531010 217592
rect 536944 217580 536972 217688
rect 603442 217676 603448 217688
rect 603500 217676 603506 217728
rect 604454 217676 604460 217728
rect 604512 217716 604518 217728
rect 614298 217716 614304 217728
rect 604512 217688 614304 217716
rect 604512 217676 604518 217688
rect 614298 217676 614304 217688
rect 614356 217676 614362 217728
rect 531004 217552 536972 217580
rect 531004 217540 531010 217552
rect 538214 217540 538220 217592
rect 538272 217580 538278 217592
rect 539134 217580 539140 217592
rect 538272 217552 539140 217580
rect 538272 217540 538278 217552
rect 539134 217540 539140 217552
rect 539192 217540 539198 217592
rect 543366 217540 543372 217592
rect 543424 217580 543430 217592
rect 606202 217580 606208 217592
rect 543424 217552 606208 217580
rect 543424 217540 543430 217552
rect 606202 217540 606208 217552
rect 606260 217540 606266 217592
rect 614114 217540 614120 217592
rect 614172 217580 614178 217592
rect 626626 217580 626632 217592
rect 614172 217552 626632 217580
rect 614172 217540 614178 217552
rect 626626 217540 626632 217552
rect 626684 217540 626690 217592
rect 115290 217404 115296 217456
rect 115348 217444 115354 217456
rect 187970 217444 187976 217456
rect 115348 217416 187976 217444
rect 115348 217404 115354 217416
rect 187970 217404 187976 217416
rect 188028 217404 188034 217456
rect 527818 217404 527824 217456
rect 527876 217444 527882 217456
rect 528462 217444 528468 217456
rect 527876 217416 528468 217444
rect 527876 217404 527882 217416
rect 528462 217404 528468 217416
rect 528520 217444 528526 217456
rect 528520 217416 598704 217444
rect 528520 217404 528526 217416
rect 168558 217308 168564 217320
rect 93826 217280 168564 217308
rect 90404 217200 90410 217252
rect 90462 217240 90468 217252
rect 93826 217240 93854 217280
rect 168558 217268 168564 217280
rect 168616 217268 168622 217320
rect 508590 217268 508596 217320
rect 508648 217308 508654 217320
rect 563008 217308 563014 217320
rect 508648 217280 563014 217308
rect 508648 217268 508654 217280
rect 563008 217268 563014 217280
rect 563066 217268 563072 217320
rect 563146 217268 563152 217320
rect 563204 217308 563210 217320
rect 572530 217308 572536 217320
rect 563204 217280 572536 217308
rect 563204 217268 563210 217280
rect 572530 217268 572536 217280
rect 572588 217268 572594 217320
rect 572668 217268 572674 217320
rect 572726 217308 572732 217320
rect 598474 217308 598480 217320
rect 572726 217280 598480 217308
rect 572726 217268 572732 217280
rect 598474 217268 598480 217280
rect 598532 217268 598538 217320
rect 90462 217212 93854 217240
rect 90462 217200 90468 217212
rect 448606 217200 448612 217252
rect 448664 217240 448670 217252
rect 449756 217240 449762 217252
rect 448664 217212 449762 217240
rect 448664 217200 448670 217212
rect 449756 217200 449762 217212
rect 449814 217200 449820 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 498286 217200 498292 217252
rect 498344 217240 498350 217252
rect 499436 217240 499442 217252
rect 498344 217212 499442 217240
rect 498344 217200 498350 217212
rect 499436 217200 499442 217212
rect 499494 217200 499500 217252
rect 506060 217132 506066 217184
rect 506118 217172 506124 217184
rect 597922 217172 597928 217184
rect 506118 217144 597928 217172
rect 506118 217132 506124 217144
rect 597922 217132 597928 217144
rect 597980 217132 597986 217184
rect 598676 217172 598704 217416
rect 603074 217404 603080 217456
rect 603132 217444 603138 217456
rect 628282 217444 628288 217456
rect 603132 217416 628288 217444
rect 603132 217404 603138 217416
rect 628282 217404 628288 217416
rect 628340 217404 628346 217456
rect 670234 217336 670240 217388
rect 670292 217376 670298 217388
rect 670602 217376 670608 217388
rect 670292 217348 670608 217376
rect 670292 217336 670298 217348
rect 670602 217336 670608 217348
rect 670660 217336 670666 217388
rect 598842 217268 598848 217320
rect 598900 217308 598906 217320
rect 622394 217308 622400 217320
rect 598900 217280 622400 217308
rect 598900 217268 598906 217280
rect 622394 217268 622400 217280
rect 622452 217268 622458 217320
rect 603074 217172 603080 217184
rect 598676 217144 603080 217172
rect 603074 217132 603080 217144
rect 603132 217132 603138 217184
rect 498608 217064 498614 217116
rect 498666 217104 498672 217116
rect 498666 217076 505094 217104
rect 498666 217064 498672 217076
rect 505066 217036 505094 217076
rect 505066 217008 574048 217036
rect 574020 216900 574048 217008
rect 574186 216996 574192 217048
rect 574244 217036 574250 217048
rect 610066 217036 610072 217048
rect 574244 217008 610072 217036
rect 574244 216996 574250 217008
rect 610066 216996 610072 217008
rect 610124 216996 610130 217048
rect 596358 216900 596364 216912
rect 574020 216872 596364 216900
rect 596358 216860 596364 216872
rect 596416 216860 596422 216912
rect 607122 216860 607128 216912
rect 607180 216900 607186 216912
rect 612274 216900 612280 216912
rect 607180 216872 612280 216900
rect 607180 216860 607186 216872
rect 612274 216860 612280 216872
rect 612332 216860 612338 216912
rect 594794 216724 594800 216776
rect 594852 216764 594858 216776
rect 613378 216764 613384 216776
rect 594852 216736 613384 216764
rect 594852 216724 594858 216736
rect 613378 216724 613384 216736
rect 613436 216724 613442 216776
rect 613562 216656 613568 216708
rect 613620 216696 613626 216708
rect 614482 216696 614488 216708
rect 613620 216668 614488 216696
rect 613620 216656 613626 216668
rect 614482 216656 614488 216668
rect 614540 216656 614546 216708
rect 648246 216656 648252 216708
rect 648304 216696 648310 216708
rect 650638 216696 650644 216708
rect 648304 216668 650644 216696
rect 648304 216656 648310 216668
rect 650638 216656 650644 216668
rect 650696 216656 650702 216708
rect 644934 215908 644940 215960
rect 644992 215948 644998 215960
rect 658918 215948 658924 215960
rect 644992 215920 658924 215948
rect 644992 215908 644998 215920
rect 658918 215908 658924 215920
rect 658976 215908 658982 215960
rect 675846 215636 675852 215688
rect 675904 215676 675910 215688
rect 676950 215676 676956 215688
rect 675904 215648 676956 215676
rect 675904 215636 675910 215648
rect 676950 215636 676956 215648
rect 677008 215636 677014 215688
rect 675846 214956 675852 215008
rect 675904 214996 675910 215008
rect 676490 214996 676496 215008
rect 675904 214968 676496 214996
rect 675904 214956 675910 214968
rect 676490 214956 676496 214968
rect 676548 214956 676554 215008
rect 574738 214820 574744 214872
rect 574796 214860 574802 214872
rect 616874 214860 616880 214872
rect 574796 214832 616880 214860
rect 574796 214820 574802 214832
rect 616874 214820 616880 214832
rect 616932 214820 616938 214872
rect 574370 214684 574376 214736
rect 574428 214724 574434 214736
rect 623314 214724 623320 214736
rect 574428 214696 623320 214724
rect 574428 214684 574434 214696
rect 623314 214684 623320 214696
rect 623372 214684 623378 214736
rect 658182 214684 658188 214736
rect 658240 214724 658246 214736
rect 665818 214724 665824 214736
rect 658240 214696 665824 214724
rect 658240 214684 658246 214696
rect 665818 214684 665824 214696
rect 665876 214684 665882 214736
rect 574554 214548 574560 214600
rect 574612 214588 574618 214600
rect 574612 214560 605834 214588
rect 574612 214548 574618 214560
rect 601786 214412 601792 214464
rect 601844 214452 601850 214464
rect 602338 214452 602344 214464
rect 601844 214424 602344 214452
rect 601844 214412 601850 214424
rect 602338 214412 602344 214424
rect 602396 214412 602402 214464
rect 604638 214412 604644 214464
rect 604696 214452 604702 214464
rect 605098 214452 605104 214464
rect 604696 214424 605104 214452
rect 604696 214412 604702 214424
rect 605098 214412 605104 214424
rect 605156 214412 605162 214464
rect 605806 214452 605834 214560
rect 607306 214548 607312 214600
rect 607364 214588 607370 214600
rect 607858 214588 607864 214600
rect 607364 214560 607864 214588
rect 607364 214548 607370 214560
rect 607858 214548 607864 214560
rect 607916 214548 607922 214600
rect 618254 214548 618260 214600
rect 618312 214588 618318 214600
rect 618898 214588 618904 214600
rect 618312 214560 618904 214588
rect 618312 214548 618318 214560
rect 618898 214548 618904 214560
rect 618956 214548 618962 214600
rect 619910 214548 619916 214600
rect 619968 214588 619974 214600
rect 620554 214588 620560 214600
rect 619968 214560 620560 214588
rect 619968 214548 619974 214560
rect 620554 214548 620560 214560
rect 620612 214548 620618 214600
rect 623958 214548 623964 214600
rect 624016 214588 624022 214600
rect 624016 214560 625154 214588
rect 624016 214548 624022 214560
rect 624418 214452 624424 214464
rect 605806 214424 624424 214452
rect 624418 214412 624424 214424
rect 624476 214412 624482 214464
rect 625126 214452 625154 214560
rect 625430 214548 625436 214600
rect 625488 214588 625494 214600
rect 626074 214588 626080 214600
rect 625488 214560 626080 214588
rect 625488 214548 625494 214560
rect 626074 214548 626080 214560
rect 626132 214548 626138 214600
rect 630030 214548 630036 214600
rect 630088 214588 630094 214600
rect 632882 214588 632888 214600
rect 630088 214560 632888 214588
rect 630088 214548 630094 214560
rect 632882 214548 632888 214560
rect 632940 214548 632946 214600
rect 646314 214548 646320 214600
rect 646372 214588 646378 214600
rect 656158 214588 656164 214600
rect 646372 214560 656164 214588
rect 646372 214548 646378 214560
rect 656158 214548 656164 214560
rect 656216 214548 656222 214600
rect 629386 214452 629392 214464
rect 625126 214424 629392 214452
rect 629386 214412 629392 214424
rect 629444 214412 629450 214464
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 41690 213976 41696 213988
rect 35860 213948 41696 213976
rect 35860 213936 35866 213948
rect 41690 213936 41696 213948
rect 41748 213936 41754 213988
rect 645854 213868 645860 213920
rect 645912 213908 645918 213920
rect 646498 213908 646504 213920
rect 645912 213880 646504 213908
rect 645912 213868 645918 213880
rect 646498 213868 646504 213880
rect 646556 213868 646562 213920
rect 648614 213868 648620 213920
rect 648672 213908 648678 213920
rect 649258 213908 649264 213920
rect 648672 213880 649264 213908
rect 648672 213868 648678 213880
rect 649258 213868 649264 213880
rect 649316 213868 649322 213920
rect 663150 213868 663156 213920
rect 663208 213908 663214 213920
rect 663702 213908 663708 213920
rect 663208 213880 663708 213908
rect 663208 213868 663214 213880
rect 663702 213868 663708 213880
rect 663760 213868 663766 213920
rect 653214 213800 653220 213852
rect 653272 213840 653278 213852
rect 654778 213840 654784 213852
rect 653272 213812 654784 213840
rect 653272 213800 653278 213812
rect 654778 213800 654784 213812
rect 654836 213800 654842 213852
rect 656526 213392 656532 213444
rect 656584 213432 656590 213444
rect 664622 213432 664628 213444
rect 656584 213404 664628 213432
rect 656584 213392 656590 213404
rect 664622 213392 664628 213404
rect 664680 213392 664686 213444
rect 643830 213324 643836 213376
rect 643888 213364 643894 213376
rect 653398 213364 653404 213376
rect 643888 213336 653404 213364
rect 643888 213324 643894 213336
rect 653398 213324 653404 213336
rect 653456 213324 653462 213376
rect 660758 213296 660764 213308
rect 654106 213268 660764 213296
rect 575474 213188 575480 213240
rect 575532 213228 575538 213240
rect 594794 213228 594800 213240
rect 575532 213200 594800 213228
rect 575532 213188 575538 213200
rect 594794 213188 594800 213200
rect 594852 213188 594858 213240
rect 645486 213188 645492 213240
rect 645544 213228 645550 213240
rect 654106 213228 654134 213268
rect 660758 213256 660764 213268
rect 660816 213256 660822 213308
rect 645544 213200 654134 213228
rect 645544 213188 645550 213200
rect 654594 213120 654600 213172
rect 654652 213160 654658 213172
rect 657538 213160 657544 213172
rect 654652 213132 657544 213160
rect 654652 213120 654658 213132
rect 657538 213120 657544 213132
rect 657596 213120 657602 213172
rect 600406 212984 600412 213036
rect 600464 213024 600470 213036
rect 601234 213024 601240 213036
rect 600464 212996 601240 213024
rect 600464 212984 600470 212996
rect 601234 212984 601240 212996
rect 601292 212984 601298 213036
rect 632698 212984 632704 213036
rect 632756 213024 632762 213036
rect 634354 213024 634360 213036
rect 632756 212996 634360 213024
rect 632756 212984 632762 212996
rect 634354 212984 634360 212996
rect 634412 212984 634418 213036
rect 654134 212916 654140 212968
rect 654192 212956 654198 212968
rect 654778 212956 654784 212968
rect 654192 212928 654784 212956
rect 654192 212916 654198 212928
rect 654778 212916 654784 212928
rect 654836 212916 654842 212968
rect 600498 212848 600504 212900
rect 600556 212888 600562 212900
rect 600866 212888 600872 212900
rect 600556 212860 600872 212888
rect 600556 212848 600562 212860
rect 600866 212848 600872 212860
rect 600924 212848 600930 212900
rect 35802 212780 35808 212832
rect 35860 212820 35866 212832
rect 39942 212820 39948 212832
rect 35860 212792 39948 212820
rect 35860 212780 35866 212792
rect 39942 212780 39948 212792
rect 40000 212780 40006 212832
rect 650454 212712 650460 212764
rect 650512 212752 650518 212764
rect 651282 212752 651288 212764
rect 650512 212724 651288 212752
rect 650512 212712 650518 212724
rect 651282 212712 651288 212724
rect 651340 212712 651346 212764
rect 664254 212712 664260 212764
rect 664312 212752 664318 212764
rect 665082 212752 665088 212764
rect 664312 212724 665088 212752
rect 664312 212712 664318 212724
rect 665082 212712 665088 212724
rect 665140 212712 665146 212764
rect 592678 212644 592684 212696
rect 592736 212684 592742 212696
rect 641714 212684 641720 212696
rect 592736 212656 641720 212684
rect 592736 212644 592742 212656
rect 641714 212644 641720 212656
rect 641772 212644 641778 212696
rect 35618 212508 35624 212560
rect 35676 212548 35682 212560
rect 39574 212548 39580 212560
rect 35676 212520 39580 212548
rect 35676 212508 35682 212520
rect 39574 212508 39580 212520
rect 39632 212508 39638 212560
rect 591298 212508 591304 212560
rect 591356 212548 591362 212560
rect 639874 212548 639880 212560
rect 591356 212520 639880 212548
rect 591356 212508 591362 212520
rect 639874 212508 639880 212520
rect 639932 212508 639938 212560
rect 578510 211148 578516 211200
rect 578568 211188 578574 211200
rect 580902 211188 580908 211200
rect 578568 211160 580908 211188
rect 578568 211148 578574 211160
rect 580902 211148 580908 211160
rect 580960 211148 580966 211200
rect 35802 209924 35808 209976
rect 35860 209964 35866 209976
rect 40402 209964 40408 209976
rect 35860 209936 40408 209964
rect 35860 209924 35866 209936
rect 40402 209924 40408 209936
rect 40460 209924 40466 209976
rect 579522 209788 579528 209840
rect 579580 209828 579586 209840
rect 582282 209828 582288 209840
rect 579580 209800 582288 209828
rect 579580 209788 579586 209800
rect 582282 209788 582288 209800
rect 582340 209788 582346 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 35802 208700 35808 208752
rect 35860 208740 35866 208752
rect 35860 208700 35894 208740
rect 35866 208672 35894 208700
rect 40034 208672 40040 208684
rect 35866 208644 40040 208672
rect 40034 208632 40040 208644
rect 40092 208632 40098 208684
rect 581638 208564 581644 208616
rect 581696 208604 581702 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652018 209516 652024 209568
rect 652076 209556 652082 209568
rect 652076 209528 654134 209556
rect 652076 209516 652082 209528
rect 654106 209080 654134 209528
rect 667750 209080 667756 209092
rect 654106 209052 667756 209080
rect 667750 209040 667756 209052
rect 667808 209040 667814 209092
rect 581696 208576 625154 208604
rect 581696 208564 581702 208576
rect 35802 208496 35808 208548
rect 35860 208536 35866 208548
rect 40586 208536 40592 208548
rect 35860 208508 40592 208536
rect 35860 208496 35866 208508
rect 40586 208496 40592 208508
rect 40644 208496 40650 208548
rect 35618 208360 35624 208412
rect 35676 208400 35682 208412
rect 41690 208400 41696 208412
rect 35676 208372 41696 208400
rect 35676 208360 35682 208372
rect 41690 208360 41696 208372
rect 41748 208360 41754 208412
rect 42058 208360 42064 208412
rect 42116 208400 42122 208412
rect 43346 208400 43352 208412
rect 42116 208372 43352 208400
rect 42116 208360 42122 208372
rect 43346 208360 43352 208372
rect 43404 208360 43410 208412
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 35802 207136 35808 207188
rect 35860 207176 35866 207188
rect 39942 207176 39948 207188
rect 35860 207148 39948 207176
rect 35860 207136 35866 207148
rect 39942 207136 39948 207148
rect 40000 207136 40006 207188
rect 580902 206864 580908 206916
rect 580960 206904 580966 206916
rect 589458 206904 589464 206916
rect 580960 206876 589464 206904
rect 580960 206864 580966 206876
rect 589458 206864 589464 206876
rect 589516 206864 589522 206916
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 582282 205504 582288 205556
rect 582340 205544 582346 205556
rect 589458 205544 589464 205556
rect 582340 205516 589464 205544
rect 582340 205504 582346 205516
rect 589458 205504 589464 205516
rect 589516 205504 589522 205556
rect 35802 204620 35808 204672
rect 35860 204660 35866 204672
rect 35860 204620 35894 204660
rect 35866 204592 35894 204620
rect 35866 204564 41414 204592
rect 41386 204524 41414 204564
rect 41506 204524 41512 204536
rect 41386 204496 41512 204524
rect 41506 204484 41512 204496
rect 41564 204484 41570 204536
rect 41690 204388 41696 204400
rect 36004 204360 41696 204388
rect 35802 204280 35808 204332
rect 35860 204320 35866 204332
rect 36004 204320 36032 204360
rect 41690 204348 41696 204360
rect 41748 204348 41754 204400
rect 35860 204292 36032 204320
rect 35860 204280 35866 204292
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 37918 202892 37924 202904
rect 35860 202864 37924 202892
rect 35860 202852 35866 202864
rect 37918 202852 37924 202864
rect 37976 202852 37982 202904
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 43254 202144 43260 202156
rect 43088 202116 43260 202144
rect 42518 201696 42524 201748
rect 42576 201736 42582 201748
rect 42886 201736 42892 201748
rect 42576 201708 42892 201736
rect 42576 201696 42582 201708
rect 42886 201696 42892 201708
rect 42944 201696 42950 201748
rect 43088 201612 43116 202116
rect 43254 202104 43260 202116
rect 43312 202104 43318 202156
rect 42702 201560 42708 201612
rect 42760 201560 42766 201612
rect 43070 201560 43076 201612
rect 43128 201560 43134 201612
rect 42720 201328 42748 201560
rect 42886 201328 42892 201340
rect 42720 201300 42892 201328
rect 42886 201288 42892 201300
rect 42944 201288 42950 201340
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 42242 190204 42248 190256
rect 42300 190244 42306 190256
rect 42886 190244 42892 190256
rect 42300 190216 42892 190244
rect 42300 190204 42306 190216
rect 42886 190204 42892 190216
rect 42944 190204 42950 190256
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 42426 187620 42432 187672
rect 42484 187660 42490 187672
rect 43070 187660 43076 187672
rect 42484 187632 43076 187660
rect 42484 187620 42490 187632
rect 43070 187620 43076 187632
rect 43128 187620 43134 187672
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 668946 184832 668952 184884
rect 669004 184872 669010 184884
rect 670694 184872 670700 184884
rect 669004 184844 670700 184872
rect 669004 184832 669010 184844
rect 670694 184832 670700 184844
rect 670752 184832 670758 184884
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 668210 177964 668216 178016
rect 668268 178004 668274 178016
rect 670786 178004 670792 178016
rect 668268 177976 670792 178004
rect 668268 177964 668274 177976
rect 670786 177964 670792 177976
rect 670844 177964 670850 178016
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 668026 175040 668032 175092
rect 668084 175080 668090 175092
rect 670418 175080 670424 175092
rect 668084 175052 670424 175080
rect 668084 175040 668090 175052
rect 670418 175040 670424 175052
rect 670476 175040 670482 175092
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 580258 171096 580264 171148
rect 580316 171136 580322 171148
rect 589458 171136 589464 171148
rect 580316 171108 589464 171136
rect 580316 171096 580322 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 667934 169668 667940 169720
rect 667992 169708 667998 169720
rect 669682 169708 669688 169720
rect 667992 169680 669688 169708
rect 667992 169668 667998 169680
rect 669682 169668 669688 169680
rect 669740 169668 669746 169720
rect 582374 168376 582380 168428
rect 582432 168416 582438 168428
rect 589458 168416 589464 168428
rect 582432 168388 589464 168416
rect 582432 168376 582438 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 578234 167288 578240 167340
rect 578292 167328 578298 167340
rect 580258 167328 580264 167340
rect 578292 167300 580264 167328
rect 578292 167288 578298 167300
rect 580258 167288 580264 167300
rect 580316 167288 580322 167340
rect 579982 167016 579988 167068
rect 580040 167056 580046 167068
rect 589458 167056 589464 167068
rect 580040 167028 589464 167056
rect 580040 167016 580046 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589642 166308 589648 166320
rect 579580 166280 589648 166308
rect 579580 166268 579586 166280
rect 589642 166268 589648 166280
rect 589700 166268 589706 166320
rect 579338 165180 579344 165232
rect 579396 165220 579402 165232
rect 582374 165220 582380 165232
rect 579396 165192 582380 165220
rect 579396 165180 579402 165192
rect 582374 165180 582380 165192
rect 582432 165180 582438 165232
rect 667934 165044 667940 165096
rect 667992 165084 667998 165096
rect 670050 165084 670056 165096
rect 667992 165056 670056 165084
rect 667992 165044 667998 165056
rect 670050 165044 670056 165056
rect 670108 165044 670114 165096
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 675846 164160 675852 164212
rect 675904 164200 675910 164212
rect 682378 164200 682384 164212
rect 675904 164172 682384 164200
rect 675904 164160 675910 164172
rect 682378 164160 682384 164172
rect 682436 164160 682442 164212
rect 578234 163616 578240 163668
rect 578292 163656 578298 163668
rect 579982 163656 579988 163668
rect 578292 163628 579988 163656
rect 578292 163616 578298 163628
rect 579982 163616 579988 163628
rect 580040 163616 580046 163668
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 578418 162664 578424 162716
rect 578476 162704 578482 162716
rect 582466 162704 582472 162716
rect 578476 162676 582472 162704
rect 578476 162664 578482 162676
rect 582466 162664 582472 162676
rect 582524 162664 582530 162716
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580718 160080 580724 160132
rect 580776 160120 580782 160132
rect 589458 160120 589464 160132
rect 580776 160092 589464 160120
rect 580776 160080 580782 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 668210 160012 668216 160064
rect 668268 160052 668274 160064
rect 670786 160052 670792 160064
rect 668268 160024 670792 160052
rect 668268 160012 668274 160024
rect 670786 160012 670792 160024
rect 670844 160012 670850 160064
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 585778 158720 585784 158772
rect 585836 158760 585842 158772
rect 589458 158760 589464 158772
rect 585836 158732 589464 158760
rect 585836 158720 585842 158732
rect 589458 158720 589464 158732
rect 589516 158720 589522 158772
rect 587158 157360 587164 157412
rect 587216 157400 587222 157412
rect 589274 157400 589280 157412
rect 587216 157372 589280 157400
rect 587216 157360 587222 157372
rect 589274 157360 589280 157372
rect 589332 157360 589338 157412
rect 668210 155524 668216 155576
rect 668268 155564 668274 155576
rect 670786 155564 670792 155576
rect 668268 155536 670792 155564
rect 668268 155524 668274 155536
rect 670786 155524 670792 155536
rect 670844 155524 670850 155576
rect 578326 154640 578332 154692
rect 578384 154680 578390 154692
rect 580534 154680 580540 154692
rect 578384 154652 580540 154680
rect 578384 154640 578390 154652
rect 580534 154640 580540 154652
rect 580592 154640 580598 154692
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 580718 152776 580724 152788
rect 578292 152748 580724 152776
rect 578292 152736 578298 152748
rect 580718 152736 580724 152748
rect 580776 152736 580782 152788
rect 580258 151784 580264 151836
rect 580316 151824 580322 151836
rect 589458 151824 589464 151836
rect 580316 151796 589464 151824
rect 580316 151784 580322 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 585778 150600 585784 150612
rect 578936 150572 585784 150600
rect 578936 150560 578942 150572
rect 585778 150560 585784 150572
rect 585836 150560 585842 150612
rect 585134 149064 585140 149116
rect 585192 149104 585198 149116
rect 589458 149104 589464 149116
rect 585192 149076 589464 149104
rect 585192 149064 585198 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 579522 148316 579528 148368
rect 579580 148356 579586 148368
rect 587158 148356 587164 148368
rect 579580 148328 587164 148356
rect 579580 148316 579586 148328
rect 587158 148316 587164 148328
rect 587216 148316 587222 148368
rect 578878 146276 578884 146328
rect 578936 146316 578942 146328
rect 585134 146316 585140 146328
rect 578936 146288 585140 146316
rect 578936 146276 578942 146288
rect 585134 146276 585140 146288
rect 585192 146276 585198 146328
rect 668762 145732 668768 145784
rect 668820 145772 668826 145784
rect 670786 145772 670792 145784
rect 668820 145744 670792 145772
rect 668820 145732 668826 145744
rect 670786 145732 670792 145744
rect 670844 145732 670850 145784
rect 584766 144916 584772 144968
rect 584824 144956 584830 144968
rect 589458 144956 589464 144968
rect 584824 144928 589464 144956
rect 584824 144916 584830 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 585962 143556 585968 143608
rect 586020 143596 586026 143608
rect 589458 143596 589464 143608
rect 586020 143568 589464 143596
rect 586020 143556 586026 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 587158 142400 587164 142452
rect 587216 142440 587222 142452
rect 589826 142440 589832 142452
rect 587216 142412 589832 142440
rect 587216 142400 587222 142412
rect 589826 142400 589832 142412
rect 589884 142400 589890 142452
rect 580442 140768 580448 140820
rect 580500 140808 580506 140820
rect 589458 140808 589464 140820
rect 580500 140780 589464 140808
rect 580500 140768 580506 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580258 140740 580264 140752
rect 578660 140712 580264 140740
rect 578660 140700 578666 140712
rect 580258 140700 580264 140712
rect 580316 140700 580322 140752
rect 583018 139408 583024 139460
rect 583076 139448 583082 139460
rect 589458 139448 589464 139460
rect 583076 139420 589464 139448
rect 583076 139408 583082 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 579522 138660 579528 138712
rect 579580 138700 579586 138712
rect 588538 138700 588544 138712
rect 579580 138672 588544 138700
rect 579580 138660 579586 138672
rect 588538 138660 588544 138672
rect 588596 138660 588602 138712
rect 579062 137300 579068 137352
rect 579120 137340 579126 137352
rect 584766 137340 584772 137352
rect 579120 137312 584772 137340
rect 579120 137300 579126 137312
rect 584766 137300 584772 137312
rect 584824 137300 584830 137352
rect 584582 136620 584588 136672
rect 584640 136660 584646 136672
rect 589458 136660 589464 136672
rect 584640 136632 589464 136660
rect 584640 136620 584646 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 580258 134512 580264 134564
rect 580316 134552 580322 134564
rect 589458 134552 589464 134564
rect 580316 134524 589464 134552
rect 580316 134512 580322 134524
rect 589458 134512 589464 134524
rect 589516 134512 589522 134564
rect 675846 133900 675852 133952
rect 675904 133940 675910 133952
rect 676490 133940 676496 133952
rect 675904 133912 676496 133940
rect 675904 133900 675910 133912
rect 676490 133900 676496 133912
rect 676548 133900 676554 133952
rect 667934 133764 667940 133816
rect 667992 133804 667998 133816
rect 669866 133804 669872 133816
rect 667992 133776 669872 133804
rect 667992 133764 667998 133776
rect 669866 133764 669872 133776
rect 669924 133764 669930 133816
rect 585778 132472 585784 132524
rect 585836 132512 585842 132524
rect 589458 132512 589464 132524
rect 585836 132484 589464 132512
rect 585836 132472 585842 132484
rect 589458 132472 589464 132484
rect 589516 132472 589522 132524
rect 581822 131248 581828 131300
rect 581880 131288 581886 131300
rect 589458 131288 589464 131300
rect 581880 131260 589464 131288
rect 581880 131248 581886 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 578878 131112 578884 131164
rect 578936 131152 578942 131164
rect 585962 131152 585968 131164
rect 578936 131124 585968 131152
rect 578936 131112 578942 131124
rect 585962 131112 585968 131124
rect 586020 131112 586026 131164
rect 668486 130772 668492 130824
rect 668544 130812 668550 130824
rect 670786 130812 670792 130824
rect 668544 130784 670792 130812
rect 668544 130772 668550 130784
rect 670786 130772 670792 130784
rect 670844 130772 670850 130824
rect 668026 129684 668032 129736
rect 668084 129724 668090 129736
rect 670142 129724 670148 129736
rect 668084 129696 670148 129724
rect 668084 129684 668090 129696
rect 670142 129684 670148 129696
rect 670200 129684 670206 129736
rect 583202 129140 583208 129192
rect 583260 129180 583266 129192
rect 590378 129180 590384 129192
rect 583260 129152 590384 129180
rect 583260 129140 583266 129152
rect 590378 129140 590384 129152
rect 590436 129140 590442 129192
rect 579522 129004 579528 129056
rect 579580 129044 579586 129056
rect 587158 129044 587164 129056
rect 579580 129016 587164 129044
rect 579580 129004 579586 129016
rect 587158 129004 587164 129016
rect 587216 129004 587222 129056
rect 579062 126964 579068 127016
rect 579120 127004 579126 127016
rect 589458 127004 589464 127016
rect 579120 126976 589464 127004
rect 579120 126964 579126 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 578326 125604 578332 125656
rect 578384 125644 578390 125656
rect 580442 125644 580448 125656
rect 578384 125616 580448 125644
rect 578384 125604 578390 125616
rect 580442 125604 580448 125616
rect 580500 125604 580506 125656
rect 675846 125400 675852 125452
rect 675904 125440 675910 125452
rect 676398 125440 676404 125452
rect 675904 125412 676404 125440
rect 675904 125400 675910 125412
rect 676398 125400 676404 125412
rect 676456 125400 676462 125452
rect 580442 124176 580448 124228
rect 580500 124216 580506 124228
rect 589458 124216 589464 124228
rect 580500 124188 589464 124216
rect 580500 124176 580506 124188
rect 589458 124176 589464 124188
rect 589516 124176 589522 124228
rect 578418 123564 578424 123616
rect 578476 123604 578482 123616
rect 583018 123604 583024 123616
rect 578476 123576 583024 123604
rect 578476 123564 578482 123576
rect 583018 123564 583024 123576
rect 583076 123564 583082 123616
rect 584398 122816 584404 122868
rect 584456 122856 584462 122868
rect 589458 122856 589464 122868
rect 584456 122828 589464 122856
rect 584456 122816 584462 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 578878 122136 578884 122188
rect 578936 122176 578942 122188
rect 584582 122176 584588 122188
rect 578936 122148 584588 122176
rect 578936 122136 578942 122148
rect 584582 122136 584588 122148
rect 584640 122136 584646 122188
rect 580626 122000 580632 122052
rect 580684 122040 580690 122052
rect 589918 122040 589924 122052
rect 580684 122012 589924 122040
rect 580684 122000 580690 122012
rect 589918 122000 589924 122012
rect 589976 122000 589982 122052
rect 587342 118668 587348 118720
rect 587400 118708 587406 118720
rect 590010 118708 590016 118720
rect 587400 118680 590016 118708
rect 587400 118668 587406 118680
rect 590010 118668 590016 118680
rect 590068 118668 590074 118720
rect 675846 118464 675852 118516
rect 675904 118504 675910 118516
rect 679618 118504 679624 118516
rect 675904 118476 679624 118504
rect 675904 118464 675910 118476
rect 679618 118464 679624 118476
rect 679676 118464 679682 118516
rect 578510 118396 578516 118448
rect 578568 118436 578574 118448
rect 580258 118436 580264 118448
rect 578568 118408 580264 118436
rect 578568 118396 578574 118408
rect 580258 118396 580264 118408
rect 580316 118396 580322 118448
rect 579522 116900 579528 116952
rect 579580 116940 579586 116952
rect 583202 116940 583208 116952
rect 579580 116912 583208 116940
rect 579580 116900 579586 116912
rect 583202 116900 583208 116912
rect 583260 116900 583266 116952
rect 668762 116832 668768 116884
rect 668820 116872 668826 116884
rect 670602 116872 670608 116884
rect 668820 116844 670608 116872
rect 668820 116832 668826 116844
rect 670602 116832 670608 116844
rect 670660 116832 670666 116884
rect 586146 115948 586152 116000
rect 586204 115988 586210 116000
rect 589458 115988 589464 116000
rect 586204 115960 589464 115988
rect 586204 115948 586210 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 583202 115200 583208 115252
rect 583260 115240 583266 115252
rect 589642 115240 589648 115252
rect 583260 115212 589648 115240
rect 583260 115200 583266 115212
rect 589642 115200 589648 115212
rect 589700 115200 589706 115252
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 583018 113160 583024 113212
rect 583076 113200 583082 113212
rect 589458 113200 589464 113212
rect 583076 113172 589464 113200
rect 583076 113160 583082 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 579522 112820 579528 112872
rect 579580 112860 579586 112872
rect 585778 112860 585784 112872
rect 579580 112832 585784 112860
rect 579580 112820 579586 112832
rect 585778 112820 585784 112832
rect 585836 112820 585842 112872
rect 585962 112412 585968 112464
rect 586020 112452 586026 112464
rect 590102 112452 590108 112464
rect 586020 112424 590108 112452
rect 586020 112412 586026 112424
rect 590102 112412 590108 112424
rect 590160 112412 590166 112464
rect 581638 110440 581644 110492
rect 581696 110480 581702 110492
rect 589458 110480 589464 110492
rect 581696 110452 589464 110480
rect 581696 110440 581702 110452
rect 589458 110440 589464 110452
rect 589516 110440 589522 110492
rect 579338 110100 579344 110152
rect 579396 110140 579402 110152
rect 581822 110140 581828 110152
rect 579396 110112 581828 110140
rect 579396 110100 579402 110112
rect 581822 110100 581828 110112
rect 581880 110100 581886 110152
rect 584582 109012 584588 109064
rect 584640 109052 584646 109064
rect 589274 109052 589280 109064
rect 584640 109024 589280 109052
rect 584640 109012 584646 109024
rect 589274 109012 589280 109024
rect 589332 109012 589338 109064
rect 667934 108808 667940 108860
rect 667992 108848 667998 108860
rect 669958 108848 669964 108860
rect 667992 108820 669964 108848
rect 667992 108808 667998 108820
rect 669958 108808 669964 108820
rect 670016 108808 670022 108860
rect 578326 108672 578332 108724
rect 578384 108712 578390 108724
rect 580626 108712 580632 108724
rect 578384 108684 580632 108712
rect 578384 108672 578390 108684
rect 580626 108672 580632 108684
rect 580684 108672 580690 108724
rect 589458 107692 589464 107704
rect 579632 107664 589464 107692
rect 578878 107584 578884 107636
rect 578936 107624 578942 107636
rect 579632 107624 579660 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 578936 107596 579660 107624
rect 578936 107584 578942 107596
rect 587158 106292 587164 106344
rect 587216 106332 587222 106344
rect 589826 106332 589832 106344
rect 587216 106304 589832 106332
rect 587216 106292 587222 106304
rect 589826 106292 589832 106304
rect 589884 106292 589890 106344
rect 668394 106156 668400 106208
rect 668452 106196 668458 106208
rect 670786 106196 670792 106208
rect 668452 106168 670792 106196
rect 668452 106156 668458 106168
rect 670786 106156 670792 106168
rect 670844 106156 670850 106208
rect 580258 104864 580264 104916
rect 580316 104904 580322 104916
rect 589458 104904 589464 104916
rect 580316 104876 589464 104904
rect 580316 104864 580322 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 668762 104660 668768 104712
rect 668820 104700 668826 104712
rect 670786 104700 670792 104712
rect 668820 104672 670792 104700
rect 668820 104660 668826 104672
rect 670786 104660 670792 104672
rect 670844 104660 670850 104712
rect 579522 103436 579528 103488
rect 579580 103476 579586 103488
rect 588538 103476 588544 103488
rect 579580 103448 588544 103476
rect 579580 103436 579586 103448
rect 588538 103436 588544 103448
rect 588596 103436 588602 103488
rect 579522 101804 579528 101856
rect 579580 101844 579586 101856
rect 584398 101844 584404 101856
rect 579580 101816 584404 101844
rect 579580 101804 579586 101816
rect 584398 101804 584404 101816
rect 584456 101804 584462 101856
rect 584398 100104 584404 100156
rect 584456 100144 584462 100156
rect 589458 100144 589464 100156
rect 584456 100116 589464 100144
rect 584456 100104 584462 100116
rect 589458 100104 589464 100116
rect 589516 100104 589522 100156
rect 579062 99356 579068 99408
rect 579120 99396 579126 99408
rect 586146 99396 586152 99408
rect 579120 99368 586152 99396
rect 579120 99356 579126 99368
rect 586146 99356 586152 99368
rect 586204 99356 586210 99408
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 578602 99220 578608 99272
rect 578660 99260 578666 99272
rect 580442 99260 580448 99272
rect 578660 99232 580448 99260
rect 578660 99220 578666 99232
rect 580442 99220 580448 99232
rect 580500 99220 580506 99272
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633434 99192 633440 99204
rect 623740 99164 633440 99192
rect 623740 99152 623746 99164
rect 633434 99152 633440 99164
rect 633492 99152 633498 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 625062 99016 625068 99068
rect 625120 99056 625126 99068
rect 636286 99056 636292 99068
rect 625120 99028 636292 99056
rect 625120 99016 625126 99028
rect 636286 99016 636292 99028
rect 636344 99016 636350 99068
rect 628282 98880 628288 98932
rect 628340 98920 628346 98932
rect 642174 98920 642180 98932
rect 628340 98892 642180 98920
rect 628340 98880 628346 98892
rect 642174 98880 642180 98892
rect 642232 98880 642238 98932
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 643646 98784 643652 98796
rect 629076 98756 643652 98784
rect 629076 98744 629082 98756
rect 643646 98744 643652 98756
rect 643704 98744 643710 98796
rect 647142 98744 647148 98796
rect 647200 98784 647206 98796
rect 661954 98784 661960 98796
rect 647200 98756 661960 98784
rect 647200 98744 647206 98756
rect 661954 98744 661960 98756
rect 662012 98744 662018 98796
rect 630490 98608 630496 98660
rect 630548 98648 630554 98660
rect 646590 98648 646596 98660
rect 630548 98620 646596 98648
rect 630548 98608 630554 98620
rect 646590 98608 646596 98620
rect 646648 98608 646654 98660
rect 631042 98200 631048 98252
rect 631100 98240 631106 98252
rect 631100 98212 634814 98240
rect 631100 98200 631106 98212
rect 634786 98172 634814 98212
rect 640702 98172 640708 98184
rect 634786 98144 640708 98172
rect 640702 98132 640708 98144
rect 640760 98132 640766 98184
rect 631980 98076 632192 98104
rect 578326 97928 578332 97980
rect 578384 97968 578390 97980
rect 587342 97968 587348 97980
rect 578384 97940 587348 97968
rect 578384 97928 578390 97940
rect 587342 97928 587348 97940
rect 587400 97928 587406 97980
rect 618714 97928 618720 97980
rect 618772 97968 618778 97980
rect 625798 97968 625804 97980
rect 618772 97940 625804 97968
rect 618772 97928 618778 97940
rect 625798 97928 625804 97940
rect 625856 97928 625862 97980
rect 629754 97928 629760 97980
rect 629812 97968 629818 97980
rect 631980 97968 632008 98076
rect 632164 98036 632192 98076
rect 645302 98036 645308 98048
rect 632164 98008 645308 98036
rect 645302 97996 645308 98008
rect 645360 97996 645366 98048
rect 629812 97940 632008 97968
rect 629812 97928 629818 97940
rect 659930 97928 659936 97980
rect 659988 97968 659994 97980
rect 665174 97968 665180 97980
rect 659988 97940 665180 97968
rect 659988 97928 659994 97940
rect 665174 97928 665180 97940
rect 665232 97928 665238 97980
rect 620186 97792 620192 97844
rect 620244 97832 620250 97844
rect 625614 97832 625620 97844
rect 620244 97804 625620 97832
rect 620244 97792 620250 97804
rect 625614 97792 625620 97804
rect 625672 97792 625678 97844
rect 627546 97792 627552 97844
rect 627604 97832 627610 97844
rect 631042 97832 631048 97844
rect 627604 97804 631048 97832
rect 627604 97792 627610 97804
rect 631042 97792 631048 97804
rect 631100 97792 631106 97844
rect 631962 97792 631968 97844
rect 632020 97832 632026 97844
rect 647510 97832 647516 97844
rect 632020 97804 647516 97832
rect 632020 97792 632026 97804
rect 647510 97792 647516 97804
rect 647568 97792 647574 97844
rect 655422 97792 655428 97844
rect 655480 97832 655486 97844
rect 662506 97832 662512 97844
rect 655480 97804 662512 97832
rect 655480 97792 655486 97804
rect 662506 97792 662512 97804
rect 662564 97792 662570 97844
rect 632698 97656 632704 97708
rect 632756 97696 632762 97708
rect 648246 97696 648252 97708
rect 632756 97668 648252 97696
rect 632756 97656 632762 97668
rect 648246 97656 648252 97668
rect 648304 97656 648310 97708
rect 651834 97656 651840 97708
rect 651892 97696 651898 97708
rect 659562 97696 659568 97708
rect 651892 97668 659568 97696
rect 651892 97656 651898 97668
rect 659562 97656 659568 97668
rect 659620 97656 659626 97708
rect 621658 97520 621664 97572
rect 621716 97560 621722 97572
rect 629294 97560 629300 97572
rect 621716 97532 629300 97560
rect 621716 97520 621722 97532
rect 629294 97520 629300 97532
rect 629352 97520 629358 97572
rect 634170 97520 634176 97572
rect 634228 97560 634234 97572
rect 634228 97532 649994 97560
rect 634228 97520 634234 97532
rect 612642 97384 612648 97436
rect 612700 97424 612706 97436
rect 618898 97424 618904 97436
rect 612700 97396 618904 97424
rect 612700 97384 612706 97396
rect 618898 97384 618904 97396
rect 618956 97384 618962 97436
rect 623130 97384 623136 97436
rect 623188 97424 623194 97436
rect 632054 97424 632060 97436
rect 623188 97396 632060 97424
rect 623188 97384 623194 97396
rect 632054 97384 632060 97396
rect 632112 97384 632118 97436
rect 633250 97384 633256 97436
rect 633308 97424 633314 97436
rect 648614 97424 648620 97436
rect 633308 97396 648620 97424
rect 633308 97384 633314 97396
rect 648614 97384 648620 97396
rect 648672 97384 648678 97436
rect 649966 97424 649994 97532
rect 650362 97520 650368 97572
rect 650420 97560 650426 97572
rect 658274 97560 658280 97572
rect 650420 97532 658280 97560
rect 650420 97520 650426 97532
rect 658274 97520 658280 97532
rect 658332 97520 658338 97572
rect 650546 97424 650552 97436
rect 649966 97396 650552 97424
rect 650546 97384 650552 97396
rect 650604 97384 650610 97436
rect 658090 97384 658096 97436
rect 658148 97424 658154 97436
rect 663058 97424 663064 97436
rect 658148 97396 663064 97424
rect 658148 97384 658154 97396
rect 663058 97384 663064 97396
rect 663116 97384 663122 97436
rect 605466 97248 605472 97300
rect 605524 97288 605530 97300
rect 611906 97288 611912 97300
rect 605524 97260 611912 97288
rect 605524 97248 605530 97260
rect 611906 97248 611912 97260
rect 611964 97248 611970 97300
rect 626074 97248 626080 97300
rect 626132 97288 626138 97300
rect 637758 97288 637764 97300
rect 626132 97260 637764 97288
rect 626132 97248 626138 97260
rect 637758 97248 637764 97260
rect 637816 97248 637822 97300
rect 643002 97248 643008 97300
rect 643060 97288 643066 97300
rect 656526 97288 656532 97300
rect 643060 97260 656532 97288
rect 643060 97248 643066 97260
rect 656526 97248 656532 97260
rect 656584 97248 656590 97300
rect 656802 97248 656808 97300
rect 656860 97288 656866 97300
rect 661402 97288 661408 97300
rect 656860 97260 661408 97288
rect 656860 97248 656866 97260
rect 661402 97248 661408 97260
rect 661460 97248 661466 97300
rect 626810 97112 626816 97164
rect 626868 97152 626874 97164
rect 639230 97152 639236 97164
rect 626868 97124 639236 97152
rect 626868 97112 626874 97124
rect 639230 97112 639236 97124
rect 639288 97112 639294 97164
rect 644290 97112 644296 97164
rect 644348 97152 644354 97164
rect 658826 97152 658832 97164
rect 644348 97124 658832 97152
rect 644348 97112 644354 97124
rect 658826 97112 658832 97124
rect 658884 97112 658890 97164
rect 624602 96976 624608 97028
rect 624660 97016 624666 97028
rect 634998 97016 635004 97028
rect 624660 96988 635004 97016
rect 624660 96976 624666 96988
rect 634998 96976 635004 96988
rect 635056 96976 635062 97028
rect 635550 96976 635556 97028
rect 635608 97016 635614 97028
rect 647694 97016 647700 97028
rect 635608 96988 647700 97016
rect 635608 96976 635614 96988
rect 647694 96976 647700 96988
rect 647752 96976 647758 97028
rect 659194 96976 659200 97028
rect 659252 97016 659258 97028
rect 663886 97016 663892 97028
rect 659252 96988 663892 97016
rect 659252 96976 659258 96988
rect 663886 96976 663892 96988
rect 663944 96976 663950 97028
rect 596174 96908 596180 96960
rect 596232 96948 596238 96960
rect 596726 96948 596732 96960
rect 596232 96920 596732 96948
rect 596232 96908 596238 96920
rect 596726 96908 596732 96920
rect 596784 96908 596790 96960
rect 597646 96908 597652 96960
rect 597704 96948 597710 96960
rect 598198 96948 598204 96960
rect 597704 96920 598204 96948
rect 597704 96908 597710 96920
rect 598198 96908 598204 96920
rect 598256 96908 598262 96960
rect 598934 96908 598940 96960
rect 598992 96948 598998 96960
rect 599670 96948 599676 96960
rect 598992 96920 599676 96948
rect 598992 96908 598998 96920
rect 599670 96908 599676 96920
rect 599728 96908 599734 96960
rect 600314 96908 600320 96960
rect 600372 96948 600378 96960
rect 601142 96948 601148 96960
rect 600372 96920 601148 96948
rect 600372 96908 600378 96920
rect 601142 96908 601148 96920
rect 601200 96908 601206 96960
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 607122 96948 607128 96960
rect 606260 96920 607128 96948
rect 606260 96908 606266 96920
rect 607122 96908 607128 96920
rect 607180 96908 607186 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 617242 96840 617248 96892
rect 617300 96880 617306 96892
rect 618162 96880 618168 96892
rect 617300 96852 618168 96880
rect 617300 96840 617306 96852
rect 618162 96840 618168 96852
rect 618220 96840 618226 96892
rect 634722 96840 634728 96892
rect 634780 96880 634786 96892
rect 650362 96880 650368 96892
rect 634780 96852 650368 96880
rect 634780 96840 634786 96852
rect 650362 96840 650368 96852
rect 650420 96840 650426 96892
rect 653950 96840 653956 96892
rect 654008 96880 654014 96892
rect 655238 96880 655244 96892
rect 654008 96852 655244 96880
rect 654008 96840 654014 96852
rect 655238 96840 655244 96852
rect 655296 96840 655302 96892
rect 656710 96840 656716 96892
rect 656768 96880 656774 96892
rect 660114 96880 660120 96892
rect 656768 96852 660120 96880
rect 656768 96840 656774 96852
rect 660114 96840 660120 96852
rect 660172 96840 660178 96892
rect 610618 96704 610624 96756
rect 610676 96744 610682 96756
rect 611262 96744 611268 96756
rect 610676 96716 611268 96744
rect 610676 96704 610682 96716
rect 611262 96704 611268 96716
rect 611320 96704 611326 96756
rect 647878 96744 647884 96756
rect 645596 96716 647884 96744
rect 640518 96568 640524 96620
rect 640576 96608 640582 96620
rect 645596 96608 645624 96716
rect 647878 96704 647884 96716
rect 647936 96704 647942 96756
rect 654778 96704 654784 96756
rect 654836 96744 654842 96756
rect 655422 96744 655428 96756
rect 654836 96716 655428 96744
rect 654836 96704 654842 96716
rect 655422 96704 655428 96716
rect 655480 96704 655486 96756
rect 656526 96704 656532 96756
rect 656584 96744 656590 96756
rect 660114 96744 660120 96756
rect 656584 96716 660120 96744
rect 656584 96704 656590 96716
rect 660114 96704 660120 96716
rect 660172 96704 660178 96756
rect 640576 96580 645624 96608
rect 640576 96568 640582 96580
rect 645762 96568 645768 96620
rect 645820 96608 645826 96620
rect 656342 96608 656348 96620
rect 645820 96580 656348 96608
rect 645820 96568 645826 96580
rect 656342 96568 656348 96580
rect 656400 96568 656406 96620
rect 639046 96432 639052 96484
rect 639104 96472 639110 96484
rect 645118 96472 645124 96484
rect 639104 96444 645124 96472
rect 639104 96432 639110 96444
rect 645118 96432 645124 96444
rect 645176 96432 645182 96484
rect 646406 96432 646412 96484
rect 646464 96472 646470 96484
rect 652018 96472 652024 96484
rect 646464 96444 652024 96472
rect 646464 96432 646470 96444
rect 652018 96432 652024 96444
rect 652076 96432 652082 96484
rect 652570 96432 652576 96484
rect 652628 96472 652634 96484
rect 665542 96472 665548 96484
rect 652628 96444 665548 96472
rect 652628 96432 652634 96444
rect 665542 96432 665548 96444
rect 665600 96432 665606 96484
rect 631226 96296 631232 96348
rect 631284 96336 631290 96348
rect 647142 96336 647148 96348
rect 631284 96308 647148 96336
rect 631284 96296 631290 96308
rect 647142 96296 647148 96308
rect 647200 96296 647206 96348
rect 648890 96296 648896 96348
rect 648948 96336 648954 96348
rect 664162 96336 664168 96348
rect 648948 96308 664168 96336
rect 648948 96296 648954 96308
rect 664162 96296 664168 96308
rect 664220 96296 664226 96348
rect 637574 96160 637580 96212
rect 637632 96200 637638 96212
rect 660666 96200 660672 96212
rect 637632 96172 660672 96200
rect 637632 96160 637638 96172
rect 660666 96160 660672 96172
rect 660724 96160 660730 96212
rect 611078 96024 611084 96076
rect 611136 96064 611142 96076
rect 622302 96064 622308 96076
rect 611136 96036 622308 96064
rect 611136 96024 611142 96036
rect 622302 96024 622308 96036
rect 622360 96024 622366 96076
rect 649902 96024 649908 96076
rect 649960 96064 649966 96076
rect 663702 96064 663708 96076
rect 649960 96036 663708 96064
rect 649960 96024 649966 96036
rect 663702 96024 663708 96036
rect 663760 96024 663766 96076
rect 644934 95956 644940 96008
rect 644992 95996 644998 96008
rect 649534 95996 649540 96008
rect 644992 95968 649540 95996
rect 644992 95956 644998 95968
rect 649534 95956 649540 95968
rect 649592 95956 649598 96008
rect 607674 95888 607680 95940
rect 607732 95928 607738 95940
rect 624970 95928 624976 95940
rect 607732 95900 624976 95928
rect 607732 95888 607738 95900
rect 624970 95888 624976 95900
rect 625028 95888 625034 95940
rect 665358 95928 665364 95940
rect 656866 95900 665364 95928
rect 643462 95820 643468 95872
rect 643520 95860 643526 95872
rect 649258 95860 649264 95872
rect 643520 95832 649264 95860
rect 643520 95820 643526 95832
rect 649258 95820 649264 95832
rect 649316 95820 649322 95872
rect 656866 95860 656894 95900
rect 665358 95888 665364 95900
rect 665416 95888 665422 95940
rect 649460 95832 656894 95860
rect 638586 95684 638592 95736
rect 638644 95724 638650 95736
rect 647326 95724 647332 95736
rect 638644 95696 647332 95724
rect 638644 95684 638650 95696
rect 647326 95684 647332 95696
rect 647384 95684 647390 95736
rect 647878 95684 647884 95736
rect 647936 95724 647942 95736
rect 649460 95724 649488 95832
rect 647936 95696 649488 95724
rect 647936 95684 647942 95696
rect 653306 95616 653312 95668
rect 653364 95656 653370 95668
rect 664346 95656 664352 95668
rect 653364 95628 664352 95656
rect 653364 95616 653370 95628
rect 664346 95616 664352 95628
rect 664404 95616 664410 95668
rect 640058 95548 640064 95600
rect 640116 95588 640122 95600
rect 647878 95588 647884 95600
rect 640116 95560 647884 95588
rect 640116 95548 640122 95560
rect 647878 95548 647884 95560
rect 647936 95548 647942 95600
rect 641530 95412 641536 95464
rect 641588 95412 641594 95464
rect 645118 95412 645124 95464
rect 645176 95452 645182 95464
rect 651834 95452 651840 95464
rect 645176 95424 651840 95452
rect 645176 95412 645182 95424
rect 651834 95412 651840 95424
rect 651892 95412 651898 95464
rect 641548 95316 641576 95412
rect 649902 95316 649908 95328
rect 641548 95288 649908 95316
rect 649902 95276 649908 95288
rect 649960 95276 649966 95328
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 626442 95180 626448 95192
rect 620980 95152 626448 95180
rect 620980 95140 620986 95152
rect 626442 95140 626448 95152
rect 626500 95140 626506 95192
rect 647694 95072 647700 95124
rect 647752 95112 647758 95124
rect 648798 95112 648804 95124
rect 647752 95084 648804 95112
rect 647752 95072 647758 95084
rect 648798 95072 648804 95084
rect 648856 95072 648862 95124
rect 579522 95004 579528 95056
rect 579580 95044 579586 95056
rect 583202 95044 583208 95056
rect 579580 95016 583208 95044
rect 579580 95004 579586 95016
rect 583202 95004 583208 95016
rect 583260 95004 583266 95056
rect 616506 95004 616512 95056
rect 616564 95044 616570 95056
rect 622946 95044 622952 95056
rect 616564 95016 622952 95044
rect 616564 95004 616570 95016
rect 622946 95004 622952 95016
rect 623004 95004 623010 95056
rect 609146 94460 609152 94512
rect 609204 94500 609210 94512
rect 620278 94500 620284 94512
rect 609204 94472 620284 94500
rect 609204 94460 609210 94472
rect 620278 94460 620284 94472
rect 620336 94460 620342 94512
rect 649534 93916 649540 93968
rect 649592 93956 649598 93968
rect 656158 93956 656164 93968
rect 649592 93928 656164 93956
rect 649592 93916 649598 93928
rect 656158 93916 656164 93928
rect 656216 93916 656222 93968
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 651282 93508 651288 93560
rect 651340 93548 651346 93560
rect 655422 93548 655428 93560
rect 651340 93520 655428 93548
rect 651340 93508 651346 93520
rect 655422 93508 655428 93520
rect 655480 93508 655486 93560
rect 578510 93440 578516 93492
rect 578568 93480 578574 93492
rect 585962 93480 585968 93492
rect 578568 93452 585968 93480
rect 578568 93440 578574 93452
rect 585962 93440 585968 93452
rect 586020 93440 586026 93492
rect 611262 93100 611268 93152
rect 611320 93140 611326 93152
rect 619266 93140 619272 93152
rect 611320 93112 619272 93140
rect 611320 93100 611326 93112
rect 619266 93100 619272 93112
rect 619324 93100 619330 93152
rect 606938 92828 606944 92880
rect 606996 92868 607002 92880
rect 610066 92868 610072 92880
rect 606996 92840 610072 92868
rect 606996 92828 607002 92840
rect 610066 92828 610072 92840
rect 610124 92828 610130 92880
rect 648614 92488 648620 92540
rect 648672 92528 648678 92540
rect 649994 92528 650000 92540
rect 648672 92500 650000 92528
rect 648672 92488 648678 92500
rect 649994 92488 650000 92500
rect 650052 92488 650058 92540
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 626442 92460 626448 92472
rect 618036 92432 626448 92460
rect 618036 92420 618042 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 647326 92352 647332 92404
rect 647384 92392 647390 92404
rect 654318 92392 654324 92404
rect 647384 92364 654324 92392
rect 647384 92352 647390 92364
rect 654318 92352 654324 92364
rect 654376 92352 654382 92404
rect 579338 91060 579344 91112
rect 579396 91100 579402 91112
rect 584582 91100 584588 91112
rect 579396 91072 584588 91100
rect 579396 91060 579402 91072
rect 584582 91060 584588 91072
rect 584640 91060 584646 91112
rect 618162 90992 618168 91044
rect 618220 91032 618226 91044
rect 626442 91032 626448 91044
rect 618220 91004 626448 91032
rect 618220 90992 618226 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 651834 90652 651840 90704
rect 651892 90692 651898 90704
rect 655422 90692 655428 90704
rect 651892 90664 655428 90692
rect 651892 90652 651898 90664
rect 655422 90652 655428 90664
rect 655480 90652 655486 90704
rect 622946 89564 622952 89616
rect 623004 89604 623010 89616
rect 625246 89604 625252 89616
rect 623004 89576 625252 89604
rect 623004 89564 623010 89576
rect 625246 89564 625252 89576
rect 625304 89564 625310 89616
rect 585134 88952 585140 89004
rect 585192 88992 585198 89004
rect 589918 88992 589924 89004
rect 585192 88964 589924 88992
rect 585192 88952 585198 88964
rect 589918 88952 589924 88964
rect 589976 88952 589982 89004
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 663886 88788 663892 88800
rect 662380 88760 663892 88788
rect 662380 88748 662386 88760
rect 663886 88748 663892 88760
rect 663944 88748 663950 88800
rect 656342 88612 656348 88664
rect 656400 88652 656406 88664
rect 657446 88652 657452 88664
rect 656400 88624 657452 88652
rect 656400 88612 656406 88624
rect 657446 88612 657452 88624
rect 657504 88612 657510 88664
rect 610066 88272 610072 88324
rect 610124 88312 610130 88324
rect 625154 88312 625160 88324
rect 610124 88284 625160 88312
rect 610124 88272 610130 88284
rect 625154 88272 625160 88284
rect 625212 88272 625218 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 622302 88136 622308 88188
rect 622360 88176 622366 88188
rect 625338 88176 625344 88188
rect 622360 88148 625344 88176
rect 622360 88136 622366 88148
rect 625338 88136 625344 88148
rect 625396 88136 625402 88188
rect 579522 88068 579528 88120
rect 579580 88108 579586 88120
rect 585134 88108 585140 88120
rect 579580 88080 585140 88108
rect 579580 88068 579586 88080
rect 585134 88068 585140 88080
rect 585192 88068 585198 88120
rect 648430 86980 648436 87032
rect 648488 87020 648494 87032
rect 662506 87020 662512 87032
rect 648488 86992 662512 87020
rect 648488 86980 648494 86992
rect 662506 86980 662512 86992
rect 662564 86980 662570 87032
rect 656710 86844 656716 86896
rect 656768 86884 656774 86896
rect 659562 86884 659568 86896
rect 656768 86856 659568 86884
rect 656768 86844 656774 86856
rect 659562 86844 659568 86856
rect 659620 86844 659626 86896
rect 649258 86708 649264 86760
rect 649316 86748 649322 86760
rect 661402 86748 661408 86760
rect 649316 86720 661408 86748
rect 649316 86708 649322 86720
rect 661402 86708 661408 86720
rect 661460 86708 661466 86760
rect 647878 86572 647884 86624
rect 647936 86612 647942 86624
rect 660114 86612 660120 86624
rect 647936 86584 660120 86612
rect 647936 86572 647942 86584
rect 660114 86572 660120 86584
rect 660172 86572 660178 86624
rect 656158 86436 656164 86488
rect 656216 86476 656222 86488
rect 660666 86476 660672 86488
rect 656216 86448 660672 86476
rect 656216 86436 656222 86448
rect 660666 86436 660672 86448
rect 660724 86436 660730 86488
rect 619266 86300 619272 86352
rect 619324 86340 619330 86352
rect 625154 86340 625160 86352
rect 619324 86312 625160 86340
rect 619324 86300 619330 86312
rect 625154 86300 625160 86312
rect 625212 86300 625218 86352
rect 652018 86300 652024 86352
rect 652076 86340 652082 86352
rect 657170 86340 657176 86352
rect 652076 86312 657176 86340
rect 652076 86300 652082 86312
rect 657170 86300 657176 86312
rect 657228 86300 657234 86352
rect 620278 85484 620284 85536
rect 620336 85524 620342 85536
rect 625338 85524 625344 85536
rect 620336 85496 625344 85524
rect 620336 85484 620342 85496
rect 625338 85484 625344 85496
rect 625396 85484 625402 85536
rect 609882 85348 609888 85400
rect 609940 85388 609946 85400
rect 609940 85360 621014 85388
rect 609940 85348 609946 85360
rect 620986 85320 621014 85360
rect 625154 85320 625160 85332
rect 620986 85292 625160 85320
rect 625154 85280 625160 85292
rect 625212 85280 625218 85332
rect 579154 84124 579160 84176
rect 579212 84164 579218 84176
rect 581638 84164 581644 84176
rect 579212 84136 581644 84164
rect 579212 84124 579218 84136
rect 581638 84124 581644 84136
rect 581696 84124 581702 84176
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 625154 84164 625160 84176
rect 608560 84136 625160 84164
rect 608560 84124 608566 84136
rect 625154 84124 625160 84136
rect 625212 84124 625218 84176
rect 579062 82356 579068 82408
rect 579120 82396 579126 82408
rect 583018 82396 583024 82408
rect 579120 82368 583024 82396
rect 579120 82356 579126 82368
rect 583018 82356 583024 82368
rect 583076 82356 583082 82408
rect 579522 82084 579528 82136
rect 579580 82124 579586 82136
rect 587158 82124 587164 82136
rect 579580 82096 587164 82124
rect 579580 82084 579586 82096
rect 587158 82084 587164 82096
rect 587216 82084 587222 82136
rect 628742 80928 628748 80980
rect 628800 80968 628806 80980
rect 642450 80968 642456 80980
rect 628800 80940 642456 80968
rect 628800 80928 628806 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 612642 80792 612648 80844
rect 612700 80832 612706 80844
rect 647418 80832 647424 80844
rect 612700 80804 647424 80832
rect 612700 80792 612706 80804
rect 647418 80792 647424 80804
rect 647476 80792 647482 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636746 80696 636752 80708
rect 595496 80668 636752 80696
rect 595496 80656 595502 80668
rect 636746 80656 636752 80668
rect 636804 80656 636810 80708
rect 629202 79976 629208 80028
rect 629260 80016 629266 80028
rect 633434 80016 633440 80028
rect 629260 79988 633440 80016
rect 629260 79976 629266 79988
rect 633434 79976 633440 79988
rect 633492 79976 633498 80028
rect 613838 79432 613844 79484
rect 613896 79472 613902 79484
rect 645946 79472 645952 79484
rect 613896 79444 645952 79472
rect 613896 79432 613902 79444
rect 645946 79432 645952 79444
rect 646004 79432 646010 79484
rect 579062 79296 579068 79348
rect 579120 79336 579126 79348
rect 588722 79336 588728 79348
rect 579120 79308 588728 79336
rect 579120 79296 579126 79308
rect 588722 79296 588728 79308
rect 588780 79296 588786 79348
rect 614022 79296 614028 79348
rect 614080 79336 614086 79348
rect 646498 79336 646504 79348
rect 614080 79308 646504 79336
rect 614080 79296 614086 79308
rect 646498 79296 646504 79308
rect 646556 79296 646562 79348
rect 633434 78072 633440 78124
rect 633492 78112 633498 78124
rect 645302 78112 645308 78124
rect 633492 78084 645308 78112
rect 633492 78072 633498 78084
rect 645302 78072 645308 78084
rect 645360 78072 645366 78124
rect 631042 77936 631048 77988
rect 631100 77976 631106 77988
rect 643094 77976 643100 77988
rect 631100 77948 643100 77976
rect 631100 77936 631106 77948
rect 643094 77936 643100 77948
rect 643152 77936 643158 77988
rect 628466 77732 628472 77784
rect 628524 77772 628530 77784
rect 632790 77772 632796 77784
rect 628524 77744 632796 77772
rect 628524 77732 628530 77744
rect 632790 77732 632796 77744
rect 632848 77732 632854 77784
rect 625798 77256 625804 77308
rect 625856 77296 625862 77308
rect 631042 77296 631048 77308
rect 625856 77268 631048 77296
rect 625856 77256 625862 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 616782 76644 616788 76696
rect 616840 76684 616846 76696
rect 646314 76684 646320 76696
rect 616840 76656 646320 76684
rect 616840 76644 616846 76656
rect 646314 76644 646320 76656
rect 646372 76644 646378 76696
rect 611998 76508 612004 76560
rect 612056 76548 612062 76560
rect 662414 76548 662420 76560
rect 612056 76520 662420 76548
rect 612056 76508 612062 76520
rect 662414 76508 662420 76520
rect 662472 76508 662478 76560
rect 578234 75828 578240 75880
rect 578292 75868 578298 75880
rect 580258 75868 580264 75880
rect 578292 75840 580264 75868
rect 578292 75828 578298 75840
rect 580258 75828 580264 75840
rect 580316 75828 580322 75880
rect 618898 75420 618904 75472
rect 618956 75460 618962 75472
rect 648614 75460 648620 75472
rect 618956 75432 648620 75460
rect 618956 75420 618962 75432
rect 648614 75420 648620 75432
rect 648672 75420 648678 75472
rect 615402 75284 615408 75336
rect 615460 75324 615466 75336
rect 646866 75324 646872 75336
rect 615460 75296 646872 75324
rect 615460 75284 615466 75296
rect 646866 75284 646872 75296
rect 646924 75284 646930 75336
rect 607122 75148 607128 75200
rect 607180 75188 607186 75200
rect 646130 75188 646136 75200
rect 607180 75160 646136 75188
rect 607180 75148 607186 75160
rect 646130 75148 646136 75160
rect 646188 75148 646194 75200
rect 578878 72428 578884 72480
rect 578936 72468 578942 72480
rect 601694 72468 601700 72480
rect 578936 72440 601700 72468
rect 578936 72428 578942 72440
rect 601694 72428 601700 72440
rect 601752 72428 601758 72480
rect 579062 71340 579068 71392
rect 579120 71380 579126 71392
rect 584398 71380 584404 71392
rect 579120 71352 584404 71380
rect 579120 71340 579126 71352
rect 584398 71340 584404 71352
rect 584456 71340 584462 71392
rect 580258 68280 580264 68332
rect 580316 68320 580322 68332
rect 604454 68320 604460 68332
rect 580316 68292 604460 68320
rect 580316 68280 580322 68292
rect 604454 68280 604460 68292
rect 604512 68280 604518 68332
rect 577498 59984 577504 60036
rect 577556 60024 577562 60036
rect 603074 60024 603080 60036
rect 577556 59996 603080 60024
rect 577556 59984 577562 59996
rect 603074 59984 603080 59996
rect 603132 59984 603138 60036
rect 576118 58624 576124 58676
rect 576176 58664 576182 58676
rect 601878 58664 601884 58676
rect 576176 58636 601884 58664
rect 576176 58624 576182 58636
rect 601878 58624 601884 58636
rect 601936 58624 601942 58676
rect 574922 57196 574928 57248
rect 574980 57236 574986 57248
rect 600314 57236 600320 57248
rect 574980 57208 600320 57236
rect 574980 57196 574986 57208
rect 600314 57196 600320 57208
rect 600372 57196 600378 57248
rect 574738 55972 574744 56024
rect 574796 56012 574802 56024
rect 598934 56012 598940 56024
rect 574796 55984 598940 56012
rect 574796 55972 574802 55984
rect 598934 55972 598940 55984
rect 598992 55972 598998 56024
rect 574554 55836 574560 55888
rect 574612 55876 574618 55888
rect 600498 55876 600504 55888
rect 574612 55848 600504 55876
rect 574612 55836 574618 55848
rect 600498 55836 600504 55848
rect 600556 55836 600562 55888
rect 464218 55372 467788 55400
rect 464218 53644 464246 55372
rect 467760 55332 467788 55372
rect 467760 55304 477494 55332
rect 477466 55196 477494 55304
rect 596450 55196 596456 55208
rect 464356 55168 471836 55196
rect 477466 55168 596456 55196
rect 464356 53644 464384 55168
rect 471808 55128 471836 55168
rect 596450 55156 596456 55168
rect 596508 55156 596514 55208
rect 471808 55100 472112 55128
rect 472084 55060 472112 55100
rect 597830 55060 597836 55072
rect 472084 55032 597836 55060
rect 597830 55020 597836 55032
rect 597888 55020 597894 55072
rect 467806 54964 471560 54992
rect 467806 54788 467834 54964
rect 471532 54924 471560 54964
rect 597646 54924 597652 54936
rect 471532 54896 471928 54924
rect 471900 54856 471928 54896
rect 471992 54896 597652 54924
rect 471992 54856 472020 54896
rect 597646 54884 597652 54896
rect 597704 54884 597710 54936
rect 471900 54828 472020 54856
rect 599118 54788 599124 54800
rect 464724 54760 467834 54788
rect 471164 54760 471836 54788
rect 464154 53592 464160 53644
rect 464212 53604 464246 53644
rect 464212 53592 464218 53604
rect 464338 53592 464344 53644
rect 464396 53592 464402 53644
rect 464522 53592 464528 53644
rect 464580 53632 464586 53644
rect 464724 53632 464752 54760
rect 471164 54584 471192 54760
rect 471808 54720 471836 54760
rect 472084 54760 599124 54788
rect 472084 54720 472112 54760
rect 599118 54748 599124 54760
rect 599176 54748 599182 54800
rect 471808 54692 472112 54720
rect 624418 54652 624424 54664
rect 472176 54624 624424 54652
rect 472176 54584 472204 54624
rect 624418 54612 624424 54624
rect 624476 54612 624482 54664
rect 465920 54556 471192 54584
rect 471256 54556 472204 54584
rect 465920 54040 465948 54556
rect 471256 54448 471284 54556
rect 625798 54516 625804 54528
rect 464908 54012 465948 54040
rect 466380 54420 471284 54448
rect 472360 54488 625804 54516
rect 464908 53644 464936 54012
rect 466380 53904 466408 54420
rect 472360 54244 472388 54488
rect 625798 54476 625804 54488
rect 625856 54476 625862 54528
rect 596174 54380 596180 54392
rect 472176 54216 472388 54244
rect 472728 54352 596180 54380
rect 472176 54040 472204 54216
rect 471946 54012 472204 54040
rect 471946 53904 471974 54012
rect 472728 53904 472756 54352
rect 596174 54340 596180 54352
rect 596232 54340 596238 54392
rect 581638 54244 581644 54256
rect 465920 53876 466408 53904
rect 467806 53876 471974 53904
rect 472360 53876 472756 53904
rect 473096 54216 581644 54244
rect 465920 53644 465948 53876
rect 467806 53768 467834 53876
rect 466104 53740 467834 53768
rect 472084 53834 472204 53836
rect 472360 53834 472388 53876
rect 472084 53808 472388 53834
rect 466104 53644 466132 53740
rect 472084 53700 472112 53808
rect 472176 53806 472388 53808
rect 473096 53700 473124 54216
rect 581638 54204 581644 54216
rect 581696 54204 581702 54256
rect 574738 54108 574744 54120
rect 471992 53672 472112 53700
rect 472820 53672 473124 53700
rect 473188 54080 574744 54108
rect 464580 53604 464752 53632
rect 464580 53592 464586 53604
rect 464890 53592 464896 53644
rect 464948 53592 464954 53644
rect 465902 53592 465908 53644
rect 465960 53592 465966 53644
rect 466086 53592 466092 53644
rect 466144 53592 466150 53644
rect 471992 53576 472020 53672
rect 472820 53576 472848 53672
rect 471974 53524 471980 53576
rect 472032 53524 472038 53576
rect 472802 53524 472808 53576
rect 472860 53524 472866 53576
rect 462222 53456 462228 53508
rect 462280 53496 462286 53508
rect 471790 53496 471796 53508
rect 462280 53468 471796 53496
rect 462280 53456 462286 53468
rect 471790 53456 471796 53468
rect 471848 53456 471854 53508
rect 461302 53320 461308 53372
rect 461360 53360 461366 53372
rect 473188 53360 473216 54080
rect 574738 54068 574744 54080
rect 574796 54068 574802 54120
rect 574554 53972 574560 53984
rect 473556 53944 574560 53972
rect 473556 53508 473584 53944
rect 574554 53932 574560 53944
rect 574612 53932 574618 53984
rect 574922 53836 574928 53848
rect 477466 53808 574928 53836
rect 473722 53592 473728 53644
rect 473780 53632 473786 53644
rect 477466 53632 477494 53808
rect 574922 53796 574928 53808
rect 574980 53796 574986 53848
rect 473780 53604 477494 53632
rect 473780 53592 473786 53604
rect 473538 53456 473544 53508
rect 473596 53456 473602 53508
rect 461360 53332 473216 53360
rect 461360 53320 461366 53332
rect 49142 53184 49148 53236
rect 49200 53224 49206 53236
rect 128998 53224 129004 53236
rect 49200 53196 129004 53224
rect 49200 53184 49206 53196
rect 128998 53184 129004 53196
rect 129056 53184 129062 53236
rect 464062 53184 464068 53236
rect 464120 53224 464126 53236
rect 471974 53224 471980 53236
rect 464120 53196 471980 53224
rect 464120 53184 464126 53196
rect 471974 53184 471980 53196
rect 472032 53184 472038 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 48958 53048 48964 53100
rect 49016 53088 49022 53100
rect 130378 53088 130384 53100
rect 49016 53060 130384 53088
rect 49016 53048 49022 53060
rect 130378 53048 130384 53060
rect 130436 53048 130442 53100
rect 459462 53048 459468 53100
rect 459520 53088 459526 53100
rect 464890 53088 464896 53100
rect 459520 53060 464896 53088
rect 459520 53048 459526 53060
rect 464890 53048 464896 53060
rect 464948 53048 464954 53100
rect 463142 52912 463148 52964
rect 463200 52952 463206 52964
rect 473722 52952 473728 52964
rect 463200 52924 473728 52952
rect 463200 52912 463206 52924
rect 473722 52912 473728 52924
rect 473780 52912 473786 52964
rect 460060 52776 460066 52828
rect 460118 52816 460124 52828
rect 466086 52816 466092 52828
rect 460118 52788 466092 52816
rect 460118 52776 460124 52788
rect 466086 52776 466092 52788
rect 466144 52776 466150 52828
rect 463602 52640 463608 52692
rect 463660 52680 463666 52692
rect 464522 52680 464528 52692
rect 463660 52652 464528 52680
rect 463660 52640 463666 52652
rect 464522 52640 464528 52652
rect 464580 52640 464586 52692
rect 465442 52640 465448 52692
rect 465500 52680 465506 52692
rect 472802 52680 472808 52692
rect 465500 52652 472808 52680
rect 465500 52640 465506 52652
rect 472802 52640 472808 52652
rect 472860 52640 472866 52692
rect 47578 51960 47584 52012
rect 47636 52000 47642 52012
rect 130562 52000 130568 52012
rect 47636 51972 130568 52000
rect 47636 51960 47642 51972
rect 130562 51960 130568 51972
rect 130620 51960 130626 52012
rect 50338 51824 50344 51876
rect 50396 51864 50402 51876
rect 129182 51864 129188 51876
rect 50396 51836 129188 51864
rect 50396 51824 50402 51836
rect 129182 51824 129188 51836
rect 129240 51824 129246 51876
rect 129550 51824 129556 51876
rect 129608 51864 129614 51876
rect 591298 51864 591304 51876
rect 129608 51836 591304 51864
rect 129608 51824 129614 51836
rect 591298 51824 591304 51836
rect 591356 51824 591362 51876
rect 128814 51688 128820 51740
rect 128872 51728 128878 51740
rect 592678 51728 592684 51740
rect 128872 51700 592684 51728
rect 128872 51688 128878 51700
rect 592678 51688 592684 51700
rect 592736 51688 592742 51740
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458174 50504 458180 50516
rect 318392 50476 458180 50504
rect 318392 50464 318398 50476
rect 458174 50464 458180 50476
rect 458232 50464 458238 50516
rect 47762 50328 47768 50380
rect 47820 50368 47826 50380
rect 130746 50368 130752 50380
rect 47820 50340 130752 50368
rect 47820 50328 47826 50340
rect 130746 50328 130752 50340
rect 130804 50328 130810 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458358 50368 458364 50380
rect 314068 50340 458364 50368
rect 314068 50328 314074 50340
rect 458358 50328 458364 50340
rect 458416 50328 458422 50380
rect 522942 50328 522948 50380
rect 523000 50368 523006 50380
rect 544010 50368 544016 50380
rect 523000 50340 544016 50368
rect 523000 50328 523006 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 50522 49104 50528 49156
rect 50580 49144 50586 49156
rect 129366 49144 129372 49156
rect 50580 49116 129372 49144
rect 50580 49104 50586 49116
rect 129366 49104 129372 49116
rect 129424 49104 129430 49156
rect 46198 48968 46204 49020
rect 46256 49008 46262 49020
rect 130930 49008 130936 49020
rect 46256 48980 130936 49008
rect 46256 48968 46262 48980
rect 130930 48968 130936 48980
rect 130988 48968 130994 49020
rect 130562 45500 130568 45552
rect 130620 45540 130626 45552
rect 132586 45540 132592 45552
rect 130620 45512 132592 45540
rect 130620 45500 130626 45512
rect 132586 45500 132592 45512
rect 132644 45500 132650 45552
rect 128998 45296 129004 45348
rect 129056 45336 129062 45348
rect 129056 45308 131206 45336
rect 129056 45296 129062 45308
rect 131178 45090 131206 45308
rect 131390 45160 131396 45212
rect 131448 45200 131454 45212
rect 133138 45200 133144 45212
rect 131448 45172 133144 45200
rect 131448 45160 131454 45172
rect 133138 45160 133144 45172
rect 133196 45160 133202 45212
rect 129550 45024 129556 45076
rect 129608 45064 129614 45076
rect 129608 45036 131068 45064
rect 129608 45024 129614 45036
rect 131040 45020 131068 45036
rect 131040 44992 131330 45020
rect 129366 44888 129372 44940
rect 129424 44928 129430 44940
rect 129424 44900 131620 44928
rect 129424 44888 129430 44900
rect 131684 44824 131790 44852
rect 128814 44752 128820 44804
rect 128872 44792 128878 44804
rect 131684 44792 131712 44824
rect 128872 44764 131712 44792
rect 128872 44752 128878 44764
rect 131868 44740 131974 44768
rect 131574 44616 131580 44668
rect 131632 44656 131638 44668
rect 131868 44656 131896 44740
rect 131632 44628 131896 44656
rect 131632 44616 131638 44628
rect 129182 44480 129188 44532
rect 129240 44520 129246 44532
rect 132144 44520 132172 44670
rect 129240 44516 131390 44520
rect 131500 44516 132172 44520
rect 129240 44492 132172 44516
rect 132236 44572 132388 44600
rect 129240 44480 129246 44492
rect 131362 44488 131528 44492
rect 43622 44276 43628 44328
rect 43680 44316 43686 44328
rect 132236 44316 132264 44572
rect 132466 44488 132526 44516
rect 132466 44328 132494 44488
rect 132586 44364 132592 44416
rect 132644 44404 132650 44416
rect 132644 44376 132756 44404
rect 132644 44364 132650 44376
rect 43680 44288 132264 44316
rect 43680 44276 43686 44288
rect 132402 44276 132408 44328
rect 132460 44288 132494 44328
rect 132460 44276 132466 44288
rect 43438 44140 43444 44192
rect 43496 44180 43502 44192
rect 131574 44180 131580 44192
rect 43496 44152 131580 44180
rect 43496 44140 43502 44152
rect 131574 44140 131580 44152
rect 131632 44140 131638 44192
rect 132972 44180 133000 44278
rect 131776 44152 133000 44180
rect 130746 44004 130752 44056
rect 130804 44044 130810 44056
rect 131776 44044 131804 44152
rect 133138 44140 133144 44192
rect 133196 44140 133202 44192
rect 130804 44016 131804 44044
rect 130804 44004 130810 44016
rect 440234 43800 440240 43852
rect 440292 43840 440298 43852
rect 441062 43840 441068 43852
rect 440292 43812 441068 43840
rect 440292 43800 440298 43812
rect 441062 43800 441068 43812
rect 441120 43800 441126 43852
rect 187326 42780 187332 42832
rect 187384 42820 187390 42832
rect 255866 42820 255872 42832
rect 187384 42792 255872 42820
rect 187384 42780 187390 42792
rect 255866 42780 255872 42792
rect 255924 42780 255930 42832
rect 307294 42712 307300 42764
rect 307352 42752 307358 42764
rect 431218 42752 431224 42764
rect 307352 42724 431224 42752
rect 307352 42712 307358 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 441062 42712 441068 42764
rect 441120 42752 441126 42764
rect 449158 42752 449164 42764
rect 441120 42724 449164 42752
rect 441120 42712 441126 42724
rect 449158 42712 449164 42724
rect 449216 42712 449222 42764
rect 453574 42712 453580 42764
rect 453632 42752 453638 42764
rect 464154 42752 464160 42764
rect 453632 42724 464160 42752
rect 453632 42712 453638 42724
rect 464154 42712 464160 42724
rect 464212 42712 464218 42764
rect 310422 42576 310428 42628
rect 310480 42616 310486 42628
rect 427078 42616 427084 42628
rect 310480 42588 427084 42616
rect 310480 42576 310486 42588
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 441246 42576 441252 42628
rect 441304 42616 441310 42628
rect 446398 42616 446404 42628
rect 441304 42588 446404 42616
rect 441304 42576 441310 42588
rect 446398 42576 446404 42588
rect 446456 42576 446462 42628
rect 454494 42440 454500 42492
rect 454552 42480 454558 42492
rect 463050 42480 463056 42492
rect 454552 42452 463056 42480
rect 454552 42440 454558 42452
rect 463050 42440 463056 42452
rect 463108 42440 463114 42492
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405182 42344 405188 42356
rect 404504 42316 405188 42344
rect 404504 42304 404510 42316
rect 405182 42304 405188 42316
rect 405240 42304 405246 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 426894 42344 426900 42356
rect 420788 42316 426900 42344
rect 420788 42304 420794 42316
rect 426894 42304 426900 42316
rect 426952 42304 426958 42356
rect 661402 42129 661408 42181
rect 661460 42129 661466 42181
rect 427078 41964 427084 42016
rect 427136 42004 427142 42016
rect 427136 41976 427814 42004
rect 427136 41964 427142 41976
rect 427786 41868 427814 41976
rect 431218 41964 431224 42016
rect 431276 42004 431282 42016
rect 441062 42004 441068 42016
rect 431276 41976 441068 42004
rect 431276 41964 431282 41976
rect 441062 41964 441068 41976
rect 441120 41964 441126 42016
rect 446398 41964 446404 42016
rect 446456 42004 446462 42016
rect 454494 42004 454500 42016
rect 446456 41976 454500 42004
rect 446456 41964 446462 41976
rect 454494 41964 454500 41976
rect 454552 41964 454558 42016
rect 441246 41868 441252 41880
rect 427786 41840 441252 41868
rect 441246 41828 441252 41840
rect 441304 41828 441310 41880
rect 449158 41828 449164 41880
rect 449216 41868 449222 41880
rect 453574 41868 453580 41880
rect 449216 41840 453580 41868
rect 449216 41828 449222 41840
rect 453574 41828 453580 41840
rect 453632 41828 453638 41880
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 426894 41420 426900 41472
rect 426952 41460 426958 41472
rect 459186 41460 459192 41472
rect 426952 41432 459192 41460
rect 426952 41420 426958 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 132500 1001920 132552 1001972
rect 133696 1001920 133748 1001972
rect 401692 992196 401744 992248
rect 404360 992196 404412 992248
rect 396080 990836 396132 990888
rect 400220 990836 400272 990888
rect 242256 989068 242308 989120
rect 245660 989068 245712 989120
rect 293960 988184 294012 988236
rect 298100 988184 298152 988236
rect 389180 987504 389232 987556
rect 391940 987504 391992 987556
rect 399760 986348 399812 986400
rect 401692 986348 401744 986400
rect 238668 985940 238720 985992
rect 242256 985940 242308 985992
rect 289728 985396 289780 985448
rect 293960 985396 294012 985448
rect 394424 983492 394476 983544
rect 396080 983492 396132 983544
rect 483020 982472 483072 982524
rect 483848 982472 483900 982524
rect 651380 959080 651432 959132
rect 677416 959080 677468 959132
rect 30104 954932 30156 954984
rect 63408 954932 63460 954984
rect 652024 896996 652076 897048
rect 676036 897064 676088 897116
rect 654784 895772 654836 895824
rect 675852 895772 675904 895824
rect 672724 895636 672776 895688
rect 676036 895636 676088 895688
rect 671068 894412 671120 894464
rect 675852 894412 675904 894464
rect 671896 894276 671948 894328
rect 676036 894276 676088 894328
rect 672540 892984 672592 893036
rect 675852 892984 675904 893036
rect 672080 892848 672132 892900
rect 676036 892848 676088 892900
rect 674840 890332 674892 890384
rect 676036 890332 676088 890384
rect 676220 890128 676272 890180
rect 676864 890128 676916 890180
rect 674380 888904 674432 888956
rect 676036 888904 676088 888956
rect 676220 888700 676272 888752
rect 677048 888700 677100 888752
rect 674656 888496 674708 888548
rect 676036 888496 676088 888548
rect 674196 887272 674248 887324
rect 676036 887272 676088 887324
rect 670884 886864 670936 886916
rect 676036 886864 676088 886916
rect 675852 886660 675904 886712
rect 676404 886660 676456 886712
rect 673092 885640 673144 885692
rect 676036 885640 676088 885692
rect 653404 880472 653456 880524
rect 675484 880472 675536 880524
rect 676036 880200 676088 880252
rect 679624 880200 679676 880252
rect 675024 879588 675076 879640
rect 677048 879588 677100 879640
rect 675116 879384 675168 879436
rect 676864 879384 676916 879436
rect 675668 879248 675720 879300
rect 678244 879248 678296 879300
rect 675852 878432 675904 878484
rect 676036 878432 676088 878484
rect 675484 877752 675536 877804
rect 675392 876732 675444 876784
rect 657544 869388 657596 869440
rect 675024 869388 675076 869440
rect 674840 869252 674892 869304
rect 675300 869252 675352 869304
rect 651472 868844 651524 868896
rect 654784 868844 654836 868896
rect 674196 868708 674248 868760
rect 675300 868708 675352 868760
rect 654140 868028 654192 868080
rect 675024 868028 675076 868080
rect 674840 867552 674892 867604
rect 675208 867552 675260 867604
rect 651472 866600 651524 866652
rect 672724 866600 672776 866652
rect 651380 865172 651432 865224
rect 653404 865172 653456 865224
rect 651472 863812 651524 863864
rect 657544 863812 657596 863864
rect 651472 862452 651524 862504
rect 654140 862452 654192 862504
rect 35808 817096 35860 817148
rect 46204 817096 46256 817148
rect 35624 816960 35676 817012
rect 60004 816960 60056 817012
rect 35808 815736 35860 815788
rect 42892 815736 42944 815788
rect 35440 815600 35492 815652
rect 44180 815600 44232 815652
rect 35624 814376 35676 814428
rect 43444 814376 43496 814428
rect 35808 814240 35860 814292
rect 45284 814240 45336 814292
rect 41328 812812 41380 812864
rect 44548 812812 44600 812864
rect 41328 811452 41380 811504
rect 43076 811452 43128 811504
rect 40960 810704 41012 810756
rect 42708 810704 42760 810756
rect 44180 810704 44232 810756
rect 62948 810704 63000 810756
rect 41328 808596 41380 808648
rect 42248 808596 42300 808648
rect 41328 807440 41380 807492
rect 43260 807440 43312 807492
rect 41144 807304 41196 807356
rect 44364 807304 44416 807356
rect 41328 806080 41380 806132
rect 50344 806080 50396 806132
rect 41144 805944 41196 805996
rect 62672 805944 62724 805996
rect 34520 802408 34572 802460
rect 41880 802408 41932 802460
rect 37924 801728 37976 801780
rect 39764 801728 39816 801780
rect 31024 801048 31076 801100
rect 42524 801048 42576 801100
rect 36544 800708 36596 800760
rect 40500 800708 40552 800760
rect 42248 799280 42300 799332
rect 42708 799280 42760 799332
rect 43628 799008 43680 799060
rect 53104 799008 53156 799060
rect 43812 797648 43864 797700
rect 57244 797648 57296 797700
rect 42248 795608 42300 795660
rect 43812 795608 43864 795660
rect 42340 793908 42392 793960
rect 44364 793908 44416 793960
rect 653404 790780 653456 790832
rect 675392 790780 675444 790832
rect 53104 790712 53156 790764
rect 62212 790712 62264 790764
rect 42616 789284 42668 789336
rect 43076 789284 43128 789336
rect 57244 789148 57296 789200
rect 62120 789148 62172 789200
rect 42708 786632 42760 786684
rect 62120 786632 62172 786684
rect 60004 786496 60056 786548
rect 62304 786496 62356 786548
rect 46204 785136 46256 785188
rect 62120 785136 62172 785188
rect 670608 784252 670660 784304
rect 675116 784252 675168 784304
rect 669228 784116 669280 784168
rect 675392 784116 675444 784168
rect 673736 782620 673788 782672
rect 675116 782620 675168 782672
rect 669044 782484 669096 782536
rect 675300 782484 675352 782536
rect 655520 781056 655572 781108
rect 675024 781056 675076 781108
rect 673920 779968 673972 780020
rect 675116 779968 675168 780020
rect 655060 778336 655112 778388
rect 674932 778336 674984 778388
rect 651472 777588 651524 777640
rect 660304 777588 660356 777640
rect 670424 776976 670476 777028
rect 675300 776976 675352 777028
rect 672724 775616 672776 775668
rect 674932 775616 674984 775668
rect 651472 775548 651524 775600
rect 669964 775548 670016 775600
rect 651380 775276 651432 775328
rect 653404 775276 653456 775328
rect 35808 774188 35860 774240
rect 41696 774188 41748 774240
rect 42064 774188 42116 774240
rect 58624 774188 58676 774240
rect 651472 774120 651524 774172
rect 655520 774120 655572 774172
rect 651472 773780 651524 773832
rect 655060 773780 655112 773832
rect 35440 773372 35492 773424
rect 41512 773372 41564 773424
rect 671436 773372 671488 773424
rect 675300 773372 675352 773424
rect 35808 773100 35860 773152
rect 41696 773168 41748 773220
rect 42064 773168 42116 773220
rect 42892 773168 42944 773220
rect 35624 772964 35676 773016
rect 41696 773032 41748 773084
rect 42064 773032 42116 773084
rect 46204 773032 46256 773084
rect 35256 772828 35308 772880
rect 41696 772828 41748 772880
rect 42064 772828 42116 772880
rect 61384 772828 61436 772880
rect 35808 771808 35860 771860
rect 39948 771808 40000 771860
rect 35624 771536 35676 771588
rect 40316 771604 40368 771656
rect 42064 771468 42116 771520
rect 45284 771468 45336 771520
rect 35808 771400 35860 771452
rect 41696 771400 41748 771452
rect 35808 770448 35860 770500
rect 40316 770448 40368 770500
rect 35440 770176 35492 770228
rect 41696 770244 41748 770296
rect 42064 770244 42116 770296
rect 43076 770244 43128 770296
rect 42064 770108 42116 770160
rect 44548 770108 44600 770160
rect 35624 770040 35676 770092
rect 41696 770040 41748 770092
rect 35808 768816 35860 768868
rect 40040 768816 40092 768868
rect 35624 768680 35676 768732
rect 41696 768680 41748 768732
rect 35808 767592 35860 767644
rect 36544 767592 36596 767644
rect 35808 766028 35860 766080
rect 39396 766028 39448 766080
rect 40040 765280 40092 765332
rect 41696 765280 41748 765332
rect 42064 765144 42116 765196
rect 42432 765144 42484 765196
rect 35808 764804 35860 764856
rect 39948 764804 40000 764856
rect 35624 764532 35676 764584
rect 41696 764600 41748 764652
rect 42064 764600 42116 764652
rect 43444 764600 43496 764652
rect 35624 763444 35676 763496
rect 39948 763444 40000 763496
rect 42064 763376 42116 763428
rect 35808 763172 35860 763224
rect 41696 763104 41748 763156
rect 60004 763172 60056 763224
rect 42064 761880 42116 761932
rect 48964 761880 49016 761932
rect 35808 761812 35860 761864
rect 41696 761812 41748 761864
rect 35164 759772 35216 759824
rect 39672 759772 39724 759824
rect 32404 759636 32456 759688
rect 41604 759636 41656 759688
rect 33784 758276 33836 758328
rect 39948 758276 40000 758328
rect 43904 755488 43956 755540
rect 62948 755488 63000 755540
rect 42616 753720 42668 753772
rect 42616 753584 42668 753636
rect 42248 749708 42300 749760
rect 42248 749164 42300 749216
rect 61384 747260 61436 747312
rect 63040 747260 63092 747312
rect 653404 746580 653456 746632
rect 675392 746580 675444 746632
rect 45284 746512 45336 746564
rect 62120 746512 62172 746564
rect 42248 745288 42300 745340
rect 42248 745084 42300 745136
rect 42800 743996 42852 744048
rect 62120 743860 62172 743912
rect 46204 743724 46256 743776
rect 62120 743724 62172 743776
rect 671804 742432 671856 742484
rect 675392 742432 675444 742484
rect 58624 742364 58676 742416
rect 62120 742364 62172 742416
rect 671620 741140 671672 741192
rect 675208 741140 675260 741192
rect 672264 739100 672316 739152
rect 675392 739100 675444 739152
rect 673552 738692 673604 738744
rect 675392 738692 675444 738744
rect 674840 738556 674892 738608
rect 675208 738556 675260 738608
rect 652024 736856 652076 736908
rect 656164 736856 656216 736908
rect 657544 735564 657596 735616
rect 675116 735972 675168 736024
rect 674012 735088 674064 735140
rect 675300 735088 675352 735140
rect 654784 734136 654836 734188
rect 675116 734544 675168 734596
rect 651472 733388 651524 733440
rect 668584 733388 668636 733440
rect 672908 732708 672960 732760
rect 675300 732708 675352 732760
rect 651472 731416 651524 731468
rect 658924 731416 658976 731468
rect 35808 731144 35860 731196
rect 41696 731076 41748 731128
rect 651380 731076 651432 731128
rect 653404 731076 653456 731128
rect 652668 730668 652720 730720
rect 661684 730668 661736 730720
rect 35808 730328 35860 730380
rect 40408 730328 40460 730380
rect 35440 730056 35492 730108
rect 41696 730056 41748 730108
rect 42064 730056 42116 730108
rect 61384 730056 61436 730108
rect 651472 729988 651524 730040
rect 657544 729988 657596 730040
rect 35624 729444 35676 729496
rect 42064 729308 42116 729360
rect 62948 729308 63000 729360
rect 41696 729240 41748 729292
rect 675300 729240 675352 729292
rect 35808 729036 35860 729088
rect 41512 729036 41564 729088
rect 675300 729036 675352 729088
rect 42064 728832 42116 728884
rect 44272 728832 44324 728884
rect 35624 728764 35676 728816
rect 41696 728764 41748 728816
rect 35440 728628 35492 728680
rect 41696 728628 41748 728680
rect 42064 728628 42116 728680
rect 44548 728628 44600 728680
rect 651472 728492 651524 728544
rect 654784 728492 654836 728544
rect 673092 728288 673144 728340
rect 670884 728084 670936 728136
rect 35808 727812 35860 727864
rect 40040 727812 40092 727864
rect 35440 727540 35492 727592
rect 41696 727608 41748 727660
rect 35808 727404 35860 727456
rect 41696 727404 41748 727456
rect 42064 727404 42116 727456
rect 43444 727404 43496 727456
rect 35624 727268 35676 727320
rect 41696 727268 41748 727320
rect 42064 727268 42116 727320
rect 43628 727268 43680 727320
rect 674840 727200 674892 727252
rect 681004 727200 681056 727252
rect 674564 726724 674616 726776
rect 683396 726724 683448 726776
rect 674380 726588 674432 726640
rect 684040 726588 684092 726640
rect 41328 726044 41380 726096
rect 41696 726044 41748 726096
rect 42064 726044 42116 726096
rect 42524 726044 42576 726096
rect 41144 725908 41196 725960
rect 41604 725908 41656 725960
rect 675300 721692 675352 721744
rect 675300 721216 675352 721268
rect 675300 720808 675352 720860
rect 675300 720468 675352 720520
rect 43628 718972 43680 719024
rect 53104 718972 53156 719024
rect 672816 717476 672868 717528
rect 673276 717476 673328 717528
rect 32404 716864 32456 716916
rect 41696 716864 41748 716916
rect 42064 716728 42116 716780
rect 42708 716728 42760 716780
rect 42064 716592 42116 716644
rect 42524 716592 42576 716644
rect 656164 716252 656216 716304
rect 673276 716252 673328 716304
rect 35164 715708 35216 715760
rect 41328 715708 41380 715760
rect 669964 715708 670016 715760
rect 673092 715708 673144 715760
rect 31668 715504 31720 715556
rect 40592 715504 40644 715556
rect 671068 715300 671120 715352
rect 673092 715300 673144 715352
rect 660304 714960 660356 715012
rect 673276 714960 673328 715012
rect 671896 714484 671948 714536
rect 673276 714484 673328 714536
rect 673276 713532 673328 713584
rect 672080 713396 672132 713448
rect 673276 713396 673328 713448
rect 672632 713260 672684 713312
rect 671068 712580 671120 712632
rect 671988 712580 672040 712632
rect 43628 712104 43680 712156
rect 51724 712104 51776 712156
rect 672448 712036 672500 712088
rect 673276 712036 673328 712088
rect 672448 711764 672500 711816
rect 673092 711764 673144 711816
rect 42248 710404 42300 710456
rect 44732 710404 44784 710456
rect 671436 709996 671488 710048
rect 673092 709996 673144 710048
rect 43628 709316 43680 709368
rect 45100 709316 45152 709368
rect 669044 709316 669096 709368
rect 673276 709316 673328 709368
rect 670608 709180 670660 709232
rect 673276 709180 673328 709232
rect 669228 708228 669280 708280
rect 673276 708228 673328 708280
rect 42248 707820 42300 707872
rect 43628 707820 43680 707872
rect 42248 707412 42300 707464
rect 42708 707412 42760 707464
rect 674656 707140 674708 707192
rect 676036 707140 676088 707192
rect 42524 706664 42576 706716
rect 42708 706460 42760 706512
rect 42248 705508 42300 705560
rect 43812 705508 43864 705560
rect 670424 705372 670476 705424
rect 673276 705372 673328 705424
rect 674288 705304 674340 705356
rect 683120 705304 683172 705356
rect 667848 705168 667900 705220
rect 673736 705236 673788 705288
rect 51724 705100 51776 705152
rect 62120 705100 62172 705152
rect 667020 703808 667072 703860
rect 673736 703808 673788 703860
rect 44732 703740 44784 703792
rect 62120 703740 62172 703792
rect 654784 701156 654836 701208
rect 673736 701156 673788 701208
rect 42708 701088 42760 701140
rect 62948 701020 63000 701072
rect 46204 698232 46256 698284
rect 62212 698232 62264 698284
rect 674288 692996 674340 693048
rect 675392 692996 675444 693048
rect 668400 692792 668452 692844
rect 673736 692792 673788 692844
rect 656440 690072 656492 690124
rect 673736 690072 673788 690124
rect 674840 688984 674892 689036
rect 675208 688984 675260 689036
rect 652760 688780 652812 688832
rect 673736 688780 673788 688832
rect 651472 688644 651524 688696
rect 657544 688644 657596 688696
rect 35808 687488 35860 687540
rect 41696 687488 41748 687540
rect 35440 687216 35492 687268
rect 651472 687216 651524 687268
rect 669964 687216 670016 687268
rect 41696 687148 41748 687200
rect 651472 687012 651524 687064
rect 654784 687012 654836 687064
rect 42064 686468 42116 686520
rect 62948 686468 63000 686520
rect 651656 686468 651708 686520
rect 667204 686468 667256 686520
rect 35624 686400 35676 686452
rect 41696 686400 41748 686452
rect 35808 686264 35860 686316
rect 41696 686264 41748 686316
rect 42064 686264 42116 686316
rect 43628 686264 43680 686316
rect 42064 686060 42116 686112
rect 44548 686060 44600 686112
rect 35440 685992 35492 686044
rect 41696 685992 41748 686044
rect 35808 685856 35860 685908
rect 41696 685856 41748 685908
rect 42064 685856 42116 685908
rect 44272 685856 44324 685908
rect 651472 685516 651524 685568
rect 656440 685516 656492 685568
rect 35808 684972 35860 685024
rect 41696 684904 41748 684956
rect 42248 684768 42300 684820
rect 45284 684768 45336 684820
rect 35624 684632 35676 684684
rect 41696 684632 41748 684684
rect 35808 684496 35860 684548
rect 41696 684496 41748 684548
rect 42064 684496 42116 684548
rect 43076 684496 43128 684548
rect 35808 683408 35860 683460
rect 41696 683408 41748 683460
rect 35624 683272 35676 683324
rect 41512 683272 41564 683324
rect 35440 683136 35492 683188
rect 41696 683068 41748 683120
rect 675484 682524 675536 682576
rect 683212 682524 683264 682576
rect 674840 682388 674892 682440
rect 683488 682388 683540 682440
rect 35624 681844 35676 681896
rect 41696 681844 41748 681896
rect 35808 681708 35860 681760
rect 41512 681708 41564 681760
rect 35808 680484 35860 680536
rect 41696 680484 41748 680536
rect 35808 679396 35860 679448
rect 41696 679396 41748 679448
rect 35808 679124 35860 679176
rect 41512 679124 41564 679176
rect 35624 678988 35676 679040
rect 41696 678988 41748 679040
rect 43996 676200 44048 676252
rect 57244 676200 57296 676252
rect 33048 674092 33100 674144
rect 41512 674092 41564 674144
rect 35164 672800 35216 672852
rect 41696 672800 41748 672852
rect 42064 672664 42116 672716
rect 42524 672664 42576 672716
rect 31024 672460 31076 672512
rect 41696 672460 41748 672512
rect 673552 671304 673604 671356
rect 668584 671100 668636 671152
rect 673552 671100 673604 671152
rect 661684 670692 661736 670744
rect 673552 670352 673604 670404
rect 670240 670216 670292 670268
rect 673552 670216 673604 670268
rect 44088 669400 44140 669452
rect 58624 669332 58676 669384
rect 658924 669332 658976 669384
rect 673552 668652 673604 668704
rect 671068 668516 671120 668568
rect 673552 668516 673604 668568
rect 671436 668176 671488 668228
rect 45652 667904 45704 667956
rect 61384 667904 61436 667956
rect 671068 667904 671120 667956
rect 673552 667904 673604 667956
rect 673552 667292 673604 667344
rect 671620 667156 671672 667208
rect 673552 667156 673604 667208
rect 42248 667020 42300 667072
rect 45652 667020 45704 667072
rect 671988 666884 672040 666936
rect 674840 666612 674892 666664
rect 676036 666612 676088 666664
rect 671896 666544 671948 666596
rect 673552 666544 673604 666596
rect 669596 665252 669648 665304
rect 673552 665252 673604 665304
rect 671712 664368 671764 664420
rect 673552 664368 673604 664420
rect 669412 663892 669464 663944
rect 673552 663892 673604 663944
rect 674840 663756 674892 663808
rect 676036 663756 676088 663808
rect 42248 663280 42300 663332
rect 42524 663076 42576 663128
rect 42248 662940 42300 662992
rect 44456 662940 44508 662992
rect 671252 661580 671304 661632
rect 674012 661580 674064 661632
rect 669228 661104 669280 661156
rect 674012 661104 674064 661156
rect 42156 661036 42208 661088
rect 43812 661036 43864 661088
rect 58624 660900 58676 660952
rect 62120 660900 62172 660952
rect 668860 660152 668912 660204
rect 674012 660152 674064 660204
rect 674840 659812 674892 659864
rect 683120 659812 683172 659864
rect 672172 659676 672224 659728
rect 674012 659676 674064 659728
rect 42524 657500 42576 657552
rect 62120 657500 62172 657552
rect 46204 656820 46256 656872
rect 62120 656820 62172 656872
rect 653404 655528 653456 655580
rect 674012 655528 674064 655580
rect 45468 655460 45520 655512
rect 62120 655460 62172 655512
rect 655520 645872 655572 645924
rect 671252 645872 671304 645924
rect 35808 644444 35860 644496
rect 41696 644444 41748 644496
rect 42064 644444 42116 644496
rect 58624 644444 58676 644496
rect 674794 643764 674846 643816
rect 35808 643492 35860 643544
rect 41144 643492 41196 643544
rect 674932 643356 674984 643408
rect 35532 643220 35584 643272
rect 41696 643288 41748 643340
rect 42064 643288 42116 643340
rect 43628 643288 43680 643340
rect 35348 643084 35400 643136
rect 41696 643084 41748 643136
rect 42064 643084 42116 643136
rect 61384 643084 61436 643136
rect 655336 643084 655388 643136
rect 671252 643084 671304 643136
rect 38568 642472 38620 642524
rect 41696 642472 41748 642524
rect 42064 642336 42116 642388
rect 62948 642336 63000 642388
rect 651472 642336 651524 642388
rect 658924 642336 658976 642388
rect 35808 642132 35860 642184
rect 39396 642132 39448 642184
rect 35440 641860 35492 641912
rect 41696 641928 41748 641980
rect 42064 641928 42116 641980
rect 43076 641928 43128 641980
rect 35624 641724 35676 641776
rect 41696 641724 41748 641776
rect 42064 641724 42116 641776
rect 45284 641724 45336 641776
rect 42064 640908 42116 640960
rect 45100 640908 45152 640960
rect 35808 640772 35860 640824
rect 40868 640568 40920 640620
rect 35624 640432 35676 640484
rect 41696 640432 41748 640484
rect 35808 640296 35860 640348
rect 41696 640296 41748 640348
rect 42064 640296 42116 640348
rect 45376 640296 45428 640348
rect 651472 640296 651524 640348
rect 668584 640296 668636 640348
rect 675208 640432 675260 640484
rect 651380 640092 651432 640144
rect 653404 640092 653456 640144
rect 675024 640092 675076 640144
rect 35808 639208 35860 639260
rect 41696 639208 41748 639260
rect 35532 639072 35584 639124
rect 39304 639072 39356 639124
rect 651656 638868 651708 638920
rect 655336 638868 655388 638920
rect 651472 638732 651524 638784
rect 655520 638732 655572 638784
rect 34428 638188 34480 638240
rect 41696 638188 41748 638240
rect 35808 637576 35860 637628
rect 36544 637576 36596 637628
rect 674472 636964 674524 637016
rect 683212 636964 683264 637016
rect 35624 636896 35676 636948
rect 40592 636896 40644 636948
rect 674288 636828 674340 636880
rect 683396 636828 683448 636880
rect 35808 636692 35860 636744
rect 40040 636556 40092 636608
rect 35808 636352 35860 636404
rect 39580 636420 39632 636472
rect 35532 636216 35584 636268
rect 39120 636148 39172 636200
rect 674932 635468 674984 635520
rect 675668 635468 675720 635520
rect 35808 634924 35860 634976
rect 40132 634924 40184 634976
rect 652024 634040 652076 634092
rect 660304 634040 660356 634092
rect 35808 633836 35860 633888
rect 40040 633700 40092 633752
rect 35808 633428 35860 633480
rect 41604 633428 41656 633480
rect 42064 633428 42116 633480
rect 60188 633428 60240 633480
rect 671528 632952 671580 633004
rect 671344 632884 671396 632936
rect 671344 632748 671396 632800
rect 671528 632612 671580 632664
rect 36544 630572 36596 630624
rect 41604 630572 41656 630624
rect 672448 629688 672500 629740
rect 673276 629688 673328 629740
rect 35164 628668 35216 628720
rect 39396 628668 39448 628720
rect 667204 626084 667256 626136
rect 673276 626084 673328 626136
rect 44180 625948 44232 626000
rect 44180 625812 44232 625864
rect 63132 625812 63184 625864
rect 669964 625404 670016 625456
rect 673276 625404 673328 625456
rect 42340 625132 42392 625184
rect 657544 625132 657596 625184
rect 673276 625132 673328 625184
rect 674288 625132 674340 625184
rect 676220 625132 676272 625184
rect 670240 624452 670292 624504
rect 672632 624452 672684 624504
rect 669412 623908 669464 623960
rect 674012 623908 674064 623960
rect 674288 623840 674340 623892
rect 676220 623840 676272 623892
rect 43996 623772 44048 623824
rect 670240 623772 670292 623824
rect 672632 623772 672684 623824
rect 671068 623228 671120 623280
rect 672632 623228 672684 623280
rect 674656 623024 674708 623076
rect 683396 623024 683448 623076
rect 42248 622820 42300 622872
rect 671896 622616 671948 622668
rect 674288 622616 674340 622668
rect 676036 622616 676088 622668
rect 674012 622548 674064 622600
rect 670424 622412 670476 622464
rect 672632 622412 672684 622464
rect 674288 622412 674340 622464
rect 676404 622412 676456 622464
rect 674288 621392 674340 621444
rect 676036 621392 676088 621444
rect 673184 621324 673236 621376
rect 674012 621324 674064 621376
rect 671436 621120 671488 621172
rect 673276 621120 673328 621172
rect 667664 620984 667716 621036
rect 674012 620984 674064 621036
rect 670884 620780 670936 620832
rect 674012 620780 674064 620832
rect 674288 620780 674340 620832
rect 676220 620780 676272 620832
rect 42248 620236 42300 620288
rect 42708 620236 42760 620288
rect 669780 620236 669832 620288
rect 674012 620236 674064 620288
rect 674288 620100 674340 620152
rect 676496 620100 676548 620152
rect 674288 619896 674340 619948
rect 676220 619896 676272 619948
rect 668400 619692 668452 619744
rect 674012 619692 674064 619744
rect 42248 619624 42300 619676
rect 43076 619624 43128 619676
rect 672448 619556 672500 619608
rect 674012 619556 674064 619608
rect 674288 619488 674340 619540
rect 676220 619488 676272 619540
rect 43812 618264 43864 618316
rect 668216 617448 668268 617500
rect 673276 617448 673328 617500
rect 42248 617312 42300 617364
rect 674288 617108 674340 617160
rect 676036 617108 676088 617160
rect 669044 616836 669096 616888
rect 674012 616836 674064 616888
rect 44180 616768 44232 616820
rect 62120 616768 62172 616820
rect 42156 616292 42208 616344
rect 42524 616292 42576 616344
rect 670608 615612 670660 615664
rect 674012 615612 674064 615664
rect 674288 615476 674340 615528
rect 683120 615476 683172 615528
rect 670608 614864 670660 614916
rect 674012 614864 674064 614916
rect 42708 614116 42760 614168
rect 62120 614116 62172 614168
rect 43260 612620 43312 612672
rect 42248 612348 42300 612400
rect 58624 612620 58676 612672
rect 62120 612620 62172 612672
rect 43766 611940 43818 611992
rect 44916 611940 44968 611992
rect 43996 611600 44048 611652
rect 44211 611532 44263 611584
rect 653404 611328 653456 611380
rect 674012 611328 674064 611380
rect 674288 611328 674340 611380
rect 675392 611328 675444 611380
rect 50160 611260 50212 611312
rect 44732 611056 44784 611108
rect 46204 610852 46256 610904
rect 44732 610716 44784 610768
rect 50160 609968 50212 610020
rect 61384 609968 61436 610020
rect 667664 608608 667716 608660
rect 674012 608608 674064 608660
rect 674288 608608 674340 608660
rect 675116 608608 675168 608660
rect 674472 603236 674524 603288
rect 675116 603236 675168 603288
rect 35808 601672 35860 601724
rect 36544 601672 36596 601724
rect 657544 600312 657596 600364
rect 674012 600448 674064 600500
rect 674288 600312 674340 600364
rect 675116 600312 675168 600364
rect 674656 599564 674708 599616
rect 675300 599564 675352 599616
rect 654784 598952 654836 599004
rect 674012 599496 674064 599548
rect 674288 599360 674340 599412
rect 675300 599360 675352 599412
rect 675300 598408 675352 598460
rect 675300 598136 675352 598188
rect 651472 597524 651524 597576
rect 669964 597524 670016 597576
rect 42892 597388 42944 597440
rect 42892 596980 42944 597032
rect 651472 596164 651524 596216
rect 664444 596164 664496 596216
rect 40132 595756 40184 595808
rect 41696 595756 41748 595808
rect 651656 595484 651708 595536
rect 653404 595484 653456 595536
rect 651472 594804 651524 594856
rect 661684 594804 661736 594856
rect 41328 594736 41380 594788
rect 41512 594736 41564 594788
rect 651472 594668 651524 594720
rect 657544 594668 657596 594720
rect 39948 594532 40000 594584
rect 41696 594532 41748 594584
rect 651472 593240 651524 593292
rect 654784 593240 654836 593292
rect 675300 592628 675352 592680
rect 683396 592628 683448 592680
rect 40960 592492 41012 592544
rect 41696 592492 41748 592544
rect 35624 590928 35676 590980
rect 41696 590928 41748 590980
rect 35808 590656 35860 590708
rect 39764 590656 39816 590708
rect 674840 590588 674892 590640
rect 682384 590588 682436 590640
rect 674288 588548 674340 588600
rect 684040 588548 684092 588600
rect 33048 587120 33100 587172
rect 41512 587120 41564 587172
rect 42064 587120 42116 587172
rect 42616 587120 42668 587172
rect 42064 586236 42116 586288
rect 35164 586168 35216 586220
rect 41696 586168 41748 586220
rect 42800 586100 42852 586152
rect 42248 586032 42300 586084
rect 33784 585896 33836 585948
rect 39856 585896 39908 585948
rect 31024 585760 31076 585812
rect 40592 585760 40644 585812
rect 42248 585556 42300 585608
rect 660304 581000 660356 581052
rect 674012 581000 674064 581052
rect 668584 579980 668636 580032
rect 674012 579980 674064 580032
rect 670240 579844 670292 579896
rect 674012 579844 674064 579896
rect 658924 579640 658976 579692
rect 673552 579640 673604 579692
rect 670792 579368 670844 579420
rect 674012 579368 674064 579420
rect 669412 579028 669464 579080
rect 674012 579028 674064 579080
rect 42248 578960 42300 579012
rect 43260 578960 43312 579012
rect 671160 578552 671212 578604
rect 674012 578552 674064 578604
rect 670424 578144 670476 578196
rect 674012 578144 674064 578196
rect 42248 577736 42300 577788
rect 42800 577736 42852 577788
rect 670240 577736 670292 577788
rect 674012 577736 674064 577788
rect 671436 577396 671488 577448
rect 674012 577396 674064 577448
rect 669412 576920 669464 576972
rect 674012 576920 674064 576972
rect 45100 575424 45152 575476
rect 62120 575424 62172 575476
rect 671620 574540 671672 574592
rect 673552 574540 673604 574592
rect 671988 574268 672040 574320
rect 673552 574268 673604 574320
rect 667480 574064 667532 574116
rect 674012 574064 674064 574116
rect 46940 573996 46992 574048
rect 62120 573996 62172 574048
rect 669596 572228 669648 572280
rect 674012 572228 674064 572280
rect 671804 571548 671856 571600
rect 674012 571548 674064 571600
rect 674472 571548 674524 571600
rect 676220 571548 676272 571600
rect 42064 570936 42116 570988
rect 42616 570936 42668 570988
rect 674840 570460 674892 570512
rect 675484 570460 675536 570512
rect 683120 570460 683172 570512
rect 671344 570392 671396 570444
rect 673552 570392 673604 570444
rect 671988 570120 672040 570172
rect 674012 570120 674064 570172
rect 669780 568556 669832 568608
rect 674012 568556 674064 568608
rect 653404 565836 653456 565888
rect 673552 565836 673604 565888
rect 665088 564408 665140 564460
rect 673552 564408 673604 564460
rect 35808 557540 35860 557592
rect 40960 557540 41012 557592
rect 35808 555024 35860 555076
rect 40500 555024 40552 555076
rect 35808 554752 35860 554804
rect 39856 554752 39908 554804
rect 657820 554752 657872 554804
rect 673552 554752 673604 554804
rect 35624 553528 35676 553580
rect 41696 553528 41748 553580
rect 35808 553392 35860 553444
rect 41328 553392 41380 553444
rect 655152 553392 655204 553444
rect 670424 553392 670476 553444
rect 651472 552644 651524 552696
rect 665824 552644 665876 552696
rect 41328 552032 41380 552084
rect 41696 552032 41748 552084
rect 675208 551760 675260 551812
rect 675208 551556 675260 551608
rect 41144 550604 41196 550656
rect 41696 550604 41748 550656
rect 42064 550604 42116 550656
rect 42984 550604 43036 550656
rect 651472 550604 651524 550656
rect 660304 550604 660356 550656
rect 651380 550332 651432 550384
rect 653404 550332 653456 550384
rect 40868 550196 40920 550248
rect 41696 550196 41748 550248
rect 651656 549856 651708 549908
rect 663064 549856 663116 549908
rect 651472 549176 651524 549228
rect 657820 549176 657872 549228
rect 675300 549448 675352 549500
rect 651472 548768 651524 548820
rect 655152 548768 655204 548820
rect 675024 548768 675076 548820
rect 41328 547884 41380 547936
rect 41696 547884 41748 547936
rect 29644 547136 29696 547188
rect 41696 547136 41748 547188
rect 675576 547136 675628 547188
rect 683212 547136 683264 547188
rect 674840 545844 674892 545896
rect 682384 545844 682436 545896
rect 673920 540880 673972 540932
rect 673736 540608 673788 540660
rect 669964 535780 670016 535832
rect 674012 535780 674064 535832
rect 674288 535712 674340 535764
rect 676036 535712 676088 535764
rect 674288 535508 674340 535560
rect 676220 535508 676272 535560
rect 664444 535440 664496 535492
rect 674012 535440 674064 535492
rect 670792 534964 670844 535016
rect 674012 534964 674064 535016
rect 674288 534896 674340 534948
rect 676036 534896 676088 534948
rect 674288 534420 674340 534472
rect 676036 534420 676088 534472
rect 670792 534352 670844 534404
rect 674012 534352 674064 534404
rect 674288 534284 674340 534336
rect 676220 534284 676272 534336
rect 661684 534216 661736 534268
rect 674012 534216 674064 534268
rect 671160 534080 671212 534132
rect 674012 534080 674064 534132
rect 674288 534080 674340 534132
rect 676036 534080 676088 534132
rect 674288 533332 674340 533384
rect 683580 533332 683632 533384
rect 671620 533060 671672 533112
rect 674012 533060 674064 533112
rect 674288 533060 674340 533112
rect 676220 533060 676272 533112
rect 674288 532924 674340 532976
rect 676036 532924 676088 532976
rect 670240 532856 670292 532908
rect 674012 532856 674064 532908
rect 674288 532788 674340 532840
rect 676404 532788 676456 532840
rect 672724 532720 672776 532772
rect 674012 532720 674064 532772
rect 674288 532176 674340 532228
rect 676404 532176 676456 532228
rect 667664 532108 667716 532160
rect 674012 532108 674064 532160
rect 674288 532040 674340 532092
rect 676220 532040 676272 532092
rect 44732 531972 44784 532024
rect 62120 531972 62172 532024
rect 674012 531972 674064 532024
rect 669412 531564 669464 531616
rect 674288 531700 674340 531752
rect 676036 531700 676088 531752
rect 671160 531428 671212 531480
rect 674012 531428 674064 531480
rect 51724 531224 51776 531276
rect 62304 531224 62356 531276
rect 42156 530680 42208 530732
rect 42708 530680 42760 530732
rect 42248 530272 42300 530324
rect 42708 530272 42760 530324
rect 667296 529932 667348 529984
rect 674012 529932 674064 529984
rect 674288 529932 674340 529984
rect 676036 529932 676088 529984
rect 674288 529320 674340 529372
rect 676220 529320 676272 529372
rect 668952 529116 669004 529168
rect 674012 529116 674064 529168
rect 674288 528980 674340 529032
rect 676220 528980 676272 529032
rect 670976 528912 671028 528964
rect 674012 528912 674064 528964
rect 672356 528708 672408 528760
rect 674012 528708 674064 528760
rect 674288 528708 674340 528760
rect 676036 528708 676088 528760
rect 44824 528572 44876 528624
rect 62120 528572 62172 528624
rect 672540 528096 672592 528148
rect 673368 528096 673420 528148
rect 47584 527076 47636 527128
rect 62120 527076 62172 527128
rect 674656 526736 674708 526788
rect 676036 526736 676088 526788
rect 674288 526328 674340 526380
rect 676036 526328 676088 526380
rect 662420 525036 662472 525088
rect 668768 525036 668820 525088
rect 674012 525036 674064 525088
rect 674288 524560 674340 524612
rect 683120 524560 683172 524612
rect 658924 521976 658976 522028
rect 662420 521976 662472 522028
rect 675484 520208 675536 520260
rect 678980 520208 679032 520260
rect 675668 518780 675720 518832
rect 677876 518780 677928 518832
rect 656164 512864 656216 512916
rect 658924 512864 658976 512916
rect 675116 503616 675168 503668
rect 679624 503616 679676 503668
rect 675300 503480 675352 503532
rect 681004 503480 681056 503532
rect 674932 500896 674984 500948
rect 681188 500896 681240 500948
rect 650644 499536 650696 499588
rect 656164 499536 656216 499588
rect 674288 494980 674340 495032
rect 674656 494980 674708 495032
rect 674288 491648 674340 491700
rect 676036 491648 676088 491700
rect 665824 491580 665876 491632
rect 674012 491580 674064 491632
rect 663064 491444 663116 491496
rect 673828 491444 673880 491496
rect 660304 491308 660356 491360
rect 674012 491308 674064 491360
rect 670792 490900 670844 490952
rect 674012 490900 674064 490952
rect 672632 489880 672684 489932
rect 673368 489880 673420 489932
rect 672448 489608 672500 489660
rect 674012 489608 674064 489660
rect 671620 489268 671672 489320
rect 674012 489268 674064 489320
rect 671160 488452 671212 488504
rect 674012 488452 674064 488504
rect 674288 486752 674340 486804
rect 676036 486752 676088 486804
rect 665088 485800 665140 485852
rect 674012 485800 674064 485852
rect 674288 485120 674340 485172
rect 676036 485120 676088 485172
rect 668584 484372 668636 484424
rect 674012 484372 674064 484424
rect 674472 483964 674524 484016
rect 676036 483964 676088 484016
rect 671804 483148 671856 483200
rect 674012 483148 674064 483200
rect 676220 482944 676272 482996
rect 677416 482944 677468 482996
rect 670424 480360 670476 480412
rect 674012 480360 674064 480412
rect 674288 480360 674340 480412
rect 683120 480360 683172 480412
rect 667480 477504 667532 477556
rect 670424 477504 670476 477556
rect 676036 476076 676088 476128
rect 680360 476076 680412 476128
rect 664444 474240 664496 474292
rect 667480 474240 667532 474292
rect 652760 467100 652812 467152
rect 664444 467100 664496 467152
rect 650828 461320 650880 461372
rect 652760 461320 652812 461372
rect 667020 456560 667072 456612
rect 667848 455948 667900 456000
rect 672172 455812 672224 455864
rect 669228 455608 669280 455660
rect 673276 455336 673328 455388
rect 673388 455200 673440 455252
rect 673506 455200 673558 455252
rect 674288 454860 674340 454912
rect 675852 454860 675904 454912
rect 672080 454792 672132 454844
rect 673046 454588 673098 454640
rect 674288 454588 674340 454640
rect 675484 454588 675536 454640
rect 672816 454452 672868 454504
rect 672954 454316 673006 454368
rect 674288 454316 674340 454368
rect 675668 454316 675720 454368
rect 672264 453908 672316 453960
rect 674288 453908 674340 453960
rect 676036 453908 676088 453960
rect 35808 429156 35860 429208
rect 41696 429156 41748 429208
rect 35808 427932 35860 427984
rect 41696 427932 41748 427984
rect 41144 424328 41196 424380
rect 41696 424328 41748 424380
rect 32772 417392 32824 417444
rect 41696 417392 41748 417444
rect 42064 417256 42116 417308
rect 42616 417256 42668 417308
rect 34520 416032 34572 416084
rect 41604 416032 41656 416084
rect 42248 406988 42300 407040
rect 42616 406988 42668 407040
rect 45284 404268 45336 404320
rect 62120 404268 62172 404320
rect 674564 403248 674616 403300
rect 676220 403248 676272 403300
rect 51448 402908 51500 402960
rect 62120 402908 62172 402960
rect 42432 402500 42484 402552
rect 42984 402500 43036 402552
rect 42432 402024 42484 402076
rect 43260 402024 43312 402076
rect 51080 400188 51132 400240
rect 62120 400188 62172 400240
rect 44824 400052 44876 400104
rect 62120 400052 62172 400104
rect 674932 398828 674984 398880
rect 676036 398828 676088 398880
rect 47768 398760 47820 398812
rect 62120 398760 62172 398812
rect 674564 396040 674616 396092
rect 676036 396040 676088 396092
rect 675208 395700 675260 395752
rect 676220 395700 676272 395752
rect 674380 394272 674432 394324
rect 676220 394272 676272 394324
rect 41328 386384 41380 386436
rect 41696 386384 41748 386436
rect 679624 386724 679676 386776
rect 675484 385976 675536 386028
rect 674840 384752 674892 384804
rect 675392 384752 675444 384804
rect 41328 382372 41380 382424
rect 41696 382372 41748 382424
rect 674380 382168 674432 382220
rect 675116 382168 675168 382220
rect 41328 379720 41380 379772
rect 41512 379720 41564 379772
rect 35808 379584 35860 379636
rect 40408 379584 40460 379636
rect 35808 378156 35860 378208
rect 41696 378156 41748 378208
rect 674380 378088 674432 378140
rect 675116 378088 675168 378140
rect 651472 373940 651524 373992
rect 657544 373940 657596 373992
rect 33968 373260 34020 373312
rect 41696 373260 41748 373312
rect 39304 371832 39356 371884
rect 41696 371832 41748 371884
rect 42064 371696 42116 371748
rect 42708 371696 42760 371748
rect 651472 370948 651524 371000
rect 654784 370948 654836 371000
rect 42340 366800 42392 366852
rect 43076 366800 43128 366852
rect 42248 364964 42300 365016
rect 42708 364964 42760 365016
rect 651012 362924 651064 362976
rect 655520 362924 655572 362976
rect 45652 361496 45704 361548
rect 62120 361496 62172 361548
rect 51080 360136 51132 360188
rect 62120 360136 62172 360188
rect 44640 357416 44692 357468
rect 62120 357416 62172 357468
rect 42248 355988 42300 356040
rect 42892 355988 42944 356040
rect 47768 355988 47820 356040
rect 62120 355988 62172 356040
rect 44640 354492 44692 354544
rect 44732 354356 44784 354408
rect 45652 354288 45704 354340
rect 45836 354152 45888 354204
rect 45468 354016 45520 354068
rect 45468 353880 45520 353932
rect 45468 353404 45520 353456
rect 45422 353132 45474 353184
rect 35808 344564 35860 344616
rect 39856 344564 39908 344616
rect 35624 343612 35676 343664
rect 40040 343612 40092 343664
rect 35808 342252 35860 342304
rect 40224 342252 40276 342304
rect 33048 341368 33100 341420
rect 40224 341368 40276 341420
rect 45468 341368 45520 341420
rect 62304 341368 62356 341420
rect 35808 341164 35860 341216
rect 40224 341164 40276 341216
rect 35808 341028 35860 341080
rect 40040 341028 40092 341080
rect 35808 339600 35860 339652
rect 37924 339600 37976 339652
rect 35532 339464 35584 339516
rect 38660 339464 38712 339516
rect 35808 335316 35860 335368
rect 40224 335316 40276 335368
rect 35808 334092 35860 334144
rect 39764 334092 39816 334144
rect 674472 331032 674524 331084
rect 675116 331032 675168 331084
rect 651380 328244 651432 328296
rect 654784 328244 654836 328296
rect 651380 325592 651432 325644
rect 653404 325592 653456 325644
rect 42432 322872 42484 322924
rect 43076 322872 43128 322924
rect 42248 321512 42300 321564
rect 42892 321512 42944 321564
rect 45468 317364 45520 317416
rect 62120 317364 62172 317416
rect 62120 314712 62172 314764
rect 45468 314644 45520 314696
rect 674380 311992 674432 312044
rect 675484 311992 675536 312044
rect 674748 309816 674800 309868
rect 675484 309816 675536 309868
rect 676220 306348 676272 306400
rect 676864 306348 676916 306400
rect 675852 304852 675904 304904
rect 676404 304852 676456 304904
rect 651380 303492 651432 303544
rect 653404 303492 653456 303544
rect 41328 300840 41380 300892
rect 41696 300840 41748 300892
rect 46388 300772 46440 300824
rect 52092 300772 52144 300824
rect 651472 300772 651524 300824
rect 658924 300772 658976 300824
rect 47584 299412 47636 299464
rect 54484 299412 54536 299464
rect 41144 299072 41196 299124
rect 41696 299072 41748 299124
rect 651472 298120 651524 298172
rect 660580 298120 660632 298172
rect 674748 297780 674800 297832
rect 675484 297780 675536 297832
rect 676036 297576 676088 297628
rect 678980 297576 679032 297628
rect 675852 297440 675904 297492
rect 678244 297440 678296 297492
rect 652208 296760 652260 296812
rect 658924 296692 658976 296744
rect 675300 296148 675352 296200
rect 41144 295468 41196 295520
rect 41696 295468 41748 295520
rect 675300 295400 675352 295452
rect 45468 295332 45520 295384
rect 62120 295332 62172 295384
rect 41328 294244 41380 294296
rect 41696 294244 41748 294296
rect 42064 294244 42116 294296
rect 42616 294244 42668 294296
rect 57428 294040 57480 294092
rect 62120 294040 62172 294092
rect 651472 293972 651524 294024
rect 664444 293972 664496 294024
rect 42064 293020 42116 293072
rect 43352 293020 43404 293072
rect 41696 292748 41748 292800
rect 41328 292680 41380 292732
rect 60372 292544 60424 292596
rect 62304 292544 62356 292596
rect 651472 292544 651524 292596
rect 660304 292544 660356 292596
rect 45468 292408 45520 292460
rect 62120 292408 62172 292460
rect 651472 289824 651524 289876
rect 663064 289824 663116 289876
rect 54484 288396 54536 288448
rect 57612 288396 57664 288448
rect 651472 288396 651524 288448
rect 672172 288396 672224 288448
rect 651472 287036 651524 287088
rect 667572 287036 667624 287088
rect 33784 286288 33836 286340
rect 41512 286288 41564 286340
rect 45468 285676 45520 285728
rect 62120 285676 62172 285728
rect 651472 285676 651524 285728
rect 667388 285676 667440 285728
rect 39948 284452 40000 284504
rect 41696 284452 41748 284504
rect 46388 284316 46440 284368
rect 63224 284316 63276 284368
rect 651472 284316 651524 284368
rect 672356 284316 672408 284368
rect 51724 282888 51776 282940
rect 62120 282888 62172 282940
rect 651472 282888 651524 282940
rect 666560 282888 666612 282940
rect 56048 281528 56100 281580
rect 62856 281528 62908 281580
rect 651472 280168 651524 280220
rect 667204 280168 667256 280220
rect 42432 280100 42484 280152
rect 43076 280100 43128 280152
rect 58624 280032 58676 280084
rect 61936 280032 61988 280084
rect 57612 278672 57664 278724
rect 61752 278672 61804 278724
rect 63500 278672 63552 278724
rect 671344 278672 671396 278724
rect 49332 278536 49384 278588
rect 60556 278536 60608 278588
rect 61936 278536 61988 278588
rect 63316 278536 63368 278588
rect 671712 278536 671764 278588
rect 650828 278400 650880 278452
rect 52092 278264 52144 278316
rect 60556 278264 60608 278316
rect 61752 278264 61804 278316
rect 651012 278264 651064 278316
rect 51908 278128 51960 278180
rect 629944 278128 629996 278180
rect 630128 278128 630180 278180
rect 650644 278128 650696 278180
rect 47768 277992 47820 278044
rect 635096 277992 635148 278044
rect 64328 277856 64380 277908
rect 637764 277856 637816 277908
rect 61936 277584 61988 277636
rect 629944 277720 629996 277772
rect 636292 277720 636344 277772
rect 630128 277584 630180 277636
rect 479984 277312 480036 277364
rect 555240 277312 555292 277364
rect 487988 277176 488040 277228
rect 565820 277176 565872 277228
rect 497924 277040 497976 277092
rect 579988 277040 580040 277092
rect 511632 276904 511684 276956
rect 600136 276904 600188 276956
rect 42248 276768 42300 276820
rect 42616 276768 42668 276820
rect 514484 276768 514536 276820
rect 603632 276768 603684 276820
rect 53288 276632 53340 276684
rect 62120 276632 62172 276684
rect 518716 276632 518768 276684
rect 609612 276632 609664 276684
rect 482836 276496 482888 276548
rect 557540 276496 557592 276548
rect 477040 276360 477092 276412
rect 550456 276360 550508 276412
rect 471612 276224 471664 276276
rect 543372 276224 543424 276276
rect 107200 275952 107252 276004
rect 163504 275952 163556 276004
rect 167552 275952 167604 276004
rect 178684 275952 178736 276004
rect 185216 275952 185268 276004
rect 221280 275952 221332 276004
rect 232504 275952 232556 276004
rect 239220 275952 239272 276004
rect 410800 275952 410852 276004
rect 455880 275952 455932 276004
rect 456064 275952 456116 276004
rect 509056 275952 509108 276004
rect 513196 275952 513248 276004
rect 601332 275952 601384 276004
rect 139124 275816 139176 275868
rect 174268 275816 174320 275868
rect 178132 275816 178184 275868
rect 216680 275816 216732 275868
rect 224224 275816 224276 275868
rect 232688 275816 232740 275868
rect 236092 275816 236144 275868
rect 250444 275816 250496 275868
rect 286876 275816 286928 275868
rect 291844 275816 291896 275868
rect 430212 275816 430264 275868
rect 484308 275816 484360 275868
rect 490564 275816 490616 275868
rect 505560 275816 505612 275868
rect 522764 275816 522816 275868
rect 615500 275816 615552 275868
rect 260932 275748 260984 275800
rect 266360 275748 266412 275800
rect 100116 275680 100168 275732
rect 159456 275680 159508 275732
rect 160468 275680 160520 275732
rect 199568 275680 199620 275732
rect 217140 275680 217192 275732
rect 224224 275680 224276 275732
rect 229008 275680 229060 275732
rect 243544 275680 243596 275732
rect 250260 275680 250312 275732
rect 259368 275680 259420 275732
rect 284576 275680 284628 275732
rect 290096 275680 290148 275732
rect 445024 275680 445076 275732
rect 498476 275680 498528 275732
rect 498844 275680 498896 275732
rect 512644 275680 512696 275732
rect 528192 275680 528244 275732
rect 622584 275680 622636 275732
rect 291660 275612 291712 275664
rect 295340 275612 295392 275664
rect 76472 275544 76524 275596
rect 86224 275544 86276 275596
rect 90732 275544 90784 275596
rect 154764 275544 154816 275596
rect 171048 275544 171100 275596
rect 211620 275544 211672 275596
rect 218336 275544 218388 275596
rect 233884 275544 233936 275596
rect 239588 275544 239640 275596
rect 255964 275544 256016 275596
rect 257344 275544 257396 275596
rect 262312 275544 262364 275596
rect 266820 275544 266872 275596
rect 276480 275544 276532 275596
rect 363880 275544 363932 275596
rect 388536 275544 388588 275596
rect 416412 275544 416464 275596
rect 462964 275544 463016 275596
rect 463148 275544 463200 275596
rect 516232 275544 516284 275596
rect 516784 275544 516836 275596
rect 526812 275544 526864 275596
rect 532332 275544 532384 275596
rect 629668 275544 629720 275596
rect 277492 275476 277544 275528
rect 285128 275476 285180 275528
rect 81256 275408 81308 275460
rect 144920 275408 144972 275460
rect 156880 275408 156932 275460
rect 96620 275272 96672 275324
rect 149612 275272 149664 275324
rect 163964 275408 164016 275460
rect 206376 275408 206428 275460
rect 221924 275408 221976 275460
rect 243728 275408 243780 275460
rect 256148 275408 256200 275460
rect 200764 275272 200816 275324
rect 214840 275272 214892 275324
rect 239404 275272 239456 275324
rect 243176 275272 243228 275324
rect 256700 275272 256752 275324
rect 285680 275408 285732 275460
rect 291292 275408 291344 275460
rect 358636 275408 358688 275460
rect 381452 275408 381504 275460
rect 386052 275408 386104 275460
rect 420460 275408 420512 275460
rect 435640 275408 435692 275460
rect 485044 275408 485096 275460
rect 485228 275408 485280 275460
rect 530400 275408 530452 275460
rect 537668 275408 537720 275460
rect 636752 275408 636804 275460
rect 269212 275340 269264 275392
rect 274640 275340 274692 275392
rect 297548 275340 297600 275392
rect 299572 275340 299624 275392
rect 299940 275340 299992 275392
rect 301136 275340 301188 275392
rect 276296 275272 276348 275324
rect 283104 275272 283156 275324
rect 290464 275272 290516 275324
rect 294144 275272 294196 275324
rect 326436 275272 326488 275324
rect 335360 275272 335412 275324
rect 371056 275272 371108 275324
rect 399208 275272 399260 275324
rect 418804 275272 418856 275324
rect 466552 275272 466604 275324
rect 467564 275272 467616 275324
rect 537484 275272 537536 275324
rect 542268 275272 542320 275324
rect 643836 275272 643888 275324
rect 269120 275204 269172 275256
rect 298744 275204 298796 275256
rect 300032 275204 300084 275256
rect 93032 275136 93084 275188
rect 152832 275136 152884 275188
rect 153384 275136 153436 275188
rect 169024 275136 169076 275188
rect 190000 275136 190052 275188
rect 222936 275136 222988 275188
rect 292856 275136 292908 275188
rect 295800 275136 295852 275188
rect 427084 275136 427136 275188
rect 477224 275136 477276 275188
rect 485044 275136 485096 275188
rect 491392 275136 491444 275188
rect 507492 275136 507544 275188
rect 594248 275136 594300 275188
rect 263232 275068 263284 275120
rect 273260 275068 273312 275120
rect 71780 275000 71832 275052
rect 141056 275000 141108 275052
rect 149796 275000 149848 275052
rect 189080 275000 189132 275052
rect 288072 275000 288124 275052
rect 292672 275000 292724 275052
rect 420552 275000 420604 275052
rect 470140 275000 470192 275052
rect 484308 275000 484360 275052
rect 485228 275000 485280 275052
rect 503444 275000 503496 275052
rect 587072 275000 587124 275052
rect 293960 274932 294012 274984
rect 296812 274932 296864 274984
rect 146208 274864 146260 274916
rect 185584 274864 185636 274916
rect 473084 274864 473136 274916
rect 544568 274864 544620 274916
rect 289268 274796 289320 274848
rect 293408 274796 293460 274848
rect 295156 274796 295208 274848
rect 297456 274796 297508 274848
rect 128544 274728 128596 274780
rect 168288 274728 168340 274780
rect 207756 274728 207808 274780
rect 210700 274728 210752 274780
rect 476764 274728 476816 274780
rect 523316 274728 523368 274780
rect 523684 274728 523736 274780
rect 533896 274728 533948 274780
rect 534724 274728 534776 274780
rect 540980 274728 541032 274780
rect 74172 274660 74224 274712
rect 76840 274660 76892 274712
rect 85948 274660 86000 274712
rect 90364 274660 90416 274712
rect 103704 274660 103756 274712
rect 104808 274660 104860 274712
rect 110788 274660 110840 274712
rect 111708 274660 111760 274712
rect 253848 274660 253900 274712
rect 256884 274660 256936 274712
rect 275100 274660 275152 274712
rect 278044 274660 278096 274712
rect 283380 274660 283432 274712
rect 289176 274660 289228 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 303436 274660 303488 274712
rect 303988 274660 304040 274712
rect 321192 274660 321244 274712
rect 328276 274660 328328 274712
rect 114376 274592 114428 274644
rect 171600 274592 171652 274644
rect 179328 274592 179380 274644
rect 214564 274592 214616 274644
rect 409788 274592 409840 274644
rect 453580 274592 453632 274644
rect 457444 274592 457496 274644
rect 480720 274592 480772 274644
rect 486792 274592 486844 274644
rect 563428 274592 563480 274644
rect 101312 274456 101364 274508
rect 160928 274456 160980 274508
rect 168748 274456 168800 274508
rect 208400 274456 208452 274508
rect 381544 274456 381596 274508
rect 392124 274456 392176 274508
rect 413836 274456 413888 274508
rect 460664 274456 460716 274508
rect 463240 274456 463292 274508
rect 484308 274456 484360 274508
rect 488356 274456 488408 274508
rect 567016 274456 567068 274508
rect 95424 274320 95476 274372
rect 157616 274320 157668 274372
rect 159272 274320 159324 274372
rect 202328 274320 202380 274372
rect 223120 274320 223172 274372
rect 247224 274320 247276 274372
rect 369124 274320 369176 274372
rect 387340 274320 387392 274372
rect 419080 274320 419132 274372
rect 467748 274320 467800 274372
rect 506204 274320 506256 274372
rect 591856 274320 591908 274372
rect 67088 274184 67140 274236
rect 130384 274184 130436 274236
rect 130844 274184 130896 274236
rect 182456 274184 182508 274236
rect 192392 274184 192444 274236
rect 224960 274184 225012 274236
rect 239220 274184 239272 274236
rect 253940 274184 253992 274236
rect 331864 274184 331916 274236
rect 337752 274184 337804 274236
rect 359464 274184 359516 274236
rect 380256 274184 380308 274236
rect 388996 274184 389048 274236
rect 425244 274184 425296 274236
rect 425704 274184 425756 274236
rect 474832 274184 474884 274236
rect 511816 274184 511868 274236
rect 598940 274184 598992 274236
rect 77668 274048 77720 274100
rect 145104 274048 145156 274100
rect 154488 274048 154540 274100
rect 198096 274048 198148 274100
rect 210056 274048 210108 274100
rect 237840 274048 237892 274100
rect 249064 274048 249116 274100
rect 265256 274048 265308 274100
rect 266360 274048 266412 274100
rect 273536 274048 273588 274100
rect 278596 274048 278648 274100
rect 285864 274048 285916 274100
rect 337752 274048 337804 274100
rect 351920 274048 351972 274100
rect 353944 274048 353996 274100
rect 369584 274048 369636 274100
rect 373264 274048 373316 274100
rect 400312 274048 400364 274100
rect 401508 274048 401560 274100
rect 442908 274048 442960 274100
rect 451188 274048 451240 274100
rect 513840 274048 513892 274100
rect 536748 274048 536800 274100
rect 634360 274048 634412 274100
rect 69388 273912 69440 273964
rect 139400 273912 139452 273964
rect 144920 273912 144972 273964
rect 147864 273912 147916 273964
rect 148600 273912 148652 273964
rect 194784 273912 194836 273964
rect 208860 273912 208912 273964
rect 237380 273912 237432 273964
rect 238484 273912 238536 273964
rect 88340 273776 88392 273828
rect 119344 273776 119396 273828
rect 120264 273776 120316 273828
rect 175280 273776 175332 273828
rect 193496 273776 193548 273828
rect 226432 273776 226484 273828
rect 271512 273912 271564 273964
rect 280344 273912 280396 273964
rect 322756 273912 322808 273964
rect 330576 273912 330628 273964
rect 335268 273912 335320 273964
rect 348332 273912 348384 273964
rect 350356 273912 350408 273964
rect 368480 273912 368532 273964
rect 377680 273912 377732 273964
rect 408592 273912 408644 273964
rect 422116 273912 422168 273964
rect 472440 273912 472492 273964
rect 474648 273912 474700 273964
rect 545764 273912 545816 273964
rect 545948 273912 546000 273964
rect 639144 273912 639196 273964
rect 258080 273776 258132 273828
rect 259368 273776 259420 273828
rect 266360 273776 266412 273828
rect 397000 273776 397052 273828
rect 435824 273776 435876 273828
rect 438124 273776 438176 273828
rect 473636 273776 473688 273828
rect 481364 273776 481416 273828
rect 556344 273776 556396 273828
rect 556804 273776 556856 273828
rect 590660 273776 590712 273828
rect 119068 273640 119120 273692
rect 173256 273640 173308 273692
rect 447784 273640 447836 273692
rect 481916 273640 481968 273692
rect 484216 273640 484268 273692
rect 559932 273640 559984 273692
rect 132040 273504 132092 273556
rect 153844 273504 153896 273556
rect 440884 273504 440936 273556
rect 471244 273504 471296 273556
rect 476028 273504 476080 273556
rect 549260 273504 549312 273556
rect 549904 273504 549956 273556
rect 583576 273504 583628 273556
rect 478696 273368 478748 273420
rect 552848 273368 552900 273420
rect 460572 273300 460624 273352
rect 461400 273300 461452 273352
rect 327724 273232 327776 273284
rect 329472 273232 329524 273284
rect 108396 273164 108448 273216
rect 165896 273164 165948 273216
rect 186412 273164 186464 273216
rect 218704 273164 218756 273216
rect 362776 273164 362828 273216
rect 385868 273164 385920 273216
rect 400036 273164 400088 273216
rect 439320 273164 439372 273216
rect 444012 273164 444064 273216
rect 503168 273164 503220 273216
rect 504180 273164 504232 273216
rect 511448 273164 511500 273216
rect 102508 273028 102560 273080
rect 162860 273028 162912 273080
rect 172244 273028 172296 273080
rect 209780 273028 209832 273080
rect 219532 273028 219584 273080
rect 244556 273028 244608 273080
rect 280988 273028 281040 273080
rect 286324 273028 286376 273080
rect 361212 273028 361264 273080
rect 384948 273028 385000 273080
rect 385684 273028 385736 273080
rect 395620 273028 395672 273080
rect 404176 273028 404228 273080
rect 446496 273028 446548 273080
rect 452292 273028 452344 273080
rect 94228 272892 94280 272944
rect 156144 272892 156196 272944
rect 166356 272892 166408 272944
rect 207296 272892 207348 272944
rect 211252 272892 211304 272944
rect 220084 272892 220136 272944
rect 220728 272892 220780 272944
rect 245752 272892 245804 272944
rect 247868 272892 247920 272944
rect 264244 272892 264296 272944
rect 333796 272892 333848 272944
rect 345940 272892 345992 272944
rect 348424 272892 348476 272944
rect 362500 272892 362552 272944
rect 365444 272892 365496 272944
rect 390928 272892 390980 272944
rect 405556 272892 405608 272944
rect 448796 272892 448848 272944
rect 455328 272892 455380 272944
rect 460572 272892 460624 272944
rect 461768 273028 461820 273080
rect 518532 273164 518584 273216
rect 515036 273028 515088 273080
rect 515404 273028 515456 273080
rect 519728 273164 519780 273216
rect 521476 273164 521528 273216
rect 614304 273164 614356 273216
rect 526812 273028 526864 273080
rect 621388 273028 621440 273080
rect 82452 272756 82504 272808
rect 148416 272756 148468 272808
rect 155684 272756 155736 272808
rect 200120 272756 200172 272808
rect 205364 272756 205416 272808
rect 234804 272756 234856 272808
rect 245384 272756 245436 272808
rect 72976 272620 73028 272672
rect 142160 272620 142212 272672
rect 142712 272620 142764 272672
rect 145564 272620 145616 272672
rect 145748 272620 145800 272672
rect 192392 272620 192444 272672
rect 197084 272620 197136 272672
rect 229100 272620 229152 272672
rect 233700 272620 233752 272672
rect 254400 272620 254452 272672
rect 262312 272756 262364 272808
rect 270960 272756 271012 272808
rect 274272 272756 274324 272808
rect 282920 272756 282972 272808
rect 325332 272756 325384 272808
rect 332968 272756 333020 272808
rect 344652 272756 344704 272808
rect 361396 272756 361448 272808
rect 362224 272756 362276 272808
rect 370320 272756 370372 272808
rect 370504 272756 370556 272808
rect 396816 272756 396868 272808
rect 406844 272756 406896 272808
rect 449992 272756 450044 272808
rect 450544 272756 450596 272808
rect 501052 272756 501104 272808
rect 504364 272756 504416 272808
rect 525616 272892 525668 272944
rect 532516 272892 532568 272944
rect 537944 272892 537996 272944
rect 538128 272892 538180 272944
rect 624976 272892 625028 272944
rect 514208 272756 514260 272808
rect 562140 272756 562192 272808
rect 562324 272756 562376 272808
rect 601148 272756 601200 272808
rect 262680 272620 262732 272672
rect 264428 272620 264480 272672
rect 276020 272620 276072 272672
rect 324044 272620 324096 272672
rect 331404 272620 331456 272672
rect 332324 272620 332376 272672
rect 343640 272620 343692 272672
rect 346216 272620 346268 272672
rect 363696 272620 363748 272672
rect 376116 272620 376168 272672
rect 406292 272620 406344 272672
rect 412272 272620 412324 272672
rect 457076 272620 457128 272672
rect 457260 272620 457312 272672
rect 459376 272620 459428 272672
rect 459560 272620 459612 272672
rect 466414 272620 466466 272672
rect 522120 272620 522172 272672
rect 529848 272620 529900 272672
rect 65892 272484 65944 272536
rect 136824 272484 136876 272536
rect 137928 272484 137980 272536
rect 116676 272348 116728 272400
rect 172520 272348 172572 272400
rect 181720 272484 181772 272536
rect 186964 272484 187016 272536
rect 195888 272484 195940 272536
rect 227904 272484 227956 272536
rect 228088 272484 228140 272536
rect 249064 272484 249116 272536
rect 254952 272484 255004 272536
rect 269304 272484 269356 272536
rect 270316 272484 270368 272536
rect 280528 272484 280580 272536
rect 329748 272484 329800 272536
rect 338856 272484 338908 272536
rect 339224 272484 339276 272536
rect 354220 272484 354272 272536
rect 354496 272484 354548 272536
rect 375564 272484 375616 272536
rect 379428 272484 379480 272536
rect 410984 272484 411036 272536
rect 416596 272484 416648 272536
rect 463884 272484 463936 272536
rect 470554 272484 470606 272536
rect 470692 272484 470744 272536
rect 532700 272484 532752 272536
rect 533712 272620 533764 272672
rect 536380 272484 536432 272536
rect 536564 272484 536616 272536
rect 538128 272484 538180 272536
rect 538680 272620 538732 272672
rect 628472 272620 628524 272672
rect 634084 272620 634136 272672
rect 640340 272620 640392 272672
rect 632060 272484 632112 272536
rect 187700 272348 187752 272400
rect 194968 272348 195020 272400
rect 227168 272348 227220 272400
rect 318708 272348 318760 272400
rect 324688 272348 324740 272400
rect 395988 272348 396040 272400
rect 434628 272348 434680 272400
rect 446864 272348 446916 272400
rect 500868 272348 500920 272400
rect 501052 272348 501104 272400
rect 509700 272348 509752 272400
rect 517428 272348 517480 272400
rect 600964 272348 601016 272400
rect 601148 272348 601200 272400
rect 635556 272348 635608 272400
rect 269120 272280 269172 272332
rect 270592 272280 270644 272332
rect 127348 272212 127400 272264
rect 179880 272212 179932 272264
rect 189080 272212 189132 272264
rect 196440 272212 196492 272264
rect 391848 272212 391900 272264
rect 428740 272212 428792 272264
rect 449716 272212 449768 272264
rect 504180 272212 504232 272264
rect 504548 272212 504600 272264
rect 507952 272212 508004 272264
rect 509700 272212 509752 272264
rect 514208 272212 514260 272264
rect 520096 272212 520148 272264
rect 610716 272212 610768 272264
rect 147404 272076 147456 272128
rect 193220 272076 193272 272128
rect 384948 272076 385000 272128
rect 418068 272076 418120 272128
rect 428464 272076 428516 272128
rect 470554 272076 470606 272128
rect 470784 272076 470836 272128
rect 124956 271940 125008 271992
rect 151084 271940 151136 271992
rect 431684 271940 431736 271992
rect 483020 272076 483072 272128
rect 547512 272076 547564 272128
rect 547696 272076 547748 272128
rect 562324 272076 562376 272128
rect 600964 272076 601016 272128
rect 607220 272076 607272 272128
rect 106004 271804 106056 271856
rect 164976 271804 165028 271856
rect 174268 271804 174320 271856
rect 189172 271804 189224 271856
rect 202972 271804 203024 271856
rect 233240 271804 233292 271856
rect 274640 271804 274692 271856
rect 279240 271804 279292 271856
rect 355324 271804 355376 271856
rect 356612 271804 356664 271856
rect 375288 271804 375340 271856
rect 403900 271804 403952 271856
rect 433156 271804 433208 271856
rect 480168 271804 480220 271856
rect 504364 271940 504416 271992
rect 504548 271940 504600 271992
rect 561956 271940 562008 271992
rect 562140 271940 562192 271992
rect 569408 271940 569460 271992
rect 484860 271804 484912 271856
rect 494704 271804 494756 271856
rect 501420 271804 501472 271856
rect 504364 271804 504416 271856
rect 578516 271804 578568 271856
rect 578884 271804 578936 271856
rect 604828 271804 604880 271856
rect 97816 271668 97868 271720
rect 158812 271668 158864 271720
rect 169852 271668 169904 271720
rect 209964 271668 210016 271720
rect 225420 271668 225472 271720
rect 228364 271668 228416 271720
rect 351184 271668 351236 271720
rect 366088 271668 366140 271720
rect 382004 271668 382056 271720
rect 414572 271668 414624 271720
rect 87144 271532 87196 271584
rect 152004 271532 152056 271584
rect 165160 271532 165212 271584
rect 205640 271532 205692 271584
rect 215944 271532 215996 271584
rect 242072 271532 242124 271584
rect 337936 271532 337988 271584
rect 350724 271532 350776 271584
rect 360844 271532 360896 271584
rect 377864 271532 377916 271584
rect 387708 271532 387760 271584
rect 421656 271668 421708 271720
rect 430396 271668 430448 271720
rect 483204 271668 483256 271720
rect 499304 271668 499356 271720
rect 582380 271668 582432 271720
rect 583024 271668 583076 271720
rect 611912 271668 611964 271720
rect 420184 271532 420236 271584
rect 431132 271532 431184 271584
rect 437204 271532 437256 271584
rect 493692 271532 493744 271584
rect 75368 271396 75420 271448
rect 142712 271396 142764 271448
rect 162676 271396 162728 271448
rect 204720 271396 204772 271448
rect 213644 271396 213696 271448
rect 240416 271396 240468 271448
rect 240784 271396 240836 271448
rect 259644 271396 259696 271448
rect 259828 271396 259880 271448
rect 272616 271396 272668 271448
rect 325516 271396 325568 271448
rect 334164 271396 334216 271448
rect 347688 271396 347740 271448
rect 364892 271396 364944 271448
rect 366364 271396 366416 271448
rect 383844 271396 383896 271448
rect 384764 271396 384816 271448
rect 419264 271396 419316 271448
rect 76840 271260 76892 271312
rect 143540 271260 143592 271312
rect 152188 271260 152240 271312
rect 197360 271260 197412 271312
rect 198280 271260 198332 271312
rect 229560 271260 229612 271312
rect 235264 271260 235316 271312
rect 255320 271260 255372 271312
rect 256700 271260 256752 271312
rect 261024 271260 261076 271312
rect 262036 271260 262088 271312
rect 274640 271260 274692 271312
rect 329564 271260 329616 271312
rect 340052 271260 340104 271312
rect 340604 271260 340656 271312
rect 355140 271260 355192 271312
rect 357164 271260 357216 271312
rect 379060 271260 379112 271312
rect 390284 271260 390336 271312
rect 426348 271396 426400 271448
rect 439964 271396 440016 271448
rect 497280 271532 497332 271584
rect 501972 271532 502024 271584
rect 585968 271532 586020 271584
rect 612004 271532 612056 271584
rect 618996 271532 619048 271584
rect 496544 271396 496596 271448
rect 504364 271396 504416 271448
rect 505008 271396 505060 271448
rect 589464 271396 589516 271448
rect 589924 271396 589976 271448
rect 633256 271396 633308 271448
rect 68192 271124 68244 271176
rect 138480 271124 138532 271176
rect 141516 271124 141568 271176
rect 189816 271124 189868 271176
rect 191196 271124 191248 271176
rect 225144 271124 225196 271176
rect 230204 271124 230256 271176
rect 252008 271124 252060 271176
rect 268016 271124 268068 271176
rect 278780 271124 278832 271176
rect 279792 271124 279844 271176
rect 287060 271124 287112 271176
rect 331128 271124 331180 271176
rect 342444 271124 342496 271176
rect 343548 271124 343600 271176
rect 360200 271124 360252 271176
rect 364156 271124 364208 271176
rect 389732 271124 389784 271176
rect 394332 271124 394384 271176
rect 432236 271260 432288 271312
rect 442908 271260 442960 271312
rect 500684 271260 500736 271312
rect 507676 271260 507728 271312
rect 593052 271260 593104 271312
rect 598204 271260 598256 271312
rect 645032 271260 645084 271312
rect 113456 270988 113508 271040
rect 169944 270988 169996 271040
rect 187424 270988 187476 271040
rect 215944 270988 215996 271040
rect 251456 270988 251508 271040
rect 266912 270988 266964 271040
rect 417424 270988 417476 271040
rect 437940 271124 437992 271176
rect 441344 271124 441396 271176
rect 445024 271124 445076 271176
rect 445668 271124 445720 271176
rect 503996 271124 504048 271176
rect 524052 271124 524104 271176
rect 617340 271124 617392 271176
rect 617524 271124 617576 271176
rect 626080 271124 626132 271176
rect 427452 270988 427504 271040
rect 479156 270988 479208 271040
rect 485044 270988 485096 271040
rect 494704 270988 494756 271040
rect 495072 270988 495124 271040
rect 575296 270988 575348 271040
rect 123760 270852 123812 270904
rect 177488 270852 177540 270904
rect 407764 270852 407816 270904
rect 440516 270852 440568 270904
rect 449164 270852 449216 270904
rect 490196 270852 490248 270904
rect 492588 270852 492640 270904
rect 571708 270852 571760 270904
rect 134432 270716 134484 270768
rect 185124 270716 185176 270768
rect 321376 270716 321428 270768
rect 327080 270716 327132 270768
rect 414664 270716 414716 270768
rect 450820 270716 450872 270768
rect 480260 270716 480312 270768
rect 486608 270716 486660 270768
rect 486976 270716 487028 270768
rect 564624 270716 564676 270768
rect 567844 270716 567896 270768
rect 597744 270716 597796 270768
rect 121460 270580 121512 270632
rect 168104 270580 168156 270632
rect 403624 270580 403676 270632
rect 433432 270580 433484 270632
rect 453304 270580 453356 270632
rect 487804 270580 487856 270632
rect 489644 270580 489696 270632
rect 568212 270580 568264 270632
rect 78864 270444 78916 270496
rect 132500 270444 132552 270496
rect 133788 270444 133840 270496
rect 136640 270444 136692 270496
rect 137008 270444 137060 270496
rect 84108 270308 84160 270360
rect 137468 270308 137520 270360
rect 137836 270444 137888 270496
rect 183652 270444 183704 270496
rect 185584 270444 185636 270496
rect 194416 270444 194468 270496
rect 200764 270444 200816 270496
rect 201868 270444 201920 270496
rect 206836 270444 206888 270496
rect 235816 270444 235868 270496
rect 278044 270444 278096 270496
rect 283840 270444 283892 270496
rect 400864 270444 400916 270496
rect 441620 270444 441672 270496
rect 456432 270444 456484 270496
rect 520280 270444 520332 270496
rect 523132 270444 523184 270496
rect 532884 270444 532936 270496
rect 186136 270308 186188 270360
rect 199936 270308 199988 270360
rect 230848 270308 230900 270360
rect 232688 270308 232740 270360
rect 248236 270308 248288 270360
rect 283104 270308 283156 270360
rect 284668 270308 284720 270360
rect 355048 270308 355100 270360
rect 376944 270308 376996 270360
rect 380532 270308 380584 270360
rect 404360 270308 404412 270360
rect 409604 270308 409656 270360
rect 454316 270308 454368 270360
rect 458824 270308 458876 270360
rect 524420 270308 524472 270360
rect 525616 270308 525668 270360
rect 619640 270444 619692 270496
rect 533528 270308 533580 270360
rect 626540 270308 626592 270360
rect 111984 270172 112036 270224
rect 168748 270172 168800 270224
rect 184848 270172 184900 270224
rect 219348 270172 219400 270224
rect 244372 270172 244424 270224
rect 262312 270172 262364 270224
rect 334348 270172 334400 270224
rect 346400 270172 346452 270224
rect 372252 270172 372304 270224
rect 397460 270172 397512 270224
rect 398748 270172 398800 270224
rect 412640 270172 412692 270224
rect 415032 270172 415084 270224
rect 460940 270172 460992 270224
rect 461400 270172 461452 270224
rect 527180 270172 527232 270224
rect 528376 270172 528428 270224
rect 623964 270172 624016 270224
rect 89628 270036 89680 270088
rect 153016 270036 153068 270088
rect 176568 270036 176620 270088
rect 211160 270036 211212 270088
rect 212448 270036 212500 270088
rect 239956 270036 240008 270088
rect 241888 270036 241940 270088
rect 260656 270036 260708 270088
rect 266176 270036 266228 270088
rect 277216 270036 277268 270088
rect 345296 270036 345348 270088
rect 358820 270036 358872 270088
rect 366640 270036 366692 270088
rect 393320 270036 393372 270088
rect 394976 270036 395028 270088
rect 408776 270036 408828 270088
rect 412456 270036 412508 270088
rect 458272 270036 458324 270088
rect 463516 270036 463568 270088
rect 530768 270036 530820 270088
rect 530952 270036 531004 270088
rect 533160 270036 533212 270088
rect 85488 269900 85540 269952
rect 149428 269900 149480 269952
rect 152832 269900 152884 269952
rect 157156 269900 157208 269952
rect 173716 269900 173768 269952
rect 212632 269900 212684 269952
rect 226616 269900 226668 269952
rect 249892 269900 249944 269952
rect 256884 269900 256936 269952
rect 268936 269900 268988 269952
rect 330208 269900 330260 269952
rect 340880 269900 340932 269952
rect 341800 269900 341852 269952
rect 357532 269900 357584 269952
rect 359188 269900 359240 269952
rect 382280 269900 382332 269952
rect 383016 269900 383068 269952
rect 411260 269900 411312 269952
rect 419632 269900 419684 269952
rect 468116 269900 468168 269952
rect 468484 269900 468536 269952
rect 538128 270036 538180 270088
rect 538312 270036 538364 270088
rect 630680 270036 630732 270088
rect 533988 269900 534040 269952
rect 537852 269900 537904 269952
rect 538036 269900 538088 269952
rect 70584 269764 70636 269816
rect 79324 269764 79376 269816
rect 80060 269764 80112 269816
rect 146392 269764 146444 269816
rect 158628 269764 158680 269816
rect 201040 269764 201092 269816
rect 201684 269764 201736 269816
rect 232504 269764 232556 269816
rect 237196 269764 237248 269816
rect 257344 269764 257396 269816
rect 258540 269764 258592 269816
rect 272248 269764 272300 269816
rect 273076 269764 273128 269816
rect 282184 269764 282236 269816
rect 326896 269764 326948 269816
rect 335544 269764 335596 269816
rect 336004 269764 336056 269816
rect 349160 269764 349212 269816
rect 351736 269764 351788 269816
rect 371240 269764 371292 269816
rect 376576 269764 376628 269816
rect 407120 269764 407172 269816
rect 417148 269764 417200 269816
rect 465080 269764 465132 269816
rect 466000 269764 466052 269816
rect 530400 269764 530452 269816
rect 122748 269628 122800 269680
rect 176200 269628 176252 269680
rect 183468 269628 183520 269680
rect 205456 269628 205508 269680
rect 392032 269628 392084 269680
rect 401692 269628 401744 269680
rect 404360 269628 404412 269680
rect 423680 269628 423732 269680
rect 423956 269628 424008 269680
rect 451372 269628 451424 269680
rect 453580 269628 453632 269680
rect 509240 269628 509292 269680
rect 538588 269764 538640 269816
rect 538772 269764 538824 269816
rect 542820 269764 542872 269816
rect 543188 269900 543240 269952
rect 640524 269900 640576 269952
rect 637580 269764 637632 269816
rect 129648 269492 129700 269544
rect 181168 269492 181220 269544
rect 204168 269492 204220 269544
rect 223488 269492 223540 269544
rect 401692 269492 401744 269544
rect 416780 269492 416832 269544
rect 424600 269492 424652 269544
rect 475016 269492 475068 269544
rect 495256 269492 495308 269544
rect 532884 269628 532936 269680
rect 616236 269628 616288 269680
rect 509884 269492 509936 269544
rect 596180 269492 596232 269544
rect 126888 269356 126940 269408
rect 178316 269356 178368 269408
rect 408408 269356 408460 269408
rect 426532 269356 426584 269408
rect 441620 269356 441672 269408
rect 458456 269356 458508 269408
rect 470968 269356 471020 269408
rect 143908 269220 143960 269272
rect 191104 269220 191156 269272
rect 282736 269220 282788 269272
rect 288808 269220 288860 269272
rect 474280 269220 474332 269272
rect 538220 269220 538272 269272
rect 538588 269356 538640 269408
rect 575480 269356 575532 269408
rect 540612 269220 540664 269272
rect 540796 269220 540848 269272
rect 543188 269220 543240 269272
rect 543372 269152 543424 269204
rect 546500 269152 546552 269204
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 42156 269016 42208 269068
rect 42892 269016 42944 269068
rect 118608 269016 118660 269068
rect 174544 269016 174596 269068
rect 175096 269016 175148 269068
rect 177672 269016 177724 269068
rect 273260 269016 273312 269068
rect 275560 269016 275612 269068
rect 436560 269016 436612 269068
rect 491668 269016 491720 269068
rect 495808 269016 495860 269068
rect 576860 269016 576912 269068
rect 115756 268880 115808 268932
rect 171232 268880 171284 268932
rect 382372 268880 382424 268932
rect 415492 268880 415544 268932
rect 433708 268880 433760 268932
rect 488540 268880 488592 268932
rect 498292 268880 498344 268932
rect 581000 268880 581052 268932
rect 188896 268812 188948 268864
rect 190460 268812 190512 268864
rect 110328 268744 110380 268796
rect 167920 268744 167972 268796
rect 168288 268744 168340 268796
rect 181996 268744 182048 268796
rect 200580 268744 200632 268796
rect 231308 268744 231360 268796
rect 387340 268744 387392 268796
rect 422300 268744 422352 268796
rect 438676 268744 438728 268796
rect 495440 268744 495492 268796
rect 500776 268744 500828 268796
rect 583760 268744 583812 268796
rect 104992 268608 105044 268660
rect 163780 268608 163832 268660
rect 176936 268608 176988 268660
rect 215116 268608 215168 268660
rect 224224 268608 224276 268660
rect 243268 268608 243320 268660
rect 352564 268608 352616 268660
rect 372620 268608 372672 268660
rect 393320 268608 393372 268660
rect 429200 268608 429252 268660
rect 441160 268608 441212 268660
rect 499580 268608 499632 268660
rect 503260 268608 503312 268660
rect 587900 268608 587952 268660
rect 99288 268472 99340 268524
rect 160468 268472 160520 268524
rect 180708 268472 180760 268524
rect 217600 268472 217652 268524
rect 231676 268472 231728 268524
rect 253204 268472 253256 268524
rect 338488 268472 338540 268524
rect 352104 268472 352156 268524
rect 367468 268472 367520 268524
rect 393504 268472 393556 268524
rect 397276 268472 397328 268524
rect 436100 268472 436152 268524
rect 446128 268472 446180 268524
rect 506480 268472 506532 268524
rect 508228 268472 508280 268524
rect 594800 268472 594852 268524
rect 92388 268336 92440 268388
rect 155500 268336 155552 268388
rect 161572 268336 161624 268388
rect 203524 268336 203576 268388
rect 210700 268336 210752 268388
rect 236644 268336 236696 268388
rect 252652 268336 252704 268388
rect 268108 268336 268160 268388
rect 348792 268336 348844 268388
rect 367100 268336 367152 268388
rect 372436 268336 372488 268388
rect 400496 268336 400548 268388
rect 402244 268336 402296 268388
rect 443092 268336 443144 268388
rect 461860 268336 461912 268388
rect 528560 268336 528612 268388
rect 541348 268336 541400 268388
rect 641720 268336 641772 268388
rect 135628 268200 135680 268252
rect 140136 268200 140188 268252
rect 140688 268200 140740 268252
rect 188620 268200 188672 268252
rect 416228 268200 416280 268252
rect 447140 268200 447192 268252
rect 493324 268200 493376 268252
rect 574100 268200 574152 268252
rect 151728 268064 151780 268116
rect 196072 268064 196124 268116
rect 422300 268064 422352 268116
rect 444380 268064 444432 268116
rect 448428 268064 448480 268116
rect 494060 268064 494112 268116
rect 527180 268064 527232 268116
rect 607404 268064 607456 268116
rect 490840 267928 490892 267980
rect 570052 267928 570104 267980
rect 276480 267724 276532 267776
rect 278044 267724 278096 267776
rect 119344 267656 119396 267708
rect 153476 267656 153528 267708
rect 153844 267656 153896 267708
rect 184480 267656 184532 267708
rect 390652 267656 390704 267708
rect 408408 267656 408460 267708
rect 422944 267656 422996 267708
rect 438124 267656 438176 267708
rect 445300 267656 445352 267708
rect 490564 267656 490616 267708
rect 509884 267656 509936 267708
rect 567844 267656 567896 267708
rect 111708 267520 111760 267572
rect 168564 267520 168616 267572
rect 169024 267520 169076 267572
rect 199384 267520 199436 267572
rect 215944 267520 215996 267572
rect 222568 267520 222620 267572
rect 353392 267520 353444 267572
rect 374460 267520 374512 267572
rect 380716 267520 380768 267572
rect 398748 267520 398800 267572
rect 404728 267520 404780 267572
rect 416228 267520 416280 267572
rect 421288 267520 421340 267572
rect 440884 267520 440936 267572
rect 450268 267520 450320 267572
rect 498844 267520 498896 267572
rect 514852 267520 514904 267572
rect 578884 267520 578936 267572
rect 86224 267384 86276 267436
rect 144736 267384 144788 267436
rect 145564 267384 145616 267436
rect 191932 267384 191984 267436
rect 199568 267384 199620 267436
rect 204352 267384 204404 267436
rect 205456 267384 205508 267436
rect 218428 267384 218480 267436
rect 233884 267384 233936 267436
rect 104808 267248 104860 267300
rect 164608 267248 164660 267300
rect 186964 267248 187016 267300
rect 219256 267248 219308 267300
rect 223488 267248 223540 267300
rect 234160 267248 234212 267300
rect 243544 267384 243596 267436
rect 251548 267384 251600 267436
rect 315304 267384 315356 267436
rect 319168 267384 319220 267436
rect 340972 267384 341024 267436
rect 355324 267384 355376 267436
rect 368296 267384 368348 267436
rect 385684 267384 385736 267436
rect 398104 267384 398156 267436
rect 417424 267384 417476 267436
rect 428740 267384 428792 267436
rect 447784 267384 447836 267436
rect 460204 267384 460256 267436
rect 516784 267384 516836 267436
rect 519820 267384 519872 267436
rect 583024 267384 583076 267436
rect 244096 267248 244148 267300
rect 321928 267248 321980 267300
rect 327724 267248 327776 267300
rect 350908 267248 350960 267300
rect 362224 267248 362276 267300
rect 371608 267248 371660 267300
rect 373264 267248 373316 267300
rect 373448 267248 373500 267300
rect 381544 267248 381596 267300
rect 383200 267248 383252 267300
rect 401692 267248 401744 267300
rect 403072 267248 403124 267300
rect 422300 267248 422352 267300
rect 432880 267248 432932 267300
rect 453304 267248 453356 267300
rect 90364 267112 90416 267164
rect 151360 267112 151412 267164
rect 168104 267112 168156 267164
rect 177028 267112 177080 267164
rect 177672 267112 177724 267164
rect 214288 267112 214340 267164
rect 220084 267112 220136 267164
rect 239128 267112 239180 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 362500 267112 362552 267164
rect 369124 267112 369176 267164
rect 373264 267112 373316 267164
rect 392032 267112 392084 267164
rect 394792 267112 394844 267164
rect 403624 267112 403676 267164
rect 413008 267112 413060 267164
rect 441620 267112 441672 267164
rect 447140 267112 447192 267164
rect 448428 267112 448480 267164
rect 452752 267112 452804 267164
rect 462964 267248 463016 267300
rect 465172 267248 465224 267300
rect 523684 267248 523736 267300
rect 524788 267248 524840 267300
rect 612004 267248 612056 267300
rect 455144 267112 455196 267164
rect 515404 267112 515456 267164
rect 517244 267112 517296 267164
rect 527180 267112 527232 267164
rect 529664 267112 529716 267164
rect 617524 267112 617576 267164
rect 79324 266976 79376 267028
rect 140136 266976 140188 267028
rect 186964 266976 187016 267028
rect 190460 266976 190512 267028
rect 224224 266976 224276 267028
rect 228364 266976 228416 267028
rect 140596 266840 140648 266892
rect 137468 266704 137520 266756
rect 150532 266840 150584 266892
rect 159456 266840 159508 266892
rect 162124 266840 162176 266892
rect 178684 266840 178736 266892
rect 209320 266840 209372 266892
rect 218704 266840 218756 266892
rect 220912 266840 220964 266892
rect 249064 266976 249116 267028
rect 250720 266976 250772 267028
rect 255964 266976 256016 267028
rect 259000 266976 259052 267028
rect 286324 266976 286376 267028
rect 287980 266976 288032 267028
rect 312820 266976 312872 267028
rect 316040 266976 316092 267028
rect 316960 266976 317012 267028
rect 321560 266976 321612 267028
rect 365812 266976 365864 267028
rect 373448 266976 373500 267028
rect 393136 266976 393188 267028
rect 420184 266976 420236 267028
rect 249064 266840 249116 266892
rect 314476 266840 314528 266892
rect 318984 266840 319036 266892
rect 332692 266840 332744 266892
rect 343824 266840 343876 266892
rect 378232 266840 378284 266892
rect 394976 266840 395028 266892
rect 427912 266840 427964 266892
rect 457444 266976 457496 267028
rect 470140 266976 470192 267028
rect 534724 266976 534776 267028
rect 539692 266976 539744 267028
rect 634084 266976 634136 267028
rect 442724 266840 442776 266892
rect 485044 266840 485096 266892
rect 499948 266840 500000 266892
rect 507860 266840 507912 266892
rect 534724 266840 534776 266892
rect 589924 266840 589976 266892
rect 151084 266704 151136 266756
rect 179512 266704 179564 266756
rect 347504 266704 347556 266756
rect 351184 266704 351236 266756
rect 388168 266704 388220 266756
rect 404360 266704 404412 266756
rect 408040 266704 408092 266756
rect 423956 266704 424008 266756
rect 434536 266704 434588 266756
rect 449164 266704 449216 266756
rect 457720 266704 457772 266756
rect 476764 266704 476816 266756
rect 485044 266704 485096 266756
rect 308680 266636 308732 266688
rect 310520 266636 310572 266688
rect 313648 266636 313700 266688
rect 317420 266636 317472 266688
rect 317788 266636 317840 266688
rect 322940 266636 322992 266688
rect 360016 266636 360068 266688
rect 366364 266636 366416 266688
rect 130384 266568 130436 266620
rect 138112 266568 138164 266620
rect 149612 266568 149664 266620
rect 159640 266568 159692 266620
rect 345112 266568 345164 266620
rect 348424 266568 348476 266620
rect 399760 266568 399812 266620
rect 407764 266568 407816 266620
rect 310336 266500 310388 266552
rect 311900 266500 311952 266552
rect 312360 266500 312412 266552
rect 314660 266500 314712 266552
rect 316132 266500 316184 266552
rect 320180 266500 320232 266552
rect 327724 266500 327776 266552
rect 331864 266500 331916 266552
rect 350080 266500 350132 266552
rect 353944 266500 353996 266552
rect 355876 266500 355928 266552
rect 360844 266500 360896 266552
rect 369952 266500 370004 266552
rect 372252 266500 372304 266552
rect 374920 266500 374972 266552
rect 380532 266500 380584 266552
rect 132500 266432 132552 266484
rect 147220 266432 147272 266484
rect 342628 266432 342680 266484
rect 345296 266432 345348 266484
rect 407212 266432 407264 266484
rect 414664 266568 414716 266620
rect 437848 266568 437900 266620
rect 447140 266568 447192 266620
rect 490012 266704 490064 266756
rect 509700 266704 509752 266756
rect 510712 266704 510764 266756
rect 511816 266704 511868 266756
rect 512368 266704 512420 266756
rect 513196 266704 513248 266756
rect 516508 266704 516560 266756
rect 517428 266704 517480 266756
rect 518992 266704 519044 266756
rect 520096 266704 520148 266756
rect 527272 266704 527324 266756
rect 528192 266704 528244 266756
rect 528928 266704 528980 266756
rect 529848 266704 529900 266756
rect 531412 266704 531464 266756
rect 532516 266704 532568 266756
rect 533068 266704 533120 266756
rect 533988 266704 534040 266756
rect 535552 266704 535604 266756
rect 536748 266704 536800 266756
rect 543004 266704 543056 266756
rect 598204 266704 598256 266756
rect 501604 266568 501656 266620
rect 504824 266568 504876 266620
rect 556804 266568 556856 266620
rect 423772 266500 423824 266552
rect 425704 266500 425756 266552
rect 426256 266500 426308 266552
rect 428464 266500 428516 266552
rect 447784 266500 447836 266552
rect 456064 266500 456116 266552
rect 491668 266432 491720 266484
rect 492588 266432 492640 266484
rect 494152 266432 494204 266484
rect 495072 266432 495124 266484
rect 502432 266432 502484 266484
rect 503444 266432 503496 266484
rect 504088 266432 504140 266484
rect 505008 266432 505060 266484
rect 506572 266432 506624 266484
rect 507676 266432 507728 266484
rect 507860 266432 507912 266484
rect 549904 266432 549956 266484
rect 163504 266364 163556 266416
rect 167092 266364 167144 266416
rect 168564 266364 168616 266416
rect 169576 266364 169628 266416
rect 211160 266364 211212 266416
rect 213460 266364 213512 266416
rect 214564 266364 214616 266416
rect 215944 266364 215996 266416
rect 239404 266364 239456 266416
rect 241612 266364 241664 266416
rect 243728 266364 243780 266416
rect 246580 266364 246632 266416
rect 250444 266364 250496 266416
rect 256516 266364 256568 266416
rect 300952 266364 301004 266416
rect 302056 266364 302108 266416
rect 303712 266364 303764 266416
rect 304540 266364 304592 266416
rect 307852 266364 307904 266416
rect 309140 266364 309192 266416
rect 309508 266364 309560 266416
rect 310704 266364 310756 266416
rect 311164 266364 311216 266416
rect 313280 266364 313332 266416
rect 320272 266364 320324 266416
rect 321376 266364 321428 266416
rect 324412 266364 324464 266416
rect 325332 266364 325384 266416
rect 328552 266364 328604 266416
rect 329748 266364 329800 266416
rect 336832 266364 336884 266416
rect 337936 266364 337988 266416
rect 346768 266364 346820 266416
rect 347688 266364 347740 266416
rect 349252 266364 349304 266416
rect 350356 266364 350408 266416
rect 357532 266364 357584 266416
rect 359464 266364 359516 266416
rect 361672 266364 361724 266416
rect 362776 266364 362828 266416
rect 369124 266364 369176 266416
rect 370504 266364 370556 266416
rect 374092 266364 374144 266416
rect 375288 266364 375340 266416
rect 379888 266364 379940 266416
rect 383016 266364 383068 266416
rect 384028 266364 384080 266416
rect 384948 266364 385000 266416
rect 386512 266364 386564 266416
rect 387708 266364 387760 266416
rect 392308 266364 392360 266416
rect 393320 266364 393372 266416
rect 398932 266364 398984 266416
rect 400036 266364 400088 266416
rect 408868 266364 408920 266416
rect 409788 266364 409840 266416
rect 411352 266364 411404 266416
rect 412272 266364 412324 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 417976 266364 418028 266416
rect 418804 266364 418856 266416
rect 425428 266364 425480 266416
rect 427084 266364 427136 266416
rect 429568 266364 429620 266416
rect 430396 266364 430448 266416
rect 432052 266364 432104 266416
rect 433156 266364 433208 266416
rect 440332 266364 440384 266416
rect 441344 266364 441396 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 444472 266364 444524 266416
rect 445668 266364 445720 266416
rect 448612 266364 448664 266416
rect 450544 266364 450596 266416
rect 454408 266364 454460 266416
rect 455328 266364 455380 266416
rect 473452 266364 473504 266416
rect 474648 266364 474700 266416
rect 475108 266364 475160 266416
rect 479524 266364 479576 266416
rect 481732 266364 481784 266416
rect 482836 266364 482888 266416
rect 483388 266364 483440 266416
rect 484216 266364 484268 266416
rect 485872 266364 485924 266416
rect 486792 266364 486844 266416
rect 487160 266296 487212 266348
rect 557724 266296 557776 266348
rect 484216 266160 484268 266212
rect 560668 266160 560720 266212
rect 482560 266024 482612 266076
rect 487160 266024 487212 266076
rect 492496 266024 492548 266076
rect 572720 266024 572772 266076
rect 513196 265888 513248 265940
rect 601700 265888 601752 265940
rect 515680 265752 515732 265804
rect 605840 265752 605892 265804
rect 209780 265616 209832 265668
rect 210700 265616 210752 265668
rect 224960 265616 225012 265668
rect 225604 265616 225656 265668
rect 280344 265616 280396 265668
rect 280988 265616 281040 265668
rect 520648 265616 520700 265668
rect 612740 265616 612792 265668
rect 479248 265480 479300 265532
rect 553400 265480 553452 265532
rect 477592 265344 477644 265396
rect 550640 265344 550692 265396
rect 469312 265208 469364 265260
rect 539968 265208 540020 265260
rect 466828 265072 466880 265124
rect 535736 265072 535788 265124
rect 64144 264460 64196 264512
rect 668952 264460 669004 264512
rect 61384 264324 61436 264376
rect 668124 264324 668176 264376
rect 55864 264188 55916 264240
rect 667940 264188 667992 264240
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 563704 259428 563756 259480
rect 675852 258680 675904 258732
rect 676404 258680 676456 258732
rect 35808 256776 35860 256828
rect 40500 256776 40552 256828
rect 553952 256708 554004 256760
rect 560944 256708 560996 256760
rect 35808 255552 35860 255604
rect 554504 255552 554556 255604
rect 558184 255552 558236 255604
rect 39580 255484 39632 255536
rect 35624 255280 35676 255332
rect 39856 255280 39908 255332
rect 35808 254056 35860 254108
rect 40224 254056 40276 254108
rect 35808 252696 35860 252748
rect 41328 252696 41380 252748
rect 35624 252560 35676 252612
rect 41696 252560 41748 252612
rect 554412 252560 554464 252612
rect 562324 252560 562376 252612
rect 35808 251200 35860 251252
rect 37924 251200 37976 251252
rect 554136 251200 554188 251252
rect 556804 251200 556856 251252
rect 35808 249908 35860 249960
rect 39764 249908 39816 249960
rect 674840 249704 674892 249756
rect 675484 249704 675536 249756
rect 675024 247936 675076 247988
rect 675392 247800 675444 247852
rect 35808 247052 35860 247104
rect 41696 247052 41748 247104
rect 559564 246304 559616 246356
rect 647240 246304 647292 246356
rect 671620 245964 671672 246016
rect 672172 245964 672224 246016
rect 553860 245624 553912 245676
rect 596824 245624 596876 245676
rect 674840 245352 674892 245404
rect 675208 245352 675260 245404
rect 553492 244264 553544 244316
rect 555424 244264 555476 244316
rect 37924 242700 37976 242752
rect 41696 242700 41748 242752
rect 42064 242632 42116 242684
rect 42708 242632 42760 242684
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553676 241476 553728 241528
rect 629944 241476 629996 241528
rect 554504 240116 554556 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 672172 236988 672224 237040
rect 671252 236852 671304 236904
rect 553768 236784 553820 236836
rect 559564 236784 559616 236836
rect 672954 236716 673006 236768
rect 671712 236512 671764 236564
rect 673184 236444 673236 236496
rect 672172 236172 672224 236224
rect 673092 236172 673144 236224
rect 671068 235900 671120 235952
rect 673414 235832 673466 235884
rect 672908 235696 672960 235748
rect 673368 234948 673420 235000
rect 673184 234812 673236 234864
rect 673460 234812 673512 234864
rect 669688 234608 669740 234660
rect 674088 234676 674140 234728
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 670240 234472 670292 234524
rect 671436 234200 671488 234252
rect 674088 234200 674140 234252
rect 652208 233860 652260 233912
rect 670884 233860 670936 233912
rect 675852 233860 675904 233912
rect 678244 233860 678296 233912
rect 672080 233248 672132 233300
rect 673184 233248 673236 233300
rect 673460 233180 673512 233232
rect 673966 233180 674018 233232
rect 670056 232976 670108 233028
rect 673000 232976 673052 233028
rect 670884 232840 670936 232892
rect 672908 232840 672960 232892
rect 663064 232636 663116 232688
rect 674380 232636 674432 232688
rect 675852 232636 675904 232688
rect 683212 232636 683264 232688
rect 660304 232500 660356 232552
rect 674564 232500 674616 232552
rect 676036 232500 676088 232552
rect 683396 232500 683448 232552
rect 156420 231548 156472 231600
rect 162676 231548 162728 231600
rect 135168 231412 135220 231464
rect 137652 231412 137704 231464
rect 155132 231412 155184 231464
rect 156972 231412 157024 231464
rect 157248 231412 157300 231464
rect 161756 231412 161808 231464
rect 662512 231412 662564 231464
rect 674840 231412 674892 231464
rect 46204 231276 46256 231328
rect 668400 231276 668452 231328
rect 92388 231140 92440 231192
rect 170772 231140 170824 231192
rect 665088 231140 665140 231192
rect 128268 231004 128320 231056
rect 195888 231004 195940 231056
rect 673184 230936 673236 230988
rect 118608 230868 118660 230920
rect 188160 230868 188212 230920
rect 674840 230800 674892 230852
rect 94504 230732 94556 230784
rect 171416 230732 171468 230784
rect 104808 230596 104860 230648
rect 179144 230596 179196 230648
rect 194416 230596 194468 230648
rect 196900 230596 196952 230648
rect 665272 230596 665324 230648
rect 439320 230528 439372 230580
rect 137652 230460 137704 230512
rect 201040 230460 201092 230512
rect 42432 230392 42484 230444
rect 43260 230392 43312 230444
rect 133788 230392 133840 230444
rect 137468 230392 137520 230444
rect 213092 230392 213144 230444
rect 261576 230392 261628 230444
rect 311992 230392 312044 230444
rect 313096 230392 313148 230444
rect 374644 230392 374696 230444
rect 376208 230392 376260 230444
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 451556 230392 451608 230444
rect 453304 230392 453356 230444
rect 476120 230392 476172 230444
rect 478604 230392 478656 230444
rect 387432 230324 387484 230376
rect 388444 230324 388496 230376
rect 398104 230324 398156 230376
rect 399392 230324 399444 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 470876 230324 470928 230376
rect 471888 230324 471940 230376
rect 493416 230324 493468 230376
rect 496360 230324 496412 230376
rect 497280 230324 497332 230376
rect 498108 230324 498160 230376
rect 510804 230324 510856 230376
rect 511908 230324 511960 230376
rect 521108 230324 521160 230376
rect 526444 230324 526496 230376
rect 530124 230324 530176 230376
rect 531136 230324 531188 230376
rect 126888 230256 126940 230308
rect 194416 230256 194468 230308
rect 194876 230256 194928 230308
rect 195428 230256 195480 230308
rect 195612 230256 195664 230308
rect 204904 230256 204956 230308
rect 206560 230256 206612 230308
rect 256424 230256 256476 230308
rect 256608 230256 256660 230308
rect 297640 230256 297692 230308
rect 297824 230256 297876 230308
rect 323400 230256 323452 230308
rect 452844 230188 452896 230240
rect 454316 230188 454368 230240
rect 468300 230188 468352 230240
rect 469128 230188 469180 230240
rect 487620 230188 487672 230240
rect 488448 230188 488500 230240
rect 95240 230120 95292 230172
rect 157616 230120 157668 230172
rect 157800 230120 157852 230172
rect 158536 230120 158588 230172
rect 162492 230120 162544 230172
rect 185584 230120 185636 230172
rect 186044 230120 186096 230172
rect 235816 230120 235868 230172
rect 240324 230120 240376 230172
rect 282184 230120 282236 230172
rect 282644 230120 282696 230172
rect 307944 230120 307996 230172
rect 308128 230120 308180 230172
rect 334992 230120 335044 230172
rect 335176 230120 335228 230172
rect 350448 230120 350500 230172
rect 444472 230120 444524 230172
rect 447692 230120 447744 230172
rect 454132 230052 454184 230104
rect 455328 230052 455380 230104
rect 82084 229984 82136 230036
rect 86224 229984 86276 230036
rect 137284 229984 137336 230036
rect 137468 229984 137520 230036
rect 156788 229984 156840 230036
rect 157432 229984 157484 230036
rect 195060 229984 195112 230036
rect 195428 229984 195480 230036
rect 215208 229984 215260 230036
rect 230480 229984 230532 230036
rect 277032 229984 277084 230036
rect 277216 229984 277268 230036
rect 302792 229984 302844 230036
rect 303252 229984 303304 230036
rect 329840 229984 329892 230036
rect 330944 229984 330996 230036
rect 355600 229984 355652 230036
rect 484400 229984 484452 230036
rect 495164 230188 495216 230240
rect 511448 230188 511500 230240
rect 517520 230188 517572 230240
rect 530768 230188 530820 230240
rect 539600 230392 539652 230444
rect 533528 230256 533580 230308
rect 538312 230256 538364 230308
rect 674676 230256 674728 230308
rect 673460 230188 673512 230240
rect 532700 230120 532752 230172
rect 547144 230120 547196 230172
rect 491484 230052 491536 230104
rect 492496 230052 492548 230104
rect 560944 230052 560996 230104
rect 568120 230052 568172 230104
rect 517244 229984 517296 230036
rect 524604 229984 524656 230036
rect 528836 229984 528888 230036
rect 533528 229984 533580 230036
rect 534632 229984 534684 230036
rect 549260 229984 549312 230036
rect 453488 229916 453540 229968
rect 455788 229916 455840 229968
rect 674452 229916 674504 229968
rect 151452 229848 151504 229900
rect 151636 229848 151688 229900
rect 157248 229848 157300 229900
rect 162308 229848 162360 229900
rect 166264 229848 166316 229900
rect 68284 229712 68336 229764
rect 144460 229712 144512 229764
rect 144828 229712 144880 229764
rect 146300 229712 146352 229764
rect 137284 229576 137336 229628
rect 156788 229712 156840 229764
rect 148140 229576 148192 229628
rect 150808 229576 150860 229628
rect 150992 229576 151044 229628
rect 153384 229576 153436 229628
rect 154396 229576 154448 229628
rect 162124 229712 162176 229764
rect 163964 229712 164016 229764
rect 225512 229848 225564 229900
rect 225696 229848 225748 229900
rect 271880 229848 271932 229900
rect 275652 229848 275704 229900
rect 311992 229848 312044 229900
rect 312636 229848 312688 229900
rect 340144 229848 340196 229900
rect 345664 229848 345716 229900
rect 360752 229848 360804 229900
rect 361212 229848 361264 229900
rect 378784 229848 378836 229900
rect 410892 229848 410944 229900
rect 417424 229848 417476 229900
rect 449624 229848 449676 229900
rect 450544 229848 450596 229900
rect 467012 229848 467064 229900
rect 474004 229848 474056 229900
rect 476672 229848 476724 229900
rect 481640 229848 481692 229900
rect 481824 229848 481876 229900
rect 493692 229848 493744 229900
rect 495992 229848 496044 229900
rect 506388 229848 506440 229900
rect 507584 229848 507636 229900
rect 516784 229848 516836 229900
rect 519176 229848 519228 229900
rect 528560 229848 528612 229900
rect 536564 229848 536616 229900
rect 559564 229848 559616 229900
rect 668584 229848 668636 229900
rect 672724 229848 672776 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 674334 229780 674386 229832
rect 173900 229712 173952 229764
rect 175924 229712 175976 229764
rect 176384 229712 176436 229764
rect 185400 229712 185452 229764
rect 185584 229712 185636 229764
rect 194876 229712 194928 229764
rect 195060 229712 195112 229764
rect 202328 229712 202380 229764
rect 204904 229712 204956 229764
rect 246120 229712 246172 229764
rect 246488 229712 246540 229764
rect 287336 229712 287388 229764
rect 287704 229712 287756 229764
rect 318248 229712 318300 229764
rect 157984 229576 158036 229628
rect 160744 229576 160796 229628
rect 160928 229576 160980 229628
rect 220360 229576 220412 229628
rect 102140 229440 102192 229492
rect 145656 229440 145708 229492
rect 146024 229372 146076 229424
rect 210056 229440 210108 229492
rect 220084 229440 220136 229492
rect 251272 229576 251324 229628
rect 251732 229576 251784 229628
rect 292488 229576 292540 229628
rect 318064 229576 318116 229628
rect 345296 229712 345348 229764
rect 351736 229712 351788 229764
rect 371056 229712 371108 229764
rect 377680 229712 377732 229764
rect 389088 229712 389140 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 457352 229712 457404 229764
rect 463884 229712 463936 229764
rect 465448 229712 465500 229764
rect 467472 229712 467524 229764
rect 469588 229712 469640 229764
rect 476764 229712 476816 229764
rect 479248 229712 479300 229764
rect 489920 229712 489972 229764
rect 492128 229712 492180 229764
rect 507124 229712 507176 229764
rect 523040 229712 523092 229764
rect 534816 229712 534868 229764
rect 538496 229712 538548 229764
rect 566832 229712 566884 229764
rect 662328 229712 662380 229764
rect 673184 229712 673236 229764
rect 509516 229644 509568 229696
rect 515496 229644 515548 229696
rect 388628 229576 388680 229628
rect 398748 229576 398800 229628
rect 526904 229576 526956 229628
rect 536104 229576 536156 229628
rect 672816 229576 672868 229628
rect 448980 229508 449032 229560
rect 451924 229508 451976 229560
rect 660948 229440 661000 229492
rect 662512 229440 662564 229492
rect 446404 229372 446456 229424
rect 448980 229372 449032 229424
rect 505652 229372 505704 229424
rect 510620 229372 510672 229424
rect 673276 229372 673328 229424
rect 110328 229304 110380 229356
rect 145840 229304 145892 229356
rect 151452 229304 151504 229356
rect 155960 229304 156012 229356
rect 123484 229168 123536 229220
rect 148140 229168 148192 229220
rect 148324 229168 148376 229220
rect 154028 229168 154080 229220
rect 154212 229168 154264 229220
rect 157800 229304 157852 229356
rect 157984 229304 158036 229356
rect 163688 229304 163740 229356
rect 166816 229304 166868 229356
rect 169116 229304 169168 229356
rect 170956 229304 171008 229356
rect 230664 229304 230716 229356
rect 413836 229304 413888 229356
rect 420000 229304 420052 229356
rect 443828 229304 443880 229356
rect 444840 229304 444892 229356
rect 472164 229304 472216 229356
rect 472992 229304 473044 229356
rect 450268 229236 450320 229288
rect 451740 229236 451792 229288
rect 495348 229236 495400 229288
rect 500224 229236 500276 229288
rect 513380 229236 513432 229288
rect 519084 229236 519136 229288
rect 162124 229168 162176 229220
rect 173900 229168 173952 229220
rect 106188 229032 106240 229084
rect 175924 229168 175976 229220
rect 180432 229168 180484 229220
rect 183376 229168 183428 229220
rect 240968 229168 241020 229220
rect 423496 229100 423548 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 450912 229100 450964 229152
rect 452752 229100 452804 229152
rect 503720 229100 503772 229152
rect 509884 229100 509936 229152
rect 515312 229100 515364 229152
rect 520924 229100 520976 229152
rect 524972 229100 525024 229152
rect 529940 229100 529992 229152
rect 179788 229032 179840 229084
rect 180064 229032 180116 229084
rect 185584 229032 185636 229084
rect 189724 229032 189776 229084
rect 100668 228896 100720 228948
rect 174636 228896 174688 228948
rect 93584 228760 93636 228812
rect 159364 228760 159416 228812
rect 162676 228760 162728 228812
rect 184848 228896 184900 228948
rect 185216 228896 185268 228948
rect 190092 228896 190144 228948
rect 192484 229032 192536 229084
rect 200396 229032 200448 229084
rect 201408 229032 201460 229084
rect 252560 229032 252612 229084
rect 257528 229032 257580 229084
rect 296352 229032 296404 229084
rect 305552 229032 305604 229084
rect 315672 229032 315724 229084
rect 326896 229032 326948 229084
rect 351092 229032 351144 229084
rect 195244 228896 195296 228948
rect 195428 228896 195480 228948
rect 246764 228896 246816 228948
rect 176108 228760 176160 228812
rect 231308 228760 231360 228812
rect 246304 228760 246356 228812
rect 253848 228896 253900 228948
rect 255228 228896 255280 228948
rect 295708 228896 295760 228948
rect 302148 228896 302200 228948
rect 331220 228896 331272 228948
rect 506388 228896 506440 228948
rect 512736 228896 512788 228948
rect 526444 228896 526496 228948
rect 544292 228896 544344 228948
rect 248236 228760 248288 228812
rect 291844 228760 291896 228812
rect 67548 228624 67600 228676
rect 146208 228624 146260 228676
rect 61384 228488 61436 228540
rect 57244 228352 57296 228404
rect 136824 228352 136876 228404
rect 137376 228488 137428 228540
rect 162308 228624 162360 228676
rect 162492 228624 162544 228676
rect 166816 228624 166868 228676
rect 166954 228624 167006 228676
rect 185400 228624 185452 228676
rect 185584 228624 185636 228676
rect 226156 228624 226208 228676
rect 226340 228624 226392 228676
rect 272524 228624 272576 228676
rect 291660 228624 291712 228676
rect 300216 228760 300268 228812
rect 300676 228760 300728 228812
rect 330484 228760 330536 228812
rect 376024 228760 376076 228812
rect 387800 228760 387852 228812
rect 478880 228760 478932 228812
rect 490380 228760 490432 228812
rect 499856 228760 499908 228812
rect 518164 228760 518216 228812
rect 518532 228760 518584 228812
rect 541624 228760 541676 228812
rect 296628 228624 296680 228676
rect 329196 228624 329248 228676
rect 336464 228624 336516 228676
rect 358820 228624 358872 228676
rect 359924 228624 359976 228676
rect 376852 228624 376904 228676
rect 485688 228624 485740 228676
rect 498292 228624 498344 228676
rect 498568 228624 498620 228676
rect 515772 228624 515824 228676
rect 517888 228624 517940 228676
rect 539416 228624 539468 228676
rect 539600 228624 539652 228676
rect 557172 228624 557224 228676
rect 147128 228488 147180 228540
rect 200396 228488 200448 228540
rect 204904 228488 204956 228540
rect 221004 228488 221056 228540
rect 112996 228216 113048 228268
rect 137192 228216 137244 228268
rect 139308 228352 139360 228404
rect 143080 228216 143132 228268
rect 143448 228216 143500 228268
rect 146024 228216 146076 228268
rect 146208 228216 146260 228268
rect 148876 228216 148928 228268
rect 153016 228352 153068 228404
rect 215852 228352 215904 228404
rect 216496 228352 216548 228404
rect 264796 228488 264848 228540
rect 272524 228488 272576 228540
rect 309876 228488 309928 228540
rect 313924 228488 313976 228540
rect 320824 228488 320876 228540
rect 325424 228488 325476 228540
rect 349160 228488 349212 228540
rect 350448 228488 350500 228540
rect 369124 228488 369176 228540
rect 371056 228488 371108 228540
rect 385224 228488 385276 228540
rect 386052 228488 386104 228540
rect 397460 228488 397512 228540
rect 224684 228352 224736 228404
rect 273812 228352 273864 228404
rect 285496 228352 285548 228404
rect 318892 228352 318944 228404
rect 330484 228352 330536 228404
rect 354956 228352 355008 228404
rect 355324 228352 355376 228404
rect 372988 228352 373040 228404
rect 373448 228352 373500 228404
rect 387156 228352 387208 228404
rect 390008 228352 390060 228404
rect 400036 228352 400088 228404
rect 205548 228216 205600 228268
rect 205916 228216 205968 228268
rect 257068 228216 257120 228268
rect 268936 228216 268988 228268
rect 306012 228216 306064 228268
rect 407764 228488 407816 228540
rect 409788 228488 409840 228540
rect 415492 228488 415544 228540
rect 485044 228488 485096 228540
rect 498660 228488 498712 228540
rect 502432 228488 502484 228540
rect 521108 228488 521160 228540
rect 527548 228488 527600 228540
rect 553216 228488 553268 228540
rect 556804 228488 556856 228540
rect 570604 228488 570656 228540
rect 402796 228352 402848 228404
rect 411628 228352 411680 228404
rect 474464 228352 474516 228404
rect 484492 228352 484544 228404
rect 490196 228352 490248 228404
rect 505192 228352 505244 228404
rect 512092 228352 512144 228404
rect 532976 228352 533028 228404
rect 537208 228352 537260 228404
rect 565636 228352 565688 228404
rect 673552 228352 673604 228404
rect 539416 228216 539468 228268
rect 540796 228216 540848 228268
rect 119988 228080 120040 228132
rect 185216 228080 185268 228132
rect 185400 228080 185452 228132
rect 126704 227944 126756 227996
rect 195244 228080 195296 228132
rect 239036 228080 239088 228132
rect 400128 228080 400180 228132
rect 415032 228012 415084 228064
rect 421932 228012 421984 228064
rect 88248 227808 88300 227860
rect 95240 227808 95292 227860
rect 133512 227808 133564 227860
rect 136640 227808 136692 227860
rect 136824 227808 136876 227860
rect 141148 227808 141200 227860
rect 141516 227808 141568 227860
rect 192484 227808 192536 227860
rect 195060 227808 195112 227860
rect 200396 227944 200448 227996
rect 210700 227944 210752 227996
rect 204904 227808 204956 227860
rect 205456 227808 205508 227860
rect 205916 227808 205968 227860
rect 210332 227808 210384 227860
rect 238392 227944 238444 227996
rect 238668 227944 238720 227996
rect 282828 227944 282880 227996
rect 416688 227876 416740 227928
rect 420644 227876 420696 227928
rect 447048 227876 447100 227928
rect 450544 227876 450596 227928
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 420644 227740 420696 227792
rect 423864 227740 423916 227792
rect 471520 227740 471572 227792
rect 479524 227740 479576 227792
rect 64788 227672 64840 227724
rect 110328 227672 110380 227724
rect 110512 227672 110564 227724
rect 182364 227672 182416 227724
rect 60648 227536 60700 227588
rect 102140 227536 102192 227588
rect 103428 227536 103480 227588
rect 175188 227536 175240 227588
rect 181536 227536 181588 227588
rect 185216 227672 185268 227724
rect 185400 227672 185452 227724
rect 192668 227672 192720 227724
rect 195244 227672 195296 227724
rect 214748 227672 214800 227724
rect 214932 227672 214984 227724
rect 262220 227672 262272 227724
rect 277032 227672 277084 227724
rect 311808 227672 311860 227724
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 184112 227536 184164 227588
rect 187516 227536 187568 227588
rect 189908 227536 189960 227588
rect 205088 227536 205140 227588
rect 205272 227536 205324 227588
rect 251916 227536 251968 227588
rect 259276 227536 259328 227588
rect 298284 227536 298336 227588
rect 301504 227536 301556 227588
rect 308588 227536 308640 227588
rect 524604 227536 524656 227588
rect 539968 227536 540020 227588
rect 96436 227400 96488 227452
rect 170772 227400 170824 227452
rect 171094 227400 171146 227452
rect 175924 227468 175976 227520
rect 185584 227400 185636 227452
rect 185768 227400 185820 227452
rect 223580 227400 223632 227452
rect 224224 227400 224276 227452
rect 241612 227400 241664 227452
rect 257896 227400 257948 227452
rect 299572 227400 299624 227452
rect 304908 227400 304960 227452
rect 333704 227400 333756 227452
rect 333888 227400 333940 227452
rect 356244 227400 356296 227452
rect 357072 227400 357124 227452
rect 374276 227400 374328 227452
rect 514024 227400 514076 227452
rect 535736 227400 535788 227452
rect 538312 227400 538364 227452
rect 556068 227400 556120 227452
rect 89628 227264 89680 227316
rect 157294 227264 157346 227316
rect 157524 227264 157576 227316
rect 176752 227264 176804 227316
rect 222476 227264 222528 227316
rect 63316 227128 63368 227180
rect 144828 227128 144880 227180
rect 150072 227128 150124 227180
rect 213276 227128 213328 227180
rect 214380 227128 214432 227180
rect 233884 227264 233936 227316
rect 235816 227264 235868 227316
rect 280252 227264 280304 227316
rect 306196 227264 306248 227316
rect 336924 227264 336976 227316
rect 340696 227264 340748 227316
rect 361396 227264 361448 227316
rect 382096 227264 382148 227316
rect 392952 227264 393004 227316
rect 224040 227128 224092 227180
rect 262864 227128 262916 227180
rect 263508 227128 263560 227180
rect 277216 227128 277268 227180
rect 281356 227128 281408 227180
rect 317604 227128 317656 227180
rect 322848 227128 322900 227180
rect 349804 227128 349856 227180
rect 355876 227128 355928 227180
rect 375564 227128 375616 227180
rect 376668 227128 376720 227180
rect 389732 227128 389784 227180
rect 393136 227128 393188 227180
rect 402612 227264 402664 227316
rect 494704 227264 494756 227316
rect 402244 227128 402296 227180
rect 408408 227128 408460 227180
rect 478604 227128 478656 227180
rect 486792 227128 486844 227180
rect 489552 227128 489604 227180
rect 504180 227128 504232 227180
rect 56508 226992 56560 227044
rect 142436 226992 142488 227044
rect 143264 226992 143316 227044
rect 204076 226992 204128 227044
rect 117228 226856 117280 226908
rect 184112 226856 184164 226908
rect 185584 226856 185636 226908
rect 205088 226856 205140 226908
rect 214380 226856 214432 226908
rect 215116 226992 215168 227044
rect 224224 226992 224276 227044
rect 218428 226856 218480 226908
rect 222476 226856 222528 226908
rect 228732 226856 228784 226908
rect 122748 226720 122800 226772
rect 185400 226720 185452 226772
rect 186136 226720 186188 226772
rect 195244 226720 195296 226772
rect 200028 226720 200080 226772
rect 205272 226720 205324 226772
rect 129556 226584 129608 226636
rect 197360 226584 197412 226636
rect 204076 226584 204128 226636
rect 208124 226584 208176 226636
rect 136548 226448 136600 226500
rect 141608 226448 141660 226500
rect 142252 226448 142304 226500
rect 202972 226448 203024 226500
rect 203524 226448 203576 226500
rect 222936 226720 222988 226772
rect 223120 226720 223172 226772
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 301504 226992 301556 227044
rect 310428 226992 310480 227044
rect 338212 226992 338264 227044
rect 338672 226992 338724 227044
rect 360108 226992 360160 227044
rect 362776 226992 362828 227044
rect 379428 226992 379480 227044
rect 391848 226992 391900 227044
rect 403532 226992 403584 227044
rect 412548 226992 412600 227044
rect 419356 226992 419408 227044
rect 486976 226992 487028 227044
rect 500960 226992 501012 227044
rect 212172 226584 212224 226636
rect 214932 226584 214984 226636
rect 219348 226584 219400 226636
rect 267372 226856 267424 226908
rect 293776 226856 293828 226908
rect 324964 226856 325016 226908
rect 510620 227264 510672 227316
rect 524420 227264 524472 227316
rect 526260 227264 526312 227316
rect 551560 227264 551612 227316
rect 506204 227128 506256 227180
rect 525984 227128 526036 227180
rect 533344 227128 533396 227180
rect 560944 227128 560996 227180
rect 505008 226992 505060 227044
rect 523040 226992 523092 227044
rect 523684 226992 523736 227044
rect 548708 226992 548760 227044
rect 555424 226992 555476 227044
rect 633716 226992 633768 227044
rect 510988 226856 511040 226908
rect 672448 226856 672500 226908
rect 673092 226856 673144 226908
rect 231032 226720 231084 226772
rect 243268 226720 243320 226772
rect 249616 226720 249668 226772
rect 290556 226720 290608 226772
rect 243452 226652 243504 226704
rect 248696 226652 248748 226704
rect 264152 226516 264204 226568
rect 269304 226516 269356 226568
rect 673276 226516 673328 226568
rect 213828 226448 213880 226500
rect 224040 226448 224092 226500
rect 351092 226448 351144 226500
rect 353024 226448 353076 226500
rect 403992 226448 404044 226500
rect 412272 226448 412324 226500
rect 474740 226448 474792 226500
rect 482744 226448 482796 226500
rect 141792 226380 141844 226432
rect 142114 226380 142166 226432
rect 271144 226380 271196 226432
rect 279608 226380 279660 226432
rect 672724 226380 672776 226432
rect 350264 226312 350316 226364
rect 351736 226312 351788 226364
rect 388536 226312 388588 226364
rect 391664 226312 391716 226364
rect 407764 226312 407816 226364
rect 408684 226312 408736 226364
rect 481640 226312 481692 226364
rect 487804 226312 487856 226364
rect 663524 226312 663576 226364
rect 665272 226312 665324 226364
rect 122564 226244 122616 226296
rect 193956 226244 194008 226296
rect 194140 226244 194192 226296
rect 244188 226244 244240 226296
rect 267004 226244 267056 226296
rect 274456 226244 274508 226296
rect 286324 226244 286376 226296
rect 289912 226244 289964 226296
rect 291016 226244 291068 226296
rect 322112 226244 322164 226296
rect 458640 226244 458692 226296
rect 462964 226244 463016 226296
rect 127624 226108 127676 226160
rect 142114 226108 142166 226160
rect 142252 226108 142304 226160
rect 209412 226108 209464 226160
rect 209688 226108 209740 226160
rect 259644 226108 259696 226160
rect 261852 226108 261904 226160
rect 300860 226108 300912 226160
rect 309048 226108 309100 226160
rect 336280 226108 336332 226160
rect 528560 226108 528612 226160
rect 542636 226108 542688 226160
rect 672604 226108 672656 226160
rect 66168 225972 66220 226024
rect 142620 225972 142672 226024
rect 142804 225972 142856 226024
rect 147588 225972 147640 226024
rect 147772 225972 147824 226024
rect 83464 225836 83516 225888
rect 156420 225836 156472 225888
rect 157340 225972 157392 226024
rect 217140 225972 217192 226024
rect 222016 225972 222068 226024
rect 269948 225972 270000 226024
rect 278412 225972 278464 226024
rect 313280 225972 313332 226024
rect 329748 225972 329800 226024
rect 353668 225972 353720 226024
rect 354588 225972 354640 226024
rect 372344 225972 372396 226024
rect 498108 225972 498160 226024
rect 514300 225972 514352 226024
rect 516600 225972 516652 226024
rect 538680 225972 538732 226024
rect 672494 225904 672546 225956
rect 183652 225836 183704 225888
rect 76564 225700 76616 225752
rect 184296 225700 184348 225752
rect 198004 225836 198056 225888
rect 204720 225700 204772 225752
rect 205088 225836 205140 225888
rect 236460 225836 236512 225888
rect 237288 225836 237340 225888
rect 240324 225836 240376 225888
rect 252468 225836 252520 225888
rect 293132 225836 293184 225888
rect 296444 225836 296496 225888
rect 327540 225836 327592 225888
rect 332232 225836 332284 225888
rect 357532 225836 357584 225888
rect 373816 225836 373868 225888
rect 377680 225836 377732 225888
rect 377864 225836 377916 225888
rect 390376 225836 390428 225888
rect 394332 225836 394384 225888
rect 403256 225836 403308 225888
rect 483756 225836 483808 225888
rect 497280 225836 497332 225888
rect 501144 225836 501196 225888
rect 519268 225836 519320 225888
rect 521752 225836 521804 225888
rect 545764 225836 545816 225888
rect 558184 225836 558236 225888
rect 571340 225836 571392 225888
rect 249340 225700 249392 225752
rect 255044 225700 255096 225752
rect 296996 225700 297048 225752
rect 315672 225700 315724 225752
rect 344652 225700 344704 225752
rect 352932 225700 352984 225752
rect 371608 225700 371660 225752
rect 371792 225700 371844 225752
rect 382740 225700 382792 225752
rect 382924 225700 382976 225752
rect 396172 225700 396224 225752
rect 488908 225700 488960 225752
rect 503628 225700 503680 225752
rect 508872 225700 508924 225752
rect 529204 225700 529256 225752
rect 535920 225700 535972 225752
rect 563980 225700 564032 225752
rect 672380 225700 672432 225752
rect 156604 225632 156656 225684
rect 671896 225632 671948 225684
rect 72424 225564 72476 225616
rect 142114 225564 142166 225616
rect 142252 225564 142304 225616
rect 147680 225564 147732 225616
rect 157340 225564 157392 225616
rect 214564 225564 214616 225616
rect 215208 225564 215260 225616
rect 266084 225564 266136 225616
rect 270040 225564 270092 225616
rect 282644 225564 282696 225616
rect 284116 225564 284168 225616
rect 320180 225564 320232 225616
rect 321376 225564 321428 225616
rect 346584 225564 346636 225616
rect 347044 225564 347096 225616
rect 367836 225564 367888 225616
rect 372528 225564 372580 225616
rect 387432 225564 387484 225616
rect 390192 225564 390244 225616
rect 401968 225564 402020 225616
rect 410984 225564 411036 225616
rect 416136 225564 416188 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 488816 225564 488868 225616
rect 494060 225564 494112 225616
rect 509516 225564 509568 225616
rect 510160 225564 510212 225616
rect 530952 225564 531004 225616
rect 531412 225564 531464 225616
rect 558276 225564 558328 225616
rect 110144 225428 110196 225480
rect 127624 225428 127676 225480
rect 125232 225292 125284 225344
rect 196164 225428 196216 225480
rect 196348 225428 196400 225480
rect 129372 225292 129424 225344
rect 199108 225292 199160 225344
rect 204720 225428 204772 225480
rect 212540 225428 212592 225480
rect 205088 225292 205140 225344
rect 208124 225292 208176 225344
rect 257712 225428 257764 225480
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 241152 225292 241204 225344
rect 286692 225292 286744 225344
rect 135076 225156 135128 225208
rect 204260 225156 204312 225208
rect 242716 225156 242768 225208
rect 285036 225156 285088 225208
rect 557632 225088 557684 225140
rect 561956 225088 562008 225140
rect 132408 225020 132460 225072
rect 201684 225020 201736 225072
rect 202696 225020 202748 225072
rect 254492 225020 254544 225072
rect 297272 225020 297324 225072
rect 305368 225020 305420 225072
rect 327724 224952 327776 225004
rect 332048 224952 332100 225004
rect 369124 224952 369176 225004
rect 373632 224952 373684 225004
rect 404176 224952 404228 225004
rect 410616 224952 410668 225004
rect 416504 224952 416556 225004
rect 422208 224952 422260 225004
rect 493692 224952 493744 225004
rect 494704 224952 494756 225004
rect 495164 224952 495216 225004
rect 567016 225020 567068 225072
rect 569132 225020 569184 225072
rect 672156 225292 672208 225344
rect 672034 225224 672086 225276
rect 563704 224952 563756 225004
rect 666468 225020 666520 225072
rect 96252 224884 96304 224936
rect 172980 224884 173032 224936
rect 102048 224748 102100 224800
rect 178500 224884 178552 224936
rect 178684 224884 178736 224936
rect 185584 224884 185636 224936
rect 185768 224884 185820 224936
rect 195244 224884 195296 224936
rect 195428 224884 195480 224936
rect 242900 224884 242952 224936
rect 274272 224884 274324 224936
rect 312452 224884 312504 224936
rect 460572 224884 460624 224936
rect 463148 224884 463200 224936
rect 630864 224952 630916 225004
rect 568856 224884 568908 224936
rect 178040 224748 178092 224800
rect 204536 224748 204588 224800
rect 204720 224748 204772 224800
rect 237748 224748 237800 224800
rect 245292 224748 245344 224800
rect 287980 224748 288032 224800
rect 319996 224748 320048 224800
rect 345940 224748 345992 224800
rect 462504 224748 462556 224800
rect 469312 224748 469364 224800
rect 506940 224748 506992 224800
rect 526720 224748 526772 224800
rect 529940 224748 529992 224800
rect 548064 224748 548116 224800
rect 548248 224748 548300 224800
rect 85488 224612 85540 224664
rect 165620 224612 165672 224664
rect 174912 224612 174964 224664
rect 178684 224612 178736 224664
rect 179328 224612 179380 224664
rect 185400 224612 185452 224664
rect 185584 224612 185636 224664
rect 235172 224612 235224 224664
rect 251088 224612 251140 224664
rect 294420 224612 294472 224664
rect 299296 224612 299348 224664
rect 331772 224612 331824 224664
rect 335176 224612 335228 224664
rect 356888 224612 356940 224664
rect 363604 224612 363656 224664
rect 368480 224612 368532 224664
rect 520464 224612 520516 224664
rect 544108 224612 544160 224664
rect 544292 224612 544344 224664
rect 545028 224612 545080 224664
rect 549260 224748 549312 224800
rect 557632 224748 557684 224800
rect 557816 224748 557868 224800
rect 562140 224748 562192 224800
rect 562324 224748 562376 224800
rect 567016 224748 567068 224800
rect 567200 224748 567252 224800
rect 572444 224884 572496 224936
rect 569224 224748 569276 224800
rect 571340 224748 571392 224800
rect 571708 224748 571760 224800
rect 616052 224748 616104 224800
rect 671820 224748 671872 224800
rect 79968 224476 80020 224528
rect 160468 224476 160520 224528
rect 161664 224476 161716 224528
rect 224868 224476 224920 224528
rect 228732 224476 228784 224528
rect 274916 224476 274968 224528
rect 275100 224476 275152 224528
rect 311164 224476 311216 224528
rect 311532 224476 311584 224528
rect 338856 224476 338908 224528
rect 346216 224476 346268 224528
rect 366548 224476 366600 224528
rect 387708 224476 387760 224528
rect 397828 224476 397880 224528
rect 456064 224476 456116 224528
rect 459744 224476 459796 224528
rect 491300 224476 491352 224528
rect 506020 224476 506072 224528
rect 515956 224476 516008 224528
rect 538864 224476 538916 224528
rect 539968 224476 540020 224528
rect 542452 224476 542504 224528
rect 542820 224476 542872 224528
rect 550640 224612 550692 224664
rect 550778 224612 550830 224664
rect 625252 224612 625304 224664
rect 666836 224612 666888 224664
rect 73712 224340 73764 224392
rect 88984 224340 89036 224392
rect 89444 224340 89496 224392
rect 167828 224340 167880 224392
rect 168288 224340 168340 224392
rect 230020 224340 230072 224392
rect 233148 224340 233200 224392
rect 277676 224340 277728 224392
rect 286692 224340 286744 224392
rect 319536 224340 319588 224392
rect 319812 224340 319864 224392
rect 347228 224340 347280 224392
rect 361212 224340 361264 224392
rect 377496 224340 377548 224392
rect 379244 224340 379296 224392
rect 393596 224340 393648 224392
rect 480536 224340 480588 224392
rect 492772 224340 492824 224392
rect 499212 224340 499264 224392
rect 516784 224340 516836 224392
rect 525616 224340 525668 224392
rect 548248 224340 548300 224392
rect 623780 224476 623832 224528
rect 667756 224408 667808 224460
rect 426440 224272 426492 224324
rect 426992 224272 427044 224324
rect 558000 224340 558052 224392
rect 625436 224340 625488 224392
rect 68928 224068 68980 224120
rect 151636 224204 151688 224256
rect 151774 224204 151826 224256
rect 155316 224204 155368 224256
rect 157248 224204 157300 224256
rect 160928 224204 160980 224256
rect 165160 224204 165212 224256
rect 227444 224204 227496 224256
rect 231676 224204 231728 224256
rect 278964 224204 279016 224256
rect 290832 224204 290884 224256
rect 323676 224204 323728 224256
rect 323952 224204 324004 224256
rect 334992 224204 335044 224256
rect 339408 224204 339460 224256
rect 88984 224068 89036 224120
rect 142114 224068 142166 224120
rect 142252 224068 142304 224120
rect 194600 224068 194652 224120
rect 195244 224068 195296 224120
rect 204628 224068 204680 224120
rect 255780 224068 255832 224120
rect 266176 224068 266228 224120
rect 303436 224068 303488 224120
rect 358084 224204 358136 224256
rect 363328 224204 363380 224256
rect 366732 224204 366784 224256
rect 381636 224204 381688 224256
rect 394516 224204 394568 224256
rect 404544 224204 404596 224256
rect 405556 224204 405608 224256
rect 414204 224204 414256 224256
rect 427912 224204 427964 224256
rect 428740 224204 428792 224256
rect 447508 224204 447560 224256
rect 448060 224204 448112 224256
rect 470232 224204 470284 224256
rect 480444 224204 480496 224256
rect 486608 224204 486660 224256
rect 500040 224204 500092 224256
rect 504456 224204 504508 224256
rect 523500 224204 523552 224256
rect 535276 224204 535328 224256
rect 557540 224136 557592 224188
rect 571708 224136 571760 224188
rect 572444 224136 572496 224188
rect 628748 224136 628800 224188
rect 362316 224068 362368 224120
rect 377404 224068 377456 224120
rect 385868 224068 385920 224120
rect 519084 224068 519136 224120
rect 535000 224068 535052 224120
rect 671482 224068 671534 224120
rect 105912 223932 105964 223984
rect 181076 223932 181128 223984
rect 201224 223932 201276 223984
rect 543004 224000 543056 224052
rect 543188 224000 543240 224052
rect 622676 224000 622728 224052
rect 205088 223932 205140 223984
rect 250628 223932 250680 223984
rect 667756 223932 667808 223984
rect 279424 223864 279476 223916
rect 284760 223864 284812 223916
rect 524420 223864 524472 223916
rect 525064 223864 525116 223916
rect 619640 223864 619692 223916
rect 108672 223796 108724 223848
rect 183836 223796 183888 223848
rect 112812 223660 112864 223712
rect 185952 223796 186004 223848
rect 186964 223796 187016 223848
rect 217784 223796 217836 223848
rect 224592 223796 224644 223848
rect 270592 223796 270644 223848
rect 667020 223796 667072 223848
rect 509516 223728 509568 223780
rect 510160 223728 510212 223780
rect 542820 223728 542872 223780
rect 543004 223728 543056 223780
rect 621572 223728 621624 223780
rect 184848 223660 184900 223712
rect 195428 223660 195480 223712
rect 195888 223660 195940 223712
rect 205088 223660 205140 223712
rect 238024 223660 238076 223712
rect 266728 223660 266780 223712
rect 505192 223592 505244 223644
rect 614948 223592 615000 223644
rect 669596 223592 669648 223644
rect 81348 223524 81400 223576
rect 153200 223524 153252 223576
rect 75828 223388 75880 223440
rect 154948 223524 155000 223576
rect 155776 223524 155828 223576
rect 159824 223524 159876 223576
rect 165620 223524 165672 223576
rect 171968 223524 172020 223576
rect 175280 223524 175332 223576
rect 176568 223524 176620 223576
rect 154212 223388 154264 223440
rect 156788 223388 156840 223440
rect 158720 223388 158772 223440
rect 181720 223388 181772 223440
rect 69572 223252 69624 223304
rect 142114 223252 142166 223304
rect 66904 223116 66956 223168
rect 146668 223252 146720 223304
rect 146944 223252 146996 223304
rect 152096 223252 152148 223304
rect 153200 223252 153252 223304
rect 155776 223252 155828 223304
rect 156420 223252 156472 223304
rect 161940 223252 161992 223304
rect 162492 223252 162544 223304
rect 186596 223524 186648 223576
rect 187332 223524 187384 223576
rect 242256 223524 242308 223576
rect 250904 223524 250956 223576
rect 291200 223524 291252 223576
rect 297916 223524 297968 223576
rect 303252 223524 303304 223576
rect 307668 223524 307720 223576
rect 335636 223524 335688 223576
rect 406752 223524 406804 223576
rect 414848 223524 414900 223576
rect 454868 223524 454920 223576
rect 460480 223524 460532 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 184664 223388 184716 223440
rect 239680 223388 239732 223440
rect 244096 223388 244148 223440
rect 286048 223388 286100 223440
rect 304724 223388 304776 223440
rect 308128 223388 308180 223440
rect 312912 223388 312964 223440
rect 342076 223456 342128 223508
rect 342812 223388 342864 223440
rect 347872 223388 347924 223440
rect 517520 223388 517572 223440
rect 531504 223388 531556 223440
rect 534816 223388 534868 223440
rect 547420 223388 547472 223440
rect 669274 223388 669326 223440
rect 336004 223320 336056 223372
rect 342260 223320 342312 223372
rect 185400 223252 185452 223304
rect 142436 223116 142488 223168
rect 144000 223116 144052 223168
rect 146576 223116 146628 223168
rect 171600 223116 171652 223168
rect 171784 223116 171836 223168
rect 185584 223116 185636 223168
rect 188896 223252 188948 223304
rect 245108 223252 245160 223304
rect 246856 223252 246908 223304
rect 288624 223252 288676 223304
rect 289728 223252 289780 223304
rect 297732 223252 297784 223304
rect 299112 223252 299164 223304
rect 328552 223252 328604 223304
rect 347228 223252 347280 223304
rect 357900 223252 357952 223304
rect 483112 223252 483164 223304
rect 496084 223252 496136 223304
rect 503352 223252 503404 223304
rect 192024 223116 192076 223168
rect 194324 223116 194376 223168
rect 199752 223116 199804 223168
rect 204260 223116 204312 223168
rect 211988 223116 212040 223168
rect 215392 223116 215444 223168
rect 216220 223116 216272 223168
rect 241336 223116 241388 223168
rect 283472 223116 283524 223168
rect 288256 223116 288308 223168
rect 321100 223116 321152 223168
rect 344652 223116 344704 223168
rect 364616 223116 364668 223168
rect 365536 223116 365588 223168
rect 379612 223116 379664 223168
rect 380072 223116 380124 223168
rect 386512 223116 386564 223168
rect 488632 223116 488684 223168
rect 502708 223116 502760 223168
rect 508228 223116 508280 223168
rect 514668 223252 514720 223304
rect 535460 223252 535512 223304
rect 561956 223252 562008 223304
rect 567844 223252 567896 223304
rect 586980 223252 587032 223304
rect 593972 223252 594024 223304
rect 71412 222980 71464 223032
rect 146944 222980 146996 223032
rect 147128 222980 147180 223032
rect 162124 222980 162176 223032
rect 162308 222980 162360 223032
rect 219716 222980 219768 223032
rect 230204 222980 230256 223032
rect 275468 222980 275520 223032
rect 278596 222980 278648 223032
rect 315028 222980 315080 223032
rect 316684 222980 316736 223032
rect 327264 222980 327316 223032
rect 328092 222980 328144 223032
rect 351460 222980 351512 223032
rect 353944 222980 353996 223032
rect 365904 222980 365956 223032
rect 366916 222980 366968 223032
rect 383844 222980 383896 223032
rect 384212 222980 384264 223032
rect 393964 222980 394016 223032
rect 493048 222980 493100 223032
rect 508596 222980 508648 223032
rect 521752 223116 521804 223168
rect 532056 223116 532108 223168
rect 559012 223116 559064 223168
rect 562324 223116 562376 223168
rect 587164 223116 587216 223168
rect 667756 223116 667808 223168
rect 527824 222980 527876 223032
rect 529480 222980 529532 223032
rect 555700 222980 555752 223032
rect 557540 222980 557592 223032
rect 559840 222980 559892 223032
rect 627092 222980 627144 223032
rect 62764 222844 62816 222896
rect 141976 222844 142028 222896
rect 142160 222844 142212 222896
rect 156604 222844 156656 222896
rect 156788 222844 156840 222896
rect 215392 222844 215444 222896
rect 215944 222844 215996 222896
rect 233332 222844 233384 222896
rect 234528 222844 234580 222896
rect 281540 222844 281592 222896
rect 282460 222844 282512 222896
rect 316316 222844 316368 222896
rect 324136 222844 324188 222896
rect 348516 222844 348568 222896
rect 349068 222844 349120 222896
rect 367192 222844 367244 222896
rect 368388 222844 368440 222896
rect 382372 222844 382424 222896
rect 383476 222844 383528 222896
rect 394884 222844 394936 222896
rect 395804 222844 395856 222896
rect 406476 222844 406528 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 479892 222844 479944 222896
rect 491944 222844 491996 222896
rect 500776 222844 500828 222896
rect 517520 222844 517572 222896
rect 519820 222844 519872 222896
rect 543372 222844 543424 222896
rect 554044 222844 554096 222896
rect 632704 222844 632756 222896
rect 651288 222844 651340 222896
rect 666468 222844 666520 222896
rect 78588 222708 78640 222760
rect 155132 222708 155184 222760
rect 155684 222708 155736 222760
rect 161940 222708 161992 222760
rect 162124 222708 162176 222760
rect 171784 222708 171836 222760
rect 171968 222708 172020 222760
rect 185400 222708 185452 222760
rect 185584 222708 185636 222760
rect 204260 222708 204312 222760
rect 204444 222708 204496 222760
rect 247408 222708 247460 222760
rect 264796 222708 264848 222760
rect 304356 222708 304408 222760
rect 543832 222708 543884 222760
rect 552388 222708 552440 222760
rect 625620 222708 625672 222760
rect 99288 222572 99340 222624
rect 87972 222436 88024 222488
rect 164976 222436 165028 222488
rect 171600 222572 171652 222624
rect 175280 222572 175332 222624
rect 197176 222572 197228 222624
rect 249984 222572 250036 222624
rect 529848 222572 529900 222624
rect 619916 222572 619968 222624
rect 176016 222504 176068 222556
rect 175648 222436 175700 222488
rect 207480 222436 207532 222488
rect 207664 222436 207716 222488
rect 258356 222436 258408 222488
rect 175832 222368 175884 222420
rect 85304 222300 85356 222352
rect 156420 222300 156472 222352
rect 194324 222300 194376 222352
rect 194508 222300 194560 222352
rect 204444 222300 204496 222352
rect 211804 222300 211856 222352
rect 228088 222300 228140 222352
rect 287888 222300 287940 222352
rect 295064 222300 295116 222352
rect 484492 222300 484544 222352
rect 562324 222436 562376 222488
rect 567844 222436 567896 222488
rect 627920 222436 627972 222488
rect 489920 222300 489972 222352
rect 491116 222300 491168 222352
rect 629852 222300 629904 222352
rect 156604 222232 156656 222284
rect 191012 222164 191064 222216
rect 482744 222164 482796 222216
rect 586980 222164 587032 222216
rect 587164 222164 587216 222216
rect 631508 222164 631560 222216
rect 97908 222096 97960 222148
rect 104348 222096 104400 222148
rect 106372 222096 106424 222148
rect 157432 222096 157484 222148
rect 172704 222096 172756 222148
rect 174084 222096 174136 222148
rect 94688 221960 94740 222012
rect 157616 221960 157668 222012
rect 104348 221824 104400 221876
rect 158352 221960 158404 222012
rect 166816 221960 166868 222012
rect 167000 221960 167052 222012
rect 169760 221960 169812 222012
rect 171784 221960 171836 222012
rect 181260 222096 181312 222148
rect 182640 222096 182692 222148
rect 191472 222096 191524 222148
rect 247592 222096 247644 222148
rect 258080 222096 258132 222148
rect 263692 222096 263744 222148
rect 270224 222096 270276 222148
rect 306380 222096 306432 222148
rect 310704 222096 310756 222148
rect 312636 222096 312688 222148
rect 331404 222096 331456 222148
rect 353760 222096 353812 222148
rect 424968 222096 425020 222148
rect 429292 222096 429344 222148
rect 452568 222096 452620 222148
rect 455604 222096 455656 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 495164 222028 495216 222080
rect 497740 222028 497792 222080
rect 515496 222028 515548 222080
rect 529848 222028 529900 222080
rect 533988 222028 534040 222080
rect 559380 222028 559432 222080
rect 559564 222028 559616 222080
rect 564808 222028 564860 222080
rect 158168 221824 158220 221876
rect 176568 221824 176620 221876
rect 231860 221960 231912 222012
rect 233700 221960 233752 222012
rect 277952 221960 278004 222012
rect 280068 221960 280120 222012
rect 313740 221960 313792 222012
rect 318248 221960 318300 222012
rect 343824 221960 343876 222012
rect 367652 221960 367704 222012
rect 380256 221960 380308 222012
rect 536104 221892 536156 221944
rect 543694 221892 543746 221944
rect 547144 221892 547196 221944
rect 556988 221892 557040 221944
rect 181260 221824 181312 221876
rect 181628 221824 181680 221876
rect 240140 221824 240192 221876
rect 263324 221824 263376 221876
rect 301228 221824 301280 221876
rect 301964 221824 302016 221876
rect 310888 221824 310940 221876
rect 313188 221824 313240 221876
rect 340420 221824 340472 221876
rect 351276 221824 351328 221876
rect 369308 221824 369360 221876
rect 509884 221824 509936 221876
rect 522580 221824 522632 221876
rect 546960 221824 547012 221876
rect 557356 221824 557408 221876
rect 562324 221892 562376 221944
rect 600596 221960 600648 222012
rect 600964 221960 601016 222012
rect 606668 221960 606720 222012
rect 80520 221688 80572 221740
rect 86224 221688 86276 221740
rect 91284 221688 91336 221740
rect 167184 221688 167236 221740
rect 167460 221688 167512 221740
rect 171416 221688 171468 221740
rect 171600 221688 171652 221740
rect 232228 221688 232280 221740
rect 239312 221688 239364 221740
rect 283656 221688 283708 221740
rect 303252 221688 303304 221740
rect 332784 221688 332836 221740
rect 357164 221688 357216 221740
rect 374644 221688 374696 221740
rect 391020 221688 391072 221740
rect 400404 221688 400456 221740
rect 475936 221688 475988 221740
rect 486148 221688 486200 221740
rect 496268 221688 496320 221740
rect 513564 221688 513616 221740
rect 524236 221688 524288 221740
rect 544292 221688 544344 221740
rect 596824 221824 596876 221876
rect 633440 221824 633492 221876
rect 562692 221688 562744 221740
rect 608600 221688 608652 221740
rect 73896 221552 73948 221604
rect 82084 221552 82136 221604
rect 86316 221552 86368 221604
rect 160836 221552 160888 221604
rect 162124 221552 162176 221604
rect 202512 221552 202564 221604
rect 59360 221416 59412 221468
rect 140780 221416 140832 221468
rect 140964 221416 141016 221468
rect 205732 221552 205784 221604
rect 208400 221552 208452 221604
rect 260840 221552 260892 221604
rect 261024 221552 261076 221604
rect 301780 221552 301832 221604
rect 308864 221552 308916 221604
rect 339684 221552 339736 221604
rect 341340 221552 341392 221604
rect 361764 221552 361816 221604
rect 369492 221552 369544 221604
rect 384028 221552 384080 221604
rect 384396 221552 384448 221604
rect 395160 221552 395212 221604
rect 400588 221552 400640 221604
rect 405832 221552 405884 221604
rect 480812 221552 480864 221604
rect 492956 221552 493008 221604
rect 497464 221552 497516 221604
rect 515128 221552 515180 221604
rect 522856 221552 522908 221604
rect 104532 221280 104584 221332
rect 106372 221280 106424 221332
rect 111156 221280 111208 221332
rect 171784 221280 171836 221332
rect 171968 221280 172020 221332
rect 226524 221416 226576 221468
rect 227904 221416 227956 221468
rect 276112 221416 276164 221468
rect 292488 221416 292540 221468
rect 326252 221416 326304 221468
rect 342168 221416 342220 221468
rect 364800 221416 364852 221468
rect 375288 221416 375340 221468
rect 390744 221416 390796 221468
rect 396816 221416 396868 221468
rect 407304 221416 407356 221468
rect 408408 221416 408460 221468
rect 416872 221416 416924 221468
rect 468944 221416 468996 221468
rect 476212 221416 476264 221468
rect 483756 221416 483808 221468
rect 533620 221552 533672 221604
rect 601792 221552 601844 221604
rect 204168 221280 204220 221332
rect 252744 221280 252796 221332
rect 266820 221280 266872 221332
rect 303804 221280 303856 221332
rect 525984 221280 526036 221332
rect 533160 221280 533212 221332
rect 546592 221416 546644 221468
rect 546960 221416 547012 221468
rect 549076 221416 549128 221468
rect 549260 221416 549312 221468
rect 600964 221416 601016 221468
rect 538312 221280 538364 221332
rect 538496 221212 538548 221264
rect 604828 221212 604880 221264
rect 138480 221144 138532 221196
rect 162124 221144 162176 221196
rect 162308 221144 162360 221196
rect 221280 221144 221332 221196
rect 222752 221144 222804 221196
rect 268292 221144 268344 221196
rect 523500 221076 523552 221128
rect 601976 221076 602028 221128
rect 124404 221008 124456 221060
rect 193404 221008 193456 221060
rect 202512 221008 202564 221060
rect 206376 221008 206428 221060
rect 219808 221008 219860 221060
rect 263048 221008 263100 221060
rect 521108 220940 521160 220992
rect 600412 220940 600464 220992
rect 600596 220940 600648 220992
rect 604644 220940 604696 220992
rect 83004 220872 83056 220924
rect 142114 220872 142166 220924
rect 142252 220872 142304 220924
rect 148324 220872 148376 220924
rect 148508 220872 148560 220924
rect 151176 220872 151228 220924
rect 158352 220872 158404 220924
rect 160652 220872 160704 220924
rect 160836 220872 160888 220924
rect 164332 220872 164384 220924
rect 164516 220872 164568 220924
rect 222292 220872 222344 220924
rect 282644 220872 282696 220924
rect 287704 220872 287756 220924
rect 456708 220872 456760 220924
rect 253848 220804 253900 220856
rect 258632 220804 258684 220856
rect 418344 220804 418396 220856
rect 424048 220804 424100 220856
rect 466092 220872 466144 220924
rect 471428 220872 471480 220924
rect 462136 220804 462188 220856
rect 517520 220804 517572 220856
rect 518532 220804 518584 220856
rect 600688 220804 600740 220856
rect 114284 220736 114336 220788
rect 146760 220736 146812 220788
rect 146944 220736 146996 220788
rect 180754 220736 180806 220788
rect 181260 220736 181312 220788
rect 190276 220736 190328 220788
rect 190414 220736 190466 220788
rect 236644 220736 236696 220788
rect 242624 220736 242676 220788
rect 246488 220736 246540 220788
rect 260196 220736 260248 220788
rect 298560 220736 298612 220788
rect 321560 220736 321612 220788
rect 324504 220736 324556 220788
rect 385224 220736 385276 220788
rect 388720 220736 388772 220788
rect 414204 220736 414256 220788
rect 418160 220736 418212 220788
rect 455328 220736 455380 220788
rect 458824 220736 458876 220788
rect 465724 220736 465776 220788
rect 469588 220736 469640 220788
rect 474004 220736 474056 220788
rect 475384 220736 475436 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 511816 220736 511868 220788
rect 101220 220600 101272 220652
rect 175464 220600 175516 220652
rect 177396 220600 177448 220652
rect 180800 220600 180852 220652
rect 181076 220600 181128 220652
rect 224224 220600 224276 220652
rect 253572 220600 253624 220652
rect 293316 220600 293368 220652
rect 302424 220600 302476 220652
rect 334072 220600 334124 220652
rect 357900 220600 357952 220652
rect 374460 220600 374512 220652
rect 500224 220600 500276 220652
rect 511816 220600 511868 220652
rect 69756 220464 69808 220516
rect 136916 220464 136968 220516
rect 137100 220464 137152 220516
rect 146944 220464 146996 220516
rect 147588 220464 147640 220516
rect 150716 220464 150768 220516
rect 150900 220464 150952 220516
rect 73068 220328 73120 220380
rect 142114 220328 142166 220380
rect 142252 220328 142304 220380
rect 144644 220328 144696 220380
rect 146760 220328 146812 220380
rect 151636 220328 151688 220380
rect 151912 220464 151964 220516
rect 211344 220464 211396 220516
rect 214104 220464 214156 220516
rect 214288 220464 214340 220516
rect 218704 220464 218756 220516
rect 223672 220464 223724 220516
rect 265164 220464 265216 220516
rect 267648 220464 267700 220516
rect 306840 220464 306892 220516
rect 338028 220464 338080 220516
rect 359004 220464 359056 220516
rect 469128 220464 469180 220516
rect 474556 220464 474608 220516
rect 488448 220464 488500 220516
rect 501880 220464 501932 220516
rect 520924 220600 520976 220652
rect 537484 220600 537536 220652
rect 531688 220464 531740 220516
rect 535736 220464 535788 220516
rect 538496 220668 538548 220720
rect 538864 220668 538916 220720
rect 544292 220668 544344 220720
rect 550640 220600 550692 220652
rect 554228 220600 554280 220652
rect 555700 220600 555752 220652
rect 608876 220600 608928 220652
rect 213644 220328 213696 220380
rect 79692 220192 79744 220244
rect 151728 220192 151780 220244
rect 151912 220192 151964 220244
rect 154028 220192 154080 220244
rect 156328 220192 156380 220244
rect 158904 220192 158956 220244
rect 164148 220192 164200 220244
rect 223856 220192 223908 220244
rect 224408 220328 224460 220380
rect 267924 220328 267976 220380
rect 273444 220328 273496 220380
rect 309232 220328 309284 220380
rect 314844 220328 314896 220380
rect 341064 220328 341116 220380
rect 342996 220328 343048 220380
rect 363420 220328 363472 220380
rect 472992 220328 473044 220380
rect 481180 220328 481232 220380
rect 496452 220328 496504 220380
rect 509332 220328 509384 220380
rect 516968 220328 517020 220380
rect 527548 220328 527600 220380
rect 531136 220328 531188 220380
rect 556528 220464 556580 220516
rect 558276 220464 558328 220516
rect 561772 220464 561824 220516
rect 561956 220464 562008 220516
rect 234160 220192 234212 220244
rect 237012 220192 237064 220244
rect 280436 220192 280488 220244
rect 283380 220192 283432 220244
rect 316316 220192 316368 220244
rect 316500 220192 316552 220244
rect 342628 220192 342680 220244
rect 348792 220192 348844 220244
rect 369952 220192 370004 220244
rect 370504 220192 370556 220244
rect 381084 220192 381136 220244
rect 388720 220192 388772 220244
rect 400956 220192 401008 220244
rect 430120 220192 430172 220244
rect 432052 220192 432104 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 473176 220192 473228 220244
rect 482008 220192 482060 220244
rect 482928 220192 482980 220244
rect 495256 220192 495308 220244
rect 501328 220192 501380 220244
rect 520188 220192 520240 220244
rect 528376 220192 528428 220244
rect 554044 220328 554096 220380
rect 554228 220328 554280 220380
rect 562324 220328 562376 220380
rect 563152 220464 563204 220516
rect 609428 220464 609480 220516
rect 566464 220328 566516 220380
rect 566832 220328 566884 220380
rect 567292 220328 567344 220380
rect 568580 220328 568632 220380
rect 569776 220328 569828 220380
rect 572674 220328 572726 220380
rect 610532 220328 610584 220380
rect 569960 220260 570012 220312
rect 548708 220192 548760 220244
rect 154396 220124 154448 220176
rect 156144 220124 156196 220176
rect 572076 220124 572128 220176
rect 611452 220192 611504 220244
rect 648620 220192 648672 220244
rect 652760 220192 652812 220244
rect 76380 220056 76432 220108
rect 152188 220056 152240 220108
rect 152372 220056 152424 220108
rect 153844 220056 153896 220108
rect 157524 220056 157576 220108
rect 214288 220056 214340 220108
rect 107844 219920 107896 219972
rect 114284 219920 114336 219972
rect 114468 219920 114520 219972
rect 121092 219784 121144 219836
rect 127624 219920 127676 219972
rect 190276 219920 190328 219972
rect 190414 219920 190466 219972
rect 213644 219920 213696 219972
rect 137100 219784 137152 219836
rect 127624 219648 127676 219700
rect 131028 219648 131080 219700
rect 197636 219784 197688 219836
rect 197820 219784 197872 219836
rect 244280 220056 244332 220108
rect 244464 220056 244516 220108
rect 288532 220056 288584 220108
rect 288716 220056 288768 220108
rect 322388 220056 322440 220108
rect 325608 220056 325660 220108
rect 352104 220056 352156 220108
rect 358820 220056 358872 220108
rect 378324 220056 378376 220108
rect 379428 220056 379480 220108
rect 392124 220056 392176 220108
rect 395988 220056 396040 220108
rect 404728 220056 404780 220108
rect 421656 220056 421708 220108
rect 426808 220056 426860 220108
rect 431960 220056 432012 220108
rect 434812 220056 434864 220108
rect 478328 220056 478380 220108
rect 489460 220056 489512 220108
rect 492496 220056 492548 220108
rect 506848 220056 506900 220108
rect 513104 220056 513156 220108
rect 534172 220056 534224 220108
rect 538128 220056 538180 220108
rect 561956 220056 562008 220108
rect 562324 219988 562376 220040
rect 607312 219988 607364 220040
rect 214748 219920 214800 219972
rect 254768 219920 254820 219972
rect 294972 219920 295024 219972
rect 325884 219920 325936 219972
rect 70584 219376 70636 219428
rect 93768 219240 93820 219292
rect 94412 219240 94464 219292
rect 109500 219376 109552 219428
rect 110420 219376 110472 219428
rect 117780 219376 117832 219428
rect 118700 219376 118752 219428
rect 123484 219512 123536 219564
rect 120264 219376 120316 219428
rect 123576 219376 123628 219428
rect 129832 219376 129884 219428
rect 130200 219376 130252 219428
rect 131856 219376 131908 219428
rect 132408 219376 132460 219428
rect 136916 219512 136968 219564
rect 142114 219648 142166 219700
rect 137652 219512 137704 219564
rect 203156 219648 203208 219700
rect 144276 219512 144328 219564
rect 208584 219648 208636 219700
rect 210516 219648 210568 219700
rect 259920 219784 259972 219836
rect 527548 219716 527600 219768
rect 548708 219852 548760 219904
rect 548892 219852 548944 219904
rect 598572 219852 598624 219904
rect 540796 219716 540848 219768
rect 606024 219852 606076 219904
rect 217140 219648 217192 219700
rect 223672 219648 223724 219700
rect 203892 219512 203944 219564
rect 214748 219512 214800 219564
rect 220452 219512 220504 219564
rect 224408 219648 224460 219700
rect 227076 219648 227128 219700
rect 272708 219648 272760 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 503628 219580 503680 219632
rect 591856 219580 591908 219632
rect 591994 219580 592046 219632
rect 620100 219716 620152 219768
rect 224224 219512 224276 219564
rect 229284 219512 229336 219564
rect 332692 219512 332744 219564
rect 337200 219512 337252 219564
rect 146760 219376 146812 219428
rect 146944 219376 146996 219428
rect 152372 219376 152424 219428
rect 152556 219376 152608 219428
rect 156236 219376 156288 219428
rect 156420 219376 156472 219428
rect 158996 219376 159048 219428
rect 159180 219376 159232 219428
rect 160008 219376 160060 219428
rect 162400 219376 162452 219428
rect 163320 219376 163372 219428
rect 163964 219376 164016 219428
rect 178040 219376 178092 219428
rect 178224 219376 178276 219428
rect 64604 219104 64656 219156
rect 66904 219104 66956 219156
rect 83832 219104 83884 219156
rect 157984 219104 158036 219156
rect 62304 218968 62356 219020
rect 72424 218968 72476 219020
rect 77208 218968 77260 219020
rect 146944 218968 146996 219020
rect 147128 218968 147180 219020
rect 156420 218968 156472 219020
rect 169116 219240 169168 219292
rect 169576 219240 169628 219292
rect 169944 219240 169996 219292
rect 170956 219240 171008 219292
rect 171416 219240 171468 219292
rect 172244 219240 172296 219292
rect 172428 219240 172480 219292
rect 173164 219240 173216 219292
rect 175740 219240 175792 219292
rect 180708 219376 180760 219428
rect 185860 219376 185912 219428
rect 186504 219376 186556 219428
rect 224408 219376 224460 219428
rect 229560 219376 229612 219428
rect 230480 219376 230532 219428
rect 237840 219376 237892 219428
rect 239312 219376 239364 219428
rect 239496 219376 239548 219428
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 241796 219376 241848 219428
rect 241980 219376 242032 219428
rect 242900 219376 242952 219428
rect 244924 219376 244976 219428
rect 272340 219376 272392 219428
rect 272708 219376 272760 219428
rect 162400 219104 162452 219156
rect 165620 219104 165672 219156
rect 165804 219104 165856 219156
rect 180064 219104 180116 219156
rect 215944 219240 215996 219292
rect 219624 219240 219676 219292
rect 264152 219240 264204 219292
rect 285864 219376 285916 219428
rect 301964 219240 302016 219292
rect 308220 219376 308272 219428
rect 309140 219376 309192 219428
rect 333704 219376 333756 219428
rect 347228 219376 347280 219428
rect 349620 219376 349672 219428
rect 350540 219376 350592 219428
rect 352104 219376 352156 219428
rect 355324 219376 355376 219428
rect 362040 219376 362092 219428
rect 367652 219376 367704 219428
rect 380256 219376 380308 219428
rect 384212 219376 384264 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 501144 219444 501196 219496
rect 596180 219444 596232 219496
rect 313924 219240 313976 219292
rect 320640 219240 320692 219292
rect 342812 219240 342864 219292
rect 419172 219240 419224 219292
rect 422668 219240 422720 219292
rect 548248 219240 548300 219292
rect 189908 219104 189960 219156
rect 190644 219104 190696 219156
rect 197820 219104 197872 219156
rect 208860 219104 208912 219156
rect 209688 219104 209740 219156
rect 218796 219104 218848 219156
rect 219348 219104 219400 219156
rect 224224 219104 224276 219156
rect 253204 219104 253256 219156
rect 265992 219104 266044 219156
rect 59820 218832 59872 218884
rect 139952 218832 140004 218884
rect 140136 218832 140188 218884
rect 162676 218968 162728 219020
rect 203524 218968 203576 219020
rect 206468 218968 206520 219020
rect 253848 218968 253900 219020
rect 259092 218968 259144 219020
rect 291660 218968 291712 219020
rect 295800 219104 295852 219156
rect 296720 219104 296772 219156
rect 314016 219104 314068 219156
rect 336004 219104 336056 219156
rect 343824 219104 343876 219156
rect 353944 219104 353996 219156
rect 542544 219104 542596 219156
rect 543004 219104 543056 219156
rect 548800 219104 548852 219156
rect 557356 219240 557408 219292
rect 560668 219240 560720 219292
rect 572536 219308 572588 219360
rect 572674 219308 572726 219360
rect 591672 219308 591724 219360
rect 591856 219308 591908 219360
rect 597744 219444 597796 219496
rect 598572 219444 598624 219496
rect 607496 219444 607548 219496
rect 297272 218968 297324 219020
rect 307392 218968 307444 219020
rect 332692 218968 332744 219020
rect 337200 218968 337252 219020
rect 345664 218968 345716 219020
rect 347228 218968 347280 219020
rect 363604 218968 363656 219020
rect 368664 218968 368716 219020
rect 377404 218968 377456 219020
rect 156788 218832 156840 218884
rect 158720 218832 158772 218884
rect 158996 218832 159048 218884
rect 171416 218832 171468 218884
rect 171784 218832 171836 218884
rect 179512 218832 179564 218884
rect 182364 218832 182416 218884
rect 189724 218832 189776 218884
rect 192852 218832 192904 218884
rect 58992 218696 59044 218748
rect 145012 218696 145064 218748
rect 146760 218696 146812 218748
rect 183744 218696 183796 218748
rect 192116 218696 192168 218748
rect 195244 218696 195296 218748
rect 198924 218832 198976 218884
rect 200028 218832 200080 218884
rect 200212 218832 200264 218884
rect 241612 218832 241664 218884
rect 241796 218832 241848 218884
rect 244924 218832 244976 218884
rect 249432 218832 249484 218884
rect 251732 218832 251784 218884
rect 252744 218832 252796 218884
rect 287888 218832 287940 218884
rect 291660 218832 291712 218884
rect 243452 218696 243504 218748
rect 251732 218696 251784 218748
rect 286324 218696 286376 218748
rect 300492 218832 300544 218884
rect 327724 218832 327776 218884
rect 340512 218832 340564 218884
rect 358084 218832 358136 218884
rect 363696 218832 363748 218884
rect 370504 218832 370556 218884
rect 376944 218832 376996 218884
rect 382740 218832 382792 218884
rect 383476 218832 383528 218884
rect 386880 218968 386932 219020
rect 398104 218968 398156 219020
rect 537484 218968 537536 219020
rect 543188 218968 543240 219020
rect 388536 218832 388588 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412548 218832 412600 218884
rect 512736 218832 512788 218884
rect 321560 218696 321612 218748
rect 327264 218696 327316 218748
rect 351092 218696 351144 218748
rect 353760 218696 353812 218748
rect 369124 218696 369176 218748
rect 370320 218696 370372 218748
rect 380072 218696 380124 218748
rect 383568 218696 383620 218748
rect 396264 218696 396316 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 429936 218696 429988 218748
rect 432696 218696 432748 218748
rect 482744 218696 482796 218748
rect 485320 218696 485372 218748
rect 513840 218696 513892 218748
rect 113640 218560 113692 218612
rect 162216 218560 162268 218612
rect 162492 218560 162544 218612
rect 171784 218560 171836 218612
rect 171968 218560 172020 218612
rect 176016 218560 176068 218612
rect 179880 218560 179932 218612
rect 210332 218560 210384 218612
rect 100392 218288 100444 218340
rect 142436 218424 142488 218476
rect 142620 218424 142672 218476
rect 143264 218424 143316 218476
rect 145104 218424 145156 218476
rect 145932 218424 145984 218476
rect 148416 218424 148468 218476
rect 148876 218424 148928 218476
rect 149244 218424 149296 218476
rect 150072 218424 150124 218476
rect 153384 218424 153436 218476
rect 186964 218424 187016 218476
rect 188712 218424 188764 218476
rect 193772 218424 193824 218476
rect 195612 218424 195664 218476
rect 198004 218424 198056 218476
rect 198280 218424 198332 218476
rect 220084 218560 220136 218612
rect 225972 218560 226024 218612
rect 267004 218560 267056 218612
rect 272340 218560 272392 218612
rect 279424 218560 279476 218612
rect 116124 218288 116176 218340
rect 117228 218288 117280 218340
rect 119436 218288 119488 218340
rect 119988 218288 120040 218340
rect 121920 218288 121972 218340
rect 122564 218288 122616 218340
rect 126060 218288 126112 218340
rect 126704 218288 126756 218340
rect 127716 218288 127768 218340
rect 128268 218288 128320 218340
rect 128544 218288 128596 218340
rect 129372 218288 129424 218340
rect 129832 218288 129884 218340
rect 132500 218288 132552 218340
rect 132684 218288 132736 218340
rect 133512 218288 133564 218340
rect 135996 218288 136048 218340
rect 136548 218288 136600 218340
rect 136916 218288 136968 218340
rect 139952 218288 140004 218340
rect 140136 218288 140188 218340
rect 170588 218288 170640 218340
rect 170772 218288 170824 218340
rect 176568 218288 176620 218340
rect 179052 218288 179104 218340
rect 196256 218288 196308 218340
rect 198096 218288 198148 218340
rect 204168 218288 204220 218340
rect 204720 218288 204772 218340
rect 207664 218288 207716 218340
rect 209688 218288 209740 218340
rect 212816 218288 212868 218340
rect 213000 218288 213052 218340
rect 224224 218424 224276 218476
rect 224408 218424 224460 218476
rect 231032 218424 231084 218476
rect 216312 218288 216364 218340
rect 238024 218424 238076 218476
rect 232872 218288 232924 218340
rect 271144 218424 271196 218476
rect 279240 218424 279292 218476
rect 305552 218560 305604 218612
rect 398472 218560 398524 218612
rect 407764 218560 407816 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 475568 218560 475620 218612
rect 482836 218560 482888 218612
rect 502708 218560 502760 218612
rect 514024 218560 514076 218612
rect 517704 218696 517756 218748
rect 518164 218696 518216 218748
rect 520004 218696 520056 218748
rect 548248 218832 548300 218884
rect 561680 218968 561732 219020
rect 563014 218968 563066 219020
rect 563152 218968 563204 219020
rect 567660 218968 567712 219020
rect 567844 218968 567896 219020
rect 574560 218968 574612 219020
rect 586980 219104 587032 219156
rect 594800 219104 594852 219156
rect 587164 218968 587216 219020
rect 548800 218832 548852 218884
rect 560484 218832 560536 218884
rect 560668 218832 560720 218884
rect 614120 218832 614172 218884
rect 548616 218696 548668 218748
rect 567844 218696 567896 218748
rect 568304 218696 568356 218748
rect 571708 218696 571760 218748
rect 571892 218696 571944 218748
rect 603080 218696 603132 218748
rect 543188 218560 543240 218612
rect 598848 218560 598900 218612
rect 294144 218424 294196 218476
rect 316684 218424 316736 218476
rect 426624 218424 426676 218476
rect 429568 218424 429620 218476
rect 500040 218424 500092 218476
rect 604460 218560 604512 218612
rect 458180 218356 458232 218408
rect 241612 218288 241664 218340
rect 246304 218288 246356 218340
rect 253204 218288 253256 218340
rect 258080 218288 258132 218340
rect 425796 218288 425848 218340
rect 428464 218288 428516 218340
rect 450728 218288 450780 218340
rect 453856 218288 453908 218340
rect 461308 218288 461360 218340
rect 497004 218288 497056 218340
rect 586980 218288 587032 218340
rect 587164 218288 587216 218340
rect 601240 218424 601292 218476
rect 670240 218424 670292 218476
rect 601056 218288 601108 218340
rect 607128 218288 607180 218340
rect 107016 218220 107068 218272
rect 55680 218152 55732 218204
rect 56508 218152 56560 218204
rect 57428 218152 57480 218204
rect 61384 218152 61436 218204
rect 66444 218152 66496 218204
rect 67548 218152 67600 218204
rect 68100 218152 68152 218204
rect 69572 218152 69624 218204
rect 75552 218152 75604 218204
rect 76564 218152 76616 218204
rect 97080 218152 97132 218204
rect 56508 218016 56560 218068
rect 57244 218016 57296 218068
rect 58164 218016 58216 218068
rect 59360 218016 59412 218068
rect 61476 218016 61528 218068
rect 62764 218016 62816 218068
rect 63960 218016 64012 218068
rect 64788 218016 64840 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 67272 218016 67324 218068
rect 68284 218016 68336 218068
rect 72240 218016 72292 218068
rect 73712 218016 73764 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 83464 218016 83516 218068
rect 84660 218016 84712 218068
rect 85304 218016 85356 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 92940 218016 92992 218068
rect 93584 218016 93636 218068
rect 95424 218016 95476 218068
rect 96252 218016 96304 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 152372 218152 152424 218204
rect 160008 218152 160060 218204
rect 162676 218152 162728 218204
rect 166632 218152 166684 218204
rect 102876 218084 102928 218136
rect 103428 218084 103480 218136
rect 103704 218084 103756 218136
rect 104808 218084 104860 218136
rect 105360 218084 105412 218136
rect 106004 218084 106056 218136
rect 111984 218084 112036 218136
rect 112812 218084 112864 218136
rect 152556 218084 152608 218136
rect 153108 218084 153160 218136
rect 155040 218084 155092 218136
rect 155684 218084 155736 218136
rect 156696 218084 156748 218136
rect 157248 218084 157300 218136
rect 170588 218016 170640 218068
rect 171968 218016 172020 218068
rect 173256 218016 173308 218068
rect 178040 218016 178092 218068
rect 178224 218016 178276 218068
rect 179328 218016 179380 218068
rect 179512 218016 179564 218068
rect 181352 218016 181404 218068
rect 184020 218016 184072 218068
rect 184664 218016 184716 218068
rect 185676 218016 185728 218068
rect 186136 218016 186188 218068
rect 188160 218016 188212 218068
rect 188896 218016 188948 218068
rect 189816 218016 189868 218068
rect 192116 218016 192168 218068
rect 192300 218016 192352 218068
rect 193036 218016 193088 218068
rect 193956 218016 194008 218068
rect 194508 218016 194560 218068
rect 194784 218016 194836 218068
rect 195888 218016 195940 218068
rect 196440 218016 196492 218068
rect 198280 218016 198332 218068
rect 200580 218152 200632 218204
rect 201500 218152 201552 218204
rect 202236 218152 202288 218204
rect 202696 218152 202748 218204
rect 203064 218152 203116 218204
rect 206284 218152 206336 218204
rect 207204 218152 207256 218204
rect 208124 218152 208176 218204
rect 211344 218152 211396 218204
rect 211804 218016 211856 218068
rect 214656 218016 214708 218068
rect 215208 218016 215260 218068
rect 215484 218016 215536 218068
rect 216496 218016 216548 218068
rect 217968 218152 218020 218204
rect 222752 218152 222804 218204
rect 222936 218152 222988 218204
rect 225604 218152 225656 218204
rect 246120 218152 246172 218204
rect 251732 218152 251784 218204
rect 328920 218152 328972 218204
rect 330484 218152 330536 218204
rect 365352 218152 365404 218204
rect 371792 218152 371844 218204
rect 374460 218152 374512 218204
rect 376024 218152 376076 218204
rect 381912 218152 381964 218204
rect 382924 218152 382976 218204
rect 401784 218152 401836 218204
rect 402796 218152 402848 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 428280 218152 428332 218204
rect 430120 218152 430172 218204
rect 433248 218152 433300 218204
rect 434720 218152 434772 218204
rect 434904 218152 434956 218204
rect 436836 218152 436888 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 491944 218152 491996 218204
rect 500960 218152 501012 218204
rect 507124 218152 507176 218204
rect 507676 218152 507728 218204
rect 513840 218152 513892 218204
rect 514024 218152 514076 218204
rect 560300 218152 560352 218204
rect 560484 218152 560536 218204
rect 563014 218152 563066 218204
rect 572674 218152 572726 218204
rect 613568 218152 613620 218204
rect 219808 218016 219860 218068
rect 221280 218016 221332 218068
rect 221832 218016 221884 218068
rect 223764 218016 223816 218068
rect 224592 218016 224644 218068
rect 225420 218016 225472 218068
rect 226156 218016 226208 218068
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233148 218016 233200 218068
rect 235356 218016 235408 218068
rect 235816 218016 235868 218068
rect 236184 218016 236236 218068
rect 237288 218016 237340 218068
rect 240324 218016 240376 218068
rect 241336 218016 241388 218068
rect 243636 218016 243688 218068
rect 244096 218016 244148 218068
rect 247776 218016 247828 218068
rect 248236 218016 248288 218068
rect 248604 218016 248656 218068
rect 249616 218016 249668 218068
rect 250260 218016 250312 218068
rect 250904 218016 250956 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 254400 218016 254452 218068
rect 255044 218016 255096 218068
rect 256056 218016 256108 218068
rect 256516 218016 256568 218068
rect 256884 218016 256936 218068
rect 257528 218016 257580 218068
rect 258540 218016 258592 218068
rect 259276 218016 259328 218068
rect 262680 218016 262732 218068
rect 263600 218016 263652 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266176 218016 266228 218068
rect 268476 218016 268528 218068
rect 268936 218016 268988 218068
rect 269304 218016 269356 218068
rect 270040 218016 270092 218068
rect 270960 218016 271012 218068
rect 272524 218016 272576 218068
rect 276756 218016 276808 218068
rect 277216 218016 277268 218068
rect 277584 218016 277636 218068
rect 278596 218016 278648 218068
rect 280896 218016 280948 218068
rect 281448 218016 281500 218068
rect 281724 218016 281776 218068
rect 282460 218016 282512 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 287520 218016 287572 218068
rect 288716 218016 288768 218068
rect 289176 218016 289228 218068
rect 289728 218016 289780 218068
rect 290004 218016 290056 218068
rect 291108 218016 291160 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 297456 218016 297508 218068
rect 297916 218016 297968 218068
rect 298284 218016 298336 218068
rect 299112 218016 299164 218068
rect 299940 218016 299992 218068
rect 300676 218016 300728 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 304080 218016 304132 218068
rect 304724 218016 304776 218068
rect 305736 218016 305788 218068
rect 306196 218016 306248 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 309876 218016 309928 218068
rect 310428 218016 310480 218068
rect 312360 218016 312412 218068
rect 312912 218016 312964 218068
rect 317328 218016 317380 218068
rect 317972 218016 318024 218068
rect 318984 218016 319036 218068
rect 319812 218016 319864 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 323124 218016 323176 218068
rect 324136 218016 324188 218068
rect 324780 218016 324832 218068
rect 325424 218016 325476 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 330576 218016 330628 218068
rect 331036 218016 331088 218068
rect 333060 218016 333112 218068
rect 333888 218016 333940 218068
rect 334716 218016 334768 218068
rect 335176 218016 335228 218068
rect 335544 218016 335596 218068
rect 338672 218016 338724 218068
rect 338856 218016 338908 218068
rect 339408 218016 339460 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 345480 218016 345532 218068
rect 347044 218016 347096 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 355416 218016 355468 218068
rect 355876 218016 355928 218068
rect 356244 218016 356296 218068
rect 356980 218016 357032 218068
rect 359556 218016 359608 218068
rect 360108 218016 360160 218068
rect 360384 218016 360436 218068
rect 361028 218016 361080 218068
rect 364524 218016 364576 218068
rect 365536 218016 365588 218068
rect 366180 218016 366232 218068
rect 366732 218016 366784 218068
rect 367836 218016 367888 218068
rect 368388 218016 368440 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373448 218016 373500 218068
rect 376116 218016 376168 218068
rect 376668 218016 376720 218068
rect 378600 218016 378652 218068
rect 379244 218016 379296 218068
rect 381084 218016 381136 218068
rect 382096 218016 382148 218068
rect 389364 218016 389416 218068
rect 390008 218016 390060 218068
rect 392676 218016 392728 218068
rect 393136 218016 393188 218068
rect 393504 218016 393556 218068
rect 394516 218016 394568 218068
rect 395160 218016 395212 218068
rect 395804 218016 395856 218068
rect 397644 218016 397696 218068
rect 400588 218016 400640 218068
rect 400956 218016 401008 218068
rect 402244 218016 402296 218068
rect 403440 218016 403492 218068
rect 403992 218016 404044 218068
rect 405096 218016 405148 218068
rect 405556 218016 405608 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 427912 218016 427964 218068
rect 429108 218016 429160 218068
rect 430580 218016 430632 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 435732 218016 435784 218068
rect 436284 218016 436336 218068
rect 436468 218016 436520 218068
rect 437480 218016 437532 218068
rect 438216 218016 438268 218068
rect 438860 218016 438912 218068
rect 439872 218016 439924 218068
rect 440332 218016 440384 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 455604 218016 455656 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 471428 218016 471480 218068
rect 472900 218016 472952 218068
rect 490380 218016 490432 218068
rect 601056 218016 601108 218068
rect 601240 218016 601292 218068
rect 563520 217948 563572 218000
rect 572168 217948 572220 218000
rect 615684 217948 615736 218000
rect 174268 217880 174320 217932
rect 523040 217812 523092 217864
rect 524236 217812 524288 217864
rect 535460 217812 535512 217864
rect 536656 217812 536708 217864
rect 533436 217676 533488 217728
rect 604000 217812 604052 217864
rect 670424 218288 670476 218340
rect 670608 218016 670660 218068
rect 675852 217948 675904 218000
rect 676772 217948 676824 218000
rect 670424 217744 670476 217796
rect 116952 217540 117004 217592
rect 189172 217540 189224 217592
rect 530952 217540 531004 217592
rect 603448 217676 603500 217728
rect 604460 217676 604512 217728
rect 614304 217676 614356 217728
rect 538220 217540 538272 217592
rect 539140 217540 539192 217592
rect 543372 217540 543424 217592
rect 606208 217540 606260 217592
rect 614120 217540 614172 217592
rect 626632 217540 626684 217592
rect 115296 217404 115348 217456
rect 187976 217404 188028 217456
rect 527824 217404 527876 217456
rect 528468 217404 528520 217456
rect 90410 217200 90462 217252
rect 168564 217268 168616 217320
rect 508596 217268 508648 217320
rect 563014 217268 563066 217320
rect 563152 217268 563204 217320
rect 572536 217268 572588 217320
rect 572674 217268 572726 217320
rect 598480 217268 598532 217320
rect 448612 217200 448664 217252
rect 449762 217200 449814 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 498292 217200 498344 217252
rect 499442 217200 499494 217252
rect 506066 217132 506118 217184
rect 597928 217132 597980 217184
rect 603080 217404 603132 217456
rect 628288 217404 628340 217456
rect 670240 217336 670292 217388
rect 670608 217336 670660 217388
rect 598848 217268 598900 217320
rect 622400 217268 622452 217320
rect 603080 217132 603132 217184
rect 498614 217064 498666 217116
rect 574192 216996 574244 217048
rect 610072 216996 610124 217048
rect 596364 216860 596416 216912
rect 607128 216860 607180 216912
rect 612280 216860 612332 216912
rect 594800 216724 594852 216776
rect 613384 216724 613436 216776
rect 613568 216656 613620 216708
rect 614488 216656 614540 216708
rect 648252 216656 648304 216708
rect 650644 216656 650696 216708
rect 644940 215908 644992 215960
rect 658924 215908 658976 215960
rect 675852 215636 675904 215688
rect 676956 215636 677008 215688
rect 675852 214956 675904 215008
rect 676496 214956 676548 215008
rect 574744 214820 574796 214872
rect 616880 214820 616932 214872
rect 574376 214684 574428 214736
rect 623320 214684 623372 214736
rect 658188 214684 658240 214736
rect 665824 214684 665876 214736
rect 574560 214548 574612 214600
rect 601792 214412 601844 214464
rect 602344 214412 602396 214464
rect 604644 214412 604696 214464
rect 605104 214412 605156 214464
rect 607312 214548 607364 214600
rect 607864 214548 607916 214600
rect 618260 214548 618312 214600
rect 618904 214548 618956 214600
rect 619916 214548 619968 214600
rect 620560 214548 620612 214600
rect 623964 214548 624016 214600
rect 624424 214412 624476 214464
rect 625436 214548 625488 214600
rect 626080 214548 626132 214600
rect 630036 214548 630088 214600
rect 632888 214548 632940 214600
rect 646320 214548 646372 214600
rect 656164 214548 656216 214600
rect 629392 214412 629444 214464
rect 35808 213936 35860 213988
rect 41696 213936 41748 213988
rect 645860 213868 645912 213920
rect 646504 213868 646556 213920
rect 648620 213868 648672 213920
rect 649264 213868 649316 213920
rect 663156 213868 663208 213920
rect 663708 213868 663760 213920
rect 653220 213800 653272 213852
rect 654784 213800 654836 213852
rect 656532 213392 656584 213444
rect 664628 213392 664680 213444
rect 643836 213324 643888 213376
rect 653404 213324 653456 213376
rect 575480 213188 575532 213240
rect 594800 213188 594852 213240
rect 645492 213188 645544 213240
rect 660764 213256 660816 213308
rect 654600 213120 654652 213172
rect 657544 213120 657596 213172
rect 600412 212984 600464 213036
rect 601240 212984 601292 213036
rect 632704 212984 632756 213036
rect 634360 212984 634412 213036
rect 654140 212916 654192 212968
rect 654784 212916 654836 212968
rect 600504 212848 600556 212900
rect 600872 212848 600924 212900
rect 35808 212780 35860 212832
rect 39948 212780 40000 212832
rect 650460 212712 650512 212764
rect 651288 212712 651340 212764
rect 664260 212712 664312 212764
rect 665088 212712 665140 212764
rect 592684 212644 592736 212696
rect 641720 212644 641772 212696
rect 35624 212508 35676 212560
rect 39580 212508 39632 212560
rect 591304 212508 591356 212560
rect 639880 212508 639932 212560
rect 578516 211148 578568 211200
rect 580908 211148 580960 211200
rect 35808 209924 35860 209976
rect 40408 209924 40460 209976
rect 579528 209788 579580 209840
rect 582288 209788 582340 209840
rect 35808 208700 35860 208752
rect 40040 208632 40092 208684
rect 581644 208564 581696 208616
rect 632152 209516 632204 209568
rect 652024 209516 652076 209568
rect 667756 209040 667808 209092
rect 35808 208496 35860 208548
rect 40592 208496 40644 208548
rect 35624 208360 35676 208412
rect 41696 208360 41748 208412
rect 42064 208360 42116 208412
rect 43352 208360 43404 208412
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 35808 207136 35860 207188
rect 39948 207136 40000 207188
rect 580908 206864 580960 206916
rect 589464 206864 589516 206916
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 582288 205504 582340 205556
rect 589464 205504 589516 205556
rect 35808 204620 35860 204672
rect 41512 204484 41564 204536
rect 35808 204280 35860 204332
rect 41696 204348 41748 204400
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 35808 202852 35860 202904
rect 37924 202852 37976 202904
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 42524 201696 42576 201748
rect 42892 201696 42944 201748
rect 43260 202104 43312 202156
rect 42708 201560 42760 201612
rect 43076 201560 43128 201612
rect 42892 201288 42944 201340
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 42248 190204 42300 190256
rect 42892 190204 42944 190256
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 42432 187620 42484 187672
rect 43076 187620 43128 187672
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 668952 184832 669004 184884
rect 670700 184832 670752 184884
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 668216 177964 668268 178016
rect 670792 177964 670844 178016
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 668032 175040 668084 175092
rect 670424 175040 670476 175092
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 580264 171096 580316 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 667940 169668 667992 169720
rect 669688 169668 669740 169720
rect 582380 168376 582432 168428
rect 589464 168376 589516 168428
rect 578240 167288 578292 167340
rect 580264 167288 580316 167340
rect 579988 167016 580040 167068
rect 589464 167016 589516 167068
rect 579528 166268 579580 166320
rect 589648 166268 589700 166320
rect 579344 165180 579396 165232
rect 582380 165180 582432 165232
rect 667940 165044 667992 165096
rect 670056 165044 670108 165096
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 675852 164160 675904 164212
rect 682384 164160 682436 164212
rect 578240 163616 578292 163668
rect 579988 163616 580040 163668
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 578424 162664 578476 162716
rect 582472 162664 582524 162716
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580724 160080 580776 160132
rect 589464 160080 589516 160132
rect 668216 160012 668268 160064
rect 670792 160012 670844 160064
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 585784 158720 585836 158772
rect 589464 158720 589516 158772
rect 587164 157360 587216 157412
rect 589280 157360 589332 157412
rect 668216 155524 668268 155576
rect 670792 155524 670844 155576
rect 578332 154640 578384 154692
rect 580540 154640 580592 154692
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 580724 152736 580776 152788
rect 580264 151784 580316 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 585784 150560 585836 150612
rect 585140 149064 585192 149116
rect 589464 149064 589516 149116
rect 579528 148316 579580 148368
rect 587164 148316 587216 148368
rect 578884 146276 578936 146328
rect 585140 146276 585192 146328
rect 668768 145732 668820 145784
rect 670792 145732 670844 145784
rect 584772 144916 584824 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 585968 143556 586020 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 587164 142400 587216 142452
rect 589832 142400 589884 142452
rect 580448 140768 580500 140820
rect 589464 140768 589516 140820
rect 578608 140700 578660 140752
rect 580264 140700 580316 140752
rect 583024 139408 583076 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 579528 138660 579580 138712
rect 588544 138660 588596 138712
rect 579068 137300 579120 137352
rect 584772 137300 584824 137352
rect 584588 136620 584640 136672
rect 589464 136620 589516 136672
rect 580264 134512 580316 134564
rect 589464 134512 589516 134564
rect 675852 133900 675904 133952
rect 676496 133900 676548 133952
rect 667940 133764 667992 133816
rect 669872 133764 669924 133816
rect 585784 132472 585836 132524
rect 589464 132472 589516 132524
rect 581828 131248 581880 131300
rect 589464 131248 589516 131300
rect 578884 131112 578936 131164
rect 585968 131112 586020 131164
rect 668492 130772 668544 130824
rect 670792 130772 670844 130824
rect 668032 129684 668084 129736
rect 670148 129684 670200 129736
rect 583208 129140 583260 129192
rect 590384 129140 590436 129192
rect 579528 129004 579580 129056
rect 587164 129004 587216 129056
rect 579068 126964 579120 127016
rect 589464 126964 589516 127016
rect 578332 125604 578384 125656
rect 580448 125604 580500 125656
rect 675852 125400 675904 125452
rect 676404 125400 676456 125452
rect 580448 124176 580500 124228
rect 589464 124176 589516 124228
rect 578424 123564 578476 123616
rect 583024 123564 583076 123616
rect 584404 122816 584456 122868
rect 589464 122816 589516 122868
rect 578884 122136 578936 122188
rect 584588 122136 584640 122188
rect 580632 122000 580684 122052
rect 589924 122000 589976 122052
rect 587348 118668 587400 118720
rect 590016 118668 590068 118720
rect 675852 118464 675904 118516
rect 679624 118464 679676 118516
rect 578516 118396 578568 118448
rect 580264 118396 580316 118448
rect 579528 116900 579580 116952
rect 583208 116900 583260 116952
rect 668768 116832 668820 116884
rect 670608 116832 670660 116884
rect 586152 115948 586204 116000
rect 589464 115948 589516 116000
rect 583208 115200 583260 115252
rect 589648 115200 589700 115252
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 583024 113160 583076 113212
rect 589464 113160 589516 113212
rect 579528 112820 579580 112872
rect 585784 112820 585836 112872
rect 585968 112412 586020 112464
rect 590108 112412 590160 112464
rect 581644 110440 581696 110492
rect 589464 110440 589516 110492
rect 579344 110100 579396 110152
rect 581828 110100 581880 110152
rect 584588 109012 584640 109064
rect 589280 109012 589332 109064
rect 667940 108808 667992 108860
rect 669964 108808 670016 108860
rect 578332 108672 578384 108724
rect 580632 108672 580684 108724
rect 578884 107584 578936 107636
rect 589464 107652 589516 107704
rect 587164 106292 587216 106344
rect 589832 106292 589884 106344
rect 668400 106156 668452 106208
rect 670792 106156 670844 106208
rect 580264 104864 580316 104916
rect 589464 104864 589516 104916
rect 668768 104660 668820 104712
rect 670792 104660 670844 104712
rect 579528 103436 579580 103488
rect 588544 103436 588596 103488
rect 579528 101804 579580 101856
rect 584404 101804 584456 101856
rect 584404 100104 584456 100156
rect 589464 100104 589516 100156
rect 579068 99356 579120 99408
rect 586152 99356 586204 99408
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 578608 99220 578660 99272
rect 580448 99220 580500 99272
rect 623688 99152 623740 99204
rect 633440 99152 633492 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 625068 99016 625120 99068
rect 636292 99016 636344 99068
rect 628288 98880 628340 98932
rect 642180 98880 642232 98932
rect 629024 98744 629076 98796
rect 643652 98744 643704 98796
rect 647148 98744 647200 98796
rect 661960 98744 662012 98796
rect 630496 98608 630548 98660
rect 646596 98608 646648 98660
rect 631048 98200 631100 98252
rect 640708 98132 640760 98184
rect 578332 97928 578384 97980
rect 587348 97928 587400 97980
rect 618720 97928 618772 97980
rect 625804 97928 625856 97980
rect 629760 97928 629812 97980
rect 645308 97996 645360 98048
rect 659936 97928 659988 97980
rect 665180 97928 665232 97980
rect 620192 97792 620244 97844
rect 625620 97792 625672 97844
rect 627552 97792 627604 97844
rect 631048 97792 631100 97844
rect 631968 97792 632020 97844
rect 647516 97792 647568 97844
rect 655428 97792 655480 97844
rect 662512 97792 662564 97844
rect 632704 97656 632756 97708
rect 648252 97656 648304 97708
rect 651840 97656 651892 97708
rect 659568 97656 659620 97708
rect 621664 97520 621716 97572
rect 629300 97520 629352 97572
rect 634176 97520 634228 97572
rect 612648 97384 612700 97436
rect 618904 97384 618956 97436
rect 623136 97384 623188 97436
rect 632060 97384 632112 97436
rect 633256 97384 633308 97436
rect 648620 97384 648672 97436
rect 650368 97520 650420 97572
rect 658280 97520 658332 97572
rect 650552 97384 650604 97436
rect 658096 97384 658148 97436
rect 663064 97384 663116 97436
rect 605472 97248 605524 97300
rect 611912 97248 611964 97300
rect 626080 97248 626132 97300
rect 637764 97248 637816 97300
rect 643008 97248 643060 97300
rect 656532 97248 656584 97300
rect 656808 97248 656860 97300
rect 661408 97248 661460 97300
rect 626816 97112 626868 97164
rect 639236 97112 639288 97164
rect 644296 97112 644348 97164
rect 658832 97112 658884 97164
rect 624608 96976 624660 97028
rect 635004 96976 635056 97028
rect 635556 96976 635608 97028
rect 647700 96976 647752 97028
rect 659200 96976 659252 97028
rect 663892 96976 663944 97028
rect 596180 96908 596232 96960
rect 596732 96908 596784 96960
rect 597652 96908 597704 96960
rect 598204 96908 598256 96960
rect 598940 96908 598992 96960
rect 599676 96908 599728 96960
rect 600320 96908 600372 96960
rect 601148 96908 601200 96960
rect 606208 96908 606260 96960
rect 607128 96908 607180 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 617248 96840 617300 96892
rect 618168 96840 618220 96892
rect 634728 96840 634780 96892
rect 650368 96840 650420 96892
rect 653956 96840 654008 96892
rect 655244 96840 655296 96892
rect 656716 96840 656768 96892
rect 660120 96840 660172 96892
rect 610624 96704 610676 96756
rect 611268 96704 611320 96756
rect 640524 96568 640576 96620
rect 647884 96704 647936 96756
rect 654784 96704 654836 96756
rect 655428 96704 655480 96756
rect 656532 96704 656584 96756
rect 660120 96704 660172 96756
rect 645768 96568 645820 96620
rect 656348 96568 656400 96620
rect 639052 96432 639104 96484
rect 645124 96432 645176 96484
rect 646412 96432 646464 96484
rect 652024 96432 652076 96484
rect 652576 96432 652628 96484
rect 665548 96432 665600 96484
rect 631232 96296 631284 96348
rect 647148 96296 647200 96348
rect 648896 96296 648948 96348
rect 664168 96296 664220 96348
rect 637580 96160 637632 96212
rect 660672 96160 660724 96212
rect 611084 96024 611136 96076
rect 622308 96024 622360 96076
rect 649908 96024 649960 96076
rect 663708 96024 663760 96076
rect 644940 95956 644992 96008
rect 649540 95956 649592 96008
rect 607680 95888 607732 95940
rect 624976 95888 625028 95940
rect 643468 95820 643520 95872
rect 649264 95820 649316 95872
rect 665364 95888 665416 95940
rect 638592 95684 638644 95736
rect 647332 95684 647384 95736
rect 647884 95684 647936 95736
rect 653312 95616 653364 95668
rect 664352 95616 664404 95668
rect 640064 95548 640116 95600
rect 647884 95548 647936 95600
rect 641536 95412 641588 95464
rect 645124 95412 645176 95464
rect 651840 95412 651892 95464
rect 649908 95276 649960 95328
rect 620928 95140 620980 95192
rect 626448 95140 626500 95192
rect 647700 95072 647752 95124
rect 648804 95072 648856 95124
rect 579528 95004 579580 95056
rect 583208 95004 583260 95056
rect 616512 95004 616564 95056
rect 622952 95004 623004 95056
rect 609152 94460 609204 94512
rect 620284 94460 620336 94512
rect 649540 93916 649592 93968
rect 656164 93916 656216 93968
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 651288 93508 651340 93560
rect 655428 93508 655480 93560
rect 578516 93440 578568 93492
rect 585968 93440 586020 93492
rect 611268 93100 611320 93152
rect 619272 93100 619324 93152
rect 606944 92828 606996 92880
rect 610072 92828 610124 92880
rect 648620 92488 648672 92540
rect 650000 92488 650052 92540
rect 617984 92420 618036 92472
rect 626448 92420 626500 92472
rect 647332 92352 647384 92404
rect 654324 92352 654376 92404
rect 579344 91060 579396 91112
rect 584588 91060 584640 91112
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 651840 90652 651892 90704
rect 655428 90652 655480 90704
rect 622952 89564 623004 89616
rect 625252 89564 625304 89616
rect 585140 88952 585192 89004
rect 589924 88952 589976 89004
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 663892 88748 663944 88800
rect 656348 88612 656400 88664
rect 657452 88612 657504 88664
rect 610072 88272 610124 88324
rect 625160 88272 625212 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 622308 88136 622360 88188
rect 625344 88136 625396 88188
rect 579528 88068 579580 88120
rect 585140 88068 585192 88120
rect 648436 86980 648488 87032
rect 662512 86980 662564 87032
rect 656716 86844 656768 86896
rect 659568 86844 659620 86896
rect 649264 86708 649316 86760
rect 661408 86708 661460 86760
rect 647884 86572 647936 86624
rect 660120 86572 660172 86624
rect 656164 86436 656216 86488
rect 660672 86436 660724 86488
rect 619272 86300 619324 86352
rect 625160 86300 625212 86352
rect 652024 86300 652076 86352
rect 657176 86300 657228 86352
rect 620284 85484 620336 85536
rect 625344 85484 625396 85536
rect 609888 85348 609940 85400
rect 625160 85280 625212 85332
rect 579160 84124 579212 84176
rect 581644 84124 581696 84176
rect 608508 84124 608560 84176
rect 625160 84124 625212 84176
rect 579068 82356 579120 82408
rect 583024 82356 583076 82408
rect 579528 82084 579580 82136
rect 587164 82084 587216 82136
rect 628748 80928 628800 80980
rect 642456 80928 642508 80980
rect 612648 80792 612700 80844
rect 647424 80792 647476 80844
rect 595444 80656 595496 80708
rect 636752 80656 636804 80708
rect 629208 79976 629260 80028
rect 633440 79976 633492 80028
rect 613844 79432 613896 79484
rect 645952 79432 646004 79484
rect 579068 79296 579120 79348
rect 588728 79296 588780 79348
rect 614028 79296 614080 79348
rect 646504 79296 646556 79348
rect 633440 78072 633492 78124
rect 645308 78072 645360 78124
rect 631048 77936 631100 77988
rect 643100 77936 643152 77988
rect 628472 77732 628524 77784
rect 632796 77732 632848 77784
rect 625804 77256 625856 77308
rect 631048 77256 631100 77308
rect 616788 76644 616840 76696
rect 646320 76644 646372 76696
rect 612004 76508 612056 76560
rect 662420 76508 662472 76560
rect 578240 75828 578292 75880
rect 580264 75828 580316 75880
rect 618904 75420 618956 75472
rect 648620 75420 648672 75472
rect 615408 75284 615460 75336
rect 646872 75284 646924 75336
rect 607128 75148 607180 75200
rect 646136 75148 646188 75200
rect 578884 72428 578936 72480
rect 601700 72428 601752 72480
rect 579068 71340 579120 71392
rect 584404 71340 584456 71392
rect 580264 68280 580316 68332
rect 604460 68280 604512 68332
rect 577504 59984 577556 60036
rect 603080 59984 603132 60036
rect 576124 58624 576176 58676
rect 601884 58624 601936 58676
rect 574928 57196 574980 57248
rect 600320 57196 600372 57248
rect 574744 55972 574796 56024
rect 598940 55972 598992 56024
rect 574560 55836 574612 55888
rect 600504 55836 600556 55888
rect 596456 55156 596508 55208
rect 597836 55020 597888 55072
rect 597652 54884 597704 54936
rect 464160 53592 464212 53644
rect 464344 53592 464396 53644
rect 464528 53592 464580 53644
rect 599124 54748 599176 54800
rect 624424 54612 624476 54664
rect 625804 54476 625856 54528
rect 596180 54340 596232 54392
rect 581644 54204 581696 54256
rect 464896 53592 464948 53644
rect 465908 53592 465960 53644
rect 466092 53592 466144 53644
rect 471980 53524 472032 53576
rect 472808 53524 472860 53576
rect 462228 53456 462280 53508
rect 471796 53456 471848 53508
rect 461308 53320 461360 53372
rect 574744 54068 574796 54120
rect 574560 53932 574612 53984
rect 473728 53592 473780 53644
rect 574928 53796 574980 53848
rect 473544 53456 473596 53508
rect 49148 53184 49200 53236
rect 129004 53184 129056 53236
rect 464068 53184 464120 53236
rect 471980 53184 472032 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 48964 53048 49016 53100
rect 130384 53048 130436 53100
rect 459468 53048 459520 53100
rect 464896 53048 464948 53100
rect 463148 52912 463200 52964
rect 473728 52912 473780 52964
rect 460066 52776 460118 52828
rect 466092 52776 466144 52828
rect 463608 52640 463660 52692
rect 464528 52640 464580 52692
rect 465448 52640 465500 52692
rect 472808 52640 472860 52692
rect 47584 51960 47636 52012
rect 130568 51960 130620 52012
rect 50344 51824 50396 51876
rect 129188 51824 129240 51876
rect 129556 51824 129608 51876
rect 591304 51824 591356 51876
rect 128820 51688 128872 51740
rect 592684 51688 592736 51740
rect 318340 50464 318392 50516
rect 458180 50464 458232 50516
rect 47768 50328 47820 50380
rect 130752 50328 130804 50380
rect 314016 50328 314068 50380
rect 458364 50328 458416 50380
rect 522948 50328 523000 50380
rect 544016 50328 544068 50380
rect 50528 49104 50580 49156
rect 129372 49104 129424 49156
rect 46204 48968 46256 49020
rect 130936 48968 130988 49020
rect 130568 45500 130620 45552
rect 132592 45500 132644 45552
rect 129004 45296 129056 45348
rect 131396 45160 131448 45212
rect 133144 45160 133196 45212
rect 129556 45024 129608 45076
rect 129372 44888 129424 44940
rect 128820 44752 128872 44804
rect 131580 44616 131632 44668
rect 129188 44480 129240 44532
rect 43628 44276 43680 44328
rect 132592 44364 132644 44416
rect 132408 44276 132460 44328
rect 43444 44140 43496 44192
rect 131580 44140 131632 44192
rect 130752 44004 130804 44056
rect 133144 44140 133196 44192
rect 440240 43800 440292 43852
rect 441068 43800 441120 43852
rect 187332 42780 187384 42832
rect 255872 42780 255924 42832
rect 307300 42712 307352 42764
rect 431224 42712 431276 42764
rect 441068 42712 441120 42764
rect 449164 42712 449216 42764
rect 453580 42712 453632 42764
rect 464160 42712 464212 42764
rect 310428 42576 310480 42628
rect 427084 42576 427136 42628
rect 441252 42576 441304 42628
rect 446404 42576 446456 42628
rect 454500 42440 454552 42492
rect 463056 42440 463108 42492
rect 404452 42304 404504 42356
rect 405188 42304 405240 42356
rect 420736 42304 420788 42356
rect 426900 42304 426952 42356
rect 661408 42129 661460 42181
rect 427084 41964 427136 42016
rect 431224 41964 431276 42016
rect 441068 41964 441120 42016
rect 446404 41964 446456 42016
rect 454500 41964 454552 42016
rect 441252 41828 441304 41880
rect 449164 41828 449216 41880
rect 453580 41828 453632 41880
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 426900 41420 426952 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 185030 1002144 185086 1002153
rect 185030 1002079 185086 1002088
rect 82174 1002008 82230 1002017
rect 81452 1001966 82174 1001994
rect 81452 997098 81480 1001966
rect 133694 1002008 133750 1002017
rect 82174 1001943 82230 1001952
rect 132500 1001972 132552 1001978
rect 133694 1001943 133696 1001952
rect 132500 1001914 132552 1001920
rect 133748 1001943 133750 1001952
rect 133696 1001914 133748 1001920
rect 81360 997070 81480 997098
rect 81360 983521 81388 997070
rect 81346 983512 81402 983521
rect 81346 983447 81402 983456
rect 132512 982569 132540 1001914
rect 185044 992234 185072 1002079
rect 483018 1002008 483074 1002017
rect 483018 1001943 483074 1001952
rect 534998 1002008 535054 1002017
rect 636198 1002008 636254 1002017
rect 535054 1001966 535500 1001994
rect 534998 1001943 535054 1001952
rect 232976 997393 233004 997628
rect 245226 997614 245700 997642
rect 232962 997384 233018 997393
rect 232962 997319 233018 997328
rect 240138 997248 240194 997257
rect 240138 997183 240194 997192
rect 184952 992206 185072 992234
rect 184952 983521 184980 992206
rect 235906 990992 235962 991001
rect 235906 990927 235962 990936
rect 235920 983793 235948 990927
rect 238668 985992 238720 985998
rect 238668 985934 238720 985940
rect 238680 984065 238708 985934
rect 238666 984056 238722 984065
rect 238666 983991 238722 984000
rect 240152 983793 240180 997183
rect 245672 989126 245700 997614
rect 285416 997393 285444 997628
rect 297850 997614 298140 997642
rect 285402 997384 285458 997393
rect 285402 997319 285458 997328
rect 292578 997384 292634 997393
rect 292578 997319 292634 997328
rect 242256 989120 242308 989126
rect 242256 989062 242308 989068
rect 245660 989120 245712 989126
rect 245660 989062 245712 989068
rect 242268 985998 242296 989062
rect 286966 988000 287022 988009
rect 286966 987935 287022 987944
rect 242256 985992 242308 985998
rect 242256 985934 242308 985940
rect 286980 983793 287008 987935
rect 289728 985448 289780 985454
rect 289728 985390 289780 985396
rect 235906 983784 235962 983793
rect 235906 983719 235962 983728
rect 240138 983784 240194 983793
rect 240138 983719 240194 983728
rect 286966 983784 287022 983793
rect 286966 983719 287022 983728
rect 184938 983512 184994 983521
rect 184938 983447 184994 983456
rect 132498 982560 132554 982569
rect 132498 982495 132554 982504
rect 289740 980937 289768 985390
rect 292592 983793 292620 997319
rect 298112 988242 298140 997614
rect 387536 997393 387564 997628
rect 399602 997614 400260 997642
rect 387522 997384 387578 997393
rect 387522 997319 387578 997328
rect 389178 990992 389234 991001
rect 389178 990927 389234 990936
rect 293960 988236 294012 988242
rect 293960 988178 294012 988184
rect 298100 988236 298152 988242
rect 298100 988178 298152 988184
rect 293972 985454 294000 988178
rect 389192 987562 389220 990927
rect 400232 990894 400260 997614
rect 404358 997384 404414 997393
rect 404358 997319 404414 997328
rect 404372 992254 404400 997319
rect 401692 992248 401744 992254
rect 401692 992190 401744 992196
rect 404360 992248 404412 992254
rect 404360 992190 404412 992196
rect 396080 990888 396132 990894
rect 396080 990830 396132 990836
rect 400220 990888 400272 990894
rect 400220 990830 400272 990836
rect 389180 987556 389232 987562
rect 389180 987498 389232 987504
rect 391940 987556 391992 987562
rect 391940 987498 391992 987504
rect 293960 985448 294012 985454
rect 293960 985390 294012 985396
rect 292578 983784 292634 983793
rect 292578 983719 292634 983728
rect 391952 983521 391980 987498
rect 396092 983550 396120 990830
rect 401704 986406 401732 992190
rect 399760 986400 399812 986406
rect 399760 986342 399812 986348
rect 401692 986400 401744 986406
rect 401692 986342 401744 986348
rect 394424 983544 394476 983550
rect 391938 983512 391994 983521
rect 391938 983447 391994 983456
rect 394422 983512 394424 983521
rect 396080 983544 396132 983550
rect 394476 983512 394478 983521
rect 399772 983521 399800 986342
rect 396080 983486 396132 983492
rect 399758 983512 399814 983521
rect 394422 983447 394478 983456
rect 399758 983447 399814 983456
rect 483032 982530 483060 1001943
rect 535472 983793 535500 1001966
rect 636198 1001943 636254 1001952
rect 636212 983793 636240 1001943
rect 535458 983784 535514 983793
rect 535458 983719 535514 983728
rect 636198 983784 636254 983793
rect 636198 983719 636254 983728
rect 483846 982560 483902 982569
rect 483020 982524 483072 982530
rect 483846 982495 483848 982504
rect 483020 982466 483072 982472
rect 483900 982495 483902 982504
rect 483848 982466 483900 982472
rect 289726 980928 289782 980937
rect 289726 980863 289782 980872
rect 30102 960256 30158 960265
rect 30102 960191 30158 960200
rect 30116 954990 30144 960191
rect 651378 959168 651434 959177
rect 651378 959103 651380 959112
rect 651432 959103 651434 959112
rect 677414 959168 677470 959177
rect 677414 959103 677416 959112
rect 651380 959074 651432 959080
rect 677468 959103 677470 959112
rect 677416 959074 677468 959080
rect 63406 959032 63462 959041
rect 63406 958967 63462 958976
rect 63420 954990 63448 958967
rect 30104 954984 30156 954990
rect 30104 954926 30156 954932
rect 63408 954984 63460 954990
rect 63408 954926 63460 954932
rect 703694 897668 703722 897804
rect 704154 897668 704182 897804
rect 704614 897668 704642 897804
rect 705074 897668 705102 897804
rect 705534 897668 705562 897804
rect 705994 897668 706022 897804
rect 706454 897668 706482 897804
rect 706914 897668 706942 897804
rect 707374 897668 707402 897804
rect 707834 897668 707862 897804
rect 708294 897668 708322 897804
rect 708754 897668 708782 897804
rect 709214 897668 709242 897804
rect 676034 897152 676090 897161
rect 676034 897087 676036 897096
rect 676088 897087 676090 897096
rect 676036 897058 676088 897064
rect 652024 897048 652076 897054
rect 652024 896990 652076 896996
rect 651472 868896 651524 868902
rect 651472 868838 651524 868844
rect 651484 868601 651512 868838
rect 651470 868592 651526 868601
rect 651470 868527 651526 868536
rect 652036 867649 652064 896990
rect 675850 896744 675906 896753
rect 675850 896679 675906 896688
rect 675864 895830 675892 896679
rect 676034 896336 676090 896345
rect 676034 896271 676090 896280
rect 654784 895824 654836 895830
rect 654784 895766 654836 895772
rect 675852 895824 675904 895830
rect 675852 895766 675904 895772
rect 653404 880524 653456 880530
rect 653404 880466 653456 880472
rect 652022 867640 652078 867649
rect 652022 867575 652078 867584
rect 651472 866652 651524 866658
rect 651472 866594 651524 866600
rect 651484 866289 651512 866594
rect 651470 866280 651526 866289
rect 651470 866215 651526 866224
rect 653416 865230 653444 880466
rect 654796 868902 654824 895766
rect 676048 895694 676076 896271
rect 672724 895688 672776 895694
rect 672724 895630 672776 895636
rect 676036 895688 676088 895694
rect 676036 895630 676088 895636
rect 671068 894464 671120 894470
rect 671068 894406 671120 894412
rect 670884 886916 670936 886922
rect 670884 886858 670936 886864
rect 657544 869440 657596 869446
rect 657544 869382 657596 869388
rect 654784 868896 654836 868902
rect 654784 868838 654836 868844
rect 654140 868080 654192 868086
rect 654140 868022 654192 868028
rect 651380 865224 651432 865230
rect 651378 865192 651380 865201
rect 653404 865224 653456 865230
rect 651432 865192 651434 865201
rect 653404 865166 653456 865172
rect 651378 865127 651434 865136
rect 651472 863864 651524 863870
rect 651470 863832 651472 863841
rect 651524 863832 651526 863841
rect 651470 863767 651526 863776
rect 654152 862510 654180 868022
rect 657556 863870 657584 869382
rect 657544 863864 657596 863870
rect 657544 863806 657596 863812
rect 651472 862504 651524 862510
rect 651472 862446 651524 862452
rect 654140 862504 654192 862510
rect 654140 862446 654192 862452
rect 651484 862345 651512 862446
rect 651470 862336 651526 862345
rect 651470 862271 651526 862280
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35622 818000 35678 818009
rect 35622 817935 35678 817944
rect 35636 817018 35664 817935
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817154 35848 817255
rect 35808 817148 35860 817154
rect 35808 817090 35860 817096
rect 46204 817148 46256 817154
rect 46204 817090 46256 817096
rect 35624 817012 35676 817018
rect 35624 816954 35676 816960
rect 35438 816912 35494 816921
rect 35438 816847 35494 816856
rect 35452 815658 35480 816847
rect 35806 816096 35862 816105
rect 35806 816031 35862 816040
rect 35820 815794 35848 816031
rect 35808 815788 35860 815794
rect 35808 815730 35860 815736
rect 42892 815788 42944 815794
rect 42892 815730 42944 815736
rect 35440 815652 35492 815658
rect 35440 815594 35492 815600
rect 35622 815280 35678 815289
rect 35622 815215 35678 815224
rect 35636 814434 35664 815215
rect 35806 814464 35862 814473
rect 35624 814428 35676 814434
rect 35806 814399 35862 814408
rect 35624 814370 35676 814376
rect 35820 814298 35848 814399
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41326 813648 41382 813657
rect 41326 813583 41382 813592
rect 41340 812870 41368 813583
rect 41328 812864 41380 812870
rect 40958 812832 41014 812841
rect 41328 812806 41380 812812
rect 40958 812767 41014 812776
rect 37922 811608 37978 811617
rect 37922 811543 37978 811552
rect 34518 811200 34574 811209
rect 34518 811135 34574 811144
rect 32586 810792 32642 810801
rect 32586 810727 32642 810736
rect 31022 809976 31078 809985
rect 31022 809911 31078 809920
rect 31036 801106 31064 809911
rect 32600 802505 32628 810727
rect 32586 802496 32642 802505
rect 34532 802466 34560 811135
rect 36542 809568 36598 809577
rect 36542 809503 36598 809512
rect 32586 802431 32642 802440
rect 34520 802460 34572 802466
rect 34520 802402 34572 802408
rect 31024 801100 31076 801106
rect 31024 801042 31076 801048
rect 36556 800766 36584 809503
rect 37936 801786 37964 811543
rect 40972 810762 41000 812767
rect 41326 812424 41382 812433
rect 41326 812359 41382 812368
rect 41142 812016 41198 812025
rect 41142 811951 41198 811960
rect 40960 810756 41012 810762
rect 40960 810698 41012 810704
rect 41156 809962 41184 811951
rect 41340 811510 41368 812359
rect 41328 811504 41380 811510
rect 41328 811446 41380 811452
rect 42708 810756 42760 810762
rect 42708 810698 42760 810704
rect 41970 810384 42026 810393
rect 41970 810319 42026 810328
rect 41786 809976 41842 809985
rect 41156 809934 41786 809962
rect 41786 809911 41842 809920
rect 41326 809160 41382 809169
rect 41326 809095 41382 809104
rect 41340 808654 41368 809095
rect 41786 808752 41842 808761
rect 41786 808687 41842 808696
rect 41328 808648 41380 808654
rect 41328 808590 41380 808596
rect 41142 808344 41198 808353
rect 41142 808279 41198 808288
rect 41156 807362 41184 808279
rect 41326 807528 41382 807537
rect 41326 807463 41328 807472
rect 41380 807463 41382 807472
rect 41328 807434 41380 807440
rect 41144 807356 41196 807362
rect 41144 807298 41196 807304
rect 41142 806712 41198 806721
rect 41142 806647 41198 806656
rect 41156 806002 41184 806647
rect 41326 806304 41382 806313
rect 41326 806239 41382 806248
rect 41340 806138 41368 806239
rect 41328 806132 41380 806138
rect 41328 806074 41380 806080
rect 41144 805996 41196 806002
rect 41144 805938 41196 805944
rect 41800 805225 41828 808687
rect 41984 805633 42012 810319
rect 42248 808648 42300 808654
rect 42248 808590 42300 808596
rect 41970 805624 42026 805633
rect 41970 805559 42026 805568
rect 41786 805216 41842 805225
rect 41786 805151 41842 805160
rect 42260 804554 42288 808590
rect 42168 804526 42288 804554
rect 41880 802460 41932 802466
rect 41880 802402 41932 802408
rect 37924 801780 37976 801786
rect 37924 801722 37976 801728
rect 39764 801780 39816 801786
rect 39764 801722 39816 801728
rect 36544 800760 36596 800766
rect 36544 800702 36596 800708
rect 39776 800601 39804 801722
rect 40500 800760 40552 800766
rect 40498 800728 40500 800737
rect 40552 800728 40554 800737
rect 40498 800663 40554 800672
rect 39762 800592 39818 800601
rect 39762 800527 39818 800536
rect 41892 800442 41920 802402
rect 42168 801009 42196 804526
rect 42720 801794 42748 810698
rect 42720 801766 42840 801794
rect 42524 801100 42576 801106
rect 42524 801042 42576 801048
rect 42154 801000 42210 801009
rect 42154 800935 42210 800944
rect 41892 800414 42288 800442
rect 42260 799459 42288 800414
rect 42182 799431 42288 799459
rect 42248 799332 42300 799338
rect 42248 799274 42300 799280
rect 42260 797619 42288 799274
rect 42182 797591 42288 797619
rect 42154 797328 42210 797337
rect 42154 797263 42210 797272
rect 42168 796960 42196 797263
rect 41786 796240 41842 796249
rect 41786 796175 41842 796184
rect 41800 795765 41828 796175
rect 42248 795660 42300 795666
rect 42248 795602 42300 795608
rect 42260 795138 42288 795602
rect 42182 795110 42288 795138
rect 41786 794880 41842 794889
rect 41786 794815 41842 794824
rect 41800 794580 41828 794815
rect 42154 794472 42210 794481
rect 42154 794407 42210 794416
rect 42168 793900 42196 794407
rect 42340 793960 42392 793966
rect 42340 793902 42392 793908
rect 42352 793302 42380 793902
rect 42182 793274 42380 793302
rect 41786 793112 41842 793121
rect 41786 793047 41842 793056
rect 41800 792744 41828 793047
rect 41786 790664 41842 790673
rect 41786 790599 41842 790608
rect 41800 790228 41828 790599
rect 42536 789630 42564 801042
rect 42812 799354 42840 801766
rect 42720 799338 42840 799354
rect 42708 799332 42840 799338
rect 42760 799326 42840 799332
rect 42708 799274 42760 799280
rect 42182 789602 42564 789630
rect 41786 789440 41842 789449
rect 41786 789375 41842 789384
rect 41800 788936 41828 789375
rect 42616 789336 42668 789342
rect 42616 789278 42668 789284
rect 42246 789168 42302 789177
rect 42246 789103 42302 789112
rect 42260 788406 42288 789103
rect 42430 788760 42486 788769
rect 42430 788695 42486 788704
rect 42182 788378 42288 788406
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 42260 786570 42288 788151
rect 42182 786542 42288 786570
rect 42444 785958 42472 788695
rect 42628 786842 42656 789278
rect 42168 785890 42196 785944
rect 42260 785930 42472 785958
rect 42536 786814 42656 786842
rect 42260 785890 42288 785930
rect 42168 785862 42288 785890
rect 42536 785278 42564 786814
rect 42708 786684 42760 786690
rect 42708 786626 42760 786632
rect 42182 785250 42564 785278
rect 42720 784802 42748 786626
rect 42536 784774 42748 784802
rect 42536 784734 42564 784774
rect 42182 784706 42564 784734
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 774752 35862 774761
rect 35806 774687 35862 774696
rect 35820 774246 35848 774687
rect 35808 774240 35860 774246
rect 35808 774182 35860 774188
rect 41696 774240 41748 774246
rect 42064 774240 42116 774246
rect 41748 774188 42064 774194
rect 41696 774182 42116 774188
rect 41708 774166 42104 774182
rect 35254 773936 35310 773945
rect 35254 773871 35310 773880
rect 35268 772886 35296 773871
rect 35622 773528 35678 773537
rect 35622 773463 35678 773472
rect 35440 773424 35492 773430
rect 35440 773366 35492 773372
rect 35452 773129 35480 773366
rect 35438 773120 35494 773129
rect 35438 773055 35494 773064
rect 35636 773022 35664 773463
rect 41512 773424 41564 773430
rect 41512 773366 41564 773372
rect 35808 773152 35860 773158
rect 35806 773120 35808 773129
rect 41524 773129 41552 773366
rect 41708 773226 42104 773242
rect 42904 773226 42932 815730
rect 44180 815652 44232 815658
rect 44180 815594 44232 815600
rect 43444 814428 43496 814434
rect 43444 814370 43496 814376
rect 43076 811504 43128 811510
rect 43076 811446 43128 811452
rect 43088 789342 43116 811446
rect 43260 807492 43312 807498
rect 43260 807434 43312 807440
rect 43076 789336 43128 789342
rect 43076 789278 43128 789284
rect 41696 773220 42116 773226
rect 41748 773214 42064 773220
rect 41696 773162 41748 773168
rect 42064 773162 42116 773168
rect 42892 773220 42944 773226
rect 42892 773162 42944 773168
rect 35860 773120 35862 773129
rect 35806 773055 35862 773064
rect 41510 773120 41566 773129
rect 41708 773090 42104 773106
rect 41510 773055 41566 773064
rect 41696 773084 42116 773090
rect 41748 773078 42064 773084
rect 41696 773026 41748 773032
rect 42064 773026 42116 773032
rect 35624 773016 35676 773022
rect 35624 772958 35676 772964
rect 35256 772880 35308 772886
rect 35256 772822 35308 772828
rect 41696 772880 41748 772886
rect 42064 772880 42116 772886
rect 41748 772828 42064 772834
rect 41696 772822 42116 772828
rect 41708 772806 42104 772822
rect 35622 772304 35678 772313
rect 35622 772239 35678 772248
rect 40314 772304 40370 772313
rect 40314 772239 40370 772248
rect 35636 771594 35664 772239
rect 35806 771896 35862 771905
rect 35806 771831 35808 771840
rect 35860 771831 35862 771840
rect 39948 771860 40000 771866
rect 35808 771802 35860 771808
rect 39948 771802 40000 771808
rect 35624 771588 35676 771594
rect 35624 771530 35676 771536
rect 39960 771497 39988 771802
rect 40328 771662 40356 772239
rect 40316 771656 40368 771662
rect 40316 771598 40368 771604
rect 42064 771520 42116 771526
rect 35806 771488 35862 771497
rect 35806 771423 35808 771432
rect 35860 771423 35862 771432
rect 39946 771488 40002 771497
rect 41708 771468 42064 771474
rect 41708 771462 42116 771468
rect 41708 771458 42104 771462
rect 39946 771423 40002 771432
rect 41696 771452 42104 771458
rect 35808 771394 35860 771400
rect 41748 771446 42104 771452
rect 41696 771394 41748 771400
rect 35438 771080 35494 771089
rect 35438 771015 35494 771024
rect 35452 770234 35480 771015
rect 35622 770672 35678 770681
rect 35622 770607 35678 770616
rect 35440 770228 35492 770234
rect 35440 770170 35492 770176
rect 35636 770098 35664 770607
rect 35808 770500 35860 770506
rect 35808 770442 35860 770448
rect 40316 770500 40368 770506
rect 40316 770442 40368 770448
rect 35820 770273 35848 770442
rect 40328 770273 40356 770442
rect 41696 770296 41748 770302
rect 35806 770264 35862 770273
rect 35806 770199 35862 770208
rect 40314 770264 40370 770273
rect 42064 770296 42116 770302
rect 41748 770244 42064 770250
rect 41696 770238 42116 770244
rect 43076 770296 43128 770302
rect 43076 770238 43128 770244
rect 41708 770222 42104 770238
rect 40314 770199 40370 770208
rect 42064 770160 42116 770166
rect 41708 770108 42064 770114
rect 41708 770102 42116 770108
rect 41708 770098 42104 770102
rect 35624 770092 35676 770098
rect 35624 770034 35676 770040
rect 41696 770092 42104 770098
rect 41748 770086 42104 770092
rect 41696 770034 41748 770040
rect 35622 769448 35678 769457
rect 35622 769383 35678 769392
rect 35636 768738 35664 769383
rect 35808 768868 35860 768874
rect 35808 768810 35860 768816
rect 40040 768868 40092 768874
rect 40040 768810 40092 768816
rect 35624 768732 35676 768738
rect 35624 768674 35676 768680
rect 35820 768641 35848 768810
rect 35806 768632 35862 768641
rect 35806 768567 35862 768576
rect 35162 768224 35218 768233
rect 35162 768159 35218 768168
rect 32402 767816 32458 767825
rect 32402 767751 32458 767760
rect 32416 759694 32444 767751
rect 33782 767000 33838 767009
rect 33782 766935 33838 766944
rect 32404 759688 32456 759694
rect 32404 759630 32456 759636
rect 33796 758334 33824 766935
rect 35176 759830 35204 768159
rect 35808 767644 35860 767650
rect 35808 767586 35860 767592
rect 36544 767644 36596 767650
rect 36544 767586 36596 767592
rect 35820 767417 35848 767586
rect 35806 767408 35862 767417
rect 35806 767343 35862 767352
rect 35806 766592 35862 766601
rect 35806 766527 35862 766536
rect 35820 766086 35848 766527
rect 35808 766080 35860 766086
rect 35808 766022 35860 766028
rect 35622 765776 35678 765785
rect 35622 765711 35678 765720
rect 35636 764590 35664 765711
rect 35808 764856 35860 764862
rect 35808 764798 35860 764804
rect 35624 764584 35676 764590
rect 35820 764561 35848 764798
rect 35624 764526 35676 764532
rect 35806 764552 35862 764561
rect 35806 764487 35862 764496
rect 35622 764144 35678 764153
rect 35622 764079 35678 764088
rect 35636 763502 35664 764079
rect 35806 763736 35862 763745
rect 35806 763671 35862 763680
rect 35624 763496 35676 763502
rect 35624 763438 35676 763444
rect 35820 763230 35848 763671
rect 35808 763224 35860 763230
rect 35808 763166 35860 763172
rect 35806 762920 35862 762929
rect 35806 762855 35862 762864
rect 35820 761870 35848 762855
rect 35808 761864 35860 761870
rect 35808 761806 35860 761812
rect 35164 759824 35216 759830
rect 35164 759766 35216 759772
rect 33784 758328 33836 758334
rect 33784 758270 33836 758276
rect 36556 757761 36584 767586
rect 39396 766080 39448 766086
rect 39396 766022 39448 766028
rect 39408 764561 39436 766022
rect 40052 765338 40080 768810
rect 41696 768732 41748 768738
rect 41696 768674 41748 768680
rect 41708 765914 41736 768674
rect 43088 765914 43116 770238
rect 41708 765886 42288 765914
rect 43088 765886 43208 765914
rect 40040 765332 40092 765338
rect 40040 765274 40092 765280
rect 41696 765332 41748 765338
rect 41696 765274 41748 765280
rect 41708 765218 41736 765274
rect 41708 765202 42104 765218
rect 41708 765196 42116 765202
rect 41708 765190 42064 765196
rect 42064 765138 42116 765144
rect 39948 764856 40000 764862
rect 39948 764798 40000 764804
rect 39394 764552 39450 764561
rect 39394 764487 39450 764496
rect 39960 764153 39988 764798
rect 41708 764658 42104 764674
rect 41696 764652 42116 764658
rect 41748 764646 42064 764652
rect 41696 764594 41748 764600
rect 42064 764594 42116 764600
rect 39946 764144 40002 764153
rect 39946 764079 40002 764088
rect 39948 763496 40000 763502
rect 39948 763438 40000 763444
rect 39960 763337 39988 763438
rect 42064 763428 42116 763434
rect 42064 763370 42116 763376
rect 39946 763328 40002 763337
rect 42076 763314 42104 763370
rect 39946 763263 40002 763272
rect 41708 763286 42104 763314
rect 41708 763162 41736 763286
rect 41696 763156 41748 763162
rect 41696 763098 41748 763104
rect 42064 761932 42116 761938
rect 42064 761874 42116 761880
rect 41696 761864 41748 761870
rect 42076 761818 42104 761874
rect 41748 761812 42104 761818
rect 41696 761806 42104 761812
rect 41708 761790 42104 761806
rect 39672 759824 39724 759830
rect 39672 759766 39724 759772
rect 39684 758033 39712 759766
rect 41604 759688 41656 759694
rect 41656 759636 41828 759642
rect 41604 759630 41828 759636
rect 41616 759614 41828 759630
rect 39948 758328 40000 758334
rect 39946 758296 39948 758305
rect 40000 758296 40002 758305
rect 39946 758231 40002 758240
rect 39670 758024 39726 758033
rect 39670 757959 39726 757968
rect 36542 757752 36598 757761
rect 36542 757687 36598 757696
rect 41800 757081 41828 759614
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 41878 756664 41934 756673
rect 41878 756599 41934 756608
rect 41892 756226 41920 756599
rect 42260 754882 42288 765886
rect 42432 765196 42484 765202
rect 42432 765138 42484 765144
rect 42444 765082 42472 765138
rect 42352 765054 42472 765082
rect 42352 763154 42380 765054
rect 42352 763126 42840 763154
rect 42614 758296 42670 758305
rect 42614 758231 42670 758240
rect 42430 758024 42486 758033
rect 42430 757959 42486 757968
rect 42168 754854 42288 754882
rect 42168 754392 42196 754854
rect 41878 754216 41934 754225
rect 41934 754174 42380 754202
rect 41878 754151 41934 754160
rect 42062 754080 42118 754089
rect 42062 754015 42118 754024
rect 42076 753780 42104 754015
rect 42154 753536 42210 753545
rect 42154 753471 42210 753480
rect 42168 753386 42196 753471
rect 42168 753358 42288 753386
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42076 751641 42104 751944
rect 42062 751632 42118 751641
rect 42062 751567 42118 751576
rect 42076 751233 42104 751369
rect 42062 751224 42118 751233
rect 42062 751159 42118 751168
rect 42260 751074 42288 753358
rect 42168 751046 42288 751074
rect 42168 750720 42196 751046
rect 42062 750408 42118 750417
rect 42062 750343 42118 750352
rect 42076 750108 42104 750343
rect 42352 749986 42380 754174
rect 42444 753522 42472 757959
rect 42628 753778 42656 758231
rect 42616 753772 42668 753778
rect 42616 753714 42668 753720
rect 42616 753636 42668 753642
rect 42616 753578 42668 753584
rect 42444 753494 42564 753522
rect 42260 749958 42380 749986
rect 42260 749766 42288 749958
rect 42248 749760 42300 749766
rect 42248 749702 42300 749708
rect 42168 749442 42196 749529
rect 42168 749414 42380 749442
rect 42352 749306 42380 749414
rect 42536 749306 42564 753494
rect 42352 749278 42564 749306
rect 42248 749216 42300 749222
rect 42248 749158 42300 749164
rect 42260 747130 42288 749158
rect 42168 747102 42288 747130
rect 42168 747048 42196 747102
rect 41786 746736 41842 746745
rect 41786 746671 41842 746680
rect 41800 746401 41828 746671
rect 42628 746594 42656 753578
rect 42812 753494 42840 763126
rect 42982 753536 43038 753545
rect 42536 746586 42656 746594
rect 42352 746566 42656 746586
rect 42720 753466 42840 753494
rect 42904 753480 42982 753494
rect 42904 753471 43038 753480
rect 42904 753466 43024 753471
rect 42352 746558 42564 746566
rect 42352 745770 42380 746558
rect 42720 745906 42748 753466
rect 42904 753001 42932 753466
rect 42890 752992 42946 753001
rect 42890 752927 42946 752936
rect 43180 746594 43208 765886
rect 42182 745742 42380 745770
rect 42444 745878 42748 745906
rect 43088 746566 43208 746594
rect 42444 745634 42472 745878
rect 42614 745784 42670 745793
rect 42614 745719 42670 745728
rect 42076 745606 42472 745634
rect 42076 745212 42104 745606
rect 42246 745512 42302 745521
rect 42628 745498 42656 745719
rect 42246 745447 42302 745456
rect 42444 745470 42656 745498
rect 42260 745346 42288 745447
rect 42248 745340 42300 745346
rect 42248 745282 42300 745288
rect 42248 745136 42300 745142
rect 42248 745078 42300 745084
rect 42260 743730 42288 745078
rect 42168 743702 42288 743730
rect 42168 743376 42196 743702
rect 42168 742750 42288 742778
rect 42168 742696 42196 742750
rect 42260 742710 42288 742750
rect 42444 742710 42472 745470
rect 42614 745104 42670 745113
rect 42614 745039 42670 745048
rect 42260 742682 42472 742710
rect 42628 742098 42656 745039
rect 42800 744048 42852 744054
rect 42182 742070 42656 742098
rect 42720 743996 42800 744002
rect 42720 743990 42852 743996
rect 42720 743974 42840 743990
rect 42720 741690 42748 743974
rect 42536 741662 42748 741690
rect 42536 741554 42564 741662
rect 42182 741526 42564 741554
rect 43088 741074 43116 746566
rect 42996 741046 43116 741074
rect 40406 732320 40462 732329
rect 40406 732255 40462 732264
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 40038 731640 40094 731649
rect 40038 731575 40094 731584
rect 35438 731368 35494 731377
rect 35438 731303 35494 731312
rect 35452 730114 35480 731303
rect 35808 731196 35860 731202
rect 35808 731138 35860 731144
rect 35820 730969 35848 731138
rect 35806 730960 35862 730969
rect 35806 730895 35862 730904
rect 35622 730552 35678 730561
rect 35622 730487 35678 730496
rect 35440 730108 35492 730114
rect 35440 730050 35492 730056
rect 35438 729736 35494 729745
rect 35438 729671 35494 729680
rect 35452 728686 35480 729671
rect 35636 729502 35664 730487
rect 35808 730380 35860 730386
rect 35808 730322 35860 730328
rect 35820 730153 35848 730322
rect 35806 730144 35862 730153
rect 35806 730079 35862 730088
rect 35624 729496 35676 729502
rect 35624 729438 35676 729444
rect 35622 729328 35678 729337
rect 35622 729263 35678 729272
rect 35636 728822 35664 729263
rect 35808 729088 35860 729094
rect 35808 729030 35860 729036
rect 35820 728929 35848 729030
rect 35806 728920 35862 728929
rect 35806 728855 35862 728864
rect 35624 728816 35676 728822
rect 35624 728758 35676 728764
rect 35440 728680 35492 728686
rect 35440 728622 35492 728628
rect 35806 728512 35862 728521
rect 35806 728447 35862 728456
rect 35438 728104 35494 728113
rect 35438 728039 35494 728048
rect 35452 727598 35480 728039
rect 35820 727870 35848 728447
rect 40052 727870 40080 731575
rect 40420 730386 40448 732255
rect 42996 731649 43024 741046
rect 42982 731640 43038 731649
rect 42982 731575 43038 731584
rect 41696 731128 41748 731134
rect 41694 731096 41696 731105
rect 41748 731096 41750 731105
rect 41694 731031 41750 731040
rect 40408 730380 40460 730386
rect 40408 730322 40460 730328
rect 41708 730114 42104 730130
rect 41696 730108 42116 730114
rect 41748 730102 42064 730108
rect 41696 730050 41748 730056
rect 42064 730050 42116 730056
rect 42064 729360 42116 729366
rect 41708 729308 42064 729314
rect 41708 729302 42116 729308
rect 41708 729298 42104 729302
rect 41696 729292 42104 729298
rect 41748 729286 42104 729292
rect 41696 729234 41748 729240
rect 41512 729088 41564 729094
rect 41512 729030 41564 729036
rect 41524 728226 41552 729030
rect 42064 728884 42116 728890
rect 42064 728826 42116 728832
rect 41696 728816 41748 728822
rect 42076 728770 42104 728826
rect 41748 728764 42104 728770
rect 41696 728758 42104 728764
rect 41708 728742 42104 728758
rect 41696 728680 41748 728686
rect 42064 728680 42116 728686
rect 41748 728628 42064 728634
rect 41696 728622 42116 728628
rect 41708 728606 42104 728622
rect 41694 728240 41750 728249
rect 41524 728198 41694 728226
rect 41694 728175 41750 728184
rect 35808 727864 35860 727870
rect 35808 727806 35860 727812
rect 40040 727864 40092 727870
rect 40040 727806 40092 727812
rect 41694 727832 41750 727841
rect 41694 727767 41750 727776
rect 43074 727832 43130 727841
rect 43074 727767 43130 727776
rect 35622 727696 35678 727705
rect 41708 727666 41736 727767
rect 35622 727631 35678 727640
rect 41696 727660 41748 727666
rect 35440 727592 35492 727598
rect 35440 727534 35492 727540
rect 35636 727326 35664 727631
rect 41696 727602 41748 727608
rect 35808 727456 35860 727462
rect 35808 727398 35860 727404
rect 41696 727456 41748 727462
rect 42064 727456 42116 727462
rect 41748 727404 42064 727410
rect 41696 727398 42116 727404
rect 35624 727320 35676 727326
rect 35820 727297 35848 727398
rect 41708 727382 42104 727398
rect 41696 727320 41748 727326
rect 35624 727262 35676 727268
rect 35806 727288 35862 727297
rect 42064 727320 42116 727326
rect 41748 727268 42064 727274
rect 41696 727262 42116 727268
rect 41708 727246 42104 727262
rect 35806 727223 35862 727232
rect 41142 726880 41198 726889
rect 41142 726815 41198 726824
rect 41156 725966 41184 726815
rect 41326 726472 41382 726481
rect 41326 726407 41382 726416
rect 41340 726102 41368 726407
rect 41328 726096 41380 726102
rect 41328 726038 41380 726044
rect 41696 726096 41748 726102
rect 42064 726096 42116 726102
rect 41748 726056 42064 726084
rect 41696 726038 41748 726044
rect 42064 726038 42116 726044
rect 42524 726096 42576 726102
rect 42524 726038 42576 726044
rect 41144 725960 41196 725966
rect 41144 725902 41196 725908
rect 41604 725960 41656 725966
rect 41604 725902 41656 725908
rect 40958 725656 41014 725665
rect 41616 725642 41644 725902
rect 41786 725656 41842 725665
rect 41616 725614 41786 725642
rect 40958 725591 41014 725600
rect 41786 725591 41842 725600
rect 32402 725248 32458 725257
rect 32402 725183 32458 725192
rect 31666 724024 31722 724033
rect 31666 723959 31722 723968
rect 31680 715562 31708 723959
rect 32416 716922 32444 725183
rect 35162 724840 35218 724849
rect 35162 724775 35218 724784
rect 32404 716916 32456 716922
rect 32404 716858 32456 716864
rect 35176 715766 35204 724775
rect 37278 724432 37334 724441
rect 37278 724367 37334 724376
rect 37292 716961 37320 724367
rect 39302 723208 39358 723217
rect 39302 723143 39358 723152
rect 37278 716952 37334 716961
rect 37278 716887 37334 716896
rect 35164 715760 35216 715766
rect 35164 715702 35216 715708
rect 31668 715556 31720 715562
rect 31668 715498 31720 715504
rect 39316 714241 39344 723143
rect 40590 715864 40646 715873
rect 40590 715799 40646 715808
rect 40604 715562 40632 715799
rect 40592 715556 40644 715562
rect 40592 715498 40644 715504
rect 40972 714921 41000 725591
rect 41786 722392 41842 722401
rect 41786 722327 41842 722336
rect 41800 718593 41828 722327
rect 41786 718584 41842 718593
rect 41786 718519 41842 718528
rect 41696 716916 41748 716922
rect 41696 716858 41748 716864
rect 41708 716802 41736 716858
rect 41708 716786 42104 716802
rect 41708 716780 42116 716786
rect 41708 716774 42064 716780
rect 42064 716722 42116 716728
rect 42536 716650 42564 726038
rect 42890 721168 42946 721177
rect 42890 721103 42946 721112
rect 42708 716780 42760 716786
rect 42708 716722 42760 716728
rect 42064 716644 42116 716650
rect 42064 716586 42116 716592
rect 42524 716644 42576 716650
rect 42524 716586 42576 716592
rect 41328 715760 41380 715766
rect 41380 715708 41552 715714
rect 41328 715702 41552 715708
rect 41340 715686 41552 715702
rect 40958 714912 41014 714921
rect 40958 714847 41014 714856
rect 39302 714232 39358 714241
rect 41524 714218 41552 715686
rect 42076 715034 42104 716586
rect 42430 715864 42486 715873
rect 42486 715822 42656 715850
rect 42430 715799 42486 715808
rect 42076 715006 42564 715034
rect 42338 714912 42394 714921
rect 42338 714854 42394 714856
rect 42260 714847 42394 714854
rect 42260 714826 42380 714847
rect 42260 714377 42288 714826
rect 42536 714762 42564 715006
rect 42352 714734 42564 714762
rect 42352 714456 42380 714734
rect 42352 714428 42472 714456
rect 42246 714368 42302 714377
rect 42246 714303 42302 714312
rect 41524 714190 42288 714218
rect 39302 714167 39358 714176
rect 42260 713062 42288 714190
rect 42444 713062 42472 714428
rect 42182 713034 42288 713062
rect 42352 713034 42472 713062
rect 42352 711226 42380 713034
rect 42182 711198 42380 711226
rect 42154 710832 42210 710841
rect 42154 710767 42210 710776
rect 42168 710561 42196 710767
rect 42248 710456 42300 710462
rect 42248 710398 42300 710404
rect 41786 709880 41842 709889
rect 41786 709815 41842 709824
rect 41800 709376 41828 709815
rect 42076 708529 42104 708696
rect 42062 708520 42118 708529
rect 42062 708455 42118 708464
rect 42260 708234 42288 710398
rect 42628 708506 42656 715822
rect 42720 714854 42748 716722
rect 42720 714826 42840 714854
rect 42168 708206 42288 708234
rect 42536 708478 42656 708506
rect 42168 708152 42196 708206
rect 42248 707872 42300 707878
rect 42248 707814 42300 707820
rect 42260 707554 42288 707814
rect 42182 707526 42288 707554
rect 42248 707464 42300 707470
rect 42248 707406 42300 707412
rect 41786 707160 41842 707169
rect 41786 707095 41842 707104
rect 41800 706860 41828 707095
rect 42260 706330 42288 707406
rect 42536 706722 42564 708478
rect 42812 707554 42840 714826
rect 42720 707526 42840 707554
rect 42720 707470 42748 707526
rect 42708 707464 42760 707470
rect 42708 707406 42760 707412
rect 42524 706716 42576 706722
rect 42524 706658 42576 706664
rect 42708 706512 42760 706518
rect 42708 706454 42760 706460
rect 42182 706302 42288 706330
rect 42430 706344 42486 706353
rect 42430 706279 42486 706288
rect 42248 705560 42300 705566
rect 42248 705502 42300 705508
rect 41786 704304 41842 704313
rect 41786 704239 41842 704248
rect 41800 703868 41828 704239
rect 42260 703746 42288 705502
rect 42076 703718 42288 703746
rect 42076 703188 42104 703718
rect 42062 703080 42118 703089
rect 42062 703015 42118 703024
rect 42076 702576 42104 703015
rect 42444 702046 42472 706279
rect 42720 705194 42748 706454
rect 42628 705166 42748 705194
rect 42628 703089 42656 705166
rect 42614 703080 42670 703089
rect 42614 703015 42670 703024
rect 42168 701978 42196 702032
rect 42260 702018 42472 702046
rect 42260 701978 42288 702018
rect 42168 701950 42288 701978
rect 42522 701856 42578 701865
rect 42352 701814 42522 701842
rect 41878 700496 41934 700505
rect 41878 700431 41934 700440
rect 41892 700165 41920 700431
rect 42352 699530 42380 701814
rect 42522 701791 42578 701800
rect 42522 701584 42578 701593
rect 42522 701519 42578 701528
rect 42182 699502 42380 699530
rect 42536 699394 42564 701519
rect 42708 701140 42760 701146
rect 42708 701082 42760 701088
rect 42352 699366 42564 699394
rect 42352 698918 42380 699366
rect 42168 698850 42196 698904
rect 42260 698890 42380 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 42720 698339 42748 701082
rect 42182 698311 42748 698339
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35438 688392 35494 688401
rect 35438 688327 35494 688336
rect 35452 687274 35480 688327
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 35820 687546 35848 687647
rect 41694 687576 41750 687585
rect 35808 687540 35860 687546
rect 41694 687511 41696 687520
rect 35808 687482 35860 687488
rect 41748 687511 41750 687520
rect 41696 687482 41748 687488
rect 35622 687304 35678 687313
rect 35440 687268 35492 687274
rect 35622 687239 35678 687248
rect 35440 687210 35492 687216
rect 35438 686896 35494 686905
rect 35438 686831 35494 686840
rect 35452 686050 35480 686831
rect 35636 686458 35664 687239
rect 41696 687200 41748 687206
rect 41694 687168 41696 687177
rect 41748 687168 41750 687177
rect 41694 687103 41750 687112
rect 42064 686520 42116 686526
rect 35806 686488 35862 686497
rect 35624 686452 35676 686458
rect 41708 686468 42064 686474
rect 41708 686462 42116 686468
rect 41708 686458 42104 686462
rect 35806 686423 35862 686432
rect 41696 686452 42104 686458
rect 35624 686394 35676 686400
rect 35820 686322 35848 686423
rect 41748 686446 42104 686452
rect 41696 686394 41748 686400
rect 41708 686322 42104 686338
rect 35808 686316 35860 686322
rect 35808 686258 35860 686264
rect 41696 686316 42116 686322
rect 41748 686310 42064 686316
rect 41696 686258 41748 686264
rect 42064 686258 42116 686264
rect 42064 686112 42116 686118
rect 35806 686080 35862 686089
rect 35440 686044 35492 686050
rect 41708 686060 42064 686066
rect 41708 686054 42116 686060
rect 41708 686050 42104 686054
rect 35806 686015 35862 686024
rect 41696 686044 42104 686050
rect 35440 685986 35492 685992
rect 35820 685914 35848 686015
rect 41748 686038 42104 686044
rect 41696 685986 41748 685992
rect 41708 685914 42104 685930
rect 35808 685908 35860 685914
rect 35808 685850 35860 685856
rect 41696 685908 42116 685914
rect 41748 685902 42064 685908
rect 41696 685850 41748 685856
rect 42064 685850 42116 685856
rect 35806 685672 35862 685681
rect 35806 685607 35862 685616
rect 35622 685264 35678 685273
rect 35622 685199 35678 685208
rect 35636 684690 35664 685199
rect 35820 685030 35848 685607
rect 35808 685024 35860 685030
rect 35808 684966 35860 684972
rect 41696 684956 41748 684962
rect 41696 684898 41748 684904
rect 35806 684856 35862 684865
rect 41708 684842 41736 684898
rect 41708 684814 42104 684842
rect 35806 684791 35862 684800
rect 35624 684684 35676 684690
rect 35624 684626 35676 684632
rect 35820 684554 35848 684791
rect 41694 684720 41750 684729
rect 41694 684655 41696 684664
rect 41748 684655 41750 684664
rect 41696 684626 41748 684632
rect 42076 684554 42104 684814
rect 42248 684820 42300 684826
rect 42248 684762 42300 684768
rect 35808 684548 35860 684554
rect 35808 684490 35860 684496
rect 41696 684548 41748 684554
rect 41696 684490 41748 684496
rect 42064 684548 42116 684554
rect 42064 684490 42116 684496
rect 35622 684448 35678 684457
rect 41708 684434 41736 684490
rect 42260 684434 42288 684762
rect 41708 684406 42288 684434
rect 35622 684383 35678 684392
rect 35438 684040 35494 684049
rect 35438 683975 35494 683984
rect 35452 683194 35480 683975
rect 35636 683330 35664 684383
rect 41694 683904 41750 683913
rect 41524 683862 41694 683890
rect 35808 683460 35860 683466
rect 35808 683402 35860 683408
rect 35624 683324 35676 683330
rect 35624 683266 35676 683272
rect 35820 683233 35848 683402
rect 41524 683330 41552 683862
rect 41694 683839 41750 683848
rect 41696 683460 41748 683466
rect 41696 683402 41748 683408
rect 41708 683346 41736 683402
rect 41512 683324 41564 683330
rect 41708 683318 41920 683346
rect 41512 683266 41564 683272
rect 35806 683224 35862 683233
rect 35440 683188 35492 683194
rect 35806 683159 35862 683168
rect 35440 683130 35492 683136
rect 41696 683120 41748 683126
rect 41694 683088 41696 683097
rect 41748 683088 41750 683097
rect 41694 683023 41750 683032
rect 35622 682816 35678 682825
rect 35622 682751 35678 682760
rect 35162 682000 35218 682009
rect 35162 681935 35218 681944
rect 33046 681592 33102 681601
rect 33046 681527 33102 681536
rect 31022 680776 31078 680785
rect 31022 680711 31078 680720
rect 31036 672518 31064 680711
rect 33060 674150 33088 681527
rect 33782 681184 33838 681193
rect 33782 681119 33838 681128
rect 33048 674144 33100 674150
rect 33048 674086 33100 674092
rect 33796 672761 33824 681119
rect 35176 672858 35204 681935
rect 35636 681902 35664 682751
rect 35806 682408 35862 682417
rect 35806 682343 35862 682352
rect 35624 681896 35676 681902
rect 35624 681838 35676 681844
rect 35820 681766 35848 682343
rect 41696 681896 41748 681902
rect 41696 681838 41748 681844
rect 35808 681760 35860 681766
rect 35808 681702 35860 681708
rect 41512 681760 41564 681766
rect 41512 681702 41564 681708
rect 41524 681034 41552 681702
rect 41708 681465 41736 681838
rect 41694 681456 41750 681465
rect 41694 681391 41750 681400
rect 41694 681048 41750 681057
rect 41524 681006 41694 681034
rect 41694 680983 41750 680992
rect 35808 680536 35860 680542
rect 35808 680478 35860 680484
rect 41696 680536 41748 680542
rect 41696 680478 41748 680484
rect 35820 680377 35848 680478
rect 35806 680368 35862 680377
rect 35806 680303 35862 680312
rect 41708 680241 41736 680478
rect 41694 680232 41750 680241
rect 41694 680167 41750 680176
rect 35806 679960 35862 679969
rect 35806 679895 35862 679904
rect 35622 679552 35678 679561
rect 35622 679487 35678 679496
rect 35636 679046 35664 679487
rect 35820 679454 35848 679895
rect 35808 679448 35860 679454
rect 41696 679448 41748 679454
rect 35808 679390 35860 679396
rect 41694 679416 41696 679425
rect 41748 679416 41750 679425
rect 41694 679351 41750 679360
rect 35808 679176 35860 679182
rect 35806 679144 35808 679153
rect 41512 679176 41564 679182
rect 35860 679144 35862 679153
rect 41512 679118 41564 679124
rect 35806 679079 35862 679088
rect 35624 679040 35676 679046
rect 35624 678982 35676 678988
rect 41524 678586 41552 679118
rect 41696 679040 41748 679046
rect 41694 679008 41696 679017
rect 41748 679008 41750 679017
rect 41694 678943 41750 678952
rect 41892 678974 41920 683318
rect 42706 681048 42762 681057
rect 42706 680983 42762 680992
rect 41892 678946 42288 678974
rect 41694 678600 41750 678609
rect 41524 678558 41694 678586
rect 41694 678535 41750 678544
rect 41512 674144 41564 674150
rect 41512 674086 41564 674092
rect 35164 672852 35216 672858
rect 35164 672794 35216 672800
rect 33782 672752 33838 672761
rect 33782 672687 33838 672696
rect 31024 672512 31076 672518
rect 31024 672454 31076 672460
rect 41524 672058 41552 674086
rect 41696 672852 41748 672858
rect 41696 672794 41748 672800
rect 41708 672738 41736 672794
rect 41708 672722 42104 672738
rect 41708 672716 42116 672722
rect 41708 672710 42064 672716
rect 42064 672658 42116 672664
rect 42260 672625 42288 678946
rect 42524 672716 42576 672722
rect 42524 672658 42576 672664
rect 42246 672616 42302 672625
rect 42536 672602 42564 672658
rect 42536 672574 42656 672602
rect 42246 672551 42302 672560
rect 41696 672512 41748 672518
rect 41748 672460 42564 672466
rect 41696 672454 42564 672460
rect 41708 672438 42564 672454
rect 41524 672030 42288 672058
rect 42168 669746 42196 669868
rect 42260 669746 42288 672030
rect 42168 669718 42288 669746
rect 41970 668536 42026 668545
rect 41970 668471 42026 668480
rect 41984 668032 42012 668471
rect 42062 667720 42118 667729
rect 42062 667655 42118 667664
rect 42076 667352 42104 667655
rect 42062 667176 42118 667185
rect 42118 667134 42472 667162
rect 42062 667111 42118 667120
rect 42248 667072 42300 667078
rect 42248 667014 42300 667020
rect 42062 666632 42118 666641
rect 42062 666567 42118 666576
rect 42076 666165 42104 666567
rect 42260 665530 42288 667014
rect 42182 665502 42288 665530
rect 41786 665136 41842 665145
rect 41786 665071 41842 665080
rect 41800 664972 41828 665071
rect 42444 664339 42472 667134
rect 42182 664311 42472 664339
rect 42536 664204 42564 672438
rect 42260 664176 42564 664204
rect 41786 664048 41842 664057
rect 41786 663983 41842 663992
rect 41800 663680 41828 663983
rect 42260 663338 42288 664176
rect 42248 663332 42300 663338
rect 42248 663274 42300 663280
rect 42628 663218 42656 672574
rect 42352 663190 42656 663218
rect 42352 663150 42380 663190
rect 42182 663122 42380 663150
rect 42524 663128 42576 663134
rect 42524 663070 42576 663076
rect 42248 662992 42300 662998
rect 42248 662934 42300 662940
rect 42260 661178 42288 662934
rect 42260 661150 42380 661178
rect 42156 661088 42208 661094
rect 42156 661030 42208 661036
rect 42168 660620 42196 661030
rect 42352 660022 42380 661150
rect 42182 659994 42380 660022
rect 42536 659371 42564 663070
rect 42182 659343 42564 659371
rect 42168 658838 42380 658866
rect 42168 658784 42196 658838
rect 42352 658798 42380 658838
rect 42720 658798 42748 680983
rect 42352 658770 42748 658798
rect 42522 658608 42578 658617
rect 42352 658566 42522 658594
rect 41800 658430 42288 658458
rect 41800 658345 41828 658430
rect 41786 658336 41842 658345
rect 41786 658271 41842 658280
rect 41786 657248 41842 657257
rect 41786 657183 41842 657192
rect 41800 656948 41828 657183
rect 42260 656350 42288 658430
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42352 655670 42380 658566
rect 42522 658543 42578 658552
rect 42524 657552 42576 657558
rect 42524 657494 42576 657500
rect 42260 655642 42380 655670
rect 42536 655126 42564 657494
rect 42182 655098 42564 655126
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 35820 644502 35848 644671
rect 35808 644496 35860 644502
rect 35808 644438 35860 644444
rect 41696 644496 41748 644502
rect 42064 644496 42116 644502
rect 41748 644446 42064 644474
rect 41696 644438 41748 644444
rect 42064 644438 42116 644444
rect 38566 644328 38622 644337
rect 38566 644263 38622 644272
rect 35346 643920 35402 643929
rect 35346 643855 35402 643864
rect 35360 643142 35388 643855
rect 35808 643544 35860 643550
rect 35530 643512 35586 643521
rect 35530 643447 35586 643456
rect 35806 643512 35808 643521
rect 35860 643512 35862 643521
rect 35806 643447 35862 643456
rect 35544 643278 35572 643447
rect 35532 643272 35584 643278
rect 35532 643214 35584 643220
rect 35348 643136 35400 643142
rect 35348 643078 35400 643084
rect 35438 642696 35494 642705
rect 35438 642631 35494 642640
rect 35806 642696 35862 642705
rect 35806 642631 35862 642640
rect 35452 641918 35480 642631
rect 35622 642288 35678 642297
rect 35622 642223 35678 642232
rect 35440 641912 35492 641918
rect 35440 641854 35492 641860
rect 35636 641782 35664 642223
rect 35820 642190 35848 642631
rect 38580 642530 38608 644263
rect 41144 643544 41196 643550
rect 41144 643486 41196 643492
rect 38568 642524 38620 642530
rect 38568 642466 38620 642472
rect 35808 642184 35860 642190
rect 35808 642126 35860 642132
rect 39396 642184 39448 642190
rect 39396 642126 39448 642132
rect 35624 641776 35676 641782
rect 35624 641718 35676 641724
rect 35806 641472 35862 641481
rect 35806 641407 35862 641416
rect 35622 641064 35678 641073
rect 35622 640999 35678 641008
rect 35636 640490 35664 640999
rect 35820 640830 35848 641407
rect 35808 640824 35860 640830
rect 35808 640766 35860 640772
rect 35806 640656 35862 640665
rect 35806 640591 35862 640600
rect 35624 640484 35676 640490
rect 35624 640426 35676 640432
rect 35820 640354 35848 640591
rect 35808 640348 35860 640354
rect 35808 640290 35860 640296
rect 39408 639849 39436 642126
rect 41156 641073 41184 643486
rect 41708 643346 42104 643362
rect 41696 643340 42116 643346
rect 41748 643334 42064 643340
rect 41696 643282 41748 643288
rect 42064 643282 42116 643288
rect 41696 643136 41748 643142
rect 42064 643136 42116 643142
rect 41748 643084 42064 643090
rect 41696 643078 42116 643084
rect 41708 643062 42104 643078
rect 41696 642524 41748 642530
rect 41748 642484 42104 642512
rect 41696 642466 41748 642472
rect 42076 642394 42104 642484
rect 42064 642388 42116 642394
rect 42064 642330 42116 642336
rect 41708 641986 42104 642002
rect 41696 641980 42116 641986
rect 41748 641974 42064 641980
rect 41696 641922 41748 641928
rect 42064 641922 42116 641928
rect 41696 641776 41748 641782
rect 42064 641776 42116 641782
rect 41748 641724 42064 641730
rect 41696 641718 42116 641724
rect 41708 641702 42104 641718
rect 41142 641064 41198 641073
rect 41142 640999 41198 641008
rect 42064 640960 42116 640966
rect 42064 640902 42116 640908
rect 42076 640778 42104 640902
rect 41708 640750 42104 640778
rect 40868 640620 40920 640626
rect 40868 640562 40920 640568
rect 40880 640257 40908 640562
rect 41708 640490 41736 640750
rect 41696 640484 41748 640490
rect 41696 640426 41748 640432
rect 41696 640348 41748 640354
rect 42064 640348 42116 640354
rect 41748 640306 42064 640334
rect 41696 640290 41748 640296
rect 42064 640290 42116 640296
rect 40866 640248 40922 640257
rect 40866 640183 40922 640192
rect 34426 639840 34482 639849
rect 34426 639775 34482 639784
rect 39394 639840 39450 639849
rect 39394 639775 39450 639784
rect 34440 638246 34468 639775
rect 35530 639432 35586 639441
rect 35530 639367 35586 639376
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 35544 639130 35572 639367
rect 35820 639266 35848 639367
rect 35808 639260 35860 639266
rect 35808 639202 35860 639208
rect 41696 639260 41748 639266
rect 41696 639202 41748 639208
rect 41708 639146 41736 639202
rect 35532 639124 35584 639130
rect 35532 639066 35584 639072
rect 39304 639124 39356 639130
rect 41708 639118 42380 639146
rect 39304 639066 39356 639072
rect 35622 638616 35678 638625
rect 35622 638551 35678 638560
rect 34428 638240 34480 638246
rect 34428 638182 34480 638188
rect 32402 637800 32458 637809
rect 32402 637735 32458 637744
rect 32416 629921 32444 637735
rect 35162 637392 35218 637401
rect 35162 637327 35218 637336
rect 32402 629912 32458 629921
rect 32402 629847 32458 629856
rect 35176 628726 35204 637327
rect 35636 636954 35664 638551
rect 35806 638208 35862 638217
rect 35806 638143 35862 638152
rect 35820 637634 35848 638143
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 36544 637628 36596 637634
rect 36544 637570 36596 637576
rect 35806 636984 35862 636993
rect 35624 636948 35676 636954
rect 35806 636919 35862 636928
rect 35624 636890 35676 636896
rect 35820 636750 35848 636919
rect 35808 636744 35860 636750
rect 35808 636686 35860 636692
rect 35530 636576 35586 636585
rect 35530 636511 35586 636520
rect 35806 636576 35862 636585
rect 35806 636511 35862 636520
rect 35544 636274 35572 636511
rect 35820 636410 35848 636511
rect 35808 636404 35860 636410
rect 35808 636346 35860 636352
rect 35532 636268 35584 636274
rect 35532 636210 35584 636216
rect 35806 635760 35862 635769
rect 35806 635695 35862 635704
rect 35820 634982 35848 635695
rect 35808 634976 35860 634982
rect 35808 634918 35860 634924
rect 35806 634536 35862 634545
rect 35806 634471 35862 634480
rect 35820 633894 35848 634471
rect 35808 633888 35860 633894
rect 35808 633830 35860 633836
rect 35806 633720 35862 633729
rect 35806 633655 35862 633664
rect 35820 633486 35848 633655
rect 35808 633480 35860 633486
rect 35808 633422 35860 633428
rect 36556 630630 36584 637570
rect 39120 636200 39172 636206
rect 39118 636168 39120 636177
rect 39172 636168 39174 636177
rect 39118 636103 39174 636112
rect 36544 630624 36596 630630
rect 36544 630566 36596 630572
rect 39316 629241 39344 639066
rect 41696 638240 41748 638246
rect 41696 638182 41748 638188
rect 40592 636948 40644 636954
rect 40592 636890 40644 636896
rect 40040 636608 40092 636614
rect 40038 636576 40040 636585
rect 40092 636576 40094 636585
rect 40038 636511 40094 636520
rect 39580 636472 39632 636478
rect 39580 636414 39632 636420
rect 39592 635769 39620 636414
rect 39578 635760 39634 635769
rect 39578 635695 39634 635704
rect 40132 634976 40184 634982
rect 40132 634918 40184 634924
rect 40144 634137 40172 634918
rect 40130 634128 40186 634137
rect 40130 634063 40186 634072
rect 40040 633752 40092 633758
rect 40040 633694 40092 633700
rect 40052 630873 40080 633694
rect 40604 632913 40632 636890
rect 41708 635066 41736 638182
rect 41708 635038 41828 635066
rect 41604 633480 41656 633486
rect 41604 633422 41656 633428
rect 41616 633321 41644 633422
rect 41602 633312 41658 633321
rect 41602 633247 41658 633256
rect 40590 632904 40646 632913
rect 40590 632839 40646 632848
rect 40038 630864 40094 630873
rect 40038 630799 40094 630808
rect 41800 630674 41828 635038
rect 42064 633480 42116 633486
rect 42064 633422 42116 633428
rect 42076 633321 42104 633422
rect 42062 633312 42118 633321
rect 42062 633247 42118 633256
rect 41800 630646 42288 630674
rect 41604 630624 41656 630630
rect 41656 630572 41828 630578
rect 41604 630566 41828 630572
rect 41616 630550 41828 630566
rect 39302 629232 39358 629241
rect 39302 629167 39358 629176
rect 35164 628720 35216 628726
rect 39396 628720 39448 628726
rect 35164 628662 35216 628668
rect 39394 628688 39396 628697
rect 39448 628688 39450 628697
rect 39394 628623 39450 628632
rect 41800 627473 41828 630550
rect 41786 627464 41842 627473
rect 41786 627399 41842 627408
rect 41786 627192 41842 627201
rect 41786 627127 41842 627136
rect 41800 626620 41828 627127
rect 42260 625274 42288 630646
rect 42352 626634 42380 639118
rect 42614 632904 42670 632913
rect 42670 632862 42840 632890
rect 42614 632839 42670 632848
rect 42614 628688 42670 628697
rect 42614 628623 42670 628632
rect 42352 626606 42564 626634
rect 42168 625246 42288 625274
rect 42168 624784 42196 625246
rect 42340 625184 42392 625190
rect 42340 625126 42392 625132
rect 42154 624608 42210 624617
rect 42154 624543 42210 624552
rect 42168 624172 42196 624543
rect 42352 623506 42380 625126
rect 42168 623478 42380 623506
rect 42168 622948 42196 623478
rect 42248 622872 42300 622878
rect 42248 622814 42300 622820
rect 42260 622554 42288 622814
rect 42260 622526 42380 622554
rect 42168 622033 42196 622336
rect 41786 622024 41842 622033
rect 41786 621959 41842 621968
rect 42154 622024 42210 622033
rect 42154 621959 42210 621968
rect 41800 621792 41828 621959
rect 42352 621126 42380 622526
rect 42182 621098 42380 621126
rect 42536 621014 42564 626606
rect 42444 620986 42564 621014
rect 41786 620800 41842 620809
rect 41786 620735 41842 620744
rect 41800 620500 41828 620735
rect 42248 620288 42300 620294
rect 42076 620236 42248 620242
rect 42076 620230 42300 620236
rect 42076 620214 42288 620230
rect 42076 619956 42104 620214
rect 42248 619676 42300 619682
rect 42248 619618 42300 619624
rect 42260 617454 42288 619618
rect 42182 617426 42288 617454
rect 42248 617364 42300 617370
rect 42248 617306 42300 617312
rect 42260 617250 42288 617306
rect 42076 617222 42288 617250
rect 42076 616828 42104 617222
rect 42444 616808 42472 620986
rect 42628 620378 42656 628623
rect 42812 627914 42840 632862
rect 42352 616780 42472 616808
rect 42536 620350 42656 620378
rect 42720 627886 42840 627914
rect 42156 616344 42208 616350
rect 42156 616286 42208 616292
rect 42168 616148 42196 616286
rect 42352 615890 42380 616780
rect 42536 616350 42564 620350
rect 42720 620294 42748 627886
rect 42708 620288 42760 620294
rect 42708 620230 42760 620236
rect 42524 616344 42576 616350
rect 42524 616286 42576 616292
rect 42168 615862 42380 615890
rect 42168 615604 42196 615862
rect 42338 615768 42394 615777
rect 42338 615703 42394 615712
rect 42352 613782 42380 615703
rect 42614 615496 42670 615505
rect 42614 615431 42670 615440
rect 42628 615346 42656 615431
rect 42182 613754 42380 613782
rect 42536 615318 42656 615346
rect 41878 613456 41934 613465
rect 41878 613391 41934 613400
rect 41892 613121 41920 613391
rect 42536 612490 42564 615318
rect 42904 614281 42932 721103
rect 43088 684729 43116 727767
rect 43074 684720 43130 684729
rect 43074 684655 43130 684664
rect 43076 684548 43128 684554
rect 43076 684490 43128 684496
rect 43088 641986 43116 684490
rect 43076 641980 43128 641986
rect 43076 641922 43128 641928
rect 43074 634128 43130 634137
rect 43074 634063 43130 634072
rect 43088 619682 43116 634063
rect 43076 619676 43128 619682
rect 43076 619618 43128 619624
rect 42890 614272 42946 614281
rect 42890 614207 42946 614216
rect 42708 614168 42760 614174
rect 42708 614110 42760 614116
rect 42182 612462 42564 612490
rect 42248 612400 42300 612406
rect 42246 612368 42248 612377
rect 42300 612368 42302 612377
rect 42246 612303 42302 612312
rect 42720 612082 42748 614110
rect 43272 612678 43300 807434
rect 43456 772313 43484 814370
rect 44192 810762 44220 815594
rect 45284 814292 45336 814298
rect 45284 814234 45336 814240
rect 44548 812864 44600 812870
rect 44548 812806 44600 812812
rect 44180 810756 44232 810762
rect 44180 810698 44232 810704
rect 44364 807356 44416 807362
rect 44364 807298 44416 807304
rect 43628 799060 43680 799066
rect 43628 799002 43680 799008
rect 43640 797337 43668 799002
rect 43812 797700 43864 797706
rect 43812 797642 43864 797648
rect 43626 797328 43682 797337
rect 43626 797263 43682 797272
rect 43824 795666 43852 797642
rect 43812 795660 43864 795666
rect 43812 795602 43864 795608
rect 44376 793966 44404 807298
rect 44364 793960 44416 793966
rect 44364 793902 44416 793908
rect 43442 772304 43498 772313
rect 43442 772239 43498 772248
rect 44270 771488 44326 771497
rect 44270 771423 44326 771432
rect 43626 770264 43682 770273
rect 43626 770199 43682 770208
rect 43444 764652 43496 764658
rect 43444 764594 43496 764600
rect 43456 753817 43484 764594
rect 43442 753808 43498 753817
rect 43442 753743 43498 753752
rect 43444 727456 43496 727462
rect 43444 727398 43496 727404
rect 43456 683913 43484 727398
rect 43640 727326 43668 770199
rect 43904 755540 43956 755546
rect 43904 755482 43956 755488
rect 43916 754089 43944 755482
rect 43902 754080 43958 754089
rect 43902 754015 43958 754024
rect 44284 728890 44312 771423
rect 44560 770166 44588 812806
rect 45098 773120 45154 773129
rect 45098 773055 45154 773064
rect 44548 770160 44600 770166
rect 44548 770102 44600 770108
rect 44454 764552 44510 764561
rect 44454 764487 44510 764496
rect 44468 753545 44496 764487
rect 44638 764144 44694 764153
rect 44638 764079 44694 764088
rect 44454 753536 44510 753545
rect 44454 753471 44510 753480
rect 44652 751233 44680 764079
rect 44914 763328 44970 763337
rect 44914 763263 44970 763272
rect 44638 751224 44694 751233
rect 44638 751159 44694 751168
rect 44272 728884 44324 728890
rect 44272 728826 44324 728832
rect 44548 728680 44600 728686
rect 44548 728622 44600 728628
rect 44270 728240 44326 728249
rect 44270 728175 44326 728184
rect 43628 727320 43680 727326
rect 43628 727262 43680 727268
rect 43810 723616 43866 723625
rect 43810 723551 43866 723560
rect 43626 720352 43682 720361
rect 43626 720287 43682 720296
rect 43640 719030 43668 720287
rect 43628 719024 43680 719030
rect 43628 718966 43680 718972
rect 43628 712156 43680 712162
rect 43628 712098 43680 712104
rect 43640 710841 43668 712098
rect 43626 710832 43682 710841
rect 43626 710767 43682 710776
rect 43628 709368 43680 709374
rect 43628 709310 43680 709316
rect 43640 707878 43668 709310
rect 43628 707872 43680 707878
rect 43628 707814 43680 707820
rect 43824 705566 43852 723551
rect 43812 705560 43864 705566
rect 43812 705502 43864 705508
rect 43628 686316 43680 686322
rect 43628 686258 43680 686264
rect 43442 683904 43498 683913
rect 43442 683839 43498 683848
rect 43442 677920 43498 677929
rect 43442 677855 43498 677864
rect 43260 612672 43312 612678
rect 43260 612614 43312 612620
rect 42536 612054 42748 612082
rect 42536 611946 42564 612054
rect 42182 611918 42564 611946
rect 43456 611153 43484 677855
rect 43640 643346 43668 686258
rect 44284 685914 44312 728175
rect 44560 686118 44588 728622
rect 44730 721576 44786 721585
rect 44730 721511 44786 721520
rect 44744 710462 44772 721511
rect 44732 710456 44784 710462
rect 44732 710398 44784 710404
rect 44730 708520 44786 708529
rect 44730 708455 44786 708464
rect 44744 703798 44772 708455
rect 44732 703792 44784 703798
rect 44732 703734 44784 703740
rect 44548 686112 44600 686118
rect 44548 686054 44600 686060
rect 44272 685908 44324 685914
rect 44272 685850 44324 685856
rect 44454 680232 44510 680241
rect 44454 680167 44510 680176
rect 44270 679416 44326 679425
rect 44270 679351 44326 679360
rect 43810 678600 43866 678609
rect 43810 678535 43866 678544
rect 43824 661094 43852 678535
rect 43994 677104 44050 677113
rect 43994 677039 44050 677048
rect 44008 676258 44036 677039
rect 43996 676252 44048 676258
rect 43996 676194 44048 676200
rect 44088 669452 44140 669458
rect 44088 669394 44140 669400
rect 44100 667729 44128 669394
rect 44086 667720 44142 667729
rect 44086 667655 44142 667664
rect 44284 666641 44312 679351
rect 44270 666632 44326 666641
rect 44270 666567 44326 666576
rect 44468 662998 44496 680167
rect 44730 679008 44786 679017
rect 44730 678943 44786 678952
rect 44744 667185 44772 678943
rect 44730 667176 44786 667185
rect 44730 667111 44786 667120
rect 44456 662992 44508 662998
rect 44456 662934 44508 662940
rect 43812 661088 43864 661094
rect 43812 661030 43864 661036
rect 43628 643340 43680 643346
rect 43628 643282 43680 643288
rect 44546 641064 44602 641073
rect 44546 640999 44602 641008
rect 44362 639840 44418 639849
rect 44362 639775 44418 639784
rect 43810 636576 43866 636585
rect 43810 636511 43866 636520
rect 43626 630864 43682 630873
rect 43626 630799 43682 630808
rect 43442 611144 43498 611153
rect 43442 611079 43498 611088
rect 43640 610745 43668 630799
rect 43824 618322 43852 636511
rect 44178 636168 44234 636177
rect 44178 636103 44234 636112
rect 43994 635760 44050 635769
rect 43994 635695 44050 635704
rect 44008 623830 44036 635695
rect 44192 626006 44220 636103
rect 44180 626000 44232 626006
rect 44180 625942 44232 625948
rect 44180 625864 44232 625870
rect 44180 625806 44232 625812
rect 44192 624617 44220 625806
rect 44178 624608 44234 624617
rect 44178 624543 44234 624552
rect 43996 623824 44048 623830
rect 43996 623766 44048 623772
rect 44178 622024 44234 622033
rect 44178 621959 44234 621968
rect 43812 618316 43864 618322
rect 43812 618258 43864 618264
rect 44192 616826 44220 621959
rect 44180 616820 44232 616826
rect 44180 616762 44232 616768
rect 44086 614272 44142 614281
rect 44086 614207 44142 614216
rect 43766 611992 43818 611998
rect 43766 611934 43818 611940
rect 43778 611833 43806 611934
rect 43764 611824 43820 611833
rect 44100 611810 44128 614207
rect 44100 611782 44251 611810
rect 43764 611759 43820 611768
rect 43996 611652 44048 611658
rect 43996 611594 44048 611600
rect 44008 611425 44036 611594
rect 44223 611590 44251 611782
rect 44211 611584 44263 611590
rect 44211 611526 44263 611532
rect 43994 611416 44050 611425
rect 43994 611351 44050 611360
rect 43626 610736 43682 610745
rect 43626 610671 43682 610680
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 40314 602032 40370 602041
rect 40314 601967 40370 601976
rect 35806 601760 35862 601769
rect 35806 601695 35808 601704
rect 35860 601695 35862 601704
rect 36544 601724 36596 601730
rect 35808 601666 35860 601672
rect 36544 601666 36596 601672
rect 35162 595810 35218 595819
rect 35162 595745 35218 595754
rect 33046 595232 33102 595241
rect 33046 595167 33102 595176
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585818 31064 594351
rect 33060 587178 33088 595167
rect 33782 593600 33838 593609
rect 33782 593535 33838 593544
rect 33048 587172 33100 587178
rect 33048 587114 33100 587120
rect 33796 585954 33824 593535
rect 35176 586226 35204 595745
rect 35622 591968 35678 591977
rect 35622 591903 35678 591912
rect 35636 590986 35664 591903
rect 35806 591560 35862 591569
rect 35806 591495 35862 591504
rect 35624 590980 35676 590986
rect 35624 590922 35676 590928
rect 35820 590714 35848 591495
rect 35808 590708 35860 590714
rect 35808 590650 35860 590656
rect 36556 589665 36584 601666
rect 39946 601352 40002 601361
rect 39946 601287 40002 601296
rect 37922 594586 37978 594595
rect 39960 594590 39988 601287
rect 40130 600944 40186 600953
rect 40130 600879 40186 600888
rect 40144 595814 40172 600879
rect 40132 595808 40184 595814
rect 40132 595750 40184 595756
rect 37922 594521 37978 594530
rect 39948 594584 40000 594590
rect 39948 594526 40000 594532
rect 36542 589656 36598 589665
rect 36542 589591 36598 589600
rect 35164 586220 35216 586226
rect 35164 586162 35216 586168
rect 33784 585948 33836 585954
rect 33784 585890 33836 585896
rect 31024 585812 31076 585818
rect 31024 585754 31076 585760
rect 37936 585177 37964 594521
rect 40328 592034 40356 601967
rect 44376 599842 44404 639775
rect 44560 600545 44588 640999
rect 44928 611998 44956 763263
rect 45112 732329 45140 773055
rect 45296 771526 45324 814234
rect 46216 785194 46244 817090
rect 60004 817012 60056 817018
rect 60004 816954 60056 816960
rect 50344 806132 50396 806138
rect 50344 806074 50396 806080
rect 46204 785188 46256 785194
rect 46204 785130 46256 785136
rect 46204 773084 46256 773090
rect 46204 773026 46256 773032
rect 45284 771520 45336 771526
rect 45284 771462 45336 771468
rect 45282 751632 45338 751641
rect 45282 751567 45338 751576
rect 45296 746570 45324 751567
rect 45284 746564 45336 746570
rect 45284 746506 45336 746512
rect 46216 743782 46244 773026
rect 48964 761932 49016 761938
rect 48964 761874 49016 761880
rect 46204 743776 46256 743782
rect 46204 743718 46256 743724
rect 45098 732320 45154 732329
rect 45098 732255 45154 732264
rect 46202 731096 46258 731105
rect 46202 731031 46258 731040
rect 45098 722800 45154 722809
rect 45098 722735 45154 722744
rect 45112 709374 45140 722735
rect 45100 709368 45152 709374
rect 45100 709310 45152 709316
rect 46216 698290 46244 731031
rect 46204 698284 46256 698290
rect 46204 698226 46256 698232
rect 45466 687576 45522 687585
rect 45466 687511 45522 687520
rect 45284 684820 45336 684826
rect 45284 684762 45336 684768
rect 45098 683088 45154 683097
rect 45098 683023 45154 683032
rect 45112 640966 45140 683023
rect 45296 641782 45324 684762
rect 45480 655518 45508 687511
rect 46202 687168 46258 687177
rect 46202 687103 46258 687112
rect 45652 667956 45704 667962
rect 45652 667898 45704 667904
rect 45664 667078 45692 667898
rect 45652 667072 45704 667078
rect 45652 667014 45704 667020
rect 46216 656878 46244 687103
rect 46204 656872 46256 656878
rect 46204 656814 46256 656820
rect 45468 655512 45520 655518
rect 45468 655454 45520 655460
rect 45284 641776 45336 641782
rect 45284 641718 45336 641724
rect 45100 640960 45152 640966
rect 45100 640902 45152 640908
rect 45376 640348 45428 640354
rect 45376 640290 45428 640296
rect 45098 640248 45154 640257
rect 45098 640183 45154 640192
rect 44916 611992 44968 611998
rect 44916 611934 44968 611940
rect 44730 611144 44786 611153
rect 44730 611079 44732 611088
rect 44784 611079 44786 611088
rect 44732 611050 44784 611056
rect 44732 610768 44784 610774
rect 44730 610736 44732 610745
rect 44784 610736 44786 610745
rect 44730 610671 44786 610680
rect 44546 600536 44602 600545
rect 44546 600471 44602 600480
rect 44638 600128 44694 600137
rect 44638 600063 44694 600072
rect 44376 599814 44496 599842
rect 44468 599729 44496 599814
rect 44454 599720 44510 599729
rect 44454 599655 44510 599664
rect 42890 597680 42946 597689
rect 42890 597615 42946 597624
rect 42904 597446 42932 597615
rect 42892 597440 42944 597446
rect 42892 597382 42944 597388
rect 42892 597032 42944 597038
rect 42892 596974 42944 596980
rect 43074 597000 43130 597009
rect 40958 596864 41014 596873
rect 40958 596799 41014 596808
rect 40972 592550 41000 596799
rect 41142 596456 41198 596465
rect 41142 596391 41198 596400
rect 40960 592544 41012 592550
rect 40960 592486 41012 592492
rect 41156 592090 41184 596391
rect 41326 595810 41382 595819
rect 41696 595808 41748 595814
rect 41326 595745 41382 595754
rect 41694 595776 41696 595785
rect 41748 595776 41750 595785
rect 41340 594794 41368 595745
rect 41694 595711 41750 595720
rect 41328 594788 41380 594794
rect 41328 594730 41380 594736
rect 41512 594788 41564 594794
rect 41512 594730 41564 594736
rect 41524 592362 41552 594730
rect 41696 594584 41748 594590
rect 41694 594552 41696 594561
rect 41748 594552 41750 594561
rect 41694 594487 41750 594496
rect 41696 592544 41748 592550
rect 41748 592492 42012 592498
rect 41696 592486 42012 592492
rect 41708 592470 42012 592486
rect 41524 592334 41920 592362
rect 41694 592104 41750 592113
rect 41156 592062 41694 592090
rect 41694 592039 41750 592048
rect 40328 592006 40448 592034
rect 39764 590708 39816 590714
rect 39764 590650 39816 590656
rect 39776 589393 39804 590650
rect 39762 589384 39818 589393
rect 39762 589319 39818 589328
rect 39856 585948 39908 585954
rect 39856 585890 39908 585896
rect 37922 585168 37978 585177
rect 37922 585103 37978 585112
rect 39868 584633 39896 585890
rect 40420 585721 40448 592006
rect 41696 590980 41748 590986
rect 41696 590922 41748 590928
rect 41708 590481 41736 590922
rect 41694 590472 41750 590481
rect 41694 590407 41750 590416
rect 41892 587194 41920 592334
rect 41984 592034 42012 592470
rect 42904 592034 42932 596974
rect 43074 596935 43130 596944
rect 41984 592006 42288 592034
rect 42904 592006 43024 592034
rect 41892 587178 42104 587194
rect 41512 587172 41564 587178
rect 41892 587172 42116 587178
rect 41892 587166 42064 587172
rect 41512 587114 41564 587120
rect 42064 587114 42116 587120
rect 40590 585984 40646 585993
rect 40590 585919 40646 585928
rect 40604 585818 40632 585919
rect 40592 585812 40644 585818
rect 40592 585754 40644 585760
rect 40406 585712 40462 585721
rect 40406 585647 40462 585656
rect 41524 585426 41552 587114
rect 42064 586288 42116 586294
rect 41708 586236 42064 586242
rect 41708 586230 42116 586236
rect 41708 586226 42104 586230
rect 41696 586220 42104 586226
rect 41748 586214 42104 586220
rect 41696 586162 41748 586168
rect 42260 586090 42288 592006
rect 42616 587172 42668 587178
rect 42616 587114 42668 587120
rect 42248 586084 42300 586090
rect 42248 586026 42300 586032
rect 42430 585984 42486 585993
rect 42430 585919 42486 585928
rect 42444 585834 42472 585919
rect 42444 585806 42564 585834
rect 42248 585608 42300 585614
rect 42300 585556 42380 585562
rect 42248 585550 42380 585556
rect 42260 585534 42380 585550
rect 41524 585398 42288 585426
rect 39854 584624 39910 584633
rect 39854 584559 39910 584568
rect 42260 583454 42288 585398
rect 42182 583426 42288 583454
rect 42352 581618 42380 585534
rect 42182 581590 42380 581618
rect 42182 580947 42288 580975
rect 42260 580281 42288 580947
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 42246 580272 42302 580281
rect 42246 580207 42302 580216
rect 41800 579768 41828 580207
rect 42536 579614 42564 585806
rect 42444 579586 42564 579614
rect 41984 578921 42012 579121
rect 42248 579012 42300 579018
rect 42248 578954 42300 578960
rect 41970 578912 42026 578921
rect 41970 578847 42026 578856
rect 42260 578626 42288 578954
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 42246 578504 42302 578513
rect 42246 578439 42302 578448
rect 42260 577946 42288 578439
rect 42182 577918 42288 577946
rect 41786 577824 41842 577833
rect 41786 577759 41842 577768
rect 42248 577788 42300 577794
rect 41800 577281 41828 577759
rect 42248 577730 42300 577736
rect 42260 576858 42288 577730
rect 42168 576830 42288 576858
rect 42444 576858 42472 579586
rect 42628 576994 42656 587114
rect 42800 586152 42852 586158
rect 42720 586100 42800 586106
rect 42720 586094 42852 586100
rect 42720 586078 42840 586094
rect 42720 577810 42748 586078
rect 42720 577794 42840 577810
rect 42720 577788 42852 577794
rect 42720 577782 42800 577788
rect 42800 577730 42852 577736
rect 42628 576966 42748 576994
rect 42444 576830 42564 576858
rect 42168 576708 42196 576830
rect 42246 575920 42302 575929
rect 42246 575855 42302 575864
rect 42260 574274 42288 575855
rect 42182 574246 42288 574274
rect 41970 573880 42026 573889
rect 41970 573815 42026 573824
rect 41984 573580 42012 573815
rect 42536 573730 42564 576830
rect 42260 573702 42564 573730
rect 42260 572982 42288 573702
rect 42720 573594 42748 576966
rect 42182 572954 42288 572982
rect 42444 573566 42748 573594
rect 42444 572438 42472 573566
rect 42614 573336 42670 573345
rect 42614 573271 42670 573280
rect 42168 572370 42196 572424
rect 42260 572410 42472 572438
rect 42260 572370 42288 572410
rect 42168 572342 42288 572370
rect 42062 571568 42118 571577
rect 42062 571503 42118 571512
rect 42076 571282 42104 571503
rect 42430 571432 42486 571441
rect 42430 571367 42486 571376
rect 42076 571254 42380 571282
rect 42064 570988 42116 570994
rect 42064 570930 42116 570936
rect 42076 570588 42104 570930
rect 41786 570208 41842 570217
rect 41786 570143 41842 570152
rect 41800 569908 41828 570143
rect 42352 569310 42380 571254
rect 42168 569242 42196 569296
rect 42260 569282 42380 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42444 568766 42472 571367
rect 42628 570994 42656 573271
rect 42616 570988 42668 570994
rect 42616 570930 42668 570936
rect 42168 568698 42196 568752
rect 42260 568738 42472 568766
rect 42260 568698 42288 568738
rect 42168 568670 42288 568698
rect 42996 567194 43024 592006
rect 42812 567166 43024 567194
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 42812 559065 42840 567166
rect 39854 559056 39910 559065
rect 39854 558991 39910 559000
rect 42798 559056 42854 559065
rect 42798 558991 42854 559000
rect 35806 558104 35862 558113
rect 35806 558039 35862 558048
rect 35820 557598 35848 558039
rect 35808 557592 35860 557598
rect 35808 557534 35860 557540
rect 35806 555656 35862 555665
rect 35806 555591 35862 555600
rect 35820 555082 35848 555591
rect 35808 555076 35860 555082
rect 35808 555018 35860 555024
rect 35806 554840 35862 554849
rect 39868 554810 39896 558991
rect 43088 558793 43116 596935
rect 44362 593192 44418 593201
rect 44362 593127 44418 593136
rect 43258 590472 43314 590481
rect 43258 590407 43314 590416
rect 43272 579018 43300 590407
rect 43442 589384 43498 589393
rect 43442 589319 43498 589328
rect 43260 579012 43312 579018
rect 43260 578954 43312 578960
rect 40498 558784 40554 558793
rect 40498 558719 40554 558728
rect 43074 558784 43130 558793
rect 43074 558719 43130 558728
rect 40512 555082 40540 558719
rect 40960 557592 41012 557598
rect 40960 557534 41012 557540
rect 40500 555076 40552 555082
rect 40500 555018 40552 555024
rect 35806 554775 35808 554784
rect 35860 554775 35862 554784
rect 39856 554804 39908 554810
rect 35808 554746 35860 554752
rect 39856 554746 39908 554752
rect 35622 554432 35678 554441
rect 35622 554367 35678 554376
rect 35636 553586 35664 554367
rect 35806 553616 35862 553625
rect 35624 553580 35676 553586
rect 35806 553551 35862 553560
rect 35624 553522 35676 553528
rect 35820 553450 35848 553551
rect 35808 553444 35860 553450
rect 35808 553386 35860 553392
rect 37922 553408 37978 553417
rect 40972 553394 41000 557534
rect 41696 553580 41748 553586
rect 41696 553522 41748 553528
rect 37922 553343 37978 553352
rect 40880 553366 41000 553394
rect 41328 553444 41380 553450
rect 41328 553386 41380 553392
rect 29642 551984 29698 551993
rect 29642 551919 29698 551928
rect 29656 547194 29684 551919
rect 29644 547188 29696 547194
rect 29644 547130 29696 547136
rect 37936 542337 37964 553343
rect 40880 550254 40908 553366
rect 41340 552514 41368 553386
rect 41708 553081 41736 553522
rect 41694 553072 41750 553081
rect 41694 553007 41750 553016
rect 43166 553072 43222 553081
rect 43166 553007 43222 553016
rect 40972 552486 41368 552514
rect 40972 550474 41000 552486
rect 41326 552392 41382 552401
rect 41326 552327 41382 552336
rect 41340 552090 41368 552327
rect 41328 552084 41380 552090
rect 41328 552026 41380 552032
rect 41696 552084 41748 552090
rect 41696 552026 41748 552032
rect 41708 551857 41736 552026
rect 41694 551848 41750 551857
rect 41694 551783 41750 551792
rect 41142 551168 41198 551177
rect 41142 551103 41198 551112
rect 41156 550662 41184 551103
rect 41144 550656 41196 550662
rect 41144 550598 41196 550604
rect 41696 550656 41748 550662
rect 42064 550656 42116 550662
rect 41748 550616 42064 550644
rect 41696 550598 41748 550604
rect 42064 550598 42116 550604
rect 42984 550656 43036 550662
rect 42984 550598 43036 550604
rect 40972 550446 41460 550474
rect 41432 550338 41460 550446
rect 41432 550310 42380 550338
rect 40868 550248 40920 550254
rect 40868 550190 40920 550196
rect 41696 550248 41748 550254
rect 42062 550216 42118 550225
rect 41748 550196 42062 550202
rect 41696 550190 42062 550196
rect 41708 550174 42062 550190
rect 42062 550151 42118 550160
rect 41786 549944 41842 549953
rect 41524 549902 41786 549930
rect 40498 549536 40554 549545
rect 40498 549471 40554 549480
rect 39210 547496 39266 547505
rect 39210 547431 39266 547440
rect 39224 543697 39252 547431
rect 40512 545329 40540 549471
rect 41326 548312 41382 548321
rect 41326 548247 41382 548256
rect 41340 547942 41368 548247
rect 41328 547936 41380 547942
rect 41328 547878 41380 547884
rect 41524 545601 41552 549902
rect 41786 549879 41842 549888
rect 41696 547936 41748 547942
rect 41696 547878 41748 547884
rect 41708 547777 41736 547878
rect 41694 547768 41750 547777
rect 41694 547703 41750 547712
rect 41696 547188 41748 547194
rect 41696 547130 41748 547136
rect 41510 545592 41566 545601
rect 41510 545527 41566 545536
rect 40498 545320 40554 545329
rect 40498 545255 40554 545264
rect 41708 543734 41736 547130
rect 42352 543734 42380 550310
rect 42798 549128 42854 549137
rect 42798 549063 42854 549072
rect 41708 543706 42288 543734
rect 42352 543706 42472 543734
rect 39210 543688 39266 543697
rect 39210 543623 39266 543632
rect 37922 542328 37978 542337
rect 37922 542263 37978 542272
rect 42260 540274 42288 543706
rect 42182 540246 42288 540274
rect 42444 538438 42472 543706
rect 42614 539608 42670 539617
rect 42614 539543 42670 539552
rect 42168 538370 42196 538424
rect 42260 538410 42472 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42430 538248 42486 538257
rect 42430 538183 42486 538192
rect 42076 537441 42104 537744
rect 42062 537432 42118 537441
rect 42062 537367 42118 537376
rect 42062 537024 42118 537033
rect 42062 536959 42118 536968
rect 42076 536588 42104 536959
rect 42444 535922 42472 538183
rect 42628 537033 42656 539543
rect 42614 537024 42670 537033
rect 42614 536959 42670 536968
rect 42812 536874 42840 549063
rect 42996 543734 43024 550598
rect 42182 535894 42472 535922
rect 42536 536846 42840 536874
rect 42904 543706 43024 543734
rect 42062 535664 42118 535673
rect 42062 535599 42118 535608
rect 42076 535364 42104 535599
rect 41786 535256 41842 535265
rect 41786 535191 41842 535200
rect 41800 534752 41828 535191
rect 42536 534086 42564 536846
rect 42706 536752 42762 536761
rect 42706 536687 42762 536696
rect 42720 535673 42748 536687
rect 42706 535664 42762 535673
rect 42706 535599 42762 535608
rect 42182 534058 42564 534086
rect 42430 533896 42486 533905
rect 42430 533831 42486 533840
rect 42444 533542 42472 533831
rect 42706 533624 42762 533633
rect 42706 533559 42762 533568
rect 42182 533514 42472 533542
rect 42246 533352 42302 533361
rect 42246 533287 42302 533296
rect 42260 531059 42288 533287
rect 42522 532672 42578 532681
rect 42522 532607 42578 532616
rect 42182 531031 42288 531059
rect 42536 530754 42564 532607
rect 42156 530732 42208 530738
rect 42156 530674 42208 530680
rect 42444 530726 42564 530754
rect 42720 530738 42748 533559
rect 42708 530732 42760 530738
rect 42168 530400 42196 530674
rect 42248 530324 42300 530330
rect 42248 530266 42300 530272
rect 42260 529771 42288 530266
rect 42182 529743 42288 529771
rect 42444 529219 42472 530726
rect 42708 530674 42760 530680
rect 42904 530618 42932 543706
rect 42720 530590 42932 530618
rect 42720 530330 42748 530590
rect 42708 530324 42760 530330
rect 42708 530266 42760 530272
rect 42614 530088 42670 530097
rect 42614 530023 42670 530032
rect 42182 529191 42472 529219
rect 42628 529122 42656 530023
rect 42444 529094 42656 529122
rect 42168 527462 42288 527490
rect 42168 527340 42196 527462
rect 42260 527354 42288 527462
rect 42444 527354 42472 529094
rect 42706 529000 42762 529009
rect 42706 528935 42762 528944
rect 42720 528850 42748 528935
rect 42260 527326 42472 527354
rect 42536 528822 42748 528850
rect 42536 526742 42564 528822
rect 42706 528728 42762 528737
rect 42706 528663 42762 528672
rect 42720 528554 42748 528663
rect 42182 526714 42564 526742
rect 42628 528526 42748 528554
rect 42628 526130 42656 528526
rect 42890 527232 42946 527241
rect 42890 527167 42946 527176
rect 42904 527082 42932 527167
rect 42536 526102 42656 526130
rect 42720 527054 42932 527082
rect 42536 526091 42564 526102
rect 42182 526063 42564 526091
rect 42720 525586 42748 527054
rect 42168 525558 42288 525586
rect 42168 525504 42196 525558
rect 42260 525518 42288 525558
rect 42536 525558 42748 525586
rect 42536 525518 42564 525558
rect 42260 525490 42564 525518
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 35806 430128 35862 430137
rect 35806 430063 35862 430072
rect 35820 429214 35848 430063
rect 35808 429208 35860 429214
rect 35808 429150 35860 429156
rect 41696 429208 41748 429214
rect 41748 429156 42196 429162
rect 41696 429150 42196 429156
rect 41708 429134 42196 429150
rect 35806 428496 35862 428505
rect 35806 428431 35862 428440
rect 35820 427990 35848 428431
rect 35808 427984 35860 427990
rect 35808 427926 35860 427932
rect 41696 427984 41748 427990
rect 41696 427926 41748 427932
rect 41708 427802 41736 427926
rect 41708 427774 42012 427802
rect 41984 426601 42012 427774
rect 42168 427145 42196 429134
rect 43180 427417 43208 553007
rect 43166 427408 43222 427417
rect 43166 427343 43222 427352
rect 42154 427136 42210 427145
rect 42154 427071 42210 427080
rect 41970 426592 42026 426601
rect 41970 426527 42026 426536
rect 42890 426592 42946 426601
rect 42890 426527 42946 426536
rect 40958 426456 41014 426465
rect 40958 426391 41014 426400
rect 39302 425640 39358 425649
rect 39302 425575 39358 425584
rect 32770 424824 32826 424833
rect 32770 424759 32826 424768
rect 32784 417450 32812 424759
rect 34518 424416 34574 424425
rect 34518 424351 34574 424360
rect 33782 424008 33838 424017
rect 33782 423943 33838 423952
rect 32772 417444 32824 417450
rect 32772 417386 32824 417392
rect 33796 414633 33824 423943
rect 34532 416090 34560 424351
rect 34520 416084 34572 416090
rect 34520 416026 34572 416032
rect 39316 415313 39344 425575
rect 40972 417761 41000 426391
rect 41142 426048 41198 426057
rect 41142 425983 41198 425992
rect 41156 424386 41184 425983
rect 41144 424380 41196 424386
rect 41144 424322 41196 424328
rect 41696 424380 41748 424386
rect 41748 424340 42012 424368
rect 41696 424322 41748 424328
rect 41786 422376 41842 422385
rect 41786 422311 41842 422320
rect 41326 419928 41382 419937
rect 41326 419863 41382 419872
rect 41340 418849 41368 419863
rect 41326 418840 41382 418849
rect 41326 418775 41382 418784
rect 41800 418577 41828 422311
rect 41786 418568 41842 418577
rect 41786 418503 41842 418512
rect 41984 418154 42012 424340
rect 42154 421560 42210 421569
rect 42154 421495 42210 421504
rect 42168 418305 42196 421495
rect 42904 420186 42932 426527
rect 43074 425232 43130 425241
rect 43074 425167 43130 425176
rect 42812 420158 42932 420186
rect 42154 418296 42210 418305
rect 42154 418231 42210 418240
rect 41984 418126 42288 418154
rect 40958 417752 41014 417761
rect 40958 417687 41014 417696
rect 41696 417444 41748 417450
rect 41696 417386 41748 417392
rect 41708 417330 41736 417386
rect 41708 417314 42104 417330
rect 41708 417308 42116 417314
rect 41708 417302 42064 417308
rect 42064 417250 42116 417256
rect 41604 416084 41656 416090
rect 41604 416026 41656 416032
rect 41616 415970 41644 416026
rect 41616 415942 41828 415970
rect 39302 415304 39358 415313
rect 39302 415239 39358 415248
rect 33782 414624 33838 414633
rect 33782 414559 33838 414568
rect 41800 413545 41828 415942
rect 41786 413536 41842 413545
rect 41786 413471 41842 413480
rect 41786 413128 41842 413137
rect 41786 413063 41842 413072
rect 41800 412624 41828 413063
rect 42260 411346 42288 418126
rect 42616 417308 42668 417314
rect 42616 417250 42668 417256
rect 42168 411318 42288 411346
rect 42168 410788 42196 411318
rect 42182 410162 42472 410190
rect 42246 409864 42302 409873
rect 42246 409799 42302 409808
rect 42260 408966 42288 409799
rect 42182 408938 42288 408966
rect 42168 408218 42196 408340
rect 42168 408190 42288 408218
rect 42062 408096 42118 408105
rect 42062 408031 42118 408040
rect 42076 407796 42104 408031
rect 42260 407130 42288 408190
rect 42444 407289 42472 410162
rect 42430 407280 42486 407289
rect 42430 407215 42486 407224
rect 41800 407017 41828 407116
rect 42260 407102 42472 407130
rect 42248 407040 42300 407046
rect 41786 407008 41842 407017
rect 42248 406982 42300 406988
rect 41786 406943 41842 406952
rect 41786 406736 41842 406745
rect 41786 406671 41842 406680
rect 41800 406504 41828 406671
rect 42260 406042 42288 406982
rect 42168 406014 42288 406042
rect 42168 405929 42196 406014
rect 42444 404977 42472 407102
rect 42628 407046 42656 417250
rect 42616 407040 42668 407046
rect 42616 406982 42668 406988
rect 42430 404968 42486 404977
rect 42430 404903 42486 404912
rect 42246 404560 42302 404569
rect 42246 404495 42302 404504
rect 42260 403458 42288 404495
rect 42182 403430 42288 403458
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42432 402552 42484 402558
rect 42432 402494 42484 402500
rect 42444 402166 42472 402494
rect 42182 402138 42472 402166
rect 42432 402076 42484 402082
rect 42432 402018 42484 402024
rect 42444 401622 42472 402018
rect 42182 401594 42472 401622
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 41786 399392 41842 399401
rect 41786 399327 41842 399336
rect 41800 399121 41828 399327
rect 41970 398848 42026 398857
rect 41970 398783 42026 398792
rect 41984 398480 42012 398783
rect 42168 395729 42196 397936
rect 42154 395720 42210 395729
rect 42154 395655 42210 395664
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41326 387152 41382 387161
rect 41326 387087 41382 387096
rect 41142 386744 41198 386753
rect 41142 386679 41198 386688
rect 41156 385937 41184 386679
rect 41340 386442 41368 387087
rect 41328 386436 41380 386442
rect 41328 386378 41380 386384
rect 41696 386436 41748 386442
rect 41748 386396 41920 386424
rect 41696 386378 41748 386384
rect 40958 385928 41014 385937
rect 40958 385863 41014 385872
rect 41142 385928 41198 385937
rect 41142 385863 41198 385872
rect 40972 382265 41000 385863
rect 41142 383072 41198 383081
rect 41142 383007 41198 383016
rect 40038 382256 40094 382265
rect 40038 382191 40094 382200
rect 40958 382256 41014 382265
rect 40958 382191 41014 382200
rect 35438 381848 35494 381857
rect 35438 381783 35494 381792
rect 33966 381032 34022 381041
rect 33966 380967 34022 380976
rect 33980 373318 34008 380967
rect 35452 374649 35480 381783
rect 39302 381440 39358 381449
rect 39302 381375 39358 381384
rect 35808 379636 35860 379642
rect 35808 379578 35860 379584
rect 35820 379409 35848 379578
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 35808 378208 35860 378214
rect 35806 378176 35808 378185
rect 35860 378176 35862 378185
rect 35806 378111 35862 378120
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 35820 376145 35848 376479
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 35438 374640 35494 374649
rect 35438 374575 35494 374584
rect 33968 373312 34020 373318
rect 33968 373254 34020 373260
rect 39316 371890 39344 381375
rect 40052 379409 40080 382191
rect 41156 381857 41184 383007
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382430 41368 382599
rect 41328 382424 41380 382430
rect 41328 382366 41380 382372
rect 41696 382424 41748 382430
rect 41696 382366 41748 382372
rect 41142 381848 41198 381857
rect 41142 381783 41198 381792
rect 41326 379808 41382 379817
rect 41326 379743 41328 379752
rect 41380 379743 41382 379752
rect 41510 379808 41566 379817
rect 41510 379743 41512 379752
rect 41328 379714 41380 379720
rect 41564 379743 41566 379752
rect 41512 379714 41564 379720
rect 40408 379636 40460 379642
rect 40408 379578 40460 379584
rect 40038 379400 40094 379409
rect 40038 379335 40094 379344
rect 40420 376961 40448 379578
rect 41708 379514 41736 382366
rect 41892 381585 41920 386396
rect 42812 385665 42840 420158
rect 43088 418154 43116 425167
rect 43088 418126 43392 418154
rect 42982 417752 43038 417761
rect 42982 417687 43038 417696
rect 42996 402558 43024 417687
rect 43364 402974 43392 418126
rect 43272 402946 43392 402974
rect 42984 402552 43036 402558
rect 42984 402494 43036 402500
rect 43272 402082 43300 402946
rect 43260 402076 43312 402082
rect 43260 402018 43312 402024
rect 42798 385656 42854 385665
rect 42798 385591 42854 385600
rect 43258 385248 43314 385257
rect 43258 385183 43314 385192
rect 41878 381576 41934 381585
rect 41878 381511 41934 381520
rect 42890 380760 42946 380769
rect 42890 380695 42946 380704
rect 41708 379486 42380 379514
rect 41696 378208 41748 378214
rect 41694 378176 41696 378185
rect 41748 378176 41750 378185
rect 41694 378111 41750 378120
rect 40406 376952 40462 376961
rect 40406 376887 40462 376896
rect 41696 373312 41748 373318
rect 41748 373260 42288 373266
rect 41696 373254 42288 373260
rect 41708 373238 42288 373254
rect 39304 371884 39356 371890
rect 39304 371826 39356 371832
rect 41696 371884 41748 371890
rect 41696 371826 41748 371832
rect 41708 371770 41736 371826
rect 41708 371754 42104 371770
rect 41708 371748 42116 371754
rect 41708 371742 42064 371748
rect 42064 371690 42116 371696
rect 42260 369458 42288 373238
rect 42182 369430 42288 369458
rect 42352 367622 42380 379486
rect 42708 371748 42760 371754
rect 42708 371690 42760 371696
rect 42182 367594 42380 367622
rect 42182 366947 42564 366975
rect 42340 366852 42392 366858
rect 42340 366794 42392 366800
rect 42352 365786 42380 366794
rect 42182 365758 42380 365786
rect 42182 365107 42472 365135
rect 42248 365016 42300 365022
rect 42248 364958 42300 364964
rect 41786 364848 41842 364857
rect 41786 364783 41842 364792
rect 41800 364548 41828 364783
rect 41786 364168 41842 364177
rect 41786 364103 41842 364112
rect 41800 363936 41828 364103
rect 42062 363624 42118 363633
rect 42062 363559 42118 363568
rect 42076 363256 42104 363559
rect 42260 362794 42288 364958
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42444 362273 42472 365107
rect 42536 363066 42564 366947
rect 42720 365022 42748 371690
rect 42708 365016 42760 365022
rect 42708 364958 42760 364964
rect 42706 363080 42762 363089
rect 42536 363038 42706 363066
rect 42706 363015 42762 363024
rect 42430 362264 42486 362273
rect 42430 362199 42486 362208
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42154 359952 42210 359961
rect 42154 359887 42210 359896
rect 42168 359584 42196 359887
rect 42430 359000 42486 359009
rect 42182 358958 42430 358986
rect 42430 358935 42486 358944
rect 41878 358728 41934 358737
rect 41878 358663 41934 358672
rect 41892 358428 41920 358663
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42904 356046 42932 380695
rect 43074 376952 43130 376961
rect 43074 376887 43130 376896
rect 43088 366858 43116 376887
rect 43076 366852 43128 366858
rect 43076 366794 43128 366800
rect 42248 356040 42300 356046
rect 42892 356040 42944 356046
rect 42248 355982 42300 355988
rect 42430 356008 42486 356017
rect 42260 355926 42288 355982
rect 42892 355982 42944 355988
rect 42430 355943 42486 355952
rect 42182 355898 42288 355926
rect 41878 355736 41934 355745
rect 41878 355671 41934 355680
rect 41892 355300 41920 355671
rect 42444 354739 42472 355943
rect 42182 354711 42472 354739
rect 43272 345545 43300 385183
rect 43456 354249 43484 589319
rect 44376 579737 44404 593127
rect 44362 579728 44418 579737
rect 44362 579663 44418 579672
rect 44652 559337 44680 600063
rect 44914 599312 44970 599321
rect 44914 599247 44970 599256
rect 44638 559328 44694 559337
rect 44638 559263 44694 559272
rect 44546 556880 44602 556889
rect 44546 556815 44602 556824
rect 44362 555248 44418 555257
rect 44362 555183 44418 555192
rect 43994 551848 44050 551857
rect 43994 551783 44050 551792
rect 43810 550760 43866 550769
rect 43810 550695 43866 550704
rect 43626 547768 43682 547777
rect 43626 547703 43682 547712
rect 43640 354793 43668 547703
rect 43824 533633 43852 550695
rect 44008 533905 44036 551783
rect 44178 548720 44234 548729
rect 44178 548655 44234 548664
rect 44192 536897 44220 548655
rect 44178 536888 44234 536897
rect 44178 536823 44234 536832
rect 43994 533896 44050 533905
rect 43994 533831 44050 533840
rect 43810 533624 43866 533633
rect 43810 533559 43866 533568
rect 44376 428097 44404 555183
rect 44560 429729 44588 556815
rect 44928 556481 44956 599247
rect 45112 598913 45140 640183
rect 45388 621014 45416 640290
rect 45296 620986 45416 621014
rect 45098 598904 45154 598913
rect 45098 598839 45154 598848
rect 45296 598097 45324 620986
rect 46204 610904 46256 610910
rect 46204 610846 46256 610852
rect 45282 598088 45338 598097
rect 45282 598023 45338 598032
rect 45098 580272 45154 580281
rect 45098 580207 45154 580216
rect 45112 575482 45140 580207
rect 45100 575476 45152 575482
rect 45100 575418 45152 575424
rect 44914 556472 44970 556481
rect 44914 556407 44970 556416
rect 45006 556064 45062 556073
rect 45006 555999 45062 556008
rect 44730 537432 44786 537441
rect 44730 537367 44786 537376
rect 44744 532030 44772 537367
rect 44732 532024 44784 532030
rect 44732 531966 44784 531972
rect 44824 528624 44876 528630
rect 44824 528566 44876 528572
rect 44836 527241 44864 528566
rect 44822 527232 44878 527241
rect 44822 527167 44878 527176
rect 44822 430944 44878 430953
rect 44822 430879 44878 430888
rect 44546 429720 44602 429729
rect 44546 429655 44602 429664
rect 44638 429312 44694 429321
rect 44638 429247 44694 429256
rect 44362 428088 44418 428097
rect 44362 428023 44418 428032
rect 44454 427680 44510 427689
rect 44454 427615 44510 427624
rect 44270 426864 44326 426873
rect 44270 426799 44326 426808
rect 43810 422784 43866 422793
rect 43810 422719 43866 422728
rect 43824 409873 43852 422719
rect 43994 421152 44050 421161
rect 43994 421087 44050 421096
rect 43810 409864 43866 409873
rect 43810 409799 43866 409808
rect 44008 408105 44036 421087
rect 43994 408096 44050 408105
rect 43994 408031 44050 408040
rect 44284 384033 44312 426799
rect 44468 384849 44496 427615
rect 44652 386481 44680 429247
rect 44836 400110 44864 430879
rect 45020 428913 45048 555999
rect 45190 551576 45246 551585
rect 45190 551511 45246 551520
rect 45204 529009 45232 551511
rect 45374 550488 45430 550497
rect 45374 550423 45430 550432
rect 45388 539617 45416 550423
rect 45374 539608 45430 539617
rect 45374 539543 45430 539552
rect 45190 529000 45246 529009
rect 45190 528935 45246 528944
rect 45006 428904 45062 428913
rect 45006 428839 45062 428848
rect 45098 423192 45154 423201
rect 45098 423127 45154 423136
rect 45112 402937 45140 423127
rect 45466 420744 45522 420753
rect 45466 420679 45522 420688
rect 45282 407280 45338 407289
rect 45282 407215 45338 407224
rect 45296 404326 45324 407215
rect 45284 404320 45336 404326
rect 45284 404262 45336 404268
rect 45098 402928 45154 402937
rect 45098 402863 45154 402872
rect 44824 400104 44876 400110
rect 44824 400046 44876 400052
rect 44638 386472 44694 386481
rect 44638 386407 44694 386416
rect 44454 384840 44510 384849
rect 44454 384775 44510 384784
rect 45098 384432 45154 384441
rect 45098 384367 45154 384376
rect 44270 384024 44326 384033
rect 44270 383959 44326 383968
rect 44914 382256 44970 382265
rect 44914 382191 44970 382200
rect 44638 380352 44694 380361
rect 44638 380287 44694 380296
rect 43810 379808 43866 379817
rect 43810 379743 43866 379752
rect 43824 359961 43852 379743
rect 43994 378176 44050 378185
rect 43994 378111 44050 378120
rect 44008 363633 44036 378111
rect 44270 377496 44326 377505
rect 44270 377431 44326 377440
rect 43994 363624 44050 363633
rect 43994 363559 44050 363568
rect 43810 359952 43866 359961
rect 43810 359887 43866 359896
rect 43626 354784 43682 354793
rect 43626 354719 43682 354728
rect 43442 354240 43498 354249
rect 43442 354175 43498 354184
rect 44284 353161 44312 377431
rect 44652 359009 44680 380287
rect 44638 359000 44694 359009
rect 44638 358935 44694 358944
rect 44640 357468 44692 357474
rect 44640 357410 44692 357416
rect 44652 356017 44680 357410
rect 44638 356008 44694 356017
rect 44638 355943 44694 355952
rect 44640 354544 44692 354550
rect 44454 354512 44510 354521
rect 44510 354492 44640 354498
rect 44510 354486 44692 354492
rect 44510 354470 44680 354486
rect 44454 354447 44510 354456
rect 44732 354408 44784 354414
rect 44732 354350 44784 354356
rect 44744 354249 44772 354350
rect 44730 354240 44786 354249
rect 44730 354175 44786 354184
rect 44270 353152 44326 353161
rect 44270 353087 44326 353096
rect 40222 345536 40278 345545
rect 40222 345471 40278 345480
rect 43258 345536 43314 345545
rect 43258 345471 43314 345480
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 35808 344616 35860 344622
rect 35808 344558 35860 344564
rect 39856 344616 39908 344622
rect 39856 344558 39908 344564
rect 35820 344321 35848 344558
rect 35806 344312 35862 344321
rect 35806 344247 35862 344256
rect 35622 343904 35678 343913
rect 35622 343839 35678 343848
rect 35636 343670 35664 343839
rect 35624 343664 35676 343670
rect 35624 343606 35676 343612
rect 33046 343496 33102 343505
rect 33046 343431 33102 343440
rect 33060 341426 33088 343431
rect 35808 342304 35860 342310
rect 35806 342272 35808 342281
rect 39868 342281 39896 344558
rect 40040 343664 40092 343670
rect 40040 343606 40092 343612
rect 35860 342272 35862 342281
rect 35806 342207 35862 342216
rect 39854 342272 39910 342281
rect 39854 342207 39910 342216
rect 40052 341873 40080 343606
rect 40236 342310 40264 345471
rect 44928 343369 44956 382191
rect 44914 343360 44970 343369
rect 44914 343295 44970 343304
rect 40224 342304 40276 342310
rect 40224 342246 40276 342252
rect 39854 341864 39910 341873
rect 39854 341799 39910 341808
rect 40038 341864 40094 341873
rect 40038 341799 40094 341808
rect 35806 341456 35862 341465
rect 33048 341420 33100 341426
rect 35806 341391 35862 341400
rect 33048 341362 33100 341368
rect 35820 341222 35848 341391
rect 35808 341216 35860 341222
rect 35808 341158 35860 341164
rect 35808 341080 35860 341086
rect 35806 341048 35808 341057
rect 35860 341048 35862 341057
rect 35806 340983 35862 340992
rect 39486 341048 39542 341057
rect 39486 340983 39542 340992
rect 35530 339824 35586 339833
rect 35530 339759 35586 339768
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35544 339522 35572 339759
rect 35820 339658 35848 339759
rect 35808 339652 35860 339658
rect 35808 339594 35860 339600
rect 37924 339652 37976 339658
rect 37924 339594 37976 339600
rect 35532 339516 35584 339522
rect 35532 339458 35584 339464
rect 35806 336152 35862 336161
rect 35806 336087 35862 336096
rect 35820 335374 35848 336087
rect 35808 335368 35860 335374
rect 35808 335310 35860 335316
rect 35806 334520 35862 334529
rect 35806 334455 35862 334464
rect 35820 334150 35848 334455
rect 35808 334144 35860 334150
rect 35808 334086 35860 334092
rect 37936 331265 37964 339594
rect 38660 339516 38712 339522
rect 38660 339458 38712 339464
rect 38672 336569 38700 339458
rect 39500 337385 39528 340983
rect 39868 340241 39896 341799
rect 40222 341456 40278 341465
rect 40222 341391 40224 341400
rect 40276 341391 40278 341400
rect 40224 341362 40276 341368
rect 40224 341216 40276 341222
rect 40224 341158 40276 341164
rect 40040 341080 40092 341086
rect 40236 341057 40264 341158
rect 45112 341057 45140 384367
rect 45282 383616 45338 383625
rect 45282 383551 45338 383560
rect 40040 341022 40092 341028
rect 40222 341048 40278 341057
rect 40052 340649 40080 341022
rect 40222 340983 40278 340992
rect 45098 341048 45154 341057
rect 45098 340983 45154 340992
rect 45296 340649 45324 383551
rect 45480 354074 45508 420679
rect 45650 363080 45706 363089
rect 45650 363015 45706 363024
rect 45664 361554 45692 363015
rect 45652 361548 45704 361554
rect 45652 361490 45704 361496
rect 45834 354784 45890 354793
rect 45834 354719 45890 354728
rect 45650 354376 45706 354385
rect 45650 354311 45652 354320
rect 45704 354311 45706 354320
rect 45652 354282 45704 354288
rect 45848 354210 45876 354719
rect 45836 354204 45888 354210
rect 45836 354146 45888 354152
rect 45468 354068 45520 354074
rect 45468 354010 45520 354016
rect 45468 353932 45520 353938
rect 45468 353874 45520 353880
rect 45480 353705 45508 353874
rect 45466 353696 45522 353705
rect 45466 353631 45522 353640
rect 45468 353456 45520 353462
rect 45466 353424 45468 353433
rect 45520 353424 45522 353433
rect 45466 353359 45522 353368
rect 45422 353184 45474 353190
rect 45420 353152 45422 353161
rect 45474 353152 45476 353161
rect 45420 353087 45476 353096
rect 45466 341456 45522 341465
rect 45466 341391 45468 341400
rect 45520 341391 45522 341400
rect 45468 341362 45520 341368
rect 40038 340640 40094 340649
rect 40038 340575 40094 340584
rect 45282 340640 45338 340649
rect 45282 340575 45338 340584
rect 39670 340232 39726 340241
rect 39670 340167 39726 340176
rect 39854 340232 39910 340241
rect 39854 340167 39910 340176
rect 39684 339833 39712 340167
rect 39670 339824 39726 339833
rect 39670 339759 39726 339768
rect 45650 339280 45706 339289
rect 45650 339215 45706 339224
rect 45466 337648 45522 337657
rect 45466 337583 45522 337592
rect 39486 337376 39542 337385
rect 39486 337311 39542 337320
rect 38658 336560 38714 336569
rect 38658 336495 38714 336504
rect 40224 335368 40276 335374
rect 40224 335310 40276 335316
rect 40236 334529 40264 335310
rect 43994 334656 44050 334665
rect 43994 334591 44050 334600
rect 44270 334656 44326 334665
rect 44270 334591 44326 334600
rect 40222 334520 40278 334529
rect 40222 334455 40278 334464
rect 43074 334520 43130 334529
rect 43074 334455 43130 334464
rect 39764 334144 39816 334150
rect 39764 334086 39816 334092
rect 39776 332897 39804 334086
rect 39762 332888 39818 332897
rect 39762 332823 39818 332832
rect 42890 332888 42946 332897
rect 42890 332823 42946 332832
rect 37922 331256 37978 331265
rect 37922 331191 37978 331200
rect 42168 325938 42196 326264
rect 42168 325910 42288 325938
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42260 324329 42288 325910
rect 42246 324320 42302 324329
rect 42246 324255 42302 324264
rect 42182 323734 42656 323762
rect 42432 322924 42484 322930
rect 42432 322866 42484 322872
rect 42444 322606 42472 322866
rect 42168 322538 42196 322592
rect 42260 322578 42472 322606
rect 42260 322538 42288 322578
rect 42168 322510 42288 322538
rect 42182 321898 42472 321926
rect 42248 321564 42300 321570
rect 42248 321506 42300 321512
rect 42260 321382 42288 321506
rect 42182 321354 42288 321382
rect 41786 321192 41842 321201
rect 41786 321127 41842 321136
rect 41800 320725 41828 321127
rect 42182 320062 42288 320090
rect 42260 319977 42288 320062
rect 41786 319968 41842 319977
rect 41786 319903 41842 319912
rect 42246 319968 42302 319977
rect 42246 319903 42302 319912
rect 41800 319532 41828 319903
rect 42444 319433 42472 321898
rect 42628 320657 42656 323734
rect 42904 321570 42932 332823
rect 43088 322930 43116 334455
rect 43076 322924 43128 322930
rect 43076 322866 43128 322872
rect 42892 321564 42944 321570
rect 42892 321506 42944 321512
rect 42614 320648 42670 320657
rect 42614 320583 42670 320592
rect 42430 319424 42486 319433
rect 42430 319359 42486 319368
rect 41786 317384 41842 317393
rect 41786 317319 41842 317328
rect 41800 317045 41828 317319
rect 42430 316432 42486 316441
rect 42182 316390 42430 316418
rect 42430 316367 42486 316376
rect 41786 316024 41842 316033
rect 41786 315959 41842 315968
rect 41800 315757 41828 315959
rect 42168 315302 42288 315330
rect 42168 315180 42196 315302
rect 42260 315194 42288 315302
rect 42260 315166 42472 315194
rect 41786 313712 41842 313721
rect 41786 313647 41842 313656
rect 41800 313344 41828 313647
rect 42444 313177 42472 315166
rect 42430 313168 42486 313177
rect 42430 313103 42486 313112
rect 42430 312896 42486 312905
rect 42430 312831 42486 312840
rect 42444 312746 42472 312831
rect 42182 312718 42472 312746
rect 42154 312624 42210 312633
rect 42154 312559 42210 312568
rect 42168 312052 42196 312559
rect 42154 311808 42210 311817
rect 42154 311743 42210 311752
rect 42168 311508 42196 311743
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41326 301608 41382 301617
rect 41326 301543 41382 301552
rect 41142 300928 41198 300937
rect 41340 300898 41368 301543
rect 41142 300863 41198 300872
rect 41328 300892 41380 300898
rect 41156 299130 41184 300863
rect 41328 300834 41380 300840
rect 41696 300892 41748 300898
rect 41748 300852 42012 300880
rect 41696 300834 41748 300840
rect 41984 299474 42012 300852
rect 41984 299446 42380 299474
rect 41144 299124 41196 299130
rect 41144 299066 41196 299072
rect 41696 299124 41748 299130
rect 41696 299066 41748 299072
rect 41708 298738 41736 299066
rect 42154 298752 42210 298761
rect 41708 298710 42154 298738
rect 42154 298687 42210 298696
rect 42352 297401 42380 299446
rect 42338 297392 42394 297401
rect 42338 297327 42394 297336
rect 43166 297120 43222 297129
rect 43166 297055 43222 297064
rect 41142 296440 41198 296449
rect 41142 296375 41198 296384
rect 41156 295526 41184 296375
rect 42798 296032 42854 296041
rect 42798 295967 42854 295976
rect 41144 295520 41196 295526
rect 41144 295462 41196 295468
rect 41696 295520 41748 295526
rect 41696 295462 41748 295468
rect 41326 295216 41382 295225
rect 41326 295151 41382 295160
rect 33782 294808 33838 294817
rect 33782 294743 33838 294752
rect 32402 293992 32458 294001
rect 32402 293927 32458 293936
rect 32416 284889 32444 293927
rect 33796 286346 33824 294743
rect 41340 294302 41368 295151
rect 41708 295066 41736 295462
rect 41708 295038 42288 295066
rect 41328 294296 41380 294302
rect 41328 294238 41380 294244
rect 41696 294296 41748 294302
rect 42064 294296 42116 294302
rect 41748 294256 42064 294284
rect 41696 294238 41748 294244
rect 42064 294238 42116 294244
rect 41326 293584 41382 293593
rect 41326 293519 41382 293528
rect 41340 292738 41368 293519
rect 42064 293072 42116 293078
rect 41708 293020 42064 293026
rect 41708 293014 42116 293020
rect 41708 292998 42104 293014
rect 41708 292806 41736 292998
rect 41696 292800 41748 292806
rect 41696 292742 41748 292748
rect 41328 292732 41380 292738
rect 41328 292674 41380 292680
rect 42260 292574 42288 295038
rect 42616 294296 42668 294302
rect 42616 294238 42668 294244
rect 42260 292546 42472 292574
rect 39946 290320 40002 290329
rect 39946 290255 40002 290264
rect 33784 286340 33836 286346
rect 33784 286282 33836 286288
rect 32402 284880 32458 284889
rect 32402 284815 32458 284824
rect 39960 284510 39988 290255
rect 41512 286340 41564 286346
rect 41512 286282 41564 286288
rect 39948 284504 40000 284510
rect 39948 284446 40000 284452
rect 41524 284322 41552 286282
rect 41696 284504 41748 284510
rect 41748 284452 42380 284458
rect 41696 284446 42380 284452
rect 41708 284430 42380 284446
rect 41524 284294 42288 284322
rect 42260 283059 42288 284294
rect 42182 283031 42288 283059
rect 42352 281874 42380 284430
rect 42182 281846 42380 281874
rect 42444 281602 42472 292546
rect 42260 281574 42472 281602
rect 42260 281466 42288 281574
rect 42168 281438 42288 281466
rect 42430 281480 42486 281489
rect 42168 281180 42196 281438
rect 42430 281415 42486 281424
rect 42444 280582 42472 281415
rect 42182 280554 42472 280582
rect 42432 280152 42484 280158
rect 42432 280094 42484 280100
rect 42168 279398 42288 279426
rect 42168 279344 42196 279398
rect 42260 279358 42288 279398
rect 42444 279358 42472 280094
rect 42260 279330 42472 279358
rect 42182 278718 42472 278746
rect 42062 278488 42118 278497
rect 42062 278423 42118 278432
rect 42076 278188 42104 278423
rect 42154 277944 42210 277953
rect 42154 277879 42210 277888
rect 42168 277508 42196 277879
rect 41786 277128 41842 277137
rect 41786 277063 41842 277072
rect 41800 276896 41828 277063
rect 42248 276820 42300 276826
rect 42248 276762 42300 276768
rect 42260 276570 42288 276762
rect 42444 276706 42472 278718
rect 42628 276826 42656 294238
rect 42812 282914 42840 295967
rect 42982 293176 43038 293185
rect 42982 293111 43038 293120
rect 42996 289814 43024 293111
rect 43180 289814 43208 297055
rect 43352 293072 43404 293078
rect 43404 293020 43576 293026
rect 43352 293014 43576 293020
rect 43364 292998 43576 293014
rect 43350 292768 43406 292777
rect 43350 292703 43406 292712
rect 43364 289814 43392 292703
rect 43548 292574 43576 292998
rect 43548 292546 43668 292574
rect 42996 289786 43116 289814
rect 43180 289786 43300 289814
rect 43364 289786 43484 289814
rect 42812 282886 42932 282914
rect 42616 276820 42668 276826
rect 42616 276762 42668 276768
rect 42444 276678 42656 276706
rect 42076 276542 42288 276570
rect 42076 276352 42104 276542
rect 42628 275913 42656 276678
rect 42614 275904 42670 275913
rect 42614 275839 42670 275848
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42168 273170 42196 273224
rect 42338 273184 42394 273193
rect 42168 273142 42338 273170
rect 42338 273119 42394 273128
rect 41786 273048 41842 273057
rect 41786 272983 41842 272992
rect 41800 272544 41828 272983
rect 41786 272368 41842 272377
rect 41786 272303 41842 272312
rect 41800 272000 41828 272303
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 41786 269784 41842 269793
rect 41786 269719 41842 269728
rect 41800 269521 41828 269719
rect 42904 269074 42932 282886
rect 43088 280158 43116 289786
rect 43076 280152 43128 280158
rect 43076 280094 43128 280100
rect 42156 269068 42208 269074
rect 42156 269010 42208 269016
rect 42892 269068 42944 269074
rect 42892 269010 42944 269016
rect 42168 268872 42196 269010
rect 42168 267753 42196 268328
rect 42154 267744 42210 267753
rect 42154 267679 42210 267688
rect 43272 263594 43300 289786
rect 43456 277953 43484 289786
rect 43442 277944 43498 277953
rect 43442 277879 43498 277888
rect 43640 273193 43668 292546
rect 43626 273184 43682 273193
rect 43626 273119 43682 273128
rect 43442 269784 43498 269793
rect 43442 269719 43498 269728
rect 43456 263594 43484 269719
rect 42996 263566 43300 263594
rect 43364 263566 43484 263594
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 40498 257136 40554 257145
rect 40498 257071 40554 257080
rect 35820 256834 35848 257071
rect 40512 256834 40540 257071
rect 35808 256828 35860 256834
rect 35808 256770 35860 256776
rect 40500 256828 40552 256834
rect 40500 256770 40552 256776
rect 42996 256329 43024 263566
rect 43364 257145 43392 263566
rect 43350 257136 43406 257145
rect 43350 257071 43406 257080
rect 35622 256320 35678 256329
rect 35622 256255 35678 256264
rect 40222 256320 40278 256329
rect 40222 256255 40278 256264
rect 42982 256320 43038 256329
rect 42982 256255 43038 256264
rect 35636 255338 35664 256255
rect 35806 255912 35862 255921
rect 35806 255847 35862 255856
rect 35820 255610 35848 255847
rect 35808 255604 35860 255610
rect 35808 255546 35860 255552
rect 39580 255536 39632 255542
rect 39578 255504 39580 255513
rect 39632 255504 39634 255513
rect 39578 255439 39634 255448
rect 35624 255332 35676 255338
rect 35624 255274 35676 255280
rect 39856 255332 39908 255338
rect 39856 255274 39908 255280
rect 39868 254289 39896 255274
rect 35806 254280 35862 254289
rect 35806 254215 35862 254224
rect 39854 254280 39910 254289
rect 39854 254215 39910 254224
rect 35820 254114 35848 254215
rect 40236 254114 40264 256255
rect 43074 255504 43130 255513
rect 43074 255439 43130 255448
rect 42890 254280 42946 254289
rect 42890 254215 42946 254224
rect 35808 254108 35860 254114
rect 35808 254050 35860 254056
rect 40224 254108 40276 254114
rect 40224 254050 40276 254056
rect 35622 253464 35678 253473
rect 35622 253399 35678 253408
rect 35636 252618 35664 253399
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 35820 252754 35848 252991
rect 35808 252748 35860 252754
rect 35808 252690 35860 252696
rect 41328 252748 41380 252754
rect 41328 252690 41380 252696
rect 35624 252612 35676 252618
rect 35624 252554 35676 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 37924 251252 37976 251258
rect 37924 251194 37976 251200
rect 35806 250608 35862 250617
rect 35806 250543 35862 250552
rect 35820 249966 35848 250543
rect 35808 249960 35860 249966
rect 35808 249902 35860 249908
rect 35806 247752 35862 247761
rect 35806 247687 35862 247696
rect 35820 247110 35848 247687
rect 35808 247104 35860 247110
rect 35808 247046 35860 247052
rect 37936 242758 37964 251194
rect 39764 249960 39816 249966
rect 39764 249902 39816 249908
rect 39776 245721 39804 249902
rect 41340 248414 41368 252690
rect 41696 252612 41748 252618
rect 41696 252554 41748 252560
rect 41708 248418 41736 252554
rect 41340 248386 41460 248414
rect 41708 248390 42380 248418
rect 39762 245712 39818 245721
rect 39762 245647 39818 245656
rect 41432 244274 41460 248386
rect 41696 247104 41748 247110
rect 41696 247046 41748 247052
rect 41708 246537 41736 247046
rect 41694 246528 41750 246537
rect 41694 246463 41750 246472
rect 41432 244246 42288 244274
rect 37924 242752 37976 242758
rect 37924 242694 37976 242700
rect 41696 242752 41748 242758
rect 41748 242700 42104 242706
rect 41696 242694 42104 242700
rect 41708 242690 42104 242694
rect 41708 242684 42116 242690
rect 41708 242678 42064 242684
rect 42064 242626 42116 242632
rect 42062 240136 42118 240145
rect 42062 240071 42118 240080
rect 42076 239836 42104 240071
rect 41984 238513 42012 238649
rect 41970 238504 42026 238513
rect 42260 238490 42288 244246
rect 41970 238439 42026 238448
rect 42168 238462 42288 238490
rect 42168 238000 42196 238462
rect 42352 238105 42380 248390
rect 42708 242684 42760 242690
rect 42708 242626 42760 242632
rect 42338 238096 42394 238105
rect 42338 238031 42394 238040
rect 41786 236600 41842 236609
rect 41786 236535 41842 236544
rect 41800 236164 41828 236535
rect 42182 234955 42380 234983
rect 41786 234696 41842 234705
rect 41786 234631 41842 234640
rect 41800 234328 41828 234631
rect 42352 233889 42380 234955
rect 42338 233880 42394 233889
rect 42338 233815 42394 233824
rect 42182 233667 42656 233695
rect 42168 233158 42288 233186
rect 42168 233104 42196 233158
rect 42260 233118 42288 233158
rect 42260 233090 42472 233118
rect 42444 232257 42472 233090
rect 42430 232248 42486 232257
rect 42430 232183 42486 232192
rect 42430 231840 42486 231849
rect 42628 231826 42656 233667
rect 42486 231798 42656 231826
rect 42430 231775 42486 231784
rect 42430 231568 42486 231577
rect 42430 231503 42486 231512
rect 42444 230670 42472 231503
rect 42182 230642 42472 230670
rect 42154 230480 42210 230489
rect 42154 230415 42210 230424
rect 42432 230444 42484 230450
rect 42168 229976 42196 230415
rect 42432 230386 42484 230392
rect 42444 229378 42472 230386
rect 42182 229350 42472 229378
rect 42720 229094 42748 242626
rect 42536 229066 42748 229094
rect 42536 228834 42564 229066
rect 42182 228806 42564 228834
rect 41970 227352 42026 227361
rect 41970 227287 42026 227296
rect 41984 226984 42012 227287
rect 42168 226358 42288 226386
rect 42168 226304 42196 226358
rect 42260 226318 42288 226358
rect 42260 226290 42656 226318
rect 42430 225720 42486 225729
rect 42182 225678 42430 225706
rect 42430 225655 42486 225664
rect 41694 224496 41750 224505
rect 41694 224431 41750 224440
rect 35530 217968 35586 217977
rect 35530 217903 35586 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35544 214305 35572 217903
rect 39946 216472 40002 216481
rect 39946 216407 40002 216416
rect 39578 216200 39634 216209
rect 39578 216135 39634 216144
rect 35530 214296 35586 214305
rect 35530 214231 35586 214240
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 35820 213994 35848 214231
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 35622 213480 35678 213489
rect 35622 213415 35678 213424
rect 35636 212566 35664 213415
rect 35806 213072 35862 213081
rect 35806 213007 35862 213016
rect 35820 212838 35848 213007
rect 35808 212832 35860 212838
rect 35808 212774 35860 212780
rect 39592 212566 39620 216135
rect 39960 212838 39988 216407
rect 41708 213994 41736 224431
rect 42168 223553 42196 225148
rect 42628 224913 42656 226290
rect 42614 224904 42670 224913
rect 42614 224839 42670 224848
rect 42154 223544 42210 223553
rect 42154 223479 42210 223488
rect 42904 216209 42932 254215
rect 43088 216481 43116 255439
rect 43442 246528 43498 246537
rect 43442 246463 43498 246472
rect 43258 245712 43314 245721
rect 43258 245647 43314 245656
rect 43272 230450 43300 245647
rect 43260 230444 43312 230450
rect 43260 230386 43312 230392
rect 43074 216472 43130 216481
rect 43074 216407 43130 216416
rect 42890 216200 42946 216209
rect 42890 216135 42946 216144
rect 43456 215294 43484 246463
rect 44008 231169 44036 334591
rect 44284 319977 44312 334591
rect 45480 325694 45508 337583
rect 45112 325666 45508 325694
rect 44270 319968 44326 319977
rect 44270 319903 44326 319912
rect 45112 316034 45140 325666
rect 45282 320648 45338 320657
rect 45282 320583 45338 320592
rect 45296 317370 45324 320583
rect 45468 317416 45520 317422
rect 45296 317364 45468 317370
rect 45296 317358 45520 317364
rect 45296 317342 45508 317358
rect 45112 316006 45324 316034
rect 45296 312905 45324 316006
rect 45468 314696 45520 314702
rect 45468 314638 45520 314644
rect 45282 312896 45338 312905
rect 45282 312831 45338 312840
rect 45480 311817 45508 314638
rect 45664 312633 45692 339215
rect 45650 312624 45706 312633
rect 45650 312559 45706 312568
rect 45466 311808 45522 311817
rect 45466 311743 45522 311752
rect 45190 300520 45246 300529
rect 45190 300455 45246 300464
rect 44362 299704 44418 299713
rect 44362 299639 44418 299648
rect 44178 299024 44234 299033
rect 44178 298959 44234 298968
rect 44192 256057 44220 298959
rect 44376 256873 44404 299639
rect 44638 298072 44694 298081
rect 44638 298007 44694 298016
rect 44362 256864 44418 256873
rect 44362 256799 44418 256808
rect 44178 256048 44234 256057
rect 44178 255983 44234 255992
rect 44652 255241 44680 298007
rect 45006 292632 45062 292641
rect 45006 292567 45062 292576
rect 45020 281489 45048 292567
rect 45204 292346 45232 300455
rect 45468 295384 45520 295390
rect 45468 295326 45520 295332
rect 45480 292641 45508 295326
rect 45466 292632 45522 292641
rect 45466 292567 45522 292576
rect 45468 292460 45520 292466
rect 45468 292402 45520 292408
rect 45480 292346 45508 292402
rect 45204 292318 45508 292346
rect 45190 291544 45246 291553
rect 45190 291479 45246 291488
rect 45006 281480 45062 281489
rect 45006 281415 45062 281424
rect 45204 278497 45232 291479
rect 45468 285728 45520 285734
rect 45468 285670 45520 285676
rect 45190 278488 45246 278497
rect 45190 278423 45246 278432
rect 45480 277394 45508 285670
rect 44836 277366 45508 277394
rect 44836 258097 44864 277366
rect 44822 258088 44878 258097
rect 44822 258023 44878 258032
rect 44638 255232 44694 255241
rect 44638 255167 44694 255176
rect 44270 254824 44326 254833
rect 44270 254759 44326 254768
rect 43994 231160 44050 231169
rect 43994 231095 44050 231104
rect 43180 215266 43484 215294
rect 41696 213988 41748 213994
rect 41696 213930 41748 213936
rect 39948 212832 40000 212838
rect 39948 212774 40000 212780
rect 35624 212560 35676 212566
rect 35624 212502 35676 212508
rect 39580 212560 39632 212566
rect 39580 212502 39632 212508
rect 35806 210216 35862 210225
rect 35806 210151 35862 210160
rect 35820 209982 35848 210151
rect 35808 209976 35860 209982
rect 35808 209918 35860 209924
rect 40408 209976 40460 209982
rect 40408 209918 40460 209924
rect 35622 209400 35678 209409
rect 35622 209335 35678 209344
rect 35636 208418 35664 209335
rect 40420 209001 40448 209918
rect 35806 208992 35862 209001
rect 35806 208927 35862 208936
rect 40406 208992 40462 209001
rect 40406 208927 40462 208936
rect 42890 208992 42946 209001
rect 42890 208927 42946 208936
rect 35820 208758 35848 208927
rect 35808 208752 35860 208758
rect 35808 208694 35860 208700
rect 40040 208684 40092 208690
rect 40040 208626 40092 208632
rect 35806 208584 35862 208593
rect 35806 208519 35808 208528
rect 35860 208519 35862 208528
rect 35808 208490 35860 208496
rect 35624 208412 35676 208418
rect 35624 208354 35676 208360
rect 40052 208185 40080 208626
rect 40592 208548 40644 208554
rect 40592 208490 40644 208496
rect 40038 208176 40094 208185
rect 40038 208111 40094 208120
rect 35806 207360 35862 207369
rect 35806 207295 35862 207304
rect 35820 207194 35848 207295
rect 35808 207188 35860 207194
rect 35808 207130 35860 207136
rect 39948 207188 40000 207194
rect 39948 207130 40000 207136
rect 35806 205320 35862 205329
rect 35806 205255 35862 205264
rect 35820 204678 35848 205255
rect 35808 204672 35860 204678
rect 35808 204614 35860 204620
rect 35806 204504 35862 204513
rect 35806 204439 35862 204448
rect 35820 204338 35848 204439
rect 35808 204332 35860 204338
rect 35808 204274 35860 204280
rect 39960 203697 39988 207130
rect 40604 206961 40632 208490
rect 41708 208418 42104 208434
rect 41696 208412 42116 208418
rect 41748 208406 42064 208412
rect 41696 208354 41748 208360
rect 42064 208354 42116 208360
rect 40590 206952 40646 206961
rect 40590 206887 40646 206896
rect 42706 206952 42762 206961
rect 42706 206887 42762 206896
rect 41512 204536 41564 204542
rect 41510 204504 41512 204513
rect 41564 204504 41566 204513
rect 41510 204439 41566 204448
rect 41696 204400 41748 204406
rect 41696 204342 41748 204348
rect 41708 204105 41736 204342
rect 41694 204096 41750 204105
rect 41694 204031 41750 204040
rect 35806 203688 35862 203697
rect 35806 203623 35862 203632
rect 39946 203688 40002 203697
rect 39946 203623 40002 203632
rect 35820 202910 35848 203623
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 37924 202904 37976 202910
rect 37924 202846 37976 202852
rect 42720 202874 42748 206887
rect 42720 202846 42840 202874
rect 37936 198801 37964 202846
rect 42812 202722 42840 202846
rect 42720 202694 42840 202722
rect 42524 201748 42576 201754
rect 42524 201690 42576 201696
rect 37922 198792 37978 198801
rect 37922 198727 37978 198736
rect 42536 197962 42564 201690
rect 42720 201618 42748 202694
rect 42904 201754 42932 208927
rect 43180 208162 43208 215266
rect 44284 212129 44312 254759
rect 44914 254008 44970 254017
rect 44914 253943 44970 253952
rect 44546 251560 44602 251569
rect 44546 251495 44602 251504
rect 44560 240145 44588 251495
rect 44730 250336 44786 250345
rect 44730 250271 44786 250280
rect 44546 240136 44602 240145
rect 44546 240071 44602 240080
rect 44744 234614 44772 250271
rect 44928 234614 44956 253943
rect 45558 252784 45614 252793
rect 45558 252719 45614 252728
rect 45098 249112 45154 249121
rect 45098 249047 45154 249056
rect 45112 234614 45140 249047
rect 44652 234586 44772 234614
rect 44836 234586 44956 234614
rect 45020 234586 45140 234614
rect 44652 230489 44680 234586
rect 44638 230480 44694 230489
rect 44638 230415 44694 230424
rect 44270 212120 44326 212129
rect 44270 212055 44326 212064
rect 44836 211313 44864 234586
rect 45020 231577 45048 234586
rect 45006 231568 45062 231577
rect 45006 231503 45062 231512
rect 45572 225729 45600 252719
rect 45834 248704 45890 248713
rect 45834 248639 45890 248648
rect 45848 231849 45876 248639
rect 46018 248296 46074 248305
rect 46018 248231 46074 248240
rect 46032 233209 46060 248231
rect 46018 233200 46074 233209
rect 46018 233135 46074 233144
rect 45834 231840 45890 231849
rect 45834 231775 45890 231784
rect 46216 231334 46244 610846
rect 46938 578232 46994 578241
rect 46938 578167 46994 578176
rect 46952 574054 46980 578167
rect 46940 574048 46992 574054
rect 46940 573990 46992 573996
rect 47582 558512 47638 558521
rect 47582 558447 47638 558456
rect 47596 527134 47624 558447
rect 47584 527128 47636 527134
rect 47584 527070 47636 527076
rect 47582 489968 47638 489977
rect 47582 489903 47638 489912
rect 46386 376136 46442 376145
rect 46386 376071 46442 376080
rect 46400 300830 46428 376071
rect 46938 338872 46994 338881
rect 46938 338807 46994 338816
rect 46952 313177 46980 338807
rect 47122 337920 47178 337929
rect 47122 337855 47178 337864
rect 47136 324329 47164 337855
rect 47122 324320 47178 324329
rect 47122 324255 47178 324264
rect 46938 313168 46994 313177
rect 46938 313103 46994 313112
rect 46388 300824 46440 300830
rect 46388 300766 46440 300772
rect 47596 299470 47624 489903
rect 47766 430536 47822 430545
rect 47766 430471 47822 430480
rect 47780 398818 47808 430471
rect 47768 398812 47820 398818
rect 47768 398754 47820 398760
rect 47766 387696 47822 387705
rect 47766 387631 47822 387640
rect 47780 356046 47808 387631
rect 47768 356040 47820 356046
rect 47768 355982 47820 355988
rect 47766 354376 47822 354385
rect 47766 354311 47822 354320
rect 47584 299464 47636 299470
rect 47584 299406 47636 299412
rect 47582 290728 47638 290737
rect 47582 290663 47638 290672
rect 46388 284368 46440 284374
rect 46388 284310 46440 284316
rect 46400 257689 46428 284310
rect 46386 257680 46442 257689
rect 46386 257615 46442 257624
rect 47214 251968 47270 251977
rect 47214 251903 47270 251912
rect 46938 251152 46994 251161
rect 46938 251087 46994 251096
rect 46204 231328 46256 231334
rect 46204 231270 46256 231276
rect 45558 225720 45614 225729
rect 45558 225655 45614 225664
rect 46952 224913 46980 251087
rect 47228 232257 47256 251903
rect 47398 247072 47454 247081
rect 47398 247007 47454 247016
rect 47412 238513 47440 247007
rect 47398 238504 47454 238513
rect 47398 238439 47454 238448
rect 47214 232248 47270 232257
rect 47214 232183 47270 232192
rect 46938 224904 46994 224913
rect 46938 224839 46994 224848
rect 44822 211304 44878 211313
rect 44822 211239 44878 211248
rect 44454 208448 44510 208457
rect 43352 208412 43404 208418
rect 44454 208383 44510 208392
rect 43352 208354 43404 208360
rect 42996 208134 43208 208162
rect 42996 202874 43024 208134
rect 43364 205634 43392 208354
rect 44178 207768 44234 207777
rect 44178 207703 44234 207712
rect 43364 205606 43944 205634
rect 43718 204504 43774 204513
rect 43718 204439 43774 204448
rect 43442 204096 43498 204105
rect 43442 204031 43498 204040
rect 43258 203688 43314 203697
rect 43258 203623 43314 203632
rect 42996 202846 43116 202874
rect 43088 201770 43116 202846
rect 43272 202162 43300 203623
rect 43260 202156 43312 202162
rect 43260 202098 43312 202104
rect 42892 201748 42944 201754
rect 43088 201742 43300 201770
rect 42892 201690 42944 201696
rect 42708 201612 42760 201618
rect 42708 201554 42760 201560
rect 43076 201612 43128 201618
rect 43076 201554 43128 201560
rect 42892 201340 42944 201346
rect 42892 201282 42944 201288
rect 42536 197934 42840 197962
rect 42430 197296 42486 197305
rect 42430 197231 42486 197240
rect 42444 196670 42472 197231
rect 42182 196642 42472 196670
rect 41970 195664 42026 195673
rect 41970 195599 42026 195608
rect 41984 195432 42012 195599
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42246 194984 42302 194993
rect 42246 194919 42302 194928
rect 41786 193488 41842 193497
rect 41786 193423 41842 193432
rect 41800 192984 41828 193423
rect 42076 191593 42104 191760
rect 42062 191584 42118 191593
rect 42062 191519 42118 191528
rect 42168 191026 42196 191148
rect 42260 191026 42288 194919
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42812 190346 42840 197934
rect 42720 190318 42840 190346
rect 42248 190256 42300 190262
rect 42248 190198 42300 190204
rect 42260 189938 42288 190198
rect 42182 189910 42288 189938
rect 42432 187672 42484 187678
rect 42246 187640 42302 187649
rect 42432 187614 42484 187620
rect 42246 187575 42302 187584
rect 42260 187459 42288 187575
rect 42182 187431 42288 187459
rect 42444 186810 42472 187614
rect 42182 186782 42472 186810
rect 41786 186416 41842 186425
rect 41786 186351 41842 186360
rect 41800 186184 41828 186351
rect 41786 186008 41842 186017
rect 41786 185943 41842 185952
rect 41800 185605 41828 185943
rect 42720 183779 42748 190318
rect 42904 190262 42932 201282
rect 42892 190256 42944 190262
rect 42892 190198 42944 190204
rect 43088 187678 43116 201554
rect 43076 187672 43128 187678
rect 43076 187614 43128 187620
rect 43272 186314 43300 201742
rect 43456 192386 43484 204031
rect 43456 192358 43576 192386
rect 43548 186314 43576 192358
rect 43732 190505 43760 204439
rect 43718 190496 43774 190505
rect 43718 190431 43774 190440
rect 43272 186286 43484 186314
rect 43548 186286 43668 186314
rect 42182 183751 42748 183779
rect 42430 183560 42486 183569
rect 42430 183495 42486 183504
rect 42246 183288 42302 183297
rect 42246 183223 42302 183232
rect 42260 183138 42288 183223
rect 42182 183110 42288 183138
rect 42444 182491 42472 183495
rect 42182 182463 42472 182491
rect 42076 180849 42104 181900
rect 42062 180840 42118 180849
rect 42062 180775 42118 180784
rect 43456 44198 43484 186286
rect 43640 44334 43668 186286
rect 43916 183569 43944 205606
rect 43902 183560 43958 183569
rect 43902 183495 43958 183504
rect 44192 183297 44220 207703
rect 44468 197305 44496 208383
rect 44638 206000 44694 206009
rect 44638 205935 44694 205944
rect 44454 197296 44510 197305
rect 44454 197231 44510 197240
rect 44652 187649 44680 205935
rect 44822 205184 44878 205193
rect 44822 205119 44878 205128
rect 44836 191593 44864 205119
rect 46202 204912 46258 204921
rect 46202 204847 46258 204856
rect 44822 191584 44878 191593
rect 44822 191519 44878 191528
rect 44638 187640 44694 187649
rect 44638 187575 44694 187584
rect 44178 183288 44234 183297
rect 44178 183223 44234 183232
rect 46216 49026 46244 204847
rect 47596 52018 47624 290663
rect 47780 278050 47808 354311
rect 47768 278044 47820 278050
rect 47768 277986 47820 277992
rect 47766 247480 47822 247489
rect 47766 247415 47822 247424
rect 47584 52012 47636 52018
rect 47584 51954 47636 51960
rect 47780 50386 47808 247415
rect 48976 53106 49004 761874
rect 50160 611312 50212 611318
rect 50160 611254 50212 611260
rect 50172 610026 50200 611254
rect 50160 610020 50212 610026
rect 50160 609962 50212 609968
rect 49330 418840 49386 418849
rect 49330 418775 49386 418784
rect 49146 334112 49202 334121
rect 49146 334047 49202 334056
rect 49160 53242 49188 334047
rect 49344 278594 49372 418775
rect 49332 278588 49384 278594
rect 49332 278530 49384 278536
rect 49148 53236 49200 53242
rect 49148 53178 49200 53184
rect 48964 53100 49016 53106
rect 48964 53042 49016 53048
rect 50356 51882 50384 806074
rect 53104 799060 53156 799066
rect 53104 799002 53156 799008
rect 53116 790770 53144 799002
rect 57244 797700 57296 797706
rect 57244 797642 57296 797648
rect 53104 790764 53156 790770
rect 53104 790706 53156 790712
rect 57256 789206 57284 797642
rect 57244 789200 57296 789206
rect 57244 789142 57296 789148
rect 60016 786554 60044 816954
rect 62948 810756 63000 810762
rect 62948 810698 63000 810704
rect 62672 805996 62724 806002
rect 62672 805938 62724 805944
rect 62212 790764 62264 790770
rect 62212 790706 62264 790712
rect 62224 790537 62252 790706
rect 62210 790528 62266 790537
rect 62210 790463 62266 790472
rect 62120 789200 62172 789206
rect 62118 789168 62120 789177
rect 62172 789168 62174 789177
rect 62118 789103 62174 789112
rect 62118 787400 62174 787409
rect 62118 787335 62174 787344
rect 62132 786690 62160 787335
rect 62120 786684 62172 786690
rect 62120 786626 62172 786632
rect 60004 786548 60056 786554
rect 60004 786490 60056 786496
rect 62304 786548 62356 786554
rect 62304 786490 62356 786496
rect 62316 786185 62344 786490
rect 62302 786176 62358 786185
rect 62302 786111 62358 786120
rect 62120 785188 62172 785194
rect 62120 785130 62172 785136
rect 62132 784961 62160 785130
rect 62118 784952 62174 784961
rect 62118 784887 62174 784896
rect 58624 774240 58676 774246
rect 58624 774182 58676 774188
rect 58636 742422 58664 774182
rect 61384 772880 61436 772886
rect 61384 772822 61436 772828
rect 60004 763224 60056 763230
rect 60004 763166 60056 763172
rect 58624 742416 58676 742422
rect 58624 742358 58676 742364
rect 53104 719024 53156 719030
rect 53104 718966 53156 718972
rect 51724 712156 51776 712162
rect 51724 712098 51776 712104
rect 51736 705158 51764 712098
rect 51724 705152 51776 705158
rect 51724 705094 51776 705100
rect 51722 538248 51778 538257
rect 51722 538183 51778 538192
rect 51736 531282 51764 538183
rect 51724 531276 51776 531282
rect 51724 531218 51776 531224
rect 51446 404968 51502 404977
rect 51446 404903 51502 404912
rect 51460 402966 51488 404903
rect 51448 402960 51500 402966
rect 51448 402902 51500 402908
rect 51080 400240 51132 400246
rect 51080 400182 51132 400188
rect 51092 395729 51120 400182
rect 51078 395720 51134 395729
rect 51078 395655 51134 395664
rect 51078 362264 51134 362273
rect 51078 362199 51134 362208
rect 51092 360194 51120 362199
rect 51080 360188 51132 360194
rect 51080 360130 51132 360136
rect 51906 353696 51962 353705
rect 51906 353631 51962 353640
rect 50526 291136 50582 291145
rect 50526 291071 50582 291080
rect 50344 51876 50396 51882
rect 50344 51818 50396 51824
rect 47768 50380 47820 50386
rect 47768 50322 47820 50328
rect 50540 49162 50568 291071
rect 51724 282940 51776 282946
rect 51724 282882 51776 282888
rect 51736 180849 51764 282882
rect 51920 278186 51948 353631
rect 52092 300824 52144 300830
rect 52092 300766 52144 300772
rect 52104 278322 52132 300766
rect 52092 278316 52144 278322
rect 52092 278258 52144 278264
rect 51908 278180 51960 278186
rect 51908 278122 51960 278128
rect 53116 264761 53144 718966
rect 57244 676252 57296 676258
rect 57244 676194 57296 676200
rect 55862 611688 55918 611697
rect 55862 611623 55918 611632
rect 54484 299464 54536 299470
rect 54484 299406 54536 299412
rect 54496 288454 54524 299406
rect 54484 288448 54536 288454
rect 54484 288390 54536 288396
rect 53288 276684 53340 276690
rect 53288 276626 53340 276632
rect 53102 264752 53158 264761
rect 53102 264687 53158 264696
rect 53300 215121 53328 276626
rect 55876 264246 55904 611623
rect 56048 281580 56100 281586
rect 56048 281522 56100 281528
rect 55864 264240 55916 264246
rect 55864 264182 55916 264188
rect 55680 218204 55732 218210
rect 55680 218146 55732 218152
rect 55692 217138 55720 218146
rect 56060 217977 56088 281522
rect 57256 278089 57284 676194
rect 58624 669384 58676 669390
rect 58624 669326 58676 669332
rect 58636 660958 58664 669326
rect 58624 660952 58676 660958
rect 58624 660894 58676 660900
rect 58624 644496 58676 644502
rect 58624 644438 58676 644444
rect 58636 612678 58664 644438
rect 58624 612672 58676 612678
rect 58624 612614 58676 612620
rect 57428 294092 57480 294098
rect 57428 294034 57480 294040
rect 57242 278080 57298 278089
rect 57242 278015 57298 278024
rect 57440 275913 57468 294034
rect 57612 288448 57664 288454
rect 57612 288390 57664 288396
rect 57624 278730 57652 288390
rect 58624 280084 58676 280090
rect 58624 280026 58676 280032
rect 57612 278724 57664 278730
rect 57612 278666 57664 278672
rect 57426 275904 57482 275913
rect 57426 275839 57482 275848
rect 57244 228404 57296 228410
rect 57244 228346 57296 228352
rect 56508 227044 56560 227050
rect 56508 226986 56560 226992
rect 56520 218210 56548 226986
rect 56508 218204 56560 218210
rect 56508 218146 56560 218152
rect 57256 218074 57284 228346
rect 58636 223553 58664 280026
rect 60016 278361 60044 763166
rect 61396 747318 61424 772822
rect 61384 747312 61436 747318
rect 61384 747254 61436 747260
rect 62120 746564 62172 746570
rect 62120 746506 62172 746512
rect 62132 746201 62160 746506
rect 62118 746192 62174 746201
rect 62118 746127 62174 746136
rect 62118 744152 62174 744161
rect 62118 744087 62174 744096
rect 62132 743918 62160 744087
rect 62120 743912 62172 743918
rect 62120 743854 62172 743860
rect 62120 743776 62172 743782
rect 62118 743744 62120 743753
rect 62172 743744 62174 743753
rect 62118 743679 62174 743688
rect 62120 742416 62172 742422
rect 62118 742384 62120 742393
rect 62172 742384 62174 742393
rect 62118 742319 62174 742328
rect 61384 730108 61436 730114
rect 61384 730050 61436 730056
rect 61396 699689 61424 730050
rect 62120 705152 62172 705158
rect 62120 705094 62172 705100
rect 62132 704449 62160 705094
rect 62118 704440 62174 704449
rect 62118 704375 62174 704384
rect 62120 703792 62172 703798
rect 62120 703734 62172 703740
rect 62132 703361 62160 703734
rect 62118 703352 62174 703361
rect 62118 703287 62174 703296
rect 61382 699680 61438 699689
rect 61382 699615 61438 699624
rect 62212 698284 62264 698290
rect 62212 698226 62264 698232
rect 62224 698057 62252 698226
rect 62210 698048 62266 698057
rect 62210 697983 62266 697992
rect 61384 667956 61436 667962
rect 61384 667898 61436 667904
rect 61396 659569 61424 667898
rect 62120 660952 62172 660958
rect 62118 660920 62120 660929
rect 62172 660920 62174 660929
rect 62118 660855 62174 660864
rect 61382 659560 61438 659569
rect 61382 659495 61438 659504
rect 62118 658336 62174 658345
rect 62118 658271 62174 658280
rect 62132 657558 62160 658271
rect 62120 657552 62172 657558
rect 62120 657494 62172 657500
rect 62120 656872 62172 656878
rect 62120 656814 62172 656820
rect 62132 656577 62160 656814
rect 62118 656568 62174 656577
rect 62118 656503 62174 656512
rect 62120 655512 62172 655518
rect 62120 655454 62172 655460
rect 62132 655353 62160 655454
rect 62118 655344 62174 655353
rect 62118 655279 62174 655288
rect 61384 643136 61436 643142
rect 61384 643078 61436 643084
rect 60188 633480 60240 633486
rect 60188 633422 60240 633428
rect 60002 278352 60058 278361
rect 60002 278287 60058 278296
rect 60200 277409 60228 633422
rect 61396 613873 61424 643078
rect 62120 616820 62172 616826
rect 62120 616762 62172 616768
rect 62132 616593 62160 616762
rect 62118 616584 62174 616593
rect 62118 616519 62174 616528
rect 62118 614680 62174 614689
rect 62118 614615 62174 614624
rect 62132 614174 62160 614615
rect 62120 614168 62172 614174
rect 62120 614110 62172 614116
rect 61382 613864 61438 613873
rect 61382 613799 61438 613808
rect 62120 612672 62172 612678
rect 62118 612640 62120 612649
rect 62172 612640 62174 612649
rect 62118 612575 62174 612584
rect 61384 610020 61436 610026
rect 61384 609962 61436 609968
rect 60372 292596 60424 292602
rect 60372 292538 60424 292544
rect 60186 277400 60242 277409
rect 60186 277335 60242 277344
rect 60384 267753 60412 292538
rect 60556 278588 60608 278594
rect 60556 278530 60608 278536
rect 60568 278322 60596 278530
rect 60556 278316 60608 278322
rect 60556 278258 60608 278264
rect 60370 267744 60426 267753
rect 60370 267679 60426 267688
rect 61396 264382 61424 609962
rect 62486 590064 62542 590073
rect 62486 589999 62542 590008
rect 62120 575476 62172 575482
rect 62120 575418 62172 575424
rect 62132 574841 62160 575418
rect 62118 574832 62174 574841
rect 62118 574767 62174 574776
rect 62120 574048 62172 574054
rect 62120 573990 62172 573996
rect 62132 573617 62160 573990
rect 62118 573608 62174 573617
rect 62118 573543 62174 573552
rect 62500 569945 62528 589999
rect 62486 569936 62542 569945
rect 62486 569871 62542 569880
rect 62486 556744 62542 556753
rect 62486 556679 62542 556688
rect 62120 532024 62172 532030
rect 62120 531966 62172 531972
rect 62132 531185 62160 531966
rect 62304 531276 62356 531282
rect 62304 531218 62356 531224
rect 62118 531176 62174 531185
rect 62118 531111 62174 531120
rect 62316 530641 62344 531218
rect 62302 530632 62358 530641
rect 62302 530567 62358 530576
rect 62120 528624 62172 528630
rect 62118 528592 62120 528601
rect 62172 528592 62174 528601
rect 62118 528527 62174 528536
rect 62500 528057 62528 556679
rect 62486 528048 62542 528057
rect 62486 527983 62542 527992
rect 62120 527128 62172 527134
rect 62118 527096 62120 527105
rect 62172 527096 62174 527105
rect 62118 527031 62174 527040
rect 62486 427136 62542 427145
rect 62486 427071 62542 427080
rect 62500 422294 62528 427071
rect 62500 422266 62620 422294
rect 62120 404320 62172 404326
rect 62120 404262 62172 404268
rect 62132 404161 62160 404262
rect 62118 404152 62174 404161
rect 62118 404087 62174 404096
rect 62592 402974 62620 422266
rect 62120 402960 62172 402966
rect 62120 402902 62172 402908
rect 62500 402946 62620 402974
rect 62132 402665 62160 402902
rect 62118 402656 62174 402665
rect 62118 402591 62174 402600
rect 62118 400616 62174 400625
rect 62118 400551 62174 400560
rect 62132 400246 62160 400551
rect 62120 400240 62172 400246
rect 62500 400217 62528 402946
rect 62120 400182 62172 400188
rect 62486 400208 62542 400217
rect 62486 400143 62542 400152
rect 62120 400104 62172 400110
rect 62120 400046 62172 400052
rect 62132 399401 62160 400046
rect 62118 399392 62174 399401
rect 62118 399327 62174 399336
rect 62120 398812 62172 398818
rect 62120 398754 62172 398760
rect 62132 398313 62160 398754
rect 62118 398304 62174 398313
rect 62118 398239 62174 398248
rect 62486 385928 62542 385937
rect 62486 385863 62542 385872
rect 62120 361548 62172 361554
rect 62120 361490 62172 361496
rect 62132 360913 62160 361490
rect 62118 360904 62174 360913
rect 62118 360839 62174 360848
rect 62120 360188 62172 360194
rect 62120 360130 62172 360136
rect 62132 359825 62160 360130
rect 62118 359816 62174 359825
rect 62118 359751 62174 359760
rect 62118 357776 62174 357785
rect 62118 357711 62174 357720
rect 62132 357474 62160 357711
rect 62120 357468 62172 357474
rect 62120 357410 62172 357416
rect 62500 357377 62528 385863
rect 62486 357368 62542 357377
rect 62486 357303 62542 357312
rect 62120 356040 62172 356046
rect 62118 356008 62120 356017
rect 62172 356008 62174 356017
rect 62118 355943 62174 355952
rect 62486 341728 62542 341737
rect 62486 341663 62542 341672
rect 62304 341420 62356 341426
rect 62304 341362 62356 341368
rect 61566 319424 61622 319433
rect 61566 319359 61622 319368
rect 61580 316033 61608 319359
rect 62120 317416 62172 317422
rect 62118 317384 62120 317393
rect 62172 317384 62174 317393
rect 62118 317319 62174 317328
rect 61566 316024 61622 316033
rect 61566 315959 61622 315968
rect 62118 314800 62174 314809
rect 62118 314735 62120 314744
rect 62172 314735 62174 314744
rect 62120 314706 62172 314712
rect 62316 314129 62344 341362
rect 62302 314120 62358 314129
rect 62302 314055 62358 314064
rect 62500 313041 62528 341663
rect 62486 313032 62542 313041
rect 62486 312967 62542 312976
rect 62486 297392 62542 297401
rect 62486 297327 62542 297336
rect 62118 295760 62174 295769
rect 62118 295695 62174 295704
rect 62132 295390 62160 295695
rect 62120 295384 62172 295390
rect 62120 295326 62172 295332
rect 62118 294128 62174 294137
rect 62118 294063 62120 294072
rect 62172 294063 62174 294072
rect 62120 294034 62172 294040
rect 62302 292768 62358 292777
rect 62302 292703 62358 292712
rect 62316 292602 62344 292703
rect 62304 292596 62356 292602
rect 62304 292538 62356 292544
rect 62118 292496 62174 292505
rect 62118 292431 62120 292440
rect 62172 292431 62174 292440
rect 62120 292402 62172 292408
rect 62500 291009 62528 297327
rect 62486 291000 62542 291009
rect 62486 290935 62542 290944
rect 62210 288552 62266 288561
rect 62210 288487 62266 288496
rect 62224 287054 62252 288487
rect 62394 287192 62450 287201
rect 62394 287127 62450 287136
rect 62224 287026 62344 287054
rect 62118 285968 62174 285977
rect 62118 285903 62174 285912
rect 62132 285734 62160 285903
rect 62120 285728 62172 285734
rect 62120 285670 62172 285676
rect 62118 283248 62174 283257
rect 62118 283183 62174 283192
rect 62132 282946 62160 283183
rect 62120 282940 62172 282946
rect 62120 282882 62172 282888
rect 62316 281058 62344 287026
rect 61948 281030 62344 281058
rect 61948 280090 61976 281030
rect 62118 280936 62174 280945
rect 62118 280871 62174 280880
rect 61936 280084 61988 280090
rect 61936 280026 61988 280032
rect 61752 278724 61804 278730
rect 61752 278666 61804 278672
rect 61764 278322 61792 278666
rect 61936 278588 61988 278594
rect 61936 278530 61988 278536
rect 61752 278316 61804 278322
rect 61752 278258 61804 278264
rect 61948 277642 61976 278530
rect 61936 277636 61988 277642
rect 61936 277578 61988 277584
rect 62132 276690 62160 280871
rect 62120 276684 62172 276690
rect 62120 276626 62172 276632
rect 62408 269793 62436 287127
rect 62394 269784 62450 269793
rect 62394 269719 62450 269728
rect 61384 264376 61436 264382
rect 61384 264318 61436 264324
rect 61384 228540 61436 228546
rect 61384 228482 61436 228488
rect 60648 227588 60700 227594
rect 60648 227530 60700 227536
rect 58622 223544 58678 223553
rect 58622 223479 58678 223488
rect 59360 221468 59412 221474
rect 59360 221410 59412 221416
rect 58992 218748 59044 218754
rect 58992 218690 59044 218696
rect 57428 218204 57480 218210
rect 57428 218146 57480 218152
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57244 218068 57296 218074
rect 57244 218010 57296 218016
rect 56046 217968 56102 217977
rect 56046 217903 56102 217912
rect 56520 217138 56548 218010
rect 57440 217274 57468 218146
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 55646 217110 55720 217138
rect 56474 217110 56548 217138
rect 57302 217246 57468 217274
rect 55646 216988 55674 217110
rect 56474 216988 56502 217110
rect 57302 216988 57330 217246
rect 58176 217138 58204 218010
rect 59004 217138 59032 218690
rect 59372 218074 59400 221410
rect 59820 218884 59872 218890
rect 59820 218826 59872 218832
rect 59360 218068 59412 218074
rect 59360 218010 59412 218016
rect 59832 217138 59860 218826
rect 60660 217274 60688 227530
rect 61396 218210 61424 228482
rect 62684 224233 62712 805938
rect 62960 787137 62988 810698
rect 653404 790832 653456 790838
rect 653404 790774 653456 790780
rect 62946 787128 63002 787137
rect 62946 787063 63002 787072
rect 651470 778424 651526 778433
rect 651470 778359 651526 778368
rect 651484 777646 651512 778359
rect 651472 777640 651524 777646
rect 651472 777582 651524 777588
rect 652022 777064 652078 777073
rect 652022 776999 652078 777008
rect 651470 776112 651526 776121
rect 651470 776047 651526 776056
rect 651484 775606 651512 776047
rect 651472 775600 651524 775606
rect 651472 775542 651524 775548
rect 651380 775328 651432 775334
rect 651378 775296 651380 775305
rect 651432 775296 651434 775305
rect 651378 775231 651434 775240
rect 651470 774208 651526 774217
rect 651470 774143 651472 774152
rect 651524 774143 651526 774152
rect 651472 774114 651524 774120
rect 651472 773832 651524 773838
rect 651472 773774 651524 773780
rect 651484 773401 651512 773774
rect 651470 773392 651526 773401
rect 651470 773327 651526 773336
rect 62948 755540 63000 755546
rect 62948 755482 63000 755488
rect 62960 747697 62988 755482
rect 62946 747688 63002 747697
rect 62946 747623 63002 747632
rect 63040 747312 63092 747318
rect 63040 747254 63092 747260
rect 63052 741849 63080 747254
rect 63038 741840 63094 741849
rect 63038 741775 63094 741784
rect 652036 736914 652064 776999
rect 653416 775334 653444 790774
rect 670608 784304 670660 784310
rect 670608 784246 670660 784252
rect 669228 784168 669280 784174
rect 669228 784110 669280 784116
rect 669044 782536 669096 782542
rect 669044 782478 669096 782484
rect 655520 781108 655572 781114
rect 655520 781050 655572 781056
rect 655060 778388 655112 778394
rect 655060 778330 655112 778336
rect 653404 775328 653456 775334
rect 653404 775270 653456 775276
rect 655072 773838 655100 778330
rect 655532 774178 655560 781050
rect 660304 777640 660356 777646
rect 660304 777582 660356 777588
rect 655520 774172 655572 774178
rect 655520 774114 655572 774120
rect 655060 773832 655112 773838
rect 655060 773774 655112 773780
rect 653404 746632 653456 746638
rect 653404 746574 653456 746580
rect 652024 736908 652076 736914
rect 652024 736850 652076 736856
rect 651470 734224 651526 734233
rect 651470 734159 651526 734168
rect 651484 733446 651512 734159
rect 651472 733440 651524 733446
rect 651472 733382 651524 733388
rect 652666 732864 652722 732873
rect 652666 732799 652722 732808
rect 651470 731776 651526 731785
rect 651470 731711 651526 731720
rect 651484 731474 651512 731711
rect 651472 731468 651524 731474
rect 651472 731410 651524 731416
rect 651380 731128 651432 731134
rect 651378 731096 651380 731105
rect 651432 731096 651434 731105
rect 651378 731031 651434 731040
rect 652680 730726 652708 732799
rect 653416 731134 653444 746574
rect 656164 736908 656216 736914
rect 656164 736850 656216 736856
rect 654784 734188 654836 734194
rect 654784 734130 654836 734136
rect 653404 731128 653456 731134
rect 653404 731070 653456 731076
rect 652668 730720 652720 730726
rect 652668 730662 652720 730668
rect 651472 730040 651524 730046
rect 651472 729982 651524 729988
rect 651484 729881 651512 729982
rect 651470 729872 651526 729881
rect 651470 729807 651526 729816
rect 62948 729360 63000 729366
rect 62948 729302 63000 729308
rect 62960 712094 62988 729302
rect 654796 728550 654824 734130
rect 651472 728544 651524 728550
rect 651470 728512 651472 728521
rect 654784 728544 654836 728550
rect 651524 728512 651526 728521
rect 654784 728486 654836 728492
rect 651470 728447 651526 728456
rect 656176 716310 656204 736850
rect 657544 735616 657596 735622
rect 657544 735558 657596 735564
rect 657556 730046 657584 735558
rect 658924 731468 658976 731474
rect 658924 731410 658976 731416
rect 657544 730040 657596 730046
rect 657544 729982 657596 729988
rect 656164 716304 656216 716310
rect 656164 716246 656216 716252
rect 62960 712066 63172 712094
rect 62946 701312 63002 701321
rect 62946 701247 63002 701256
rect 62960 701078 62988 701247
rect 62948 701072 63000 701078
rect 62948 701014 63000 701020
rect 63144 700913 63172 712066
rect 654784 701208 654836 701214
rect 654784 701150 654836 701156
rect 63130 700904 63186 700913
rect 63130 700839 63186 700848
rect 651470 689480 651526 689489
rect 651470 689415 651526 689424
rect 651484 688702 651512 689415
rect 652760 688832 652812 688838
rect 651654 688800 651710 688809
rect 652760 688774 652812 688780
rect 651654 688735 651710 688744
rect 651472 688696 651524 688702
rect 651472 688638 651524 688644
rect 651470 687440 651526 687449
rect 651470 687375 651526 687384
rect 651484 687274 651512 687375
rect 651472 687268 651524 687274
rect 651472 687210 651524 687216
rect 651472 687064 651524 687070
rect 651472 687006 651524 687012
rect 651484 686769 651512 687006
rect 651470 686760 651526 686769
rect 651470 686695 651526 686704
rect 651668 686526 651696 688735
rect 62948 686520 63000 686526
rect 62948 686462 63000 686468
rect 651656 686520 651708 686526
rect 651656 686462 651708 686468
rect 62960 657665 62988 686462
rect 651472 685568 651524 685574
rect 651472 685510 651524 685516
rect 651484 685273 651512 685510
rect 651470 685264 651526 685273
rect 651470 685199 651526 685208
rect 652574 684448 652630 684457
rect 652772 684434 652800 688774
rect 654796 687070 654824 701150
rect 656440 690124 656492 690130
rect 656440 690066 656492 690072
rect 654784 687064 654836 687070
rect 654784 687006 654836 687012
rect 656452 685574 656480 690066
rect 657544 688696 657596 688702
rect 657544 688638 657596 688644
rect 656440 685568 656492 685574
rect 656440 685510 656492 685516
rect 652630 684406 652800 684434
rect 652574 684383 652630 684392
rect 62946 657656 63002 657665
rect 62946 657591 63002 657600
rect 653404 655580 653456 655586
rect 653404 655522 653456 655528
rect 651470 643240 651526 643249
rect 651470 643175 651526 643184
rect 651484 642394 651512 643175
rect 62948 642388 63000 642394
rect 62948 642330 63000 642336
rect 651472 642388 651524 642394
rect 651472 642330 651524 642336
rect 62960 612105 62988 642330
rect 652022 641880 652078 641889
rect 652022 641815 652078 641824
rect 651470 640792 651526 640801
rect 651470 640727 651526 640736
rect 651484 640354 651512 640727
rect 651472 640348 651524 640354
rect 651472 640290 651524 640296
rect 651380 640144 651432 640150
rect 651378 640112 651380 640121
rect 651432 640112 651434 640121
rect 651378 640047 651434 640056
rect 651656 638920 651708 638926
rect 651656 638862 651708 638868
rect 651472 638784 651524 638790
rect 651472 638726 651524 638732
rect 651484 638625 651512 638726
rect 651470 638616 651526 638625
rect 651470 638551 651526 638560
rect 651668 638217 651696 638862
rect 651654 638208 651710 638217
rect 651654 638143 651710 638152
rect 652036 634098 652064 641815
rect 653416 640150 653444 655522
rect 655520 645924 655572 645930
rect 655520 645866 655572 645872
rect 655336 643136 655388 643142
rect 655336 643078 655388 643084
rect 653404 640144 653456 640150
rect 653404 640086 653456 640092
rect 655348 638926 655376 643078
rect 655336 638920 655388 638926
rect 655336 638862 655388 638868
rect 655532 638790 655560 645866
rect 655520 638784 655572 638790
rect 655520 638726 655572 638732
rect 652024 634092 652076 634098
rect 652024 634034 652076 634040
rect 63132 625864 63184 625870
rect 63132 625806 63184 625812
rect 63144 618089 63172 625806
rect 657556 625190 657584 688638
rect 658936 669390 658964 731410
rect 660316 715018 660344 777582
rect 668584 733440 668636 733446
rect 668584 733382 668636 733388
rect 661684 730720 661736 730726
rect 661684 730662 661736 730668
rect 660304 715012 660356 715018
rect 660304 714954 660356 714960
rect 661696 670750 661724 730662
rect 667848 705220 667900 705226
rect 667848 705162 667900 705168
rect 667020 703860 667072 703866
rect 667020 703802 667072 703808
rect 661684 670744 661736 670750
rect 661684 670686 661736 670692
rect 658924 669384 658976 669390
rect 658924 669326 658976 669332
rect 658924 642388 658976 642394
rect 658924 642330 658976 642336
rect 657544 625184 657596 625190
rect 657544 625126 657596 625132
rect 63130 618080 63186 618089
rect 63130 618015 63186 618024
rect 62946 612096 63002 612105
rect 62946 612031 63002 612040
rect 64142 611416 64198 611425
rect 64142 611351 64198 611360
rect 653404 611380 653456 611386
rect 63314 595776 63370 595785
rect 63314 595711 63370 595720
rect 63130 594144 63186 594153
rect 63130 594079 63186 594088
rect 62946 590744 63002 590753
rect 62946 590679 63002 590688
rect 62960 287054 62988 590679
rect 63144 568585 63172 594079
rect 63328 571169 63356 595711
rect 63314 571160 63370 571169
rect 63314 571095 63370 571104
rect 63130 568576 63186 568585
rect 63130 568511 63186 568520
rect 63314 550216 63370 550225
rect 63314 550151 63370 550160
rect 63328 525745 63356 550151
rect 63314 525736 63370 525745
rect 63314 525671 63370 525680
rect 63314 381576 63370 381585
rect 63314 381511 63370 381520
rect 63328 354521 63356 381511
rect 63314 354512 63370 354521
rect 63314 354447 63370 354456
rect 63130 341456 63186 341465
rect 63130 341391 63186 341400
rect 63144 311817 63172 341391
rect 63406 332616 63462 332625
rect 63406 332551 63462 332560
rect 63130 311808 63186 311817
rect 63130 311743 63186 311752
rect 63130 298752 63186 298761
rect 63130 298687 63186 298696
rect 63144 289785 63172 298687
rect 63130 289776 63186 289785
rect 63130 289711 63186 289720
rect 62960 287026 63080 287054
rect 63052 282914 63080 287026
rect 63222 284608 63278 284617
rect 63222 284543 63278 284552
rect 63236 284374 63264 284543
rect 63224 284368 63276 284374
rect 63224 284310 63276 284316
rect 63052 282886 63356 282914
rect 62854 282160 62910 282169
rect 62854 282095 62910 282104
rect 62868 281586 62896 282095
rect 62856 281580 62908 281586
rect 62856 281522 62908 281528
rect 63130 280392 63186 280401
rect 63130 280327 63186 280336
rect 62946 278896 63002 278905
rect 62946 278831 63002 278840
rect 62960 273254 62988 278831
rect 62960 273226 63080 273254
rect 63052 229094 63080 273226
rect 62960 229066 63080 229094
rect 62670 224224 62726 224233
rect 62670 224159 62726 224168
rect 62960 223553 62988 229066
rect 63144 224505 63172 280327
rect 63328 278594 63356 282886
rect 63420 278746 63448 332551
rect 63420 278730 63540 278746
rect 63420 278724 63552 278730
rect 63420 278718 63500 278724
rect 63500 278666 63552 278672
rect 63316 278588 63368 278594
rect 63316 278530 63368 278536
rect 64156 264518 64184 611351
rect 653404 611322 653456 611328
rect 651470 597952 651526 597961
rect 651470 597887 651526 597896
rect 651484 597582 651512 597887
rect 651472 597576 651524 597582
rect 651472 597518 651524 597524
rect 651470 596728 651526 596737
rect 651470 596663 651526 596672
rect 651484 596222 651512 596663
rect 651472 596216 651524 596222
rect 651472 596158 651524 596164
rect 653416 595542 653444 611322
rect 657544 600364 657596 600370
rect 657544 600306 657596 600312
rect 654784 599004 654836 599010
rect 654784 598946 654836 598952
rect 651656 595536 651708 595542
rect 651656 595478 651708 595484
rect 653404 595536 653456 595542
rect 653404 595478 653456 595484
rect 651470 595368 651526 595377
rect 651470 595303 651526 595312
rect 651484 594862 651512 595303
rect 651668 595105 651696 595478
rect 651654 595096 651710 595105
rect 651654 595031 651710 595040
rect 651472 594856 651524 594862
rect 651472 594798 651524 594804
rect 651472 594720 651524 594726
rect 651472 594662 651524 594668
rect 651484 594153 651512 594662
rect 651470 594144 651526 594153
rect 651470 594079 651526 594088
rect 654796 593298 654824 598946
rect 657556 594726 657584 600306
rect 657544 594720 657596 594726
rect 657544 594662 657596 594668
rect 651472 593292 651524 593298
rect 651472 593234 651524 593240
rect 654784 593292 654836 593298
rect 654784 593234 654836 593240
rect 651484 592929 651512 593234
rect 651470 592920 651526 592929
rect 651470 592855 651526 592864
rect 658936 579698 658964 642330
rect 660304 634092 660356 634098
rect 660304 634034 660356 634040
rect 660316 581058 660344 634034
rect 664444 596216 664496 596222
rect 664444 596158 664496 596164
rect 661684 594856 661736 594862
rect 661684 594798 661736 594804
rect 660304 581052 660356 581058
rect 660304 580994 660356 581000
rect 658924 579692 658976 579698
rect 658924 579634 658976 579640
rect 653404 565888 653456 565894
rect 653404 565830 653456 565836
rect 651470 553480 651526 553489
rect 651470 553415 651526 553424
rect 651484 552702 651512 553415
rect 651472 552696 651524 552702
rect 651472 552638 651524 552644
rect 651654 552120 651710 552129
rect 651654 552055 651710 552064
rect 651470 551168 651526 551177
rect 651470 551103 651526 551112
rect 651484 550662 651512 551103
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 651380 550384 651432 550390
rect 651378 550352 651380 550361
rect 651432 550352 651434 550361
rect 651378 550287 651434 550296
rect 651668 549914 651696 552055
rect 653416 550390 653444 565830
rect 657820 554804 657872 554810
rect 657820 554746 657872 554752
rect 655152 553444 655204 553450
rect 655152 553386 655204 553392
rect 653404 550384 653456 550390
rect 653404 550326 653456 550332
rect 651656 549908 651708 549914
rect 651656 549850 651708 549856
rect 651470 549264 651526 549273
rect 651470 549199 651472 549208
rect 651524 549199 651526 549208
rect 651472 549170 651524 549176
rect 655164 548826 655192 553386
rect 657832 549234 657860 554746
rect 660304 550656 660356 550662
rect 660304 550598 660356 550604
rect 657820 549228 657872 549234
rect 657820 549170 657872 549176
rect 651472 548820 651524 548826
rect 651472 548762 651524 548768
rect 655152 548820 655204 548826
rect 655152 548762 655204 548768
rect 651484 548457 651512 548762
rect 651470 548448 651526 548457
rect 651470 548383 651526 548392
rect 658924 522028 658976 522034
rect 658924 521970 658976 521976
rect 658936 512922 658964 521970
rect 656164 512916 656216 512922
rect 656164 512858 656216 512864
rect 658924 512916 658976 512922
rect 658924 512858 658976 512864
rect 656176 499594 656204 512858
rect 650644 499588 650696 499594
rect 650644 499530 650696 499536
rect 656164 499588 656216 499594
rect 656164 499530 656216 499536
rect 64326 353424 64382 353433
rect 64326 353359 64382 353368
rect 64340 277914 64368 353359
rect 650656 278186 650684 499530
rect 660316 491366 660344 550598
rect 661696 534274 661724 594798
rect 663064 549908 663116 549914
rect 663064 549850 663116 549856
rect 661684 534268 661736 534274
rect 661684 534210 661736 534216
rect 662420 525088 662472 525094
rect 662420 525030 662472 525036
rect 662432 522034 662460 525030
rect 662420 522028 662472 522034
rect 662420 521970 662472 521976
rect 663076 491502 663104 549850
rect 664456 535498 664484 596158
rect 665088 564460 665140 564466
rect 665088 564402 665140 564408
rect 664444 535492 664496 535498
rect 664444 535434 664496 535440
rect 663064 491496 663116 491502
rect 663064 491438 663116 491444
rect 660304 491360 660356 491366
rect 660304 491302 660356 491308
rect 665100 485858 665128 564402
rect 665824 552696 665876 552702
rect 665824 552638 665876 552644
rect 665836 491638 665864 552638
rect 665824 491632 665876 491638
rect 665824 491574 665876 491580
rect 665088 485852 665140 485858
rect 665088 485794 665140 485800
rect 664444 474292 664496 474298
rect 664444 474234 664496 474240
rect 664456 467158 664484 474234
rect 652760 467152 652812 467158
rect 652760 467094 652812 467100
rect 664444 467152 664496 467158
rect 664444 467094 664496 467100
rect 652772 461378 652800 467094
rect 650828 461372 650880 461378
rect 650828 461314 650880 461320
rect 652760 461372 652812 461378
rect 652760 461314 652812 461320
rect 650840 278458 650868 461314
rect 667032 456618 667060 703802
rect 667662 698320 667718 698329
rect 667662 698255 667718 698264
rect 667204 686520 667256 686526
rect 667204 686462 667256 686468
rect 667216 626142 667244 686462
rect 667478 645824 667534 645833
rect 667478 645759 667534 645768
rect 667204 626136 667256 626142
rect 667204 626078 667256 626084
rect 667294 600944 667350 600953
rect 667294 600879 667350 600888
rect 667308 529990 667336 600879
rect 667492 574122 667520 645759
rect 667676 621042 667704 698255
rect 667664 621036 667716 621042
rect 667664 620978 667716 620984
rect 667664 608660 667716 608666
rect 667664 608602 667716 608608
rect 667480 574116 667532 574122
rect 667480 574058 667532 574064
rect 667676 532166 667704 608602
rect 667664 532160 667716 532166
rect 667664 532102 667716 532108
rect 667296 529984 667348 529990
rect 667296 529926 667348 529932
rect 667480 477556 667532 477562
rect 667480 477498 667532 477504
rect 667492 474298 667520 477498
rect 667480 474292 667532 474298
rect 667480 474234 667532 474240
rect 667020 456612 667072 456618
rect 667020 456554 667072 456560
rect 667860 456006 667888 705162
rect 668400 692844 668452 692850
rect 668400 692786 668452 692792
rect 668214 687848 668270 687857
rect 668214 687783 668270 687792
rect 668228 617506 668256 687783
rect 668412 619750 668440 692786
rect 668596 671158 668624 733382
rect 668858 730144 668914 730153
rect 668858 730079 668914 730088
rect 668584 671152 668636 671158
rect 668584 671094 668636 671100
rect 668872 660210 668900 730079
rect 669056 709374 669084 782478
rect 669044 709368 669096 709374
rect 669044 709310 669096 709316
rect 669240 708286 669268 784110
rect 670424 777028 670476 777034
rect 670424 776970 670476 776976
rect 669964 775600 670016 775606
rect 669964 775542 670016 775548
rect 669594 735720 669650 735729
rect 669594 735655 669650 735664
rect 669410 728784 669466 728793
rect 669410 728719 669466 728728
rect 669228 708280 669280 708286
rect 669228 708222 669280 708228
rect 669042 689480 669098 689489
rect 669042 689415 669098 689424
rect 668860 660204 668912 660210
rect 668860 660146 668912 660152
rect 668584 640348 668636 640354
rect 668584 640290 668636 640296
rect 668400 619744 668452 619750
rect 668400 619686 668452 619692
rect 668216 617500 668268 617506
rect 668216 617442 668268 617448
rect 668596 580038 668624 640290
rect 669056 616894 669084 689415
rect 669424 663950 669452 728719
rect 669608 665310 669636 735655
rect 669976 715766 670004 775542
rect 669964 715760 670016 715766
rect 669964 715702 670016 715708
rect 670436 705430 670464 776970
rect 670620 709238 670648 784246
rect 670896 728142 670924 886858
rect 670884 728136 670936 728142
rect 670884 728078 670936 728084
rect 671080 715358 671108 894406
rect 671896 894328 671948 894334
rect 671896 894270 671948 894276
rect 671436 773424 671488 773430
rect 671436 773366 671488 773372
rect 671250 733816 671306 733825
rect 671250 733751 671306 733760
rect 671068 715352 671120 715358
rect 671068 715294 671120 715300
rect 671068 712632 671120 712638
rect 671068 712574 671120 712580
rect 670608 709232 670660 709238
rect 670608 709174 670660 709180
rect 670424 705424 670476 705430
rect 670424 705366 670476 705372
rect 670882 695872 670938 695881
rect 670882 695807 670938 695816
rect 669964 687268 670016 687274
rect 669964 687210 670016 687216
rect 669778 685808 669834 685817
rect 669778 685743 669834 685752
rect 669596 665304 669648 665310
rect 669596 665246 669648 665252
rect 669412 663944 669464 663950
rect 669412 663886 669464 663892
rect 669228 661156 669280 661162
rect 669228 661098 669280 661104
rect 669044 616888 669096 616894
rect 669044 616830 669096 616836
rect 668766 594824 668822 594833
rect 668766 594759 668822 594768
rect 668584 580032 668636 580038
rect 668584 579974 668636 579980
rect 668582 562320 668638 562329
rect 668582 562255 668638 562264
rect 668596 484430 668624 562255
rect 668780 525094 668808 594759
rect 668950 593464 669006 593473
rect 668950 593399 669006 593408
rect 668964 529174 668992 593399
rect 668952 529168 669004 529174
rect 668952 529110 669004 529116
rect 668768 525088 668820 525094
rect 668768 525030 668820 525036
rect 668584 484424 668636 484430
rect 668584 484366 668636 484372
rect 667848 456000 667900 456006
rect 667848 455942 667900 455948
rect 669240 455666 669268 661098
rect 669594 644328 669650 644337
rect 669594 644263 669650 644272
rect 669412 623960 669464 623966
rect 669412 623902 669464 623908
rect 669424 579086 669452 623902
rect 669412 579080 669464 579086
rect 669412 579022 669464 579028
rect 669412 576972 669464 576978
rect 669412 576914 669464 576920
rect 669424 531622 669452 576914
rect 669608 572286 669636 644263
rect 669792 620294 669820 685743
rect 669976 625462 670004 687210
rect 670606 685536 670662 685545
rect 670606 685471 670662 685480
rect 670240 670268 670292 670274
rect 670240 670210 670292 670216
rect 669964 625456 670016 625462
rect 669964 625398 670016 625404
rect 670252 624510 670280 670210
rect 670240 624504 670292 624510
rect 670240 624446 670292 624452
rect 670240 623824 670292 623830
rect 670240 623766 670292 623772
rect 669780 620288 669832 620294
rect 669780 620230 669832 620236
rect 669964 597576 670016 597582
rect 669964 597518 670016 597524
rect 669596 572280 669648 572286
rect 669596 572222 669648 572228
rect 669780 568608 669832 568614
rect 669780 568550 669832 568556
rect 669412 531616 669464 531622
rect 669412 531558 669464 531564
rect 669228 455660 669280 455666
rect 669228 455602 669280 455608
rect 669792 455433 669820 568550
rect 669976 535838 670004 597518
rect 670252 579902 670280 623766
rect 670424 622464 670476 622470
rect 670424 622406 670476 622412
rect 670240 579896 670292 579902
rect 670240 579838 670292 579844
rect 670436 578202 670464 622406
rect 670620 615670 670648 685471
rect 670896 620838 670924 695807
rect 671080 668574 671108 712574
rect 671068 668568 671120 668574
rect 671068 668510 671120 668516
rect 671068 667956 671120 667962
rect 671068 667898 671120 667904
rect 671080 623286 671108 667898
rect 671264 661638 671292 733751
rect 671448 710054 671476 773366
rect 671908 746594 671936 894270
rect 672540 893036 672592 893042
rect 672540 892978 672592 892984
rect 672080 892900 672132 892906
rect 672080 892842 672132 892848
rect 671908 746566 672028 746594
rect 671804 742484 671856 742490
rect 671804 742426 671856 742432
rect 671620 741192 671672 741198
rect 671620 741134 671672 741140
rect 671436 710048 671488 710054
rect 671436 709990 671488 709996
rect 671436 668228 671488 668234
rect 671436 668170 671488 668176
rect 671252 661632 671304 661638
rect 671252 661574 671304 661580
rect 671448 654134 671476 668170
rect 671632 667214 671660 741134
rect 671816 736934 671844 742426
rect 672000 736934 672028 746566
rect 671724 736906 671844 736934
rect 671908 736906 672028 736934
rect 671724 692774 671752 736906
rect 671908 714542 671936 736906
rect 671896 714536 671948 714542
rect 671896 714478 671948 714484
rect 672092 713454 672120 892842
rect 672264 739152 672316 739158
rect 672264 739094 672316 739100
rect 672080 713448 672132 713454
rect 672080 713390 672132 713396
rect 671986 713280 672042 713289
rect 671986 713215 672042 713224
rect 672000 712638 672028 713215
rect 671988 712632 672040 712638
rect 671988 712574 672040 712580
rect 671986 712464 672042 712473
rect 671986 712399 672042 712408
rect 671724 692746 671844 692774
rect 671620 667208 671672 667214
rect 671620 667150 671672 667156
rect 671816 667026 671844 692746
rect 671724 666998 671844 667026
rect 671724 664426 671752 666998
rect 672000 666942 672028 712399
rect 671988 666936 672040 666942
rect 671988 666878 672040 666884
rect 671896 666596 671948 666602
rect 671896 666538 671948 666544
rect 671712 664420 671764 664426
rect 671712 664362 671764 664368
rect 671908 654134 671936 666538
rect 672276 664057 672304 739094
rect 672552 713697 672580 892978
rect 672736 866658 672764 895630
rect 675850 895520 675906 895529
rect 675850 895455 675906 895464
rect 675864 894470 675892 895455
rect 676034 894704 676090 894713
rect 676034 894639 676090 894648
rect 675852 894464 675904 894470
rect 675852 894406 675904 894412
rect 676048 894334 676076 894639
rect 676036 894328 676088 894334
rect 676036 894270 676088 894276
rect 675850 893888 675906 893897
rect 675850 893823 675906 893832
rect 675864 893042 675892 893823
rect 676034 893072 676090 893081
rect 675852 893036 675904 893042
rect 676034 893007 676090 893016
rect 675852 892978 675904 892984
rect 676048 892906 676076 893007
rect 676036 892900 676088 892906
rect 676036 892842 676088 892848
rect 676034 892664 676090 892673
rect 676090 892622 676444 892650
rect 676034 892599 676090 892608
rect 676034 891440 676090 891449
rect 676034 891375 676090 891384
rect 675298 891032 675354 891041
rect 675298 890967 675354 890976
rect 674840 890384 674892 890390
rect 674840 890326 674892 890332
rect 674380 888956 674432 888962
rect 674380 888898 674432 888904
rect 674196 887324 674248 887330
rect 674196 887266 674248 887272
rect 673092 885692 673144 885698
rect 673092 885634 673144 885640
rect 672724 866652 672776 866658
rect 672724 866594 672776 866600
rect 672724 775668 672776 775674
rect 672724 775610 672776 775616
rect 672736 717614 672764 775610
rect 672908 732760 672960 732766
rect 672908 732702 672960 732708
rect 672920 724514 672948 732702
rect 673104 728346 673132 885634
rect 674208 868766 674236 887266
rect 674392 869530 674420 888898
rect 674656 888548 674708 888554
rect 674656 888490 674708 888496
rect 674668 872174 674696 888490
rect 674852 874721 674880 890326
rect 675024 879640 675076 879646
rect 674944 879588 675024 879594
rect 674944 879582 675076 879588
rect 674944 879566 675064 879582
rect 674944 876194 674972 879566
rect 675116 879436 675168 879442
rect 675116 879378 675168 879384
rect 675128 879074 675156 879378
rect 675312 879074 675340 890967
rect 676048 890390 676076 891375
rect 676036 890384 676088 890390
rect 676036 890326 676088 890332
rect 676034 890216 676090 890225
rect 676090 890186 676260 890202
rect 676090 890180 676272 890186
rect 676090 890174 676220 890180
rect 676034 890151 676090 890160
rect 676220 890122 676272 890128
rect 676034 889400 676090 889409
rect 676090 889358 676260 889386
rect 676034 889335 676090 889344
rect 676034 888992 676090 889001
rect 676034 888927 676036 888936
rect 676088 888927 676090 888936
rect 676036 888898 676088 888904
rect 676232 888758 676260 889358
rect 676220 888752 676272 888758
rect 676220 888694 676272 888700
rect 676034 888584 676090 888593
rect 676034 888519 676036 888528
rect 676088 888519 676090 888528
rect 676036 888490 676088 888496
rect 676034 887360 676090 887369
rect 676034 887295 676036 887304
rect 676088 887295 676090 887304
rect 676036 887266 676088 887272
rect 676034 886952 676090 886961
rect 676034 886887 676036 886896
rect 676088 886887 676090 886896
rect 676036 886858 676088 886864
rect 676416 886718 676444 892622
rect 679622 891848 679678 891857
rect 679622 891783 679678 891792
rect 676864 890180 676916 890186
rect 676864 890122 676916 890128
rect 675852 886712 675904 886718
rect 675852 886654 675904 886660
rect 676404 886712 676456 886718
rect 676404 886654 676456 886660
rect 675484 880524 675536 880530
rect 675484 880466 675536 880472
rect 675036 879046 675156 879074
rect 675220 879046 675340 879074
rect 675036 877010 675064 879046
rect 675220 877169 675248 879046
rect 675496 878084 675524 880466
rect 675668 879300 675720 879306
rect 675668 879242 675720 879248
rect 675680 878529 675708 879242
rect 675666 878520 675722 878529
rect 675864 878490 675892 886654
rect 676034 885728 676090 885737
rect 676034 885663 676036 885672
rect 676088 885663 676090 885672
rect 676036 885634 676088 885640
rect 676036 880252 676088 880258
rect 676036 880194 676088 880200
rect 676048 878490 676076 880194
rect 676876 879442 676904 890122
rect 678242 889808 678298 889817
rect 678242 889743 678298 889752
rect 677048 888752 677100 888758
rect 677048 888694 677100 888700
rect 677060 879646 677088 888694
rect 677048 879640 677100 879646
rect 677048 879582 677100 879588
rect 676864 879436 676916 879442
rect 676864 879378 676916 879384
rect 678256 879306 678284 889743
rect 679636 880258 679664 891783
rect 681002 890624 681058 890633
rect 681002 890559 681058 890568
rect 681016 880705 681044 890559
rect 683118 888176 683174 888185
rect 683118 888111 683174 888120
rect 681002 880696 681058 880705
rect 681002 880631 681058 880640
rect 683132 880433 683160 888111
rect 683118 880424 683174 880433
rect 683118 880359 683174 880368
rect 679624 880252 679676 880258
rect 679624 880194 679676 880200
rect 678244 879300 678296 879306
rect 678244 879242 678296 879248
rect 675666 878455 675722 878464
rect 675852 878484 675904 878490
rect 675852 878426 675904 878432
rect 676036 878484 676088 878490
rect 676036 878426 676088 878432
rect 675484 877804 675536 877810
rect 675484 877746 675536 877752
rect 675496 877540 675524 877746
rect 675206 877160 675262 877169
rect 675206 877095 675262 877104
rect 675036 876982 675432 877010
rect 675404 876860 675432 876982
rect 675392 876784 675444 876790
rect 675392 876726 675444 876732
rect 675404 876248 675432 876726
rect 674944 876166 675064 876194
rect 674838 874712 674894 874721
rect 674838 874647 674894 874656
rect 675036 873202 675064 876166
rect 675482 874712 675538 874721
rect 675482 874647 675538 874656
rect 675496 874412 675524 874647
rect 675574 874168 675630 874177
rect 675574 874103 675630 874112
rect 675588 873868 675616 874103
rect 675036 873174 675418 873202
rect 675758 873080 675814 873089
rect 675758 873015 675814 873024
rect 675022 872808 675078 872817
rect 675022 872743 675078 872752
rect 674668 872146 674880 872174
rect 674392 869502 674696 869530
rect 674668 869122 674696 869502
rect 674852 869310 674880 872146
rect 675036 869530 675064 872743
rect 675772 872576 675800 873015
rect 675390 870496 675446 870505
rect 675390 870431 675446 870440
rect 675404 870060 675432 870431
rect 675036 869502 675418 869530
rect 675024 869440 675076 869446
rect 675024 869382 675076 869388
rect 674840 869304 674892 869310
rect 674840 869246 674892 869252
rect 674668 869094 674880 869122
rect 674196 868760 674248 868766
rect 674196 868702 674248 868708
rect 674852 867610 674880 869094
rect 675036 868170 675064 869382
rect 675300 869304 675352 869310
rect 675300 869246 675352 869252
rect 675312 868889 675340 869246
rect 675312 868861 675418 868889
rect 675300 868760 675352 868766
rect 675300 868702 675352 868708
rect 675312 868238 675340 868702
rect 675312 868210 675418 868238
rect 675036 868142 675248 868170
rect 675024 868080 675076 868086
rect 675024 868022 675076 868028
rect 674840 867604 674892 867610
rect 674840 867546 674892 867552
rect 675036 865858 675064 868022
rect 675220 867694 675248 868142
rect 675220 867666 675418 867694
rect 675208 867604 675260 867610
rect 675208 867546 675260 867552
rect 675220 867049 675248 867546
rect 675220 867021 675418 867049
rect 675036 865830 675418 865858
rect 675298 865736 675354 865745
rect 675298 865671 675354 865680
rect 675312 863818 675340 865671
rect 675758 865464 675814 865473
rect 675758 865399 675814 865408
rect 675772 865195 675800 865399
rect 675666 865056 675722 865065
rect 675666 864991 675722 865000
rect 675680 864552 675708 864991
rect 675312 863790 675432 863818
rect 675404 863328 675432 863790
rect 675392 790832 675444 790838
rect 675392 790774 675444 790780
rect 675404 788868 675432 790774
rect 675772 788089 675800 788324
rect 675758 788080 675814 788089
rect 675758 788015 675814 788024
rect 675128 787665 675418 787693
rect 675128 786729 675156 787665
rect 675404 786729 675432 787032
rect 675114 786720 675170 786729
rect 675114 786655 675170 786664
rect 675390 786720 675446 786729
rect 675390 786655 675446 786664
rect 674852 785182 675418 785210
rect 673736 782672 673788 782678
rect 673736 782614 673788 782620
rect 673274 777472 673330 777481
rect 673274 777407 673330 777416
rect 673092 728340 673144 728346
rect 673092 728282 673144 728288
rect 672920 724486 673040 724514
rect 672644 717586 672764 717614
rect 672644 714490 672672 717586
rect 672816 717528 672868 717534
rect 672816 717470 672868 717476
rect 672644 714462 672764 714490
rect 672538 713688 672594 713697
rect 672538 713623 672594 713632
rect 672736 713538 672764 714462
rect 672460 713510 672764 713538
rect 672460 712094 672488 713510
rect 672632 713312 672684 713318
rect 672632 713254 672684 713260
rect 672448 712088 672500 712094
rect 672448 712030 672500 712036
rect 672448 711816 672500 711822
rect 672448 711758 672500 711764
rect 672460 670041 672488 711758
rect 672446 670032 672502 670041
rect 672446 669967 672502 669976
rect 672644 669497 672672 713254
rect 672828 708393 672856 717470
rect 673012 715850 673040 724486
rect 673288 717534 673316 777407
rect 673552 738744 673604 738750
rect 673552 738686 673604 738692
rect 673564 736934 673592 738686
rect 673564 736906 673684 736934
rect 673458 734360 673514 734369
rect 673458 734295 673514 734304
rect 673472 732850 673500 734295
rect 673472 732822 673592 732850
rect 673564 727274 673592 732822
rect 673472 727246 673592 727274
rect 673276 717528 673328 717534
rect 673276 717470 673328 717476
rect 673274 716544 673330 716553
rect 673274 716479 673330 716488
rect 673288 716310 673316 716479
rect 673276 716304 673328 716310
rect 673276 716246 673328 716252
rect 673274 716136 673330 716145
rect 673274 716071 673330 716080
rect 672920 715822 673040 715850
rect 672920 708642 672948 715822
rect 673092 715760 673144 715766
rect 673090 715728 673092 715737
rect 673144 715728 673146 715737
rect 673090 715663 673146 715672
rect 673092 715352 673144 715358
rect 673090 715320 673092 715329
rect 673144 715320 673146 715329
rect 673090 715255 673146 715264
rect 673090 715048 673146 715057
rect 673288 715018 673316 716071
rect 673090 714983 673146 714992
rect 673276 715012 673328 715018
rect 673104 711822 673132 714983
rect 673276 714954 673328 714960
rect 673276 714536 673328 714542
rect 673274 714504 673276 714513
rect 673328 714504 673330 714513
rect 673274 714439 673330 714448
rect 673274 714096 673330 714105
rect 673274 714031 673330 714040
rect 673288 713590 673316 714031
rect 673276 713584 673328 713590
rect 673276 713526 673328 713532
rect 673276 713448 673328 713454
rect 673276 713390 673328 713396
rect 673288 712881 673316 713390
rect 673274 712872 673330 712881
rect 673274 712807 673330 712816
rect 673276 712088 673328 712094
rect 673276 712030 673328 712036
rect 673092 711816 673144 711822
rect 673092 711758 673144 711764
rect 673288 711657 673316 712030
rect 673274 711648 673330 711657
rect 673274 711583 673330 711592
rect 673274 710424 673330 710433
rect 673274 710359 673330 710368
rect 673092 710048 673144 710054
rect 673090 710016 673092 710025
rect 673144 710016 673146 710025
rect 673090 709951 673146 709960
rect 673288 709374 673316 710359
rect 673276 709368 673328 709374
rect 673276 709310 673328 709316
rect 673276 709232 673328 709238
rect 673274 709200 673276 709209
rect 673328 709200 673330 709209
rect 673274 709135 673330 709144
rect 673274 708792 673330 708801
rect 673274 708727 673330 708736
rect 672920 708614 673040 708642
rect 672814 708384 672870 708393
rect 672814 708319 672870 708328
rect 673012 705194 673040 708614
rect 673288 708286 673316 708727
rect 673276 708280 673328 708286
rect 673276 708222 673328 708228
rect 673276 705424 673328 705430
rect 673274 705392 673276 705401
rect 673328 705392 673330 705401
rect 673274 705327 673330 705336
rect 672920 705166 673040 705194
rect 672630 669488 672686 669497
rect 672630 669423 672686 669432
rect 672262 664048 672318 664057
rect 672262 663983 672318 663992
rect 672920 662969 672948 705166
rect 673274 696960 673330 696969
rect 673274 696895 673330 696904
rect 673090 686216 673146 686225
rect 673090 686151 673146 686160
rect 673104 683114 673132 686151
rect 673104 683086 673224 683114
rect 672906 662960 672962 662969
rect 672906 662895 672962 662904
rect 672172 659728 672224 659734
rect 672172 659670 672224 659676
rect 671448 654106 671568 654134
rect 671252 645924 671304 645930
rect 671252 645866 671304 645872
rect 671264 645561 671292 645866
rect 671250 645552 671306 645561
rect 671250 645487 671306 645496
rect 671252 643136 671304 643142
rect 671252 643078 671304 643084
rect 671264 641481 671292 643078
rect 671250 641472 671306 641481
rect 671250 641407 671306 641416
rect 671540 640334 671568 654106
rect 671724 654106 671936 654134
rect 672184 654134 672212 659670
rect 672184 654106 672304 654134
rect 671724 649994 671752 654106
rect 671986 652488 672042 652497
rect 671986 652423 672042 652432
rect 671724 649966 671936 649994
rect 671710 647864 671766 647873
rect 671710 647799 671766 647808
rect 671540 640306 671660 640334
rect 671342 638616 671398 638625
rect 671342 638551 671398 638560
rect 671356 632942 671384 638551
rect 671632 633026 671660 640306
rect 671540 633010 671660 633026
rect 671528 633004 671660 633010
rect 671580 632998 671660 633004
rect 671528 632946 671580 632952
rect 671344 632936 671396 632942
rect 671344 632878 671396 632884
rect 671344 632800 671396 632806
rect 671344 632742 671396 632748
rect 671356 627994 671384 632742
rect 671528 632664 671580 632670
rect 671528 632606 671580 632612
rect 671356 627966 671476 627994
rect 671448 624209 671476 627966
rect 671540 627914 671568 632606
rect 671540 627886 671660 627914
rect 671434 624200 671490 624209
rect 671434 624135 671490 624144
rect 671068 623280 671120 623286
rect 671068 623222 671120 623228
rect 671436 621172 671488 621178
rect 671436 621114 671488 621120
rect 670884 620832 670936 620838
rect 670884 620774 670936 620780
rect 670608 615664 670660 615670
rect 670608 615606 670660 615612
rect 670608 614916 670660 614922
rect 670608 614858 670660 614864
rect 670424 578196 670476 578202
rect 670424 578138 670476 578144
rect 670240 577788 670292 577794
rect 670240 577730 670292 577736
rect 669964 535832 670016 535838
rect 669964 535774 670016 535780
rect 670252 532914 670280 577730
rect 670424 553444 670476 553450
rect 670424 553386 670476 553392
rect 670436 551585 670464 553386
rect 670422 551576 670478 551585
rect 670422 551511 670478 551520
rect 670422 549672 670478 549681
rect 670422 549607 670478 549616
rect 670240 532908 670292 532914
rect 670240 532850 670292 532856
rect 670436 480418 670464 549607
rect 670424 480412 670476 480418
rect 670424 480354 670476 480360
rect 670436 477562 670464 480354
rect 670424 477556 670476 477562
rect 670424 477498 670476 477504
rect 669778 455424 669834 455433
rect 669778 455359 669834 455368
rect 670620 455161 670648 614858
rect 670974 607744 671030 607753
rect 670974 607679 671030 607688
rect 670792 579420 670844 579426
rect 670792 579362 670844 579368
rect 670804 535022 670832 579362
rect 670792 535016 670844 535022
rect 670792 534958 670844 534964
rect 670792 534404 670844 534410
rect 670792 534346 670844 534352
rect 670804 490958 670832 534346
rect 670988 528970 671016 607679
rect 671160 578604 671212 578610
rect 671160 578546 671212 578552
rect 671172 534138 671200 578546
rect 671448 577454 671476 621114
rect 671436 577448 671488 577454
rect 671436 577390 671488 577396
rect 671632 574598 671660 627886
rect 671724 611354 671752 647799
rect 671908 622674 671936 649966
rect 672000 622826 672028 652423
rect 672276 640334 672304 654106
rect 672814 649224 672870 649233
rect 672814 649159 672870 649168
rect 672184 640306 672304 640334
rect 672000 622798 672120 622826
rect 671896 622668 671948 622674
rect 671896 622610 671948 622616
rect 672092 622418 672120 622798
rect 672000 622390 672120 622418
rect 671724 611326 671844 611354
rect 671620 574592 671672 574598
rect 671620 574534 671672 574540
rect 671816 571606 671844 611326
rect 672000 574326 672028 622390
rect 671988 574320 672040 574326
rect 671988 574262 672040 574268
rect 671804 571600 671856 571606
rect 671804 571542 671856 571548
rect 671344 570444 671396 570450
rect 671344 570386 671396 570392
rect 671160 534132 671212 534138
rect 671160 534074 671212 534080
rect 671160 531480 671212 531486
rect 671160 531422 671212 531428
rect 670976 528964 671028 528970
rect 670976 528906 671028 528912
rect 670792 490952 670844 490958
rect 670792 490894 670844 490900
rect 671172 488510 671200 531422
rect 671160 488504 671212 488510
rect 671160 488446 671212 488452
rect 670606 455152 670662 455161
rect 670606 455087 670662 455096
rect 657542 403336 657598 403345
rect 657542 403271 657598 403280
rect 652022 400888 652078 400897
rect 652022 400823 652078 400832
rect 651472 373992 651524 373998
rect 651472 373934 651524 373940
rect 651484 373289 651512 373934
rect 651470 373280 651526 373289
rect 651470 373215 651526 373224
rect 652036 372201 652064 400823
rect 652206 396672 652262 396681
rect 652206 396607 652262 396616
rect 652220 373969 652248 396607
rect 654782 382936 654838 382945
rect 654782 382871 654838 382880
rect 652206 373960 652262 373969
rect 652206 373895 652262 373904
rect 652022 372192 652078 372201
rect 652022 372127 652078 372136
rect 654796 371006 654824 382871
rect 657556 373998 657584 403271
rect 670514 392592 670570 392601
rect 670514 392527 670570 392536
rect 657544 373992 657596 373998
rect 657544 373934 657596 373940
rect 651472 371000 651524 371006
rect 651472 370942 651524 370948
rect 654784 371000 654836 371006
rect 654784 370942 654836 370948
rect 651484 370705 651512 370942
rect 651470 370696 651526 370705
rect 651470 370631 651526 370640
rect 655518 366344 655574 366353
rect 655518 366279 655574 366288
rect 655532 362982 655560 366279
rect 651012 362976 651064 362982
rect 651012 362918 651064 362924
rect 655520 362976 655572 362982
rect 655520 362918 655572 362924
rect 650828 278452 650880 278458
rect 650828 278394 650880 278400
rect 651024 278322 651052 362918
rect 654782 358592 654838 358601
rect 654782 358527 654838 358536
rect 652022 356688 652078 356697
rect 652022 356623 652078 356632
rect 651380 328296 651432 328302
rect 651380 328238 651432 328244
rect 651392 328137 651420 328238
rect 651378 328128 651434 328137
rect 651378 328063 651434 328072
rect 652036 326913 652064 356623
rect 652390 351112 652446 351121
rect 652390 351047 652446 351056
rect 652404 329769 652432 351047
rect 653402 338736 653458 338745
rect 653402 338671 653458 338680
rect 652390 329760 652446 329769
rect 652390 329695 652446 329704
rect 652022 326904 652078 326913
rect 652022 326839 652078 326848
rect 651378 325680 651434 325689
rect 653416 325650 653444 338671
rect 654796 328302 654824 358527
rect 669410 347304 669466 347313
rect 669410 347239 669466 347248
rect 654784 328296 654836 328302
rect 654784 328238 654836 328244
rect 651378 325615 651380 325624
rect 651432 325615 651434 325624
rect 653404 325644 653456 325650
rect 651380 325586 651432 325592
rect 653404 325586 653456 325592
rect 653402 313304 653458 313313
rect 653402 313239 653458 313248
rect 652298 309904 652354 309913
rect 652298 309839 652354 309848
rect 651380 303544 651432 303550
rect 651380 303486 651432 303492
rect 651392 303385 651420 303486
rect 651378 303376 651434 303385
rect 651378 303311 651434 303320
rect 652312 302161 652340 309839
rect 653416 303550 653444 313239
rect 658922 311944 658978 311953
rect 658922 311879 658978 311888
rect 653404 303544 653456 303550
rect 653404 303486 653456 303492
rect 652298 302152 652354 302161
rect 652298 302087 652354 302096
rect 658936 300830 658964 311879
rect 651472 300824 651524 300830
rect 651472 300766 651524 300772
rect 658924 300824 658976 300830
rect 658924 300766 658976 300772
rect 651484 300665 651512 300766
rect 651470 300656 651526 300665
rect 651470 300591 651526 300600
rect 651470 298752 651526 298761
rect 651470 298687 651526 298696
rect 651484 298178 651512 298687
rect 651472 298172 651524 298178
rect 651472 298114 651524 298120
rect 660580 298172 660632 298178
rect 660580 298114 660632 298120
rect 652390 297528 652446 297537
rect 652390 297463 652446 297472
rect 652206 296848 652262 296857
rect 652206 296783 652208 296792
rect 652260 296783 652262 296792
rect 652208 296754 652260 296760
rect 652404 296714 652432 297463
rect 652312 296686 652432 296714
rect 658924 296744 658976 296750
rect 658924 296686 658976 296692
rect 651654 295352 651710 295361
rect 651654 295287 651710 295296
rect 651470 294264 651526 294273
rect 651470 294199 651526 294208
rect 651484 294030 651512 294199
rect 651472 294024 651524 294030
rect 651472 293966 651524 293972
rect 651470 293040 651526 293049
rect 651470 292975 651526 292984
rect 651484 292602 651512 292975
rect 651472 292596 651524 292602
rect 651472 292538 651524 292544
rect 651668 291825 651696 295287
rect 651654 291816 651710 291825
rect 651654 291751 651710 291760
rect 652114 291544 652170 291553
rect 652114 291479 652170 291488
rect 651470 290456 651526 290465
rect 651470 290391 651526 290400
rect 651484 289882 651512 290391
rect 651472 289876 651524 289882
rect 651472 289818 651524 289824
rect 651654 289232 651710 289241
rect 651654 289167 651710 289176
rect 651470 288688 651526 288697
rect 651470 288623 651526 288632
rect 651484 288454 651512 288623
rect 651472 288448 651524 288454
rect 651472 288390 651524 288396
rect 651668 287745 651696 289167
rect 651654 287736 651710 287745
rect 651654 287671 651710 287680
rect 651470 287464 651526 287473
rect 651470 287399 651526 287408
rect 651484 287094 651512 287399
rect 651472 287088 651524 287094
rect 651472 287030 651524 287036
rect 652128 287054 652156 291479
rect 652312 287054 652340 296686
rect 652128 287026 652248 287054
rect 652312 287026 652616 287054
rect 651470 285968 651526 285977
rect 651470 285903 651526 285912
rect 651484 285734 651512 285903
rect 651472 285728 651524 285734
rect 651472 285670 651524 285676
rect 651470 284744 651526 284753
rect 651470 284679 651526 284688
rect 651484 284374 651512 284679
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 651470 283384 651526 283393
rect 651470 283319 651526 283328
rect 651484 282946 651512 283319
rect 651472 282940 651524 282946
rect 651472 282882 651524 282888
rect 652022 282160 652078 282169
rect 652022 282095 652078 282104
rect 651470 280936 651526 280945
rect 651470 280871 651526 280880
rect 651484 280226 651512 280871
rect 651472 280220 651524 280226
rect 651472 280162 651524 280168
rect 651012 278316 651064 278322
rect 651012 278258 651064 278264
rect 629944 278180 629996 278186
rect 629944 278122 629996 278128
rect 630128 278180 630180 278186
rect 630128 278122 630180 278128
rect 650644 278180 650696 278186
rect 650644 278122 650696 278128
rect 64328 277908 64380 277914
rect 64328 277850 64380 277856
rect 65904 272542 65932 278052
rect 67100 274242 67128 278052
rect 67088 274236 67140 274242
rect 67088 274178 67140 274184
rect 65892 272536 65944 272542
rect 65892 272478 65944 272484
rect 68204 271182 68232 278052
rect 69400 273970 69428 278052
rect 69388 273964 69440 273970
rect 69388 273906 69440 273912
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 70596 269822 70624 278052
rect 71792 275058 71820 278052
rect 71780 275052 71832 275058
rect 71780 274994 71832 275000
rect 72988 272678 73016 278052
rect 74184 274718 74212 278052
rect 74172 274712 74224 274718
rect 74172 274654 74224 274660
rect 72976 272672 73028 272678
rect 72976 272614 73028 272620
rect 75380 271454 75408 278052
rect 76484 275602 76512 278052
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 76840 274712 76892 274718
rect 76840 274654 76892 274660
rect 75368 271448 75420 271454
rect 75368 271390 75420 271396
rect 76852 271318 76880 274654
rect 77680 274106 77708 278052
rect 77668 274100 77720 274106
rect 77668 274042 77720 274048
rect 76840 271312 76892 271318
rect 76840 271254 76892 271260
rect 78876 270502 78904 278052
rect 78864 270496 78916 270502
rect 78864 270438 78916 270444
rect 80072 269822 80100 278052
rect 81268 275466 81296 278052
rect 81256 275460 81308 275466
rect 81256 275402 81308 275408
rect 82464 272814 82492 278052
rect 83674 278038 84148 278066
rect 84778 278038 85528 278066
rect 82452 272808 82504 272814
rect 82452 272750 82504 272756
rect 84120 270366 84148 278038
rect 84108 270360 84160 270366
rect 84108 270302 84160 270308
rect 85500 269958 85528 278038
rect 85960 274718 85988 278052
rect 86224 275596 86276 275602
rect 86224 275538 86276 275544
rect 85948 274712 86000 274718
rect 85948 274654 86000 274660
rect 85488 269952 85540 269958
rect 85488 269894 85540 269900
rect 70584 269816 70636 269822
rect 70584 269758 70636 269764
rect 79324 269816 79376 269822
rect 79324 269758 79376 269764
rect 80060 269816 80112 269822
rect 80060 269758 80112 269764
rect 79336 267034 79364 269758
rect 86236 267442 86264 275538
rect 87156 271590 87184 278052
rect 88352 273834 88380 278052
rect 89562 278038 89668 278066
rect 88340 273828 88392 273834
rect 88340 273770 88392 273776
rect 87144 271584 87196 271590
rect 87144 271526 87196 271532
rect 89640 270094 89668 278038
rect 90744 275602 90772 278052
rect 91862 278038 92428 278066
rect 90732 275596 90784 275602
rect 90732 275538 90784 275544
rect 90364 274712 90416 274718
rect 90364 274654 90416 274660
rect 89628 270088 89680 270094
rect 89628 270030 89680 270036
rect 86224 267436 86276 267442
rect 86224 267378 86276 267384
rect 90376 267170 90404 274654
rect 92400 268394 92428 278038
rect 93044 275194 93072 278052
rect 93032 275188 93084 275194
rect 93032 275130 93084 275136
rect 94240 272950 94268 278052
rect 95436 274378 95464 278052
rect 96632 275330 96660 278052
rect 96620 275324 96672 275330
rect 96620 275266 96672 275272
rect 95424 274372 95476 274378
rect 95424 274314 95476 274320
rect 94228 272944 94280 272950
rect 94228 272886 94280 272892
rect 97828 271726 97856 278052
rect 99038 278038 99328 278066
rect 97816 271720 97868 271726
rect 97816 271662 97868 271668
rect 99300 268530 99328 278038
rect 100128 275738 100156 278052
rect 100116 275732 100168 275738
rect 100116 275674 100168 275680
rect 101324 274514 101352 278052
rect 101312 274508 101364 274514
rect 101312 274450 101364 274456
rect 102520 273086 102548 278052
rect 103716 274718 103744 278052
rect 104912 277394 104940 278052
rect 104912 277366 105032 277394
rect 103704 274712 103756 274718
rect 103704 274654 103756 274660
rect 104808 274712 104860 274718
rect 104808 274654 104860 274660
rect 102508 273080 102560 273086
rect 102508 273022 102560 273028
rect 99288 268524 99340 268530
rect 99288 268466 99340 268472
rect 92388 268388 92440 268394
rect 92388 268330 92440 268336
rect 104820 267306 104848 274654
rect 105004 268666 105032 277366
rect 106016 271862 106044 278052
rect 107212 276010 107240 278052
rect 107200 276004 107252 276010
rect 107200 275946 107252 275952
rect 108408 273222 108436 278052
rect 109618 278038 110368 278066
rect 108396 273216 108448 273222
rect 108396 273158 108448 273164
rect 106004 271856 106056 271862
rect 106004 271798 106056 271804
rect 110340 268802 110368 278038
rect 110800 274718 110828 278052
rect 110788 274712 110840 274718
rect 110788 274654 110840 274660
rect 111708 274712 111760 274718
rect 111708 274654 111760 274660
rect 110328 268796 110380 268802
rect 110328 268738 110380 268744
rect 104992 268660 105044 268666
rect 104992 268602 105044 268608
rect 111720 267578 111748 274654
rect 111996 270230 112024 278052
rect 113206 278038 113496 278066
rect 113468 271046 113496 278038
rect 114388 274650 114416 278052
rect 115506 278038 115796 278066
rect 114376 274644 114428 274650
rect 114376 274586 114428 274592
rect 113456 271040 113508 271046
rect 113456 270982 113508 270988
rect 111984 270224 112036 270230
rect 111984 270166 112036 270172
rect 115768 268938 115796 278038
rect 116688 272406 116716 278052
rect 117898 278038 118648 278066
rect 116676 272400 116728 272406
rect 116676 272342 116728 272348
rect 118620 269074 118648 278038
rect 119080 273698 119108 278052
rect 120276 273834 120304 278052
rect 119344 273828 119396 273834
rect 119344 273770 119396 273776
rect 120264 273828 120316 273834
rect 120264 273770 120316 273776
rect 119068 273692 119120 273698
rect 119068 273634 119120 273640
rect 118608 269068 118660 269074
rect 118608 269010 118660 269016
rect 115756 268932 115808 268938
rect 115756 268874 115808 268880
rect 119356 267714 119384 273770
rect 121472 270638 121500 278052
rect 122590 278038 122788 278066
rect 121460 270632 121512 270638
rect 121460 270574 121512 270580
rect 122760 269686 122788 278038
rect 123772 270910 123800 278052
rect 124968 271998 124996 278052
rect 126178 278038 126928 278066
rect 124956 271992 125008 271998
rect 124956 271934 125008 271940
rect 123760 270904 123812 270910
rect 123760 270846 123812 270852
rect 122748 269680 122800 269686
rect 122748 269622 122800 269628
rect 126900 269414 126928 278038
rect 127360 272270 127388 278052
rect 128556 274786 128584 278052
rect 128544 274780 128596 274786
rect 128544 274722 128596 274728
rect 127348 272264 127400 272270
rect 127348 272206 127400 272212
rect 129660 269550 129688 278052
rect 130856 274242 130884 278052
rect 130384 274236 130436 274242
rect 130384 274178 130436 274184
rect 130844 274236 130896 274242
rect 130844 274178 130896 274184
rect 129648 269544 129700 269550
rect 129648 269486 129700 269492
rect 126888 269408 126940 269414
rect 126888 269350 126940 269356
rect 119344 267708 119396 267714
rect 119344 267650 119396 267656
rect 111708 267572 111760 267578
rect 111708 267514 111760 267520
rect 104808 267300 104860 267306
rect 104808 267242 104860 267248
rect 90364 267164 90416 267170
rect 90364 267106 90416 267112
rect 79324 267028 79376 267034
rect 79324 266970 79376 266976
rect 130396 266626 130424 274178
rect 132052 273562 132080 278052
rect 133262 278038 133828 278066
rect 132040 273556 132092 273562
rect 132040 273498 132092 273504
rect 133800 270502 133828 278038
rect 134444 270774 134472 278052
rect 134432 270768 134484 270774
rect 134432 270710 134484 270716
rect 132500 270496 132552 270502
rect 132500 270438 132552 270444
rect 133788 270496 133840 270502
rect 133788 270438 133840 270444
rect 130384 266620 130436 266626
rect 130384 266562 130436 266568
rect 132512 266490 132540 270438
rect 135640 268258 135668 278052
rect 136850 278038 137048 278066
rect 136824 272536 136876 272542
rect 136824 272478 136876 272484
rect 136640 270496 136692 270502
rect 136638 270464 136640 270473
rect 136692 270464 136694 270473
rect 136638 270399 136694 270408
rect 135628 268252 135680 268258
rect 135628 268194 135680 268200
rect 132500 266484 132552 266490
rect 132500 266426 132552 266432
rect 64144 264512 64196 264518
rect 64144 264454 64196 264460
rect 136836 264330 136864 272478
rect 137020 270502 137048 278038
rect 137940 272542 137968 278052
rect 139136 275874 139164 278052
rect 140346 278038 140728 278066
rect 139124 275868 139176 275874
rect 139124 275810 139176 275816
rect 139400 273964 139452 273970
rect 139400 273906 139452 273912
rect 137928 272536 137980 272542
rect 137928 272478 137980 272484
rect 138480 271176 138532 271182
rect 138480 271118 138532 271124
rect 137008 270496 137060 270502
rect 137836 270496 137888 270502
rect 137008 270438 137060 270444
rect 137834 270464 137836 270473
rect 137888 270464 137890 270473
rect 137834 270399 137890 270408
rect 137468 270360 137520 270366
rect 137468 270302 137520 270308
rect 137480 266762 137508 270302
rect 137468 266756 137520 266762
rect 137468 266698 137520 266704
rect 138112 266620 138164 266626
rect 138112 266562 138164 266568
rect 136836 264302 137310 264330
rect 138124 264316 138152 266562
rect 138492 264330 138520 271118
rect 139412 264330 139440 273906
rect 140700 268258 140728 278038
rect 141056 275052 141108 275058
rect 141056 274994 141108 275000
rect 140136 268252 140188 268258
rect 140136 268194 140188 268200
rect 140688 268252 140740 268258
rect 140688 268194 140740 268200
rect 140148 267034 140176 268194
rect 140136 267028 140188 267034
rect 140136 266970 140188 266976
rect 140596 266892 140648 266898
rect 140596 266834 140648 266840
rect 138492 264302 138966 264330
rect 139412 264302 139794 264330
rect 140608 264316 140636 266834
rect 141068 264330 141096 274994
rect 141528 271182 141556 278052
rect 142724 272678 142752 278052
rect 142160 272672 142212 272678
rect 142160 272614 142212 272620
rect 142712 272672 142764 272678
rect 142712 272614 142764 272620
rect 141516 271176 141568 271182
rect 141516 271118 141568 271124
rect 142172 264330 142200 272614
rect 142712 271448 142764 271454
rect 142712 271390 142764 271396
rect 142724 264330 142752 271390
rect 143540 271312 143592 271318
rect 143540 271254 143592 271260
rect 143552 264330 143580 271254
rect 143920 269278 143948 278052
rect 145130 278038 145788 278066
rect 144920 275460 144972 275466
rect 144920 275402 144972 275408
rect 144932 273970 144960 275402
rect 145104 274100 145156 274106
rect 145104 274042 145156 274048
rect 144920 273964 144972 273970
rect 144920 273906 144972 273912
rect 143908 269272 143960 269278
rect 143908 269214 143960 269220
rect 144736 267436 144788 267442
rect 144736 267378 144788 267384
rect 141068 264302 141450 264330
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143552 264302 143934 264330
rect 144748 264316 144776 267378
rect 145116 264330 145144 274042
rect 145760 272678 145788 278038
rect 146220 274922 146248 278052
rect 146208 274916 146260 274922
rect 146208 274858 146260 274864
rect 145564 272672 145616 272678
rect 145564 272614 145616 272620
rect 145748 272672 145800 272678
rect 145748 272614 145800 272620
rect 145576 267442 145604 272614
rect 147416 272134 147444 278052
rect 148612 273970 148640 278052
rect 149612 275324 149664 275330
rect 149612 275266 149664 275272
rect 147864 273964 147916 273970
rect 147864 273906 147916 273912
rect 148600 273964 148652 273970
rect 148600 273906 148652 273912
rect 147404 272128 147456 272134
rect 147404 272070 147456 272076
rect 146392 269816 146444 269822
rect 146392 269758 146444 269764
rect 145564 267436 145616 267442
rect 145564 267378 145616 267384
rect 145116 264302 145590 264330
rect 146404 264316 146432 269758
rect 147220 266484 147272 266490
rect 147220 266426 147272 266432
rect 147232 264316 147260 266426
rect 147876 264330 147904 273906
rect 148416 272808 148468 272814
rect 148416 272750 148468 272756
rect 148428 264330 148456 272750
rect 149428 269952 149480 269958
rect 149428 269894 149480 269900
rect 149440 264330 149468 269894
rect 149624 266626 149652 275266
rect 149808 275058 149836 278052
rect 151018 278038 151768 278066
rect 149796 275052 149848 275058
rect 149796 274994 149848 275000
rect 151084 271992 151136 271998
rect 151084 271934 151136 271940
rect 150532 266892 150584 266898
rect 150532 266834 150584 266840
rect 149612 266620 149664 266626
rect 149612 266562 149664 266568
rect 147876 264302 148074 264330
rect 148428 264302 148902 264330
rect 149440 264302 149730 264330
rect 150544 264316 150572 266834
rect 151096 266762 151124 271934
rect 151740 268122 151768 278038
rect 152004 271584 152056 271590
rect 152004 271526 152056 271532
rect 151728 268116 151780 268122
rect 151728 268058 151780 268064
rect 151360 267164 151412 267170
rect 151360 267106 151412 267112
rect 151084 266756 151136 266762
rect 151084 266698 151136 266704
rect 151372 264316 151400 267106
rect 152016 264330 152044 271526
rect 152200 271318 152228 278052
rect 153396 275194 153424 278052
rect 152832 275188 152884 275194
rect 152832 275130 152884 275136
rect 153384 275188 153436 275194
rect 153384 275130 153436 275136
rect 152188 271312 152240 271318
rect 152188 271254 152240 271260
rect 152844 269958 152872 275130
rect 154500 274106 154528 278052
rect 154764 275596 154816 275602
rect 154764 275538 154816 275544
rect 154488 274100 154540 274106
rect 154488 274042 154540 274048
rect 153844 273556 153896 273562
rect 153844 273498 153896 273504
rect 153016 270088 153068 270094
rect 153016 270030 153068 270036
rect 152832 269952 152884 269958
rect 152832 269894 152884 269900
rect 152016 264302 152214 264330
rect 153028 264316 153056 270030
rect 153856 267714 153884 273498
rect 154776 267734 154804 275538
rect 155696 272814 155724 278052
rect 156892 275466 156920 278052
rect 158102 278038 158668 278066
rect 156880 275460 156932 275466
rect 156880 275402 156932 275408
rect 157616 274372 157668 274378
rect 157616 274314 157668 274320
rect 156144 272944 156196 272950
rect 156144 272886 156196 272892
rect 155684 272808 155736 272814
rect 155684 272750 155736 272756
rect 155500 268388 155552 268394
rect 155500 268330 155552 268336
rect 153476 267708 153528 267714
rect 153476 267650 153528 267656
rect 153844 267708 153896 267714
rect 153844 267650 153896 267656
rect 154684 267706 154804 267734
rect 153488 264330 153516 267650
rect 153488 264302 153870 264330
rect 154684 264316 154712 267706
rect 155512 264316 155540 268330
rect 156156 264330 156184 272886
rect 157156 269952 157208 269958
rect 157156 269894 157208 269900
rect 156156 264302 156354 264330
rect 157168 264316 157196 269894
rect 157628 264330 157656 274314
rect 158640 269822 158668 278038
rect 159284 274378 159312 278052
rect 160480 275738 160508 278052
rect 159456 275732 159508 275738
rect 159456 275674 159508 275680
rect 160468 275732 160520 275738
rect 160468 275674 160520 275680
rect 159272 274372 159324 274378
rect 159272 274314 159324 274320
rect 158812 271720 158864 271726
rect 158812 271662 158864 271668
rect 158628 269816 158680 269822
rect 158628 269758 158680 269764
rect 157628 264302 158010 264330
rect 158824 264316 158852 271662
rect 159468 266898 159496 275674
rect 160928 274508 160980 274514
rect 160928 274450 160980 274456
rect 160468 268524 160520 268530
rect 160468 268466 160520 268472
rect 159456 266892 159508 266898
rect 159456 266834 159508 266840
rect 159640 266620 159692 266626
rect 159640 266562 159692 266568
rect 159652 264316 159680 266562
rect 160480 264316 160508 268466
rect 160940 264330 160968 274450
rect 161584 268394 161612 278052
rect 162780 277394 162808 278052
rect 162688 277366 162808 277394
rect 162688 271454 162716 277366
rect 163504 276004 163556 276010
rect 163504 275946 163556 275952
rect 162860 273080 162912 273086
rect 162860 273022 162912 273028
rect 162676 271448 162728 271454
rect 162676 271390 162728 271396
rect 161572 268388 161624 268394
rect 161572 268330 161624 268336
rect 162124 266892 162176 266898
rect 162124 266834 162176 266840
rect 160940 264302 161322 264330
rect 162136 264316 162164 266834
rect 162872 264330 162900 273022
rect 163516 266422 163544 275946
rect 163976 275466 164004 278052
rect 163964 275460 164016 275466
rect 163964 275402 164016 275408
rect 164976 271856 165028 271862
rect 164976 271798 165028 271804
rect 163780 268660 163832 268666
rect 163780 268602 163832 268608
rect 163504 266416 163556 266422
rect 163504 266358 163556 266364
rect 162872 264302 162978 264330
rect 163792 264316 163820 268602
rect 164608 267300 164660 267306
rect 164608 267242 164660 267248
rect 164620 264316 164648 267242
rect 164988 264330 165016 271798
rect 165172 271590 165200 278052
rect 165896 273216 165948 273222
rect 165896 273158 165948 273164
rect 165160 271584 165212 271590
rect 165160 271526 165212 271532
rect 165908 264330 165936 273158
rect 166368 272950 166396 278052
rect 167564 276010 167592 278052
rect 167552 276004 167604 276010
rect 167552 275946 167604 275952
rect 168288 274780 168340 274786
rect 168288 274722 168340 274728
rect 166356 272944 166408 272950
rect 166356 272886 166408 272892
rect 168104 270632 168156 270638
rect 168104 270574 168156 270580
rect 167920 268796 167972 268802
rect 167920 268738 167972 268744
rect 167092 266416 167144 266422
rect 167092 266358 167144 266364
rect 164988 264302 165462 264330
rect 165908 264302 166290 264330
rect 167104 264316 167132 266358
rect 167932 264316 167960 268738
rect 168116 267170 168144 270574
rect 168300 268802 168328 274722
rect 168760 274514 168788 278052
rect 169024 275188 169076 275194
rect 169024 275130 169076 275136
rect 168748 274508 168800 274514
rect 168748 274450 168800 274456
rect 168748 270224 168800 270230
rect 168748 270166 168800 270172
rect 168288 268796 168340 268802
rect 168288 268738 168340 268744
rect 168564 267572 168616 267578
rect 168564 267514 168616 267520
rect 168104 267164 168156 267170
rect 168104 267106 168156 267112
rect 168576 266422 168604 267514
rect 168564 266416 168616 266422
rect 168564 266358 168616 266364
rect 168760 264316 168788 270166
rect 169036 267578 169064 275130
rect 169864 271726 169892 278052
rect 171060 275602 171088 278052
rect 171048 275596 171100 275602
rect 171048 275538 171100 275544
rect 171600 274644 171652 274650
rect 171600 274586 171652 274592
rect 169852 271720 169904 271726
rect 169852 271662 169904 271668
rect 169944 271040 169996 271046
rect 169944 270982 169996 270988
rect 169024 267572 169076 267578
rect 169024 267514 169076 267520
rect 169576 266416 169628 266422
rect 169576 266358 169628 266364
rect 169588 264316 169616 266358
rect 169956 264330 169984 270982
rect 171232 268932 171284 268938
rect 171232 268874 171284 268880
rect 169956 264302 170430 264330
rect 171244 264316 171272 268874
rect 171612 264330 171640 274586
rect 172256 273086 172284 278052
rect 173466 278038 173756 278066
rect 174662 278038 175136 278066
rect 175858 278038 176608 278066
rect 173256 273692 173308 273698
rect 173256 273634 173308 273640
rect 172244 273080 172296 273086
rect 172244 273022 172296 273028
rect 172520 272400 172572 272406
rect 172520 272342 172572 272348
rect 172532 264330 172560 272342
rect 173268 264330 173296 273634
rect 173728 269958 173756 278038
rect 174268 275868 174320 275874
rect 174268 275810 174320 275816
rect 174280 271862 174308 275810
rect 174268 271856 174320 271862
rect 174268 271798 174320 271804
rect 173716 269952 173768 269958
rect 173716 269894 173768 269900
rect 175108 269074 175136 278038
rect 175280 273828 175332 273834
rect 175280 273770 175332 273776
rect 174544 269068 174596 269074
rect 174544 269010 174596 269016
rect 175096 269068 175148 269074
rect 175096 269010 175148 269016
rect 171612 264302 172086 264330
rect 172532 264302 172914 264330
rect 173268 264302 173742 264330
rect 174556 264316 174584 269010
rect 175292 264330 175320 273770
rect 176580 270094 176608 278038
rect 176568 270088 176620 270094
rect 176568 270030 176620 270036
rect 176200 269680 176252 269686
rect 176200 269622 176252 269628
rect 175292 264302 175398 264330
rect 176212 264316 176240 269622
rect 176948 268666 176976 278052
rect 178144 275874 178172 278052
rect 178684 276004 178736 276010
rect 178684 275946 178736 275952
rect 178132 275868 178184 275874
rect 178132 275810 178184 275816
rect 177488 270904 177540 270910
rect 177488 270846 177540 270852
rect 176936 268660 176988 268666
rect 176936 268602 176988 268608
rect 177028 267164 177080 267170
rect 177028 267106 177080 267112
rect 177040 264316 177068 267106
rect 177500 264330 177528 270846
rect 178316 269408 178368 269414
rect 178316 269350 178368 269356
rect 177672 269068 177724 269074
rect 177672 269010 177724 269016
rect 177684 267170 177712 269010
rect 177672 267164 177724 267170
rect 177672 267106 177724 267112
rect 178328 264330 178356 269350
rect 178696 266898 178724 275946
rect 179340 274650 179368 278052
rect 180550 278038 180748 278066
rect 179328 274644 179380 274650
rect 179328 274586 179380 274592
rect 179880 272264 179932 272270
rect 179880 272206 179932 272212
rect 178684 266892 178736 266898
rect 178684 266834 178736 266840
rect 179512 266756 179564 266762
rect 179512 266698 179564 266704
rect 177500 264302 177882 264330
rect 178328 264302 178710 264330
rect 179524 264316 179552 266698
rect 179892 264330 179920 272206
rect 180720 268530 180748 278038
rect 181732 272542 181760 278052
rect 182942 278038 183508 278066
rect 184138 278038 184888 278066
rect 182456 274236 182508 274242
rect 182456 274178 182508 274184
rect 181720 272536 181772 272542
rect 181720 272478 181772 272484
rect 181168 269544 181220 269550
rect 181168 269486 181220 269492
rect 180708 268524 180760 268530
rect 180708 268466 180760 268472
rect 179892 264302 180366 264330
rect 181180 264316 181208 269486
rect 181996 268796 182048 268802
rect 181996 268738 182048 268744
rect 182008 264316 182036 268738
rect 182468 264330 182496 274178
rect 183480 269686 183508 278038
rect 183652 270496 183704 270502
rect 183652 270438 183704 270444
rect 183468 269680 183520 269686
rect 183468 269622 183520 269628
rect 182468 264302 182850 264330
rect 183664 264316 183692 270438
rect 184860 270230 184888 278038
rect 185228 276010 185256 278052
rect 185216 276004 185268 276010
rect 185216 275946 185268 275952
rect 185584 274916 185636 274922
rect 185584 274858 185636 274864
rect 185124 270768 185176 270774
rect 185124 270710 185176 270716
rect 184848 270224 184900 270230
rect 184848 270166 184900 270172
rect 184480 267708 184532 267714
rect 184480 267650 184532 267656
rect 184492 264316 184520 267650
rect 185136 264330 185164 270710
rect 185596 270502 185624 274858
rect 186424 273222 186452 278052
rect 187436 278038 187634 278066
rect 186412 273216 186464 273222
rect 186412 273158 186464 273164
rect 186964 272536 187016 272542
rect 186964 272478 187016 272484
rect 185584 270496 185636 270502
rect 185584 270438 185636 270444
rect 186136 270360 186188 270366
rect 186136 270302 186188 270308
rect 185136 264302 185334 264330
rect 186148 264316 186176 270302
rect 186976 267306 187004 272478
rect 187436 271046 187464 278038
rect 188816 277394 188844 278052
rect 188816 277366 188936 277394
rect 187700 272400 187752 272406
rect 187700 272342 187752 272348
rect 187424 271040 187476 271046
rect 187424 270982 187476 270988
rect 186964 267300 187016 267306
rect 186964 267242 187016 267248
rect 186964 267028 187016 267034
rect 186964 266970 187016 266976
rect 186976 264316 187004 266970
rect 187712 264330 187740 272342
rect 188908 268870 188936 277366
rect 190012 275194 190040 278052
rect 190000 275188 190052 275194
rect 190000 275130 190052 275136
rect 189080 275052 189132 275058
rect 189080 274994 189132 275000
rect 189092 272270 189120 274994
rect 189080 272264 189132 272270
rect 189080 272206 189132 272212
rect 189172 271856 189224 271862
rect 189172 271798 189224 271804
rect 188896 268864 188948 268870
rect 188896 268806 188948 268812
rect 188620 268252 188672 268258
rect 188620 268194 188672 268200
rect 187712 264302 187818 264330
rect 188632 264316 188660 268194
rect 189184 264330 189212 271798
rect 191208 271182 191236 278052
rect 192404 274242 192432 278052
rect 192392 274236 192444 274242
rect 192392 274178 192444 274184
rect 193508 273834 193536 278052
rect 194718 278038 195008 278066
rect 194784 273964 194836 273970
rect 194784 273906 194836 273912
rect 193496 273828 193548 273834
rect 193496 273770 193548 273776
rect 192392 272672 192444 272678
rect 192392 272614 192444 272620
rect 189816 271176 189868 271182
rect 189816 271118 189868 271124
rect 191196 271176 191248 271182
rect 191196 271118 191248 271124
rect 189828 264330 189856 271118
rect 191104 269272 191156 269278
rect 191104 269214 191156 269220
rect 190460 268864 190512 268870
rect 190460 268806 190512 268812
rect 190472 267034 190500 268806
rect 190460 267028 190512 267034
rect 190460 266970 190512 266976
rect 189184 264302 189474 264330
rect 189828 264302 190302 264330
rect 191116 264316 191144 269214
rect 191932 267436 191984 267442
rect 191932 267378 191984 267384
rect 191944 264316 191972 267378
rect 192404 264330 192432 272614
rect 193220 272128 193272 272134
rect 193220 272070 193272 272076
rect 193232 264330 193260 272070
rect 194416 270496 194468 270502
rect 194416 270438 194468 270444
rect 192404 264302 192786 264330
rect 193232 264302 193614 264330
rect 194428 264316 194456 270438
rect 194796 264330 194824 273906
rect 194980 272406 195008 278038
rect 195900 272542 195928 278052
rect 197096 272678 197124 278052
rect 198096 274100 198148 274106
rect 198096 274042 198148 274048
rect 197084 272672 197136 272678
rect 197084 272614 197136 272620
rect 195888 272536 195940 272542
rect 195888 272478 195940 272484
rect 194968 272400 195020 272406
rect 194968 272342 195020 272348
rect 196440 272264 196492 272270
rect 196440 272206 196492 272212
rect 196072 268116 196124 268122
rect 196072 268058 196124 268064
rect 194796 264302 195270 264330
rect 196084 264316 196112 268058
rect 196452 264330 196480 272206
rect 197360 271312 197412 271318
rect 197360 271254 197412 271260
rect 197372 264330 197400 271254
rect 198108 264330 198136 274042
rect 198292 271318 198320 278052
rect 199502 278038 199976 278066
rect 199568 275732 199620 275738
rect 199568 275674 199620 275680
rect 198280 271312 198332 271318
rect 198280 271254 198332 271260
rect 199384 267572 199436 267578
rect 199384 267514 199436 267520
rect 196452 264302 196926 264330
rect 197372 264302 197754 264330
rect 198108 264302 198582 264330
rect 199396 264316 199424 267514
rect 199580 267442 199608 275674
rect 199948 270366 199976 278038
rect 200120 272808 200172 272814
rect 200120 272750 200172 272756
rect 199936 270360 199988 270366
rect 199936 270302 199988 270308
rect 199568 267436 199620 267442
rect 199568 267378 199620 267384
rect 200132 264330 200160 272750
rect 200592 268802 200620 278052
rect 201788 277394 201816 278052
rect 201696 277366 201816 277394
rect 200764 275324 200816 275330
rect 200764 275266 200816 275272
rect 200776 270502 200804 275266
rect 200764 270496 200816 270502
rect 200764 270438 200816 270444
rect 201696 269822 201724 277366
rect 202328 274372 202380 274378
rect 202328 274314 202380 274320
rect 201868 270496 201920 270502
rect 201868 270438 201920 270444
rect 201040 269816 201092 269822
rect 201040 269758 201092 269764
rect 201684 269816 201736 269822
rect 201684 269758 201736 269764
rect 200580 268796 200632 268802
rect 200580 268738 200632 268744
rect 200132 264302 200238 264330
rect 201052 264316 201080 269758
rect 201880 264316 201908 270438
rect 202340 264330 202368 274314
rect 202984 271862 203012 278052
rect 202972 271856 203024 271862
rect 202972 271798 203024 271804
rect 204180 269550 204208 278052
rect 205376 272814 205404 278052
rect 206586 278038 206876 278066
rect 206376 275460 206428 275466
rect 206376 275402 206428 275408
rect 205364 272808 205416 272814
rect 205364 272750 205416 272756
rect 205640 271584 205692 271590
rect 205640 271526 205692 271532
rect 204720 271448 204772 271454
rect 204720 271390 204772 271396
rect 204168 269544 204220 269550
rect 204168 269486 204220 269492
rect 203524 268388 203576 268394
rect 203524 268330 203576 268336
rect 202340 264302 202722 264330
rect 203536 264316 203564 268330
rect 204352 267436 204404 267442
rect 204352 267378 204404 267384
rect 204364 264316 204392 267378
rect 204732 264330 204760 271390
rect 205456 269680 205508 269686
rect 205456 269622 205508 269628
rect 205468 267442 205496 269622
rect 205456 267436 205508 267442
rect 205456 267378 205508 267384
rect 205652 264330 205680 271526
rect 206388 264330 206416 275402
rect 206848 270502 206876 278038
rect 207768 274786 207796 278052
rect 207756 274780 207808 274786
rect 207756 274722 207808 274728
rect 208400 274508 208452 274514
rect 208400 274450 208452 274456
rect 207296 272944 207348 272950
rect 207296 272886 207348 272892
rect 206836 270496 206888 270502
rect 206836 270438 206888 270444
rect 207308 264330 207336 272886
rect 208412 264330 208440 274450
rect 208872 273970 208900 278052
rect 210068 274106 210096 278052
rect 210700 274780 210752 274786
rect 210700 274722 210752 274728
rect 210056 274100 210108 274106
rect 210056 274042 210108 274048
rect 208860 273964 208912 273970
rect 208860 273906 208912 273912
rect 209780 273080 209832 273086
rect 209780 273022 209832 273028
rect 209320 266892 209372 266898
rect 209320 266834 209372 266840
rect 204732 264302 205206 264330
rect 205652 264302 206034 264330
rect 206388 264302 206862 264330
rect 207308 264302 207690 264330
rect 208412 264302 208518 264330
rect 209332 264316 209360 266834
rect 209792 265674 209820 273022
rect 209964 271720 210016 271726
rect 209964 271662 210016 271668
rect 209780 265668 209832 265674
rect 209780 265610 209832 265616
rect 209976 264330 210004 271662
rect 210712 268394 210740 274722
rect 211264 272950 211292 278052
rect 211620 275596 211672 275602
rect 211620 275538 211672 275544
rect 211252 272944 211304 272950
rect 211252 272886 211304 272892
rect 211160 270088 211212 270094
rect 211160 270030 211212 270036
rect 210700 268388 210752 268394
rect 210700 268330 210752 268336
rect 211172 266422 211200 270030
rect 211160 266416 211212 266422
rect 211160 266358 211212 266364
rect 210700 265668 210752 265674
rect 210700 265610 210752 265616
rect 210712 264330 210740 265610
rect 211632 264330 211660 275538
rect 212460 270094 212488 278052
rect 213656 271454 213684 278052
rect 214852 275330 214880 278052
rect 214840 275324 214892 275330
rect 214840 275266 214892 275272
rect 214564 274644 214616 274650
rect 214564 274586 214616 274592
rect 213644 271448 213696 271454
rect 213644 271390 213696 271396
rect 212448 270088 212500 270094
rect 212448 270030 212500 270036
rect 212632 269952 212684 269958
rect 212632 269894 212684 269900
rect 209976 264302 210174 264330
rect 210712 264302 211002 264330
rect 211632 264302 211830 264330
rect 212644 264316 212672 269894
rect 214288 267164 214340 267170
rect 214288 267106 214340 267112
rect 213460 266416 213512 266422
rect 213460 266358 213512 266364
rect 213472 264316 213500 266358
rect 214300 264316 214328 267106
rect 214576 266422 214604 274586
rect 215956 271590 215984 278052
rect 216680 275868 216732 275874
rect 216680 275810 216732 275816
rect 215944 271584 215996 271590
rect 215944 271526 215996 271532
rect 215944 271040 215996 271046
rect 215944 270982 215996 270988
rect 215116 268660 215168 268666
rect 215116 268602 215168 268608
rect 214564 266416 214616 266422
rect 214564 266358 214616 266364
rect 215128 264316 215156 268602
rect 215956 267578 215984 270982
rect 215944 267572 215996 267578
rect 215944 267514 215996 267520
rect 215944 266416 215996 266422
rect 215944 266358 215996 266364
rect 215956 264316 215984 266358
rect 216692 264330 216720 275810
rect 217152 275738 217180 278052
rect 217140 275732 217192 275738
rect 217140 275674 217192 275680
rect 218348 275602 218376 278052
rect 218336 275596 218388 275602
rect 218336 275538 218388 275544
rect 218704 273216 218756 273222
rect 218704 273158 218756 273164
rect 217600 268524 217652 268530
rect 217600 268466 217652 268472
rect 216692 264302 216798 264330
rect 217612 264316 217640 268466
rect 218428 267436 218480 267442
rect 218428 267378 218480 267384
rect 218440 264316 218468 267378
rect 218716 266898 218744 273158
rect 219544 273086 219572 278052
rect 219532 273080 219584 273086
rect 219532 273022 219584 273028
rect 220740 272950 220768 278052
rect 221280 276004 221332 276010
rect 221280 275946 221332 275952
rect 220084 272944 220136 272950
rect 220084 272886 220136 272892
rect 220728 272944 220780 272950
rect 220728 272886 220780 272892
rect 219348 270224 219400 270230
rect 219348 270166 219400 270172
rect 219360 267458 219388 270166
rect 219360 267430 219664 267458
rect 219256 267300 219308 267306
rect 219256 267242 219308 267248
rect 218704 266892 218756 266898
rect 218704 266834 218756 266840
rect 219268 264316 219296 267242
rect 219636 264330 219664 267430
rect 220096 267170 220124 272886
rect 220084 267164 220136 267170
rect 220084 267106 220136 267112
rect 220912 266892 220964 266898
rect 220912 266834 220964 266840
rect 219636 264302 220110 264330
rect 220924 264316 220952 266834
rect 221292 264330 221320 275946
rect 221936 275466 221964 278052
rect 221924 275460 221976 275466
rect 221924 275402 221976 275408
rect 222936 275188 222988 275194
rect 222936 275130 222988 275136
rect 222568 267572 222620 267578
rect 222568 267514 222620 267520
rect 221292 264302 221766 264330
rect 222580 264316 222608 267514
rect 222948 264330 222976 275130
rect 223132 274378 223160 278052
rect 224236 275874 224264 278052
rect 224224 275868 224276 275874
rect 224224 275810 224276 275816
rect 224224 275732 224276 275738
rect 224224 275674 224276 275680
rect 223120 274372 223172 274378
rect 223120 274314 223172 274320
rect 223488 269544 223540 269550
rect 223488 269486 223540 269492
rect 223500 267306 223528 269486
rect 224236 268666 224264 275674
rect 224960 274236 225012 274242
rect 224960 274178 225012 274184
rect 224224 268660 224276 268666
rect 224224 268602 224276 268608
rect 223488 267300 223540 267306
rect 223488 267242 223540 267248
rect 224224 267028 224276 267034
rect 224224 266970 224276 266976
rect 222948 264302 223422 264330
rect 224236 264316 224264 266970
rect 224972 265674 225000 274178
rect 225432 271726 225460 278052
rect 226432 273828 226484 273834
rect 226432 273770 226484 273776
rect 225420 271720 225472 271726
rect 225420 271662 225472 271668
rect 225144 271176 225196 271182
rect 225144 271118 225196 271124
rect 224960 265668 225012 265674
rect 224960 265610 225012 265616
rect 225156 265554 225184 271118
rect 225604 265668 225656 265674
rect 225604 265610 225656 265616
rect 225064 265526 225184 265554
rect 225064 264316 225092 265526
rect 225616 264330 225644 265610
rect 226444 264330 226472 273770
rect 226628 269958 226656 278052
rect 227838 278038 228128 278066
rect 228100 272542 228128 278038
rect 229020 275738 229048 278052
rect 229008 275732 229060 275738
rect 229008 275674 229060 275680
rect 229100 272672 229152 272678
rect 229100 272614 229152 272620
rect 227904 272536 227956 272542
rect 227904 272478 227956 272484
rect 228088 272536 228140 272542
rect 228088 272478 228140 272484
rect 227168 272400 227220 272406
rect 227168 272342 227220 272348
rect 226616 269952 226668 269958
rect 226616 269894 226668 269900
rect 227180 264330 227208 272342
rect 227916 264330 227944 272478
rect 228364 271720 228416 271726
rect 228364 271662 228416 271668
rect 228376 267034 228404 271662
rect 228364 267028 228416 267034
rect 228364 266970 228416 266976
rect 229112 264330 229140 272614
rect 229560 271312 229612 271318
rect 229560 271254 229612 271260
rect 229572 264330 229600 271254
rect 230216 271182 230244 278052
rect 231334 278038 231716 278066
rect 230204 271176 230256 271182
rect 230204 271118 230256 271124
rect 230848 270360 230900 270366
rect 230848 270302 230900 270308
rect 225616 264302 225906 264330
rect 226444 264302 226734 264330
rect 227180 264302 227562 264330
rect 227916 264302 228390 264330
rect 229112 264302 229218 264330
rect 229572 264302 230046 264330
rect 230860 264316 230888 270302
rect 231308 268796 231360 268802
rect 231308 268738 231360 268744
rect 231320 264330 231348 268738
rect 231688 268530 231716 278038
rect 232516 276010 232544 278052
rect 232504 276004 232556 276010
rect 232504 275946 232556 275952
rect 232688 275868 232740 275874
rect 232688 275810 232740 275816
rect 232700 270366 232728 275810
rect 233712 272678 233740 278052
rect 234922 278038 235304 278066
rect 233884 275596 233936 275602
rect 233884 275538 233936 275544
rect 233700 272672 233752 272678
rect 233700 272614 233752 272620
rect 233240 271856 233292 271862
rect 233240 271798 233292 271804
rect 232688 270360 232740 270366
rect 232688 270302 232740 270308
rect 232504 269816 232556 269822
rect 232504 269758 232556 269764
rect 231676 268524 231728 268530
rect 231676 268466 231728 268472
rect 231320 264302 231702 264330
rect 232516 264316 232544 269758
rect 233252 264330 233280 271798
rect 233896 267442 233924 275538
rect 234804 272808 234856 272814
rect 234804 272750 234856 272756
rect 233884 267436 233936 267442
rect 233884 267378 233936 267384
rect 234160 267300 234212 267306
rect 234160 267242 234212 267248
rect 233252 264302 233358 264330
rect 234172 264316 234200 267242
rect 234816 264330 234844 272750
rect 235276 271318 235304 278038
rect 236104 275874 236132 278052
rect 236092 275868 236144 275874
rect 236092 275810 236144 275816
rect 235264 271312 235316 271318
rect 235264 271254 235316 271260
rect 235816 270496 235868 270502
rect 235816 270438 235868 270444
rect 234816 264302 235014 264330
rect 235828 264316 235856 270438
rect 237208 269822 237236 278052
rect 237840 274100 237892 274106
rect 237840 274042 237892 274048
rect 237380 273964 237432 273970
rect 237380 273906 237432 273912
rect 237196 269816 237248 269822
rect 237196 269758 237248 269764
rect 236644 268388 236696 268394
rect 236644 268330 236696 268336
rect 236656 264316 236684 268330
rect 237392 264330 237420 273906
rect 237852 264330 237880 274042
rect 238496 273970 238524 278052
rect 239220 276004 239272 276010
rect 239220 275946 239272 275952
rect 239232 274242 239260 275946
rect 239600 275602 239628 278052
rect 239588 275596 239640 275602
rect 239588 275538 239640 275544
rect 239404 275324 239456 275330
rect 239404 275266 239456 275272
rect 239220 274236 239272 274242
rect 239220 274178 239272 274184
rect 238484 273964 238536 273970
rect 238484 273906 238536 273912
rect 239128 267164 239180 267170
rect 239128 267106 239180 267112
rect 237392 264302 237498 264330
rect 237852 264302 238326 264330
rect 239140 264316 239168 267106
rect 239416 266422 239444 275266
rect 240796 271454 240824 278052
rect 241992 277394 242020 278052
rect 241900 277366 242020 277394
rect 240416 271448 240468 271454
rect 240416 271390 240468 271396
rect 240784 271448 240836 271454
rect 240784 271390 240836 271396
rect 239956 270088 240008 270094
rect 239956 270030 240008 270036
rect 239404 266416 239456 266422
rect 239404 266358 239456 266364
rect 239968 264316 239996 270030
rect 240428 264330 240456 271390
rect 241900 270094 241928 277366
rect 243188 275330 243216 278052
rect 243544 275732 243596 275738
rect 243544 275674 243596 275680
rect 243176 275324 243228 275330
rect 243176 275266 243228 275272
rect 242072 271584 242124 271590
rect 242072 271526 242124 271532
rect 241888 270088 241940 270094
rect 241888 270030 241940 270036
rect 241612 266416 241664 266422
rect 241612 266358 241664 266364
rect 240428 264302 240810 264330
rect 241624 264316 241652 266358
rect 242084 264330 242112 271526
rect 243268 268660 243320 268666
rect 243268 268602 243320 268608
rect 242084 264302 242466 264330
rect 243280 264316 243308 268602
rect 243556 267442 243584 275674
rect 243728 275460 243780 275466
rect 243728 275402 243780 275408
rect 243544 267436 243596 267442
rect 243544 267378 243596 267384
rect 243740 266422 243768 275402
rect 244384 270230 244412 278052
rect 245396 278038 245502 278066
rect 246790 278038 246988 278066
rect 244556 273080 244608 273086
rect 244556 273022 244608 273028
rect 244372 270224 244424 270230
rect 244372 270166 244424 270172
rect 244096 267300 244148 267306
rect 244096 267242 244148 267248
rect 243728 266416 243780 266422
rect 243728 266358 243780 266364
rect 244108 264316 244136 267242
rect 244568 264330 244596 273022
rect 245396 272814 245424 278038
rect 245752 272944 245804 272950
rect 245752 272886 245804 272892
rect 245384 272808 245436 272814
rect 245384 272750 245436 272756
rect 244568 264302 244950 264330
rect 245764 264316 245792 272886
rect 246960 267170 246988 278038
rect 247224 274372 247276 274378
rect 247224 274314 247276 274320
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 246580 266416 246632 266422
rect 246580 266358 246632 266364
rect 246592 264316 246620 266358
rect 247236 264330 247264 274314
rect 247880 272950 247908 278052
rect 249076 274106 249104 278052
rect 250272 275738 250300 278052
rect 250444 275868 250496 275874
rect 250444 275810 250496 275816
rect 250260 275732 250312 275738
rect 250260 275674 250312 275680
rect 249064 274100 249116 274106
rect 249064 274042 249116 274048
rect 247868 272944 247920 272950
rect 247868 272886 247920 272892
rect 249064 272536 249116 272542
rect 249064 272478 249116 272484
rect 248236 270360 248288 270366
rect 248236 270302 248288 270308
rect 247236 264302 247434 264330
rect 248248 264316 248276 270302
rect 249076 267034 249104 272478
rect 249892 269952 249944 269958
rect 249892 269894 249944 269900
rect 249064 267028 249116 267034
rect 249064 266970 249116 266976
rect 249064 266892 249116 266898
rect 249064 266834 249116 266840
rect 249076 264316 249104 266834
rect 249904 264316 249932 269894
rect 250456 266422 250484 275810
rect 251468 271046 251496 278052
rect 252008 271176 252060 271182
rect 252008 271118 252060 271124
rect 251456 271040 251508 271046
rect 251456 270982 251508 270988
rect 251548 267436 251600 267442
rect 251548 267378 251600 267384
rect 250720 267028 250772 267034
rect 250720 266970 250772 266976
rect 250444 266416 250496 266422
rect 250444 266358 250496 266364
rect 250732 264316 250760 266970
rect 251560 264316 251588 267378
rect 252020 264330 252048 271118
rect 252664 268394 252692 278052
rect 253860 274718 253888 278052
rect 253848 274712 253900 274718
rect 253848 274654 253900 274660
rect 253940 274236 253992 274242
rect 253940 274178 253992 274184
rect 253204 268524 253256 268530
rect 253204 268466 253256 268472
rect 252652 268388 252704 268394
rect 252652 268330 252704 268336
rect 252020 264302 252402 264330
rect 253216 264316 253244 268466
rect 253952 264330 253980 274178
rect 254400 272672 254452 272678
rect 254400 272614 254452 272620
rect 254412 264330 254440 272614
rect 254964 272542 254992 278052
rect 255964 275596 256016 275602
rect 255964 275538 256016 275544
rect 254952 272536 255004 272542
rect 254952 272478 255004 272484
rect 255320 271312 255372 271318
rect 255320 271254 255372 271260
rect 255332 264330 255360 271254
rect 255976 267034 256004 275538
rect 256160 275466 256188 278052
rect 257356 275602 257384 278052
rect 257344 275596 257396 275602
rect 257344 275538 257396 275544
rect 256148 275460 256200 275466
rect 256148 275402 256200 275408
rect 256700 275324 256752 275330
rect 256700 275266 256752 275272
rect 256712 271318 256740 275266
rect 256884 274712 256936 274718
rect 256884 274654 256936 274660
rect 256700 271312 256752 271318
rect 256700 271254 256752 271260
rect 256896 269958 256924 274654
rect 258080 273828 258132 273834
rect 258080 273770 258132 273776
rect 256884 269952 256936 269958
rect 256884 269894 256936 269900
rect 257344 269816 257396 269822
rect 257344 269758 257396 269764
rect 255964 267028 256016 267034
rect 255964 266970 256016 266976
rect 256516 266416 256568 266422
rect 256516 266358 256568 266364
rect 253952 264302 254058 264330
rect 254412 264302 254886 264330
rect 255332 264302 255714 264330
rect 256528 264316 256556 266358
rect 257356 264316 257384 269758
rect 258092 264330 258120 273770
rect 258552 269822 258580 278052
rect 259748 277394 259776 278052
rect 259748 277366 259868 277394
rect 259368 275732 259420 275738
rect 259368 275674 259420 275680
rect 259380 273834 259408 275674
rect 259368 273828 259420 273834
rect 259368 273770 259420 273776
rect 259840 271454 259868 277366
rect 260944 275806 260972 278052
rect 260932 275800 260984 275806
rect 260932 275742 260984 275748
rect 259644 271448 259696 271454
rect 259644 271390 259696 271396
rect 259828 271448 259880 271454
rect 259828 271390 259880 271396
rect 258540 269816 258592 269822
rect 258540 269758 258592 269764
rect 259000 267028 259052 267034
rect 259000 266970 259052 266976
rect 258092 264302 258198 264330
rect 259012 264316 259040 266970
rect 259656 264330 259684 271390
rect 262048 271318 262076 278052
rect 262312 275596 262364 275602
rect 262312 275538 262364 275544
rect 262324 272814 262352 275538
rect 263244 275126 263272 278052
rect 263232 275120 263284 275126
rect 263232 275062 263284 275068
rect 264244 272944 264296 272950
rect 264244 272886 264296 272892
rect 262312 272808 262364 272814
rect 262312 272750 262364 272756
rect 262680 272672 262732 272678
rect 262680 272614 262732 272620
rect 261024 271312 261076 271318
rect 261024 271254 261076 271260
rect 262036 271312 262088 271318
rect 262036 271254 262088 271260
rect 260656 270088 260708 270094
rect 260656 270030 260708 270036
rect 259656 264302 259854 264330
rect 260668 264316 260696 270030
rect 261036 264330 261064 271254
rect 262312 270224 262364 270230
rect 262312 270166 262364 270172
rect 261036 264302 261510 264330
rect 262324 264316 262352 270166
rect 262692 264330 262720 272614
rect 264256 267734 264284 272886
rect 264440 272678 264468 278052
rect 265650 278038 266216 278066
rect 265256 274100 265308 274106
rect 265256 274042 265308 274048
rect 264428 272672 264480 272678
rect 264428 272614 264480 272620
rect 264256 267706 264376 267734
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 262692 264302 263166 264330
rect 263980 264316 264008 267106
rect 264348 264330 264376 267706
rect 265268 264330 265296 274042
rect 266188 270094 266216 278038
rect 266360 275800 266412 275806
rect 266360 275742 266412 275748
rect 266372 274106 266400 275742
rect 266832 275602 266860 278052
rect 266820 275596 266872 275602
rect 266820 275538 266872 275544
rect 266360 274100 266412 274106
rect 266360 274042 266412 274048
rect 266360 273828 266412 273834
rect 266360 273770 266412 273776
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 266372 264330 266400 273770
rect 268028 271182 268056 278052
rect 269224 275398 269252 278052
rect 269212 275392 269264 275398
rect 269212 275334 269264 275340
rect 269120 275256 269172 275262
rect 269120 275198 269172 275204
rect 269132 272338 269160 275198
rect 270328 272542 270356 278052
rect 271524 273970 271552 278052
rect 272734 278038 273116 278066
rect 273930 278038 274312 278066
rect 271512 273964 271564 273970
rect 271512 273906 271564 273912
rect 270960 272808 271012 272814
rect 270960 272750 271012 272756
rect 269304 272536 269356 272542
rect 269304 272478 269356 272484
rect 270316 272536 270368 272542
rect 270316 272478 270368 272484
rect 269120 272332 269172 272338
rect 269120 272274 269172 272280
rect 268016 271176 268068 271182
rect 268016 271118 268068 271124
rect 266912 271040 266964 271046
rect 266912 270982 266964 270988
rect 266924 264330 266952 270982
rect 268936 269952 268988 269958
rect 268936 269894 268988 269900
rect 268108 268388 268160 268394
rect 268108 268330 268160 268336
rect 264348 264302 264822 264330
rect 265268 264302 265650 264330
rect 266372 264302 266478 264330
rect 266924 264302 267306 264330
rect 268120 264316 268148 268330
rect 268948 264316 268976 269894
rect 269316 264330 269344 272478
rect 270592 272332 270644 272338
rect 270592 272274 270644 272280
rect 269316 264302 269790 264330
rect 270604 264316 270632 272274
rect 270972 264330 271000 272750
rect 272616 271448 272668 271454
rect 272616 271390 272668 271396
rect 272248 269816 272300 269822
rect 272248 269758 272300 269764
rect 270972 264302 271446 264330
rect 272260 264316 272288 269758
rect 272628 264330 272656 271390
rect 273088 269822 273116 278038
rect 273260 275120 273312 275126
rect 273260 275062 273312 275068
rect 273076 269816 273128 269822
rect 273076 269758 273128 269764
rect 273272 269074 273300 275062
rect 273536 274100 273588 274106
rect 273536 274042 273588 274048
rect 273260 269068 273312 269074
rect 273260 269010 273312 269016
rect 273548 264330 273576 274042
rect 274284 272814 274312 278038
rect 274640 275392 274692 275398
rect 274640 275334 274692 275340
rect 274272 272808 274324 272814
rect 274272 272750 274324 272756
rect 274652 271862 274680 275334
rect 275112 274718 275140 278052
rect 276308 275330 276336 278052
rect 276480 275596 276532 275602
rect 276480 275538 276532 275544
rect 276296 275324 276348 275330
rect 276296 275266 276348 275272
rect 275100 274712 275152 274718
rect 275100 274654 275152 274660
rect 276020 272672 276072 272678
rect 276020 272614 276072 272620
rect 274640 271856 274692 271862
rect 274640 271798 274692 271804
rect 274640 271312 274692 271318
rect 274640 271254 274692 271260
rect 274652 264330 274680 271254
rect 275560 269068 275612 269074
rect 275560 269010 275612 269016
rect 272628 264302 273102 264330
rect 273548 264302 273930 264330
rect 274652 264302 274758 264330
rect 275572 264316 275600 269010
rect 276032 264330 276060 272614
rect 276492 267782 276520 275538
rect 277504 275534 277532 278052
rect 277492 275528 277544 275534
rect 277492 275470 277544 275476
rect 278044 274712 278096 274718
rect 278044 274654 278096 274660
rect 278056 270502 278084 274654
rect 278608 274106 278636 278052
rect 278596 274100 278648 274106
rect 278596 274042 278648 274048
rect 279240 271856 279292 271862
rect 279240 271798 279292 271804
rect 278780 271176 278832 271182
rect 278780 271118 278832 271124
rect 278044 270496 278096 270502
rect 278044 270438 278096 270444
rect 277216 270088 277268 270094
rect 277216 270030 277268 270036
rect 276480 267776 276532 267782
rect 276480 267718 276532 267724
rect 276032 264302 276414 264330
rect 277228 264316 277256 270030
rect 278044 267776 278096 267782
rect 278044 267718 278096 267724
rect 278056 264316 278084 267718
rect 278792 264330 278820 271118
rect 279252 264330 279280 271798
rect 279804 271182 279832 278052
rect 280344 273964 280396 273970
rect 280344 273906 280396 273912
rect 279792 271176 279844 271182
rect 279792 271118 279844 271124
rect 280356 265674 280384 273906
rect 281000 273086 281028 278052
rect 282210 278038 282776 278066
rect 280988 273080 281040 273086
rect 280988 273022 281040 273028
rect 280528 272536 280580 272542
rect 280528 272478 280580 272484
rect 280344 265668 280396 265674
rect 280344 265610 280396 265616
rect 278792 264302 278898 264330
rect 279252 264302 279726 264330
rect 280540 264316 280568 272478
rect 282184 269816 282236 269822
rect 282184 269758 282236 269764
rect 280988 265668 281040 265674
rect 280988 265610 281040 265616
rect 281000 264330 281028 265610
rect 281000 264302 281382 264330
rect 282196 264316 282224 269758
rect 282748 269278 282776 278038
rect 283104 275324 283156 275330
rect 283104 275266 283156 275272
rect 282920 272808 282972 272814
rect 282920 272750 282972 272756
rect 282736 269272 282788 269278
rect 282736 269214 282788 269220
rect 282932 264330 282960 272750
rect 283116 270366 283144 275266
rect 283392 274718 283420 278052
rect 284588 275738 284616 278052
rect 284576 275732 284628 275738
rect 284576 275674 284628 275680
rect 285128 275528 285180 275534
rect 285128 275470 285180 275476
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283840 270496 283892 270502
rect 283840 270438 283892 270444
rect 283104 270360 283156 270366
rect 283104 270302 283156 270308
rect 282932 264302 283038 264330
rect 283852 264316 283880 270438
rect 284668 270360 284720 270366
rect 284668 270302 284720 270308
rect 284680 264316 284708 270302
rect 285140 264330 285168 275470
rect 285692 275466 285720 278052
rect 286888 275874 286916 278052
rect 286876 275868 286928 275874
rect 286876 275810 286928 275816
rect 285680 275460 285732 275466
rect 285680 275402 285732 275408
rect 288084 275058 288112 278052
rect 288072 275052 288124 275058
rect 288072 274994 288124 275000
rect 289280 274854 289308 278052
rect 290096 275732 290148 275738
rect 290096 275674 290148 275680
rect 289268 274848 289320 274854
rect 289268 274790 289320 274796
rect 289176 274712 289228 274718
rect 289176 274654 289228 274660
rect 285864 274100 285916 274106
rect 285864 274042 285916 274048
rect 285876 264330 285904 274042
rect 286324 273080 286376 273086
rect 286324 273022 286376 273028
rect 286336 267034 286364 273022
rect 287060 271176 287112 271182
rect 287060 271118 287112 271124
rect 286324 267028 286376 267034
rect 286324 266970 286376 266976
rect 287072 264330 287100 271118
rect 288808 269272 288860 269278
rect 288808 269214 288860 269220
rect 287980 267028 288032 267034
rect 287980 266970 288032 266976
rect 285140 264302 285522 264330
rect 285876 264302 286350 264330
rect 287072 264302 287178 264330
rect 287992 264316 288020 266970
rect 288820 264316 288848 269214
rect 289188 264330 289216 274654
rect 290108 264330 290136 275674
rect 290476 275330 290504 278052
rect 291672 275670 291700 278052
rect 291844 275868 291896 275874
rect 291844 275810 291896 275816
rect 291660 275664 291712 275670
rect 291660 275606 291712 275612
rect 291292 275460 291344 275466
rect 291292 275402 291344 275408
rect 290464 275324 290516 275330
rect 290464 275266 290516 275272
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291304 264316 291332 275402
rect 291856 264330 291884 275810
rect 292868 275194 292896 278052
rect 292856 275188 292908 275194
rect 292856 275130 292908 275136
rect 292672 275052 292724 275058
rect 292672 274994 292724 275000
rect 292684 264330 292712 274994
rect 293972 274990 294000 278052
rect 294144 275324 294196 275330
rect 294144 275266 294196 275272
rect 293960 274984 294012 274990
rect 293960 274926 294012 274932
rect 293408 274848 293460 274854
rect 293408 274790 293460 274796
rect 293420 264330 293448 274790
rect 294156 264330 294184 275266
rect 295168 274854 295196 278052
rect 295340 275664 295392 275670
rect 295340 275606 295392 275612
rect 295156 274848 295208 274854
rect 295156 274790 295208 274796
rect 295352 264330 295380 275606
rect 295800 275188 295852 275194
rect 295800 275130 295852 275136
rect 295812 264330 295840 275130
rect 296364 274718 296392 278052
rect 297560 275398 297588 278052
rect 297548 275392 297600 275398
rect 297548 275334 297600 275340
rect 298756 275262 298784 278052
rect 299952 275398 299980 278052
rect 300964 278038 301070 278066
rect 302266 278038 302464 278066
rect 299572 275392 299624 275398
rect 299572 275334 299624 275340
rect 299940 275392 299992 275398
rect 299940 275334 299992 275340
rect 298744 275256 298796 275262
rect 298744 275198 298796 275204
rect 296812 274984 296864 274990
rect 296812 274926 296864 274932
rect 296352 274712 296404 274718
rect 296352 274654 296404 274660
rect 296824 264330 296852 274926
rect 297456 274848 297508 274854
rect 297456 274790 297508 274796
rect 297468 264330 297496 274790
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 298388 264330 298416 274654
rect 291856 264302 292146 264330
rect 292684 264302 292974 264330
rect 293420 264302 293802 264330
rect 294156 264302 294630 264330
rect 295352 264302 295458 264330
rect 295812 264302 296286 264330
rect 296824 264302 297114 264330
rect 297468 264302 297942 264330
rect 298388 264302 298770 264330
rect 299584 264316 299612 275334
rect 300032 275256 300084 275262
rect 300032 275198 300084 275204
rect 300044 264330 300072 275198
rect 300964 266422 300992 278038
rect 301136 275392 301188 275398
rect 301136 275334 301188 275340
rect 300952 266416 301004 266422
rect 300952 266358 301004 266364
rect 301148 264330 301176 275334
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300044 264302 300426 264330
rect 301148 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 278038
rect 303448 274718 303476 278052
rect 303724 278038 304658 278066
rect 305012 278038 305854 278066
rect 306392 278038 307050 278066
rect 307772 278038 308154 278066
rect 309152 278038 309350 278066
rect 303436 274712 303488 274718
rect 303436 274654 303488 274660
rect 303724 266422 303752 278038
rect 303988 274712 304040 274718
rect 303988 274654 304040 274660
rect 303712 266416 303764 266422
rect 303712 266358 303764 266364
rect 304000 264330 304028 274654
rect 304540 266416 304592 266422
rect 304540 266358 304592 266364
rect 302436 264302 302910 264330
rect 303738 264302 304028 264330
rect 304552 264316 304580 266358
rect 305012 264330 305040 278038
rect 306392 266370 306420 278038
rect 307772 267734 307800 278038
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266688 308732 266694
rect 308680 266630 308732 266636
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266630
rect 309152 266422 309180 278038
rect 310532 266694 310560 278052
rect 310716 278038 311742 278066
rect 311912 278038 312938 278066
rect 313292 278038 314134 278066
rect 314672 278038 315238 278066
rect 316052 278038 316434 278066
rect 317432 278038 317630 278066
rect 318826 278038 319024 278066
rect 310520 266688 310572 266694
rect 310520 266630 310572 266636
rect 310336 266552 310388 266558
rect 310336 266494 310388 266500
rect 309140 266416 309192 266422
rect 309140 266358 309192 266364
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309520 264316 309548 266358
rect 310348 264316 310376 266494
rect 310716 266422 310744 278038
rect 311912 266558 311940 278038
rect 312820 267028 312872 267034
rect 312820 266970 312872 266976
rect 311900 266552 311952 266558
rect 311900 266494 311952 266500
rect 312360 266552 312412 266558
rect 312360 266494 312412 266500
rect 310704 266416 310756 266422
rect 310704 266358 310756 266364
rect 311164 266416 311216 266422
rect 311164 266358 311216 266364
rect 311176 264316 311204 266358
rect 312372 264330 312400 266494
rect 312018 264302 312400 264330
rect 312832 264316 312860 266970
rect 313292 266422 313320 278038
rect 314476 266892 314528 266898
rect 314476 266834 314528 266840
rect 313648 266688 313700 266694
rect 313648 266630 313700 266636
rect 313280 266416 313332 266422
rect 313280 266358 313332 266364
rect 313660 264316 313688 266630
rect 314488 264316 314516 266834
rect 314672 266558 314700 278038
rect 315304 267436 315356 267442
rect 315304 267378 315356 267384
rect 314660 266552 314712 266558
rect 314660 266494 314712 266500
rect 315316 264316 315344 267378
rect 316052 267034 316080 278038
rect 316040 267028 316092 267034
rect 316040 266970 316092 266976
rect 316960 267028 317012 267034
rect 316960 266970 317012 266976
rect 316132 266552 316184 266558
rect 316132 266494 316184 266500
rect 316144 264316 316172 266494
rect 316972 264316 317000 266970
rect 317432 266694 317460 278038
rect 318708 272400 318760 272406
rect 318708 272342 318760 272348
rect 318720 267734 318748 272342
rect 318628 267706 318748 267734
rect 317420 266688 317472 266694
rect 317420 266630 317472 266636
rect 317788 266688 317840 266694
rect 317788 266630 317840 266636
rect 317800 264316 317828 266630
rect 318628 264316 318656 267706
rect 318996 266898 319024 278038
rect 319180 278038 320022 278066
rect 320192 278038 321218 278066
rect 321572 278038 322414 278066
rect 322952 278038 323518 278066
rect 319180 267442 319208 278038
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319168 267436 319220 267442
rect 319168 267378 319220 267384
rect 318984 266892 319036 266898
rect 318984 266834 319036 266840
rect 319456 264316 319484 269078
rect 320192 266558 320220 278038
rect 321192 274712 321244 274718
rect 321192 274654 321244 274660
rect 321204 267734 321232 274654
rect 321376 270768 321428 270774
rect 321376 270710 321428 270716
rect 321112 267706 321232 267734
rect 320180 266552 320232 266558
rect 320180 266494 320232 266500
rect 320272 266416 320324 266422
rect 320272 266358 320324 266364
rect 320284 264316 320312 266358
rect 321112 264316 321140 267706
rect 321388 266422 321416 270710
rect 321572 267034 321600 278038
rect 322756 273964 322808 273970
rect 322756 273906 322808 273912
rect 321928 267300 321980 267306
rect 321928 267242 321980 267248
rect 321560 267028 321612 267034
rect 321560 266970 321612 266976
rect 321376 266416 321428 266422
rect 321376 266358 321428 266364
rect 321940 264316 321968 267242
rect 322768 264316 322796 273906
rect 322952 266694 322980 278038
rect 324044 272672 324096 272678
rect 324044 272614 324096 272620
rect 322940 266688 322992 266694
rect 322940 266630 322992 266636
rect 324056 264330 324084 272614
rect 324700 272406 324728 278052
rect 325712 278038 325910 278066
rect 325332 272808 325384 272814
rect 325332 272750 325384 272756
rect 324688 272400 324740 272406
rect 324688 272342 324740 272348
rect 325344 266422 325372 272750
rect 325516 271448 325568 271454
rect 325516 271390 325568 271396
rect 324412 266416 324464 266422
rect 324412 266358 324464 266364
rect 325332 266416 325384 266422
rect 325332 266358 325384 266364
rect 323610 264302 324084 264330
rect 324424 264316 324452 266358
rect 325528 264330 325556 271390
rect 325712 269142 325740 278038
rect 326436 275324 326488 275330
rect 326436 275266 326488 275272
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 275266
rect 327092 270774 327120 278052
rect 328288 274718 328316 278052
rect 328276 274712 328328 274718
rect 328276 274654 328328 274660
rect 329484 273290 329512 278052
rect 330588 273970 330616 278052
rect 331416 278038 331798 278066
rect 330576 273964 330628 273970
rect 330576 273906 330628 273912
rect 327724 273284 327776 273290
rect 327724 273226 327776 273232
rect 329472 273284 329524 273290
rect 329472 273226 329524 273232
rect 327080 270768 327132 270774
rect 327080 270710 327132 270716
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269758
rect 327736 267306 327764 273226
rect 331416 272678 331444 278038
rect 331864 274236 331916 274242
rect 331864 274178 331916 274184
rect 331404 272672 331456 272678
rect 331404 272614 331456 272620
rect 329748 272536 329800 272542
rect 329748 272478 329800 272484
rect 329564 271312 329616 271318
rect 329564 271254 329616 271260
rect 327724 267300 327776 267306
rect 327724 267242 327776 267248
rect 327724 266552 327776 266558
rect 327724 266494 327776 266500
rect 327736 264316 327764 266494
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 328564 264316 328592 266358
rect 329576 264330 329604 271254
rect 329760 266422 329788 272478
rect 331128 271176 331180 271182
rect 331128 271118 331180 271124
rect 330208 269952 330260 269958
rect 330208 269894 330260 269900
rect 329748 266416 329800 266422
rect 329748 266358 329800 266364
rect 329406 264302 329604 264330
rect 330220 264316 330248 269894
rect 331140 267734 331168 271118
rect 331048 267706 331168 267734
rect 331048 264316 331076 267706
rect 331876 266558 331904 274178
rect 332980 272814 333008 278052
rect 333796 272944 333848 272950
rect 333796 272886 333848 272892
rect 332968 272808 333020 272814
rect 332968 272750 333020 272756
rect 332324 272672 332376 272678
rect 332324 272614 332376 272620
rect 331864 266552 331916 266558
rect 331864 266494 331916 266500
rect 332336 264330 332364 272614
rect 332692 266892 332744 266898
rect 332692 266834 332744 266840
rect 331890 264302 332364 264330
rect 332704 264316 332732 266834
rect 333808 264330 333836 272886
rect 334176 271454 334204 278052
rect 335372 275330 335400 278052
rect 335556 278038 336582 278066
rect 335360 275324 335412 275330
rect 335360 275266 335412 275272
rect 335268 273964 335320 273970
rect 335268 273906 335320 273912
rect 334164 271448 334216 271454
rect 334164 271390 334216 271396
rect 334348 270224 334400 270230
rect 334348 270166 334400 270172
rect 333546 264302 333836 264330
rect 334360 264316 334388 270166
rect 335280 267734 335308 273906
rect 335556 269822 335584 278038
rect 337764 274242 337792 278052
rect 337752 274236 337804 274242
rect 337752 274178 337804 274184
rect 337752 274100 337804 274106
rect 337752 274042 337804 274048
rect 335544 269816 335596 269822
rect 335544 269758 335596 269764
rect 336004 269816 336056 269822
rect 336004 269758 336056 269764
rect 335188 267706 335308 267734
rect 335188 264316 335216 267706
rect 336016 264316 336044 269758
rect 337764 267734 337792 274042
rect 338868 272542 338896 278052
rect 338856 272536 338908 272542
rect 338856 272478 338908 272484
rect 339224 272536 339276 272542
rect 339224 272478 339276 272484
rect 337936 271584 337988 271590
rect 337936 271526 337988 271532
rect 337672 267706 337792 267734
rect 336832 266416 336884 266422
rect 336832 266358 336884 266364
rect 336844 264316 336872 266358
rect 337672 264316 337700 267706
rect 337948 266422 337976 271526
rect 338488 268524 338540 268530
rect 338488 268466 338540 268472
rect 337936 266416 337988 266422
rect 337936 266358 337988 266364
rect 338500 264316 338528 268466
rect 339236 264330 339264 272478
rect 340064 271318 340092 278052
rect 340892 278038 341274 278066
rect 340052 271312 340104 271318
rect 340052 271254 340104 271260
rect 340604 271312 340656 271318
rect 340604 271254 340656 271260
rect 340616 264330 340644 271254
rect 340892 269958 340920 278038
rect 342456 271182 342484 278052
rect 343652 272678 343680 278052
rect 343836 278038 344862 278066
rect 343640 272672 343692 272678
rect 343640 272614 343692 272620
rect 342444 271176 342496 271182
rect 342444 271118 342496 271124
rect 343548 271176 343600 271182
rect 343548 271118 343600 271124
rect 340880 269952 340932 269958
rect 340880 269894 340932 269900
rect 341800 269952 341852 269958
rect 341800 269894 341852 269900
rect 340972 267436 341024 267442
rect 340972 267378 341024 267384
rect 339236 264302 339342 264330
rect 340170 264302 340644 264330
rect 340984 264316 341012 267378
rect 341812 264316 341840 269894
rect 343560 267734 343588 271118
rect 343468 267706 343588 267734
rect 342628 266484 342680 266490
rect 342628 266426 342680 266432
rect 342640 264316 342668 266426
rect 343468 264316 343496 267706
rect 343836 266898 343864 278038
rect 345952 272950 345980 278052
rect 346412 278038 347162 278066
rect 345940 272944 345992 272950
rect 345940 272886 345992 272892
rect 344652 272808 344704 272814
rect 344652 272750 344704 272756
rect 343824 266892 343876 266898
rect 343824 266834 343876 266840
rect 344664 264330 344692 272750
rect 346216 272672 346268 272678
rect 346216 272614 346268 272620
rect 345296 270088 345348 270094
rect 345296 270030 345348 270036
rect 345112 266620 345164 266626
rect 345112 266562 345164 266568
rect 344310 264302 344692 264330
rect 345124 264316 345152 266562
rect 345308 266490 345336 270030
rect 345296 266484 345348 266490
rect 345296 266426 345348 266432
rect 346228 264330 346256 272614
rect 346412 270230 346440 278038
rect 348344 273970 348372 278052
rect 349172 278038 349554 278066
rect 348332 273964 348384 273970
rect 348332 273906 348384 273912
rect 348424 272944 348476 272950
rect 348424 272886 348476 272892
rect 347688 271448 347740 271454
rect 347688 271390 347740 271396
rect 346400 270224 346452 270230
rect 346400 270166 346452 270172
rect 347504 266756 347556 266762
rect 347504 266698 347556 266704
rect 346768 266416 346820 266422
rect 346768 266358 346820 266364
rect 345966 264302 346256 264330
rect 346780 264316 346808 266358
rect 347516 264330 347544 266698
rect 347700 266422 347728 271390
rect 348436 266626 348464 272886
rect 349172 269822 349200 278038
rect 350356 273964 350408 273970
rect 350356 273906 350408 273912
rect 349160 269816 349212 269822
rect 349160 269758 349212 269764
rect 348792 268388 348844 268394
rect 348792 268330 348844 268336
rect 348424 266620 348476 266626
rect 348424 266562 348476 266568
rect 347688 266416 347740 266422
rect 347688 266358 347740 266364
rect 348804 264330 348832 268330
rect 350080 266552 350132 266558
rect 350080 266494 350132 266500
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 347516 264302 347622 264330
rect 348450 264302 348832 264330
rect 349264 264316 349292 266358
rect 350092 264316 350120 266494
rect 350368 266422 350396 273906
rect 350736 271590 350764 278052
rect 351932 274106 351960 278052
rect 352116 278038 353142 278066
rect 351920 274100 351972 274106
rect 351920 274042 351972 274048
rect 351184 271720 351236 271726
rect 351184 271662 351236 271668
rect 350724 271584 350776 271590
rect 350724 271526 350776 271532
rect 350908 267300 350960 267306
rect 350908 267242 350960 267248
rect 350356 266416 350408 266422
rect 350356 266358 350408 266364
rect 350920 264316 350948 267242
rect 351196 266762 351224 271662
rect 351736 269816 351788 269822
rect 351736 269758 351788 269764
rect 351184 266756 351236 266762
rect 351184 266698 351236 266704
rect 351748 264316 351776 269758
rect 352116 268530 352144 278038
rect 353944 274100 353996 274106
rect 353944 274042 353996 274048
rect 352564 268660 352616 268666
rect 352564 268602 352616 268608
rect 352104 268524 352156 268530
rect 352104 268466 352156 268472
rect 352576 264316 352604 268602
rect 353392 267572 353444 267578
rect 353392 267514 353444 267520
rect 353404 264316 353432 267514
rect 353956 266558 353984 274042
rect 354232 272542 354260 278052
rect 355152 278038 355442 278066
rect 354220 272536 354272 272542
rect 354220 272478 354272 272484
rect 354496 272536 354548 272542
rect 354496 272478 354548 272484
rect 353944 266552 353996 266558
rect 353944 266494 353996 266500
rect 354508 264330 354536 272478
rect 355152 271318 355180 278038
rect 356624 271862 356652 278052
rect 357544 278038 357834 278066
rect 358832 278038 359030 278066
rect 355324 271856 355376 271862
rect 355324 271798 355376 271804
rect 356612 271856 356664 271862
rect 356612 271798 356664 271804
rect 355140 271312 355192 271318
rect 355140 271254 355192 271260
rect 355048 270360 355100 270366
rect 355048 270302 355100 270308
rect 354246 264302 354536 264330
rect 355060 264316 355088 270302
rect 355336 267442 355364 271798
rect 357164 271312 357216 271318
rect 357164 271254 357216 271260
rect 355324 267436 355376 267442
rect 355324 267378 355376 267384
rect 355876 266552 355928 266558
rect 355876 266494 355928 266500
rect 355888 264316 355916 266494
rect 357176 264330 357204 271254
rect 357544 269958 357572 278038
rect 358636 275460 358688 275466
rect 358636 275402 358688 275408
rect 357532 269952 357584 269958
rect 357532 269894 357584 269900
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 356730 264302 357204 264330
rect 357544 264316 357572 266358
rect 358648 264330 358676 275402
rect 358832 270094 358860 278038
rect 359464 274236 359516 274242
rect 359464 274178 359516 274184
rect 358820 270088 358872 270094
rect 358820 270030 358872 270036
rect 359188 269952 359240 269958
rect 359188 269894 359240 269900
rect 358386 264302 358676 264330
rect 359200 264316 359228 269894
rect 359476 266422 359504 274178
rect 360212 271182 360240 278052
rect 361212 273080 361264 273086
rect 361212 273022 361264 273028
rect 360844 271584 360896 271590
rect 360844 271526 360896 271532
rect 360200 271176 360252 271182
rect 360200 271118 360252 271124
rect 360016 266688 360068 266694
rect 360016 266630 360068 266636
rect 359464 266416 359516 266422
rect 359464 266358 359516 266364
rect 360028 264316 360056 266630
rect 360856 266558 360884 271526
rect 360844 266552 360896 266558
rect 360844 266494 360896 266500
rect 361224 264330 361252 273022
rect 361408 272814 361436 278052
rect 362512 272950 362540 278052
rect 362776 273216 362828 273222
rect 362776 273158 362828 273164
rect 362500 272944 362552 272950
rect 362500 272886 362552 272892
rect 361396 272808 361448 272814
rect 361396 272750 361448 272756
rect 362224 272808 362276 272814
rect 362224 272750 362276 272756
rect 362236 267306 362264 272750
rect 362224 267300 362276 267306
rect 362224 267242 362276 267248
rect 362500 267164 362552 267170
rect 362500 267106 362552 267112
rect 361672 266416 361724 266422
rect 361672 266358 361724 266364
rect 360870 264302 361252 264330
rect 361684 264316 361712 266358
rect 362512 264316 362540 267106
rect 362788 266422 362816 273158
rect 363708 272678 363736 278052
rect 363880 275596 363932 275602
rect 363880 275538 363932 275544
rect 363696 272672 363748 272678
rect 363696 272614 363748 272620
rect 363892 267734 363920 275538
rect 364904 271454 364932 278052
rect 365444 272944 365496 272950
rect 365444 272886 365496 272892
rect 364892 271448 364944 271454
rect 364892 271390 364944 271396
rect 364156 271176 364208 271182
rect 364156 271118 364208 271124
rect 363800 267706 363920 267734
rect 362776 266416 362828 266422
rect 362776 266358 362828 266364
rect 363800 264330 363828 267706
rect 363354 264302 363828 264330
rect 364168 264316 364196 271118
rect 365456 264330 365484 272886
rect 366100 271726 366128 278052
rect 367112 278038 367310 278066
rect 366088 271720 366140 271726
rect 366088 271662 366140 271668
rect 366364 271448 366416 271454
rect 366364 271390 366416 271396
rect 365812 267028 365864 267034
rect 365812 266970 365864 266976
rect 365010 264302 365484 264330
rect 365824 264316 365852 266970
rect 366376 266694 366404 271390
rect 366640 270088 366692 270094
rect 366640 270030 366692 270036
rect 366364 266688 366416 266694
rect 366364 266630 366416 266636
rect 366652 264316 366680 270030
rect 367112 268394 367140 278038
rect 368492 273970 368520 278052
rect 369124 274372 369176 274378
rect 369124 274314 369176 274320
rect 368480 273964 368532 273970
rect 368480 273906 368532 273912
rect 367468 268524 367520 268530
rect 367468 268466 367520 268472
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 367480 264316 367508 268466
rect 368296 267436 368348 267442
rect 368296 267378 368348 267384
rect 368308 264316 368336 267378
rect 369136 267170 369164 274314
rect 369596 274106 369624 278052
rect 370332 278038 370806 278066
rect 371252 278038 372002 278066
rect 372632 278038 373198 278066
rect 369584 274100 369636 274106
rect 369584 274042 369636 274048
rect 370332 272814 370360 278038
rect 371056 275324 371108 275330
rect 371056 275266 371108 275272
rect 370320 272808 370372 272814
rect 370320 272750 370372 272756
rect 370504 272808 370556 272814
rect 370504 272750 370556 272756
rect 369124 267164 369176 267170
rect 369124 267106 369176 267112
rect 369952 266552 370004 266558
rect 369952 266494 370004 266500
rect 369124 266416 369176 266422
rect 369124 266358 369176 266364
rect 369136 264316 369164 266358
rect 369964 264316 369992 266494
rect 370516 266422 370544 272750
rect 370504 266416 370556 266422
rect 370504 266358 370556 266364
rect 371068 264330 371096 275266
rect 371252 269822 371280 278038
rect 372252 270224 372304 270230
rect 372252 270166 372304 270172
rect 371240 269816 371292 269822
rect 371240 269758 371292 269764
rect 371608 267300 371660 267306
rect 371608 267242 371660 267248
rect 370806 264302 371096 264330
rect 371620 264316 371648 267242
rect 372264 266558 372292 270166
rect 372632 268666 372660 278038
rect 374380 277394 374408 278052
rect 374380 277366 374500 277394
rect 373264 274100 373316 274106
rect 373264 274042 373316 274048
rect 372620 268660 372672 268666
rect 372620 268602 372672 268608
rect 372436 268388 372488 268394
rect 372436 268330 372488 268336
rect 372252 266552 372304 266558
rect 372252 266494 372304 266500
rect 372448 264316 372476 268330
rect 373276 267306 373304 274042
rect 374472 267578 374500 277366
rect 375576 272542 375604 278052
rect 376786 278038 376984 278066
rect 376116 272672 376168 272678
rect 376116 272614 376168 272620
rect 375564 272536 375616 272542
rect 375564 272478 375616 272484
rect 375288 271856 375340 271862
rect 375288 271798 375340 271804
rect 374460 267572 374512 267578
rect 374460 267514 374512 267520
rect 373264 267300 373316 267306
rect 373264 267242 373316 267248
rect 373448 267300 373500 267306
rect 373448 267242 373500 267248
rect 373264 267164 373316 267170
rect 373264 267106 373316 267112
rect 373276 264316 373304 267106
rect 373460 267034 373488 267242
rect 373448 267028 373500 267034
rect 373448 266970 373500 266976
rect 374920 266552 374972 266558
rect 374920 266494 374972 266500
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 266494
rect 375300 266422 375328 271798
rect 375288 266416 375340 266422
rect 375288 266358 375340 266364
rect 376128 264330 376156 272614
rect 376956 270366 376984 278038
rect 377680 273964 377732 273970
rect 377680 273906 377732 273912
rect 376944 270360 376996 270366
rect 376944 270302 376996 270308
rect 376576 269816 376628 269822
rect 376576 269758 376628 269764
rect 375774 264302 376156 264330
rect 376588 264316 376616 269758
rect 377692 264330 377720 273906
rect 377876 271590 377904 278052
rect 377864 271584 377916 271590
rect 377864 271526 377916 271532
rect 379072 271318 379100 278052
rect 380268 274242 380296 278052
rect 381464 275466 381492 278052
rect 382292 278038 382674 278066
rect 381452 275460 381504 275466
rect 381452 275402 381504 275408
rect 381544 274508 381596 274514
rect 381544 274450 381596 274456
rect 380256 274236 380308 274242
rect 380256 274178 380308 274184
rect 379428 272536 379480 272542
rect 379428 272478 379480 272484
rect 379060 271312 379112 271318
rect 379060 271254 379112 271260
rect 378232 266892 378284 266898
rect 378232 266834 378284 266840
rect 377430 264302 377720 264330
rect 378244 264316 378272 266834
rect 379440 264330 379468 272478
rect 380532 270360 380584 270366
rect 380532 270302 380584 270308
rect 380544 266558 380572 270302
rect 380716 267572 380768 267578
rect 380716 267514 380768 267520
rect 380532 266552 380584 266558
rect 380532 266494 380584 266500
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379468 264330
rect 379900 264316 379928 266358
rect 380728 264316 380756 267514
rect 381556 267306 381584 274450
rect 382004 271720 382056 271726
rect 382004 271662 382056 271668
rect 381544 267300 381596 267306
rect 381544 267242 381596 267248
rect 382016 264330 382044 271662
rect 382292 269958 382320 278038
rect 383856 271454 383884 278052
rect 385052 274666 385080 278052
rect 384960 274638 385080 274666
rect 385880 278038 386170 278066
rect 384960 273086 384988 274638
rect 385880 273222 385908 278038
rect 386052 275460 386104 275466
rect 386052 275402 386104 275408
rect 385868 273216 385920 273222
rect 385868 273158 385920 273164
rect 384948 273080 385000 273086
rect 384948 273022 385000 273028
rect 385684 273080 385736 273086
rect 385684 273022 385736 273028
rect 384948 272128 385000 272134
rect 384948 272070 385000 272076
rect 383844 271448 383896 271454
rect 383844 271390 383896 271396
rect 384764 271448 384816 271454
rect 384764 271390 384816 271396
rect 382280 269952 382332 269958
rect 382280 269894 382332 269900
rect 383016 269952 383068 269958
rect 383016 269894 383068 269900
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 383028 266422 383056 269894
rect 383200 267300 383252 267306
rect 383200 267242 383252 267248
rect 383016 266416 383068 266422
rect 383016 266358 383068 266364
rect 383212 264316 383240 267242
rect 384028 266416 384080 266422
rect 384028 266358 384080 266364
rect 384040 264316 384068 266358
rect 384776 264330 384804 271390
rect 384960 266422 384988 272070
rect 385696 267442 385724 273022
rect 385684 267436 385736 267442
rect 385684 267378 385736 267384
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 386064 264330 386092 275402
rect 387352 274378 387380 278052
rect 388548 275602 388576 278052
rect 388536 275596 388588 275602
rect 388536 275538 388588 275544
rect 387340 274372 387392 274378
rect 387340 274314 387392 274320
rect 388996 274236 389048 274242
rect 388996 274178 389048 274184
rect 387708 271584 387760 271590
rect 387708 271526 387760 271532
rect 387340 268796 387392 268802
rect 387340 268738 387392 268744
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 384776 264302 384882 264330
rect 385710 264302 386092 264330
rect 386524 264316 386552 266358
rect 387352 264316 387380 268738
rect 387720 266422 387748 271526
rect 388168 266756 388220 266762
rect 388168 266698 388220 266704
rect 387708 266416 387760 266422
rect 387708 266358 387760 266364
rect 388180 264316 388208 266698
rect 389008 264316 389036 274178
rect 389744 271182 389772 278052
rect 390940 272950 390968 278052
rect 392136 274514 392164 278052
rect 392124 274508 392176 274514
rect 392124 274450 392176 274456
rect 390928 272944 390980 272950
rect 390928 272886 390980 272892
rect 391848 272264 391900 272270
rect 391848 272206 391900 272212
rect 390284 271312 390336 271318
rect 390284 271254 390336 271260
rect 389732 271176 389784 271182
rect 389732 271118 389784 271124
rect 390296 264330 390324 271254
rect 390652 267708 390704 267714
rect 390652 267650 390704 267656
rect 389850 264302 390324 264330
rect 390664 264316 390692 267650
rect 391860 264330 391888 272206
rect 393332 270094 393360 278052
rect 393516 278038 394450 278066
rect 393320 270088 393372 270094
rect 393320 270030 393372 270036
rect 392032 269680 392084 269686
rect 392032 269622 392084 269628
rect 392044 267170 392072 269622
rect 393320 268660 393372 268666
rect 393320 268602 393372 268608
rect 392032 267164 392084 267170
rect 392032 267106 392084 267112
rect 393136 267028 393188 267034
rect 393136 266970 393188 266976
rect 392308 266416 392360 266422
rect 392308 266358 392360 266364
rect 391506 264302 391888 264330
rect 392320 264316 392348 266358
rect 393148 264316 393176 266970
rect 393332 266422 393360 268602
rect 393516 268530 393544 278038
rect 395632 273086 395660 278052
rect 395620 273080 395672 273086
rect 395620 273022 395672 273028
rect 396828 272814 396856 278052
rect 397472 278038 398038 278066
rect 397000 273828 397052 273834
rect 397000 273770 397052 273776
rect 396816 272808 396868 272814
rect 396816 272750 396868 272756
rect 395988 272400 396040 272406
rect 395988 272342 396040 272348
rect 394332 271176 394384 271182
rect 394332 271118 394384 271124
rect 393504 268524 393556 268530
rect 393504 268466 393556 268472
rect 393320 266416 393372 266422
rect 393320 266358 393372 266364
rect 394344 264330 394372 271118
rect 394976 270088 395028 270094
rect 394976 270030 395028 270036
rect 394792 267164 394844 267170
rect 394792 267106 394844 267112
rect 393990 264302 394372 264330
rect 394804 264316 394832 267106
rect 394988 266898 395016 270030
rect 394976 266892 395028 266898
rect 394976 266834 395028 266840
rect 396000 264330 396028 272342
rect 397012 267734 397040 273770
rect 397472 270230 397500 278038
rect 399220 275330 399248 278052
rect 399208 275324 399260 275330
rect 399208 275266 399260 275272
rect 400324 274106 400352 278052
rect 400508 278038 401534 278066
rect 401704 278038 402730 278066
rect 400312 274100 400364 274106
rect 400312 274042 400364 274048
rect 400036 273216 400088 273222
rect 400036 273158 400088 273164
rect 397460 270224 397512 270230
rect 397460 270166 397512 270172
rect 398748 270224 398800 270230
rect 398748 270166 398800 270172
rect 397276 268524 397328 268530
rect 397276 268466 397328 268472
rect 396920 267706 397040 267734
rect 396920 264330 396948 267706
rect 395646 264302 396028 264330
rect 396474 264302 396948 264330
rect 397288 264316 397316 268466
rect 398760 267578 398788 270166
rect 398748 267572 398800 267578
rect 398748 267514 398800 267520
rect 398104 267436 398156 267442
rect 398104 267378 398156 267384
rect 398116 264316 398144 267378
rect 399760 266620 399812 266626
rect 399760 266562 399812 266568
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 266562
rect 400048 266422 400076 273158
rect 400508 268394 400536 278038
rect 401508 274100 401560 274106
rect 401508 274042 401560 274048
rect 400864 270496 400916 270502
rect 400864 270438 400916 270444
rect 400496 268388 400548 268394
rect 400496 268330 400548 268336
rect 400036 266416 400088 266422
rect 400036 266358 400088 266364
rect 400876 264330 400904 270438
rect 401520 267734 401548 274042
rect 401704 269686 401732 278038
rect 403912 271862 403940 278052
rect 404372 278038 405122 278066
rect 404176 273080 404228 273086
rect 404176 273022 404228 273028
rect 403900 271856 403952 271862
rect 403900 271798 403952 271804
rect 403624 270632 403676 270638
rect 403624 270574 403676 270580
rect 401692 269680 401744 269686
rect 401692 269622 401744 269628
rect 401692 269544 401744 269550
rect 401692 269486 401744 269492
rect 400614 264302 400904 264330
rect 401428 267706 401548 267734
rect 401428 264316 401456 267706
rect 401704 267306 401732 269486
rect 402244 268388 402296 268394
rect 402244 268330 402296 268336
rect 401692 267300 401744 267306
rect 401692 267242 401744 267248
rect 402256 264316 402284 268330
rect 403072 267300 403124 267306
rect 403072 267242 403124 267248
rect 403084 264316 403112 267242
rect 403636 267170 403664 270574
rect 403624 267164 403676 267170
rect 403624 267106 403676 267112
rect 404188 264330 404216 273022
rect 404372 270366 404400 278038
rect 405556 272944 405608 272950
rect 405556 272886 405608 272892
rect 404360 270360 404412 270366
rect 404360 270302 404412 270308
rect 404360 269680 404412 269686
rect 404360 269622 404412 269628
rect 404372 266762 404400 269622
rect 404728 267572 404780 267578
rect 404728 267514 404780 267520
rect 404360 266756 404412 266762
rect 404360 266698 404412 266704
rect 403926 264302 404216 264330
rect 404740 264316 404768 267514
rect 405568 264316 405596 272886
rect 406304 272678 406332 278052
rect 407132 278038 407514 278066
rect 406844 272808 406896 272814
rect 406844 272750 406896 272756
rect 406292 272672 406344 272678
rect 406292 272614 406344 272620
rect 406856 264330 406884 272750
rect 407132 269822 407160 278038
rect 408604 273970 408632 278052
rect 408788 278038 409814 278066
rect 408592 273964 408644 273970
rect 408592 273906 408644 273912
rect 407764 270904 407816 270910
rect 407764 270846 407816 270852
rect 407120 269816 407172 269822
rect 407120 269758 407172 269764
rect 407776 266626 407804 270846
rect 408788 270094 408816 278038
rect 410800 276004 410852 276010
rect 410800 275946 410852 275952
rect 409788 274644 409840 274650
rect 409788 274586 409840 274592
rect 409604 270360 409656 270366
rect 409604 270302 409656 270308
rect 408776 270088 408828 270094
rect 408776 270030 408828 270036
rect 408408 269408 408460 269414
rect 408408 269350 408460 269356
rect 408420 267714 408448 269350
rect 408408 267708 408460 267714
rect 408408 267650 408460 267656
rect 408040 266756 408092 266762
rect 408040 266698 408092 266704
rect 407764 266620 407816 266626
rect 407764 266562 407816 266568
rect 407212 266484 407264 266490
rect 407212 266426 407264 266432
rect 406410 264302 406884 264330
rect 407224 264316 407252 266426
rect 408052 264316 408080 266698
rect 408868 266416 408920 266422
rect 408868 266358 408920 266364
rect 408880 264316 408908 266358
rect 409616 264330 409644 270302
rect 409800 266422 409828 274586
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410812 264330 410840 275946
rect 410996 272542 411024 278052
rect 411272 278038 412206 278066
rect 412652 278038 413402 278066
rect 410984 272536 411036 272542
rect 410984 272478 411036 272484
rect 411272 269958 411300 278038
rect 412272 272672 412324 272678
rect 412272 272614 412324 272620
rect 411260 269952 411312 269958
rect 411260 269894 411312 269900
rect 412284 266422 412312 272614
rect 412652 270230 412680 278038
rect 413836 274508 413888 274514
rect 413836 274450 413888 274456
rect 412640 270224 412692 270230
rect 412640 270166 412692 270172
rect 412456 270088 412508 270094
rect 412456 270030 412508 270036
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 412272 266416 412324 266422
rect 412272 266358 412324 266364
rect 409616 264302 409722 264330
rect 410550 264302 410840 264330
rect 411364 264316 411392 266358
rect 412468 264330 412496 270030
rect 413008 267164 413060 267170
rect 413008 267106 413060 267112
rect 412206 264302 412496 264330
rect 413020 264316 413048 267106
rect 413848 264316 413876 274450
rect 414584 271726 414612 278052
rect 415504 278038 415794 278066
rect 416792 278038 416898 278066
rect 414572 271720 414624 271726
rect 414572 271662 414624 271668
rect 414664 270768 414716 270774
rect 414664 270710 414716 270716
rect 414676 266626 414704 270710
rect 415032 270224 415084 270230
rect 415032 270166 415084 270172
rect 414664 266620 414716 266626
rect 414664 266562 414716 266568
rect 415044 264330 415072 270166
rect 415504 268938 415532 278038
rect 416412 275596 416464 275602
rect 416412 275538 416464 275544
rect 415492 268932 415544 268938
rect 415492 268874 415544 268880
rect 416228 268252 416280 268258
rect 416228 268194 416280 268200
rect 416240 267578 416268 268194
rect 416228 267572 416280 267578
rect 416228 267514 416280 267520
rect 416424 266422 416452 275538
rect 416596 272536 416648 272542
rect 416596 272478 416648 272484
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 414690 264302 415072 264330
rect 415504 264316 415532 266358
rect 416608 264330 416636 272478
rect 416792 269550 416820 278038
rect 418080 272134 418108 278052
rect 418804 275324 418856 275330
rect 418804 275266 418856 275272
rect 418068 272128 418120 272134
rect 418068 272070 418120 272076
rect 417424 271040 417476 271046
rect 417424 270982 417476 270988
rect 417148 269816 417200 269822
rect 417148 269758 417200 269764
rect 416780 269544 416832 269550
rect 416780 269486 416832 269492
rect 416346 264302 416636 264330
rect 417160 264316 417188 269758
rect 417436 267442 417464 270982
rect 417424 267436 417476 267442
rect 417424 267378 417476 267384
rect 418816 266422 418844 275266
rect 419080 274372 419132 274378
rect 419080 274314 419132 274320
rect 417976 266416 418028 266422
rect 417976 266358 418028 266364
rect 418804 266416 418856 266422
rect 418804 266358 418856 266364
rect 417988 264316 418016 266358
rect 419092 264330 419120 274314
rect 419276 271454 419304 278052
rect 420472 275466 420500 278052
rect 420460 275460 420512 275466
rect 420460 275402 420512 275408
rect 420552 275052 420604 275058
rect 420552 274994 420604 275000
rect 420184 271584 420236 271590
rect 420184 271526 420236 271532
rect 419264 271448 419316 271454
rect 419264 271390 419316 271396
rect 419632 269952 419684 269958
rect 419632 269894 419684 269900
rect 418830 264302 419120 264330
rect 419644 264316 419672 269894
rect 420196 267034 420224 271526
rect 420564 267734 420592 274994
rect 421668 271726 421696 278052
rect 422312 278038 422878 278066
rect 423692 278038 423982 278066
rect 422116 273964 422168 273970
rect 422116 273906 422168 273912
rect 421656 271720 421708 271726
rect 421656 271662 421708 271668
rect 420472 267706 420592 267734
rect 420184 267028 420236 267034
rect 420184 266970 420236 266976
rect 420472 264316 420500 267706
rect 421288 267572 421340 267578
rect 421288 267514 421340 267520
rect 421300 264316 421328 267514
rect 422128 264316 422156 273906
rect 422312 268802 422340 278038
rect 423692 269686 423720 278038
rect 425256 274242 425284 278052
rect 425244 274236 425296 274242
rect 425244 274178 425296 274184
rect 425704 274236 425756 274242
rect 425704 274178 425756 274184
rect 423680 269680 423732 269686
rect 423680 269622 423732 269628
rect 423956 269680 424008 269686
rect 423956 269622 424008 269628
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 422300 268116 422352 268122
rect 422300 268058 422352 268064
rect 422312 267306 422340 268058
rect 422944 267708 422996 267714
rect 422944 267650 422996 267656
rect 422300 267300 422352 267306
rect 422300 267242 422352 267248
rect 422956 264316 422984 267650
rect 423968 266762 423996 269622
rect 424600 269544 424652 269550
rect 424600 269486 424652 269492
rect 423956 266756 424008 266762
rect 423956 266698 424008 266704
rect 423772 266552 423824 266558
rect 423772 266494 423824 266500
rect 423784 264316 423812 266494
rect 424612 264316 424640 269486
rect 425716 266558 425744 274178
rect 426360 271454 426388 278052
rect 426544 278038 427570 278066
rect 426348 271448 426400 271454
rect 426348 271390 426400 271396
rect 426544 269414 426572 278038
rect 427084 275188 427136 275194
rect 427084 275130 427136 275136
rect 426532 269408 426584 269414
rect 426532 269350 426584 269356
rect 425704 266552 425756 266558
rect 425704 266494 425756 266500
rect 426256 266552 426308 266558
rect 426256 266494 426308 266500
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426268 264316 426296 266494
rect 427096 266422 427124 275130
rect 428752 272270 428780 278052
rect 429212 278038 429962 278066
rect 428740 272264 428792 272270
rect 428740 272206 428792 272212
rect 428464 272128 428516 272134
rect 428464 272070 428516 272076
rect 427452 271040 427504 271046
rect 427452 270982 427504 270988
rect 427084 266416 427136 266422
rect 427084 266358 427136 266364
rect 427464 264330 427492 270982
rect 427912 266892 427964 266898
rect 427912 266834 427964 266840
rect 427110 264302 427492 264330
rect 427924 264316 427952 266834
rect 428476 266558 428504 272070
rect 429212 268666 429240 278038
rect 430212 275868 430264 275874
rect 430212 275810 430264 275816
rect 429200 268660 429252 268666
rect 429200 268602 429252 268608
rect 428740 267436 428792 267442
rect 428740 267378 428792 267384
rect 428464 266552 428516 266558
rect 428464 266494 428516 266500
rect 428752 264316 428780 267378
rect 429568 266416 429620 266422
rect 429568 266358 429620 266364
rect 429580 264316 429608 266358
rect 430224 264330 430252 275810
rect 430396 271720 430448 271726
rect 430396 271662 430448 271668
rect 430408 266422 430436 271662
rect 431144 271590 431172 278052
rect 431684 271992 431736 271998
rect 431684 271934 431736 271940
rect 431132 271584 431184 271590
rect 431132 271526 431184 271532
rect 430396 266416 430448 266422
rect 430396 266358 430448 266364
rect 431696 264330 431724 271934
rect 432248 271318 432276 278052
rect 433156 271856 433208 271862
rect 433156 271798 433208 271804
rect 432236 271312 432288 271318
rect 432236 271254 432288 271260
rect 432880 267300 432932 267306
rect 432880 267242 432932 267248
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 430224 264302 430422 264330
rect 431250 264302 431724 264330
rect 432064 264316 432092 266358
rect 432892 264316 432920 267242
rect 433168 266422 433196 271798
rect 433444 270638 433472 278052
rect 434640 272406 434668 278052
rect 435640 275460 435692 275466
rect 435640 275402 435692 275408
rect 434628 272400 434680 272406
rect 434628 272342 434680 272348
rect 433432 270632 433484 270638
rect 433432 270574 433484 270580
rect 433708 268932 433760 268938
rect 433708 268874 433760 268880
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 433720 264316 433748 268874
rect 434536 266756 434588 266762
rect 434536 266698 434588 266704
rect 434548 264316 434576 266698
rect 435652 264330 435680 275402
rect 435836 273834 435864 278052
rect 436112 278038 437046 278066
rect 437952 278038 438242 278066
rect 435824 273828 435876 273834
rect 435824 273770 435876 273776
rect 436112 268530 436140 278038
rect 437204 271584 437256 271590
rect 437204 271526 437256 271532
rect 436560 269068 436612 269074
rect 436560 269010 436612 269016
rect 436100 268524 436152 268530
rect 436100 268466 436152 268472
rect 436572 264330 436600 269010
rect 437216 264330 437244 271526
rect 437952 271182 437980 278038
rect 438124 273828 438176 273834
rect 438124 273770 438176 273776
rect 437940 271176 437992 271182
rect 437940 271118 437992 271124
rect 438136 267714 438164 273770
rect 439332 273222 439360 278052
rect 439320 273216 439372 273222
rect 439320 273158 439372 273164
rect 439964 271448 440016 271454
rect 439964 271390 440016 271396
rect 438676 268796 438728 268802
rect 438676 268738 438728 268744
rect 438124 267708 438176 267714
rect 438124 267650 438176 267656
rect 437848 266620 437900 266626
rect 437848 266562 437900 266568
rect 435390 264302 435680 264330
rect 436218 264302 436600 264330
rect 437046 264302 437244 264330
rect 437860 264316 437888 266562
rect 438688 264316 438716 268738
rect 439976 264330 440004 271390
rect 440528 270910 440556 278052
rect 441724 277394 441752 278052
rect 441632 277366 441752 277394
rect 440884 273556 440936 273562
rect 440884 273498 440936 273504
rect 440516 270904 440568 270910
rect 440516 270846 440568 270852
rect 440896 267578 440924 273498
rect 441344 271176 441396 271182
rect 441344 271118 441396 271124
rect 441160 268660 441212 268666
rect 441160 268602 441212 268608
rect 440884 267572 440936 267578
rect 440884 267514 440936 267520
rect 440332 266416 440384 266422
rect 440332 266358 440384 266364
rect 439530 264302 440004 264330
rect 440344 264316 440372 266358
rect 441172 264316 441200 268602
rect 441356 266422 441384 271118
rect 441632 270502 441660 277366
rect 442920 274106 442948 278052
rect 443104 278038 444130 278066
rect 444392 278038 445326 278066
rect 442908 274100 442960 274106
rect 442908 274042 442960 274048
rect 442908 271312 442960 271318
rect 442908 271254 442960 271260
rect 441620 270496 441672 270502
rect 441620 270438 441672 270444
rect 441620 269408 441672 269414
rect 441620 269350 441672 269356
rect 441632 267170 441660 269350
rect 441620 267164 441672 267170
rect 441620 267106 441672 267112
rect 442724 266892 442776 266898
rect 442724 266834 442776 266840
rect 441344 266416 441396 266422
rect 441344 266358 441396 266364
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 266834
rect 442920 266422 442948 271254
rect 443104 268394 443132 278038
rect 444012 273216 444064 273222
rect 444012 273158 444064 273164
rect 443092 268388 443144 268394
rect 443092 268330 443144 268336
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 444024 264330 444052 273158
rect 444392 268122 444420 278038
rect 445024 275732 445076 275738
rect 445024 275674 445076 275680
rect 445036 271182 445064 275674
rect 446508 273086 446536 278052
rect 447152 278038 447626 278066
rect 446496 273080 446548 273086
rect 446496 273022 446548 273028
rect 446864 272400 446916 272406
rect 446864 272342 446916 272348
rect 445024 271176 445076 271182
rect 445024 271118 445076 271124
rect 445668 271176 445720 271182
rect 445668 271118 445720 271124
rect 444380 268116 444432 268122
rect 444380 268058 444432 268064
rect 445300 267708 445352 267714
rect 445300 267650 445352 267656
rect 444472 266416 444524 266422
rect 444472 266358 444524 266364
rect 442736 264302 442842 264330
rect 443670 264302 444052 264330
rect 444484 264316 444512 266358
rect 445312 264316 445340 267650
rect 445680 266422 445708 271118
rect 446128 268524 446180 268530
rect 446128 268466 446180 268472
rect 445668 266416 445720 266422
rect 445668 266358 445720 266364
rect 446140 264316 446168 268466
rect 446876 264330 446904 272342
rect 447152 268258 447180 278038
rect 447784 273692 447836 273698
rect 447784 273634 447836 273640
rect 447140 268252 447192 268258
rect 447140 268194 447192 268200
rect 447796 267442 447824 273634
rect 448808 272950 448836 278052
rect 448796 272944 448848 272950
rect 448796 272886 448848 272892
rect 450004 272814 450032 278052
rect 450832 278038 451214 278066
rect 451384 278038 452410 278066
rect 449992 272808 450044 272814
rect 449992 272750 450044 272756
rect 450544 272808 450596 272814
rect 450544 272750 450596 272756
rect 449716 272264 449768 272270
rect 449716 272206 449768 272212
rect 449164 270904 449216 270910
rect 449164 270846 449216 270852
rect 448428 268116 448480 268122
rect 448428 268058 448480 268064
rect 447784 267436 447836 267442
rect 447784 267378 447836 267384
rect 448440 267170 448468 268058
rect 447140 267164 447192 267170
rect 447140 267106 447192 267112
rect 448428 267164 448480 267170
rect 448428 267106 448480 267112
rect 447152 266626 447180 267106
rect 449176 266762 449204 270846
rect 449164 266756 449216 266762
rect 449164 266698 449216 266704
rect 447140 266620 447192 266626
rect 447140 266562 447192 266568
rect 447784 266552 447836 266558
rect 447784 266494 447836 266500
rect 446876 264302 446982 264330
rect 447796 264316 447824 266494
rect 448612 266416 448664 266422
rect 448612 266358 448664 266364
rect 448624 264316 448652 266358
rect 449728 264330 449756 272206
rect 450268 267572 450320 267578
rect 450268 267514 450320 267520
rect 449466 264302 449756 264330
rect 450280 264316 450308 267514
rect 450556 266422 450584 272750
rect 450832 270774 450860 278038
rect 451188 274100 451240 274106
rect 451188 274042 451240 274048
rect 450820 270768 450872 270774
rect 450820 270710 450872 270716
rect 451200 267734 451228 274042
rect 451384 269686 451412 278038
rect 453592 274650 453620 278052
rect 454328 278038 454710 278066
rect 453580 274644 453632 274650
rect 453580 274586 453632 274592
rect 452292 273080 452344 273086
rect 452292 273022 452344 273028
rect 451372 269680 451424 269686
rect 451372 269622 451424 269628
rect 451108 267706 451228 267734
rect 450544 266416 450596 266422
rect 450544 266358 450596 266364
rect 451108 264316 451136 267706
rect 452304 264330 452332 273022
rect 453304 270632 453356 270638
rect 453304 270574 453356 270580
rect 453316 267306 453344 270574
rect 454328 270366 454356 278038
rect 455892 276010 455920 278052
rect 455880 276004 455932 276010
rect 455880 275946 455932 275952
rect 456064 276004 456116 276010
rect 456064 275946 456116 275952
rect 455328 272944 455380 272950
rect 455328 272886 455380 272892
rect 454316 270360 454368 270366
rect 454316 270302 454368 270308
rect 453580 269680 453632 269686
rect 453580 269622 453632 269628
rect 453304 267300 453356 267306
rect 453304 267242 453356 267248
rect 452752 267164 452804 267170
rect 452752 267106 452804 267112
rect 451950 264302 452332 264330
rect 452764 264316 452792 267106
rect 453592 264316 453620 269622
rect 455144 267164 455196 267170
rect 455144 267106 455196 267112
rect 454408 266416 454460 266422
rect 454408 266358 454460 266364
rect 454420 264316 454448 266358
rect 455156 264330 455184 267106
rect 455340 266422 455368 272886
rect 456076 266558 456104 275946
rect 457088 272678 457116 278052
rect 457444 274644 457496 274650
rect 457444 274586 457496 274592
rect 457076 272672 457128 272678
rect 457076 272614 457128 272620
rect 457260 272672 457312 272678
rect 457260 272614 457312 272620
rect 456432 270496 456484 270502
rect 456432 270438 456484 270444
rect 456064 266552 456116 266558
rect 456064 266494 456116 266500
rect 455328 266416 455380 266422
rect 455328 266358 455380 266364
rect 456444 264330 456472 270438
rect 457272 264330 457300 272614
rect 457456 267034 457484 274586
rect 458284 270094 458312 278052
rect 458468 278038 459494 278066
rect 458272 270088 458324 270094
rect 458272 270030 458324 270036
rect 458468 269414 458496 278038
rect 460676 274514 460704 278052
rect 460952 278038 461886 278066
rect 460664 274508 460716 274514
rect 460664 274450 460716 274456
rect 460572 273352 460624 273358
rect 460572 273294 460624 273300
rect 460584 272950 460612 273294
rect 460572 272944 460624 272950
rect 460572 272886 460624 272892
rect 459376 272672 459428 272678
rect 459374 272640 459376 272649
rect 459560 272672 459612 272678
rect 459428 272640 459430 272649
rect 459560 272614 459612 272620
rect 459374 272575 459430 272584
rect 458824 270360 458876 270366
rect 458824 270302 458876 270308
rect 458456 269408 458508 269414
rect 458456 269350 458508 269356
rect 457444 267028 457496 267034
rect 457444 266970 457496 266976
rect 457720 266756 457772 266762
rect 457720 266698 457772 266704
rect 455156 264302 455262 264330
rect 456090 264302 456472 264330
rect 456918 264302 457300 264330
rect 457732 264316 457760 266698
rect 458836 264330 458864 270302
rect 459572 267730 459600 272614
rect 460952 270230 460980 278038
rect 462976 275602 463004 278052
rect 463896 278038 464186 278066
rect 465092 278038 465382 278066
rect 462964 275596 463016 275602
rect 462964 275538 463016 275544
rect 463148 275596 463200 275602
rect 463148 275538 463200 275544
rect 463160 274666 463188 275538
rect 462976 274638 463188 274666
rect 461400 273352 461452 273358
rect 461400 273294 461452 273300
rect 461412 273170 461440 273294
rect 461412 273142 461808 273170
rect 461780 273086 461808 273142
rect 461768 273080 461820 273086
rect 461768 273022 461820 273028
rect 460940 270224 460992 270230
rect 460940 270166 460992 270172
rect 461400 270224 461452 270230
rect 461400 270166 461452 270172
rect 458574 264302 458864 264330
rect 459388 267702 459600 267730
rect 459388 264316 459416 267702
rect 460204 267436 460256 267442
rect 460204 267378 460256 267384
rect 460216 264316 460244 267378
rect 461412 264330 461440 270166
rect 461860 268388 461912 268394
rect 461860 268330 461912 268336
rect 461058 264302 461440 264330
rect 461872 264316 461900 268330
rect 462976 267306 463004 274638
rect 463240 274508 463292 274514
rect 463240 274450 463292 274456
rect 463252 273254 463280 274450
rect 463160 273226 463280 273254
rect 462964 267300 463016 267306
rect 462964 267242 463016 267248
rect 463160 264330 463188 273226
rect 463896 272542 463924 278038
rect 463884 272536 463936 272542
rect 463884 272478 463936 272484
rect 464710 272368 464766 272377
rect 464710 272303 464766 272312
rect 463516 270088 463568 270094
rect 463516 270030 463568 270036
rect 462714 264302 463188 264330
rect 463528 264316 463556 270030
rect 464724 264330 464752 272303
rect 465092 269822 465120 278038
rect 466564 275330 466592 278052
rect 466552 275324 466604 275330
rect 466552 275266 466604 275272
rect 467564 275324 467616 275330
rect 467564 275266 467616 275272
rect 466414 272672 466466 272678
rect 466090 272640 466146 272649
rect 466146 272620 466414 272626
rect 466146 272614 466466 272620
rect 466146 272598 466454 272614
rect 466090 272575 466146 272584
rect 465080 269816 465132 269822
rect 465080 269758 465132 269764
rect 466000 269816 466052 269822
rect 466000 269758 466052 269764
rect 465172 267300 465224 267306
rect 465172 267242 465224 267248
rect 464370 264302 464752 264330
rect 465184 264316 465212 267242
rect 466012 264316 466040 269758
rect 466828 265124 466880 265130
rect 466828 265066 466880 265072
rect 466840 264316 466868 265066
rect 467576 264330 467604 275266
rect 467760 274378 467788 278052
rect 468128 278038 468970 278066
rect 467748 274372 467800 274378
rect 467748 274314 467800 274320
rect 468128 269958 468156 278038
rect 470152 275058 470180 278052
rect 470140 275052 470192 275058
rect 470140 274994 470192 275000
rect 471256 273562 471284 278052
rect 471612 276276 471664 276282
rect 471612 276218 471664 276224
rect 471244 273556 471296 273562
rect 471244 273498 471296 273504
rect 470554 272536 470606 272542
rect 470692 272536 470744 272542
rect 470554 272478 470606 272484
rect 470690 272504 470692 272513
rect 470744 272504 470746 272513
rect 470566 272354 470594 272478
rect 470690 272439 470746 272448
rect 470566 272326 470640 272354
rect 470612 272218 470640 272326
rect 470612 272190 470824 272218
rect 470796 272134 470824 272190
rect 470554 272128 470606 272134
rect 470784 272128 470836 272134
rect 470606 272076 470640 272082
rect 470554 272070 470640 272076
rect 470784 272070 470836 272076
rect 470566 272054 470640 272070
rect 470612 271969 470640 272054
rect 470598 271960 470654 271969
rect 470598 271895 470654 271904
rect 468116 269952 468168 269958
rect 468116 269894 468168 269900
rect 468484 269952 468536 269958
rect 468484 269894 468536 269900
rect 467576 264302 467682 264330
rect 468496 264316 468524 269894
rect 470968 269408 471020 269414
rect 470968 269350 471020 269356
rect 470140 267028 470192 267034
rect 470140 266970 470192 266976
rect 469312 265260 469364 265266
rect 469312 265202 469364 265208
rect 469324 264316 469352 265202
rect 470152 264316 470180 266970
rect 470980 264316 471008 269350
rect 471624 264330 471652 276218
rect 472452 273970 472480 278052
rect 473084 274916 473136 274922
rect 473084 274858 473136 274864
rect 472440 273964 472492 273970
rect 472440 273906 472492 273912
rect 473096 264330 473124 274858
rect 473648 273834 473676 278052
rect 474844 274242 474872 278052
rect 475028 278038 476054 278066
rect 474832 274236 474884 274242
rect 474832 274178 474884 274184
rect 474648 273964 474700 273970
rect 474648 273906 474700 273912
rect 473636 273828 473688 273834
rect 473636 273770 473688 273776
rect 474280 269272 474332 269278
rect 474280 269214 474332 269220
rect 473452 266416 473504 266422
rect 473452 266358 473504 266364
rect 471624 264302 471822 264330
rect 472650 264302 473124 264330
rect 473464 264316 473492 266358
rect 474292 264316 474320 269214
rect 474660 266422 474688 273906
rect 475028 269550 475056 278038
rect 477040 276412 477092 276418
rect 477040 276354 477092 276360
rect 476764 274780 476816 274786
rect 476764 274722 476816 274728
rect 476028 273556 476080 273562
rect 476028 273498 476080 273504
rect 475016 269544 475068 269550
rect 475016 269486 475068 269492
rect 476040 267734 476068 273498
rect 475948 267706 476068 267734
rect 474648 266416 474700 266422
rect 474648 266358 474700 266364
rect 475108 266416 475160 266422
rect 475108 266358 475160 266364
rect 475120 264316 475148 266358
rect 475948 264316 475976 267706
rect 476776 266762 476804 274722
rect 476764 266756 476816 266762
rect 476764 266698 476816 266704
rect 477052 264330 477080 276354
rect 477236 275194 477264 278052
rect 478064 278038 478354 278066
rect 479168 278038 479550 278066
rect 477224 275188 477276 275194
rect 477224 275130 477276 275136
rect 478064 271969 478092 278038
rect 478696 273420 478748 273426
rect 478696 273362 478748 273368
rect 478050 271960 478106 271969
rect 478050 271895 478106 271904
rect 477592 265396 477644 265402
rect 477592 265338 477644 265344
rect 476790 264302 477080 264330
rect 477604 264316 477632 265338
rect 478708 264330 478736 273362
rect 479168 271046 479196 278038
rect 479984 277364 480036 277370
rect 479984 277306 480036 277312
rect 479522 271960 479578 271969
rect 479522 271895 479578 271904
rect 479156 271040 479208 271046
rect 479156 270982 479208 270988
rect 479536 266422 479564 271895
rect 479524 266416 479576 266422
rect 479524 266358 479576 266364
rect 479248 265532 479300 265538
rect 479248 265474 479300 265480
rect 478446 264302 478736 264330
rect 479260 264316 479288 265474
rect 479996 264330 480024 277306
rect 480732 274650 480760 278052
rect 480720 274644 480772 274650
rect 480720 274586 480772 274592
rect 481364 273828 481416 273834
rect 481364 273770 481416 273776
rect 480168 271856 480220 271862
rect 480220 271804 480300 271810
rect 480168 271798 480300 271804
rect 480180 271782 480300 271798
rect 480272 270774 480300 271782
rect 480260 270768 480312 270774
rect 480260 270710 480312 270716
rect 481376 264330 481404 273770
rect 481928 273698 481956 278052
rect 483124 277394 483152 278052
rect 483124 277366 483244 277394
rect 482836 276548 482888 276554
rect 482836 276490 482888 276496
rect 481916 273692 481968 273698
rect 481916 273634 481968 273640
rect 482848 266422 482876 276490
rect 483020 272128 483072 272134
rect 483020 272070 483072 272076
rect 483032 271969 483060 272070
rect 483018 271960 483074 271969
rect 483018 271895 483074 271904
rect 483216 271726 483244 277366
rect 484320 275874 484348 278052
rect 484872 278038 485530 278066
rect 484308 275868 484360 275874
rect 484308 275810 484360 275816
rect 484308 275052 484360 275058
rect 484308 274994 484360 275000
rect 484320 274514 484348 274994
rect 484308 274508 484360 274514
rect 484308 274450 484360 274456
rect 484216 273692 484268 273698
rect 484216 273634 484268 273640
rect 483204 271720 483256 271726
rect 483204 271662 483256 271668
rect 484228 266422 484256 273634
rect 484872 271862 484900 278038
rect 485044 275460 485096 275466
rect 485044 275402 485096 275408
rect 485228 275460 485280 275466
rect 485228 275402 485280 275408
rect 485056 275194 485084 275402
rect 485044 275188 485096 275194
rect 485044 275130 485096 275136
rect 485240 275058 485268 275402
rect 485228 275052 485280 275058
rect 485228 274994 485280 275000
rect 484860 271856 484912 271862
rect 484860 271798 484912 271804
rect 485044 271040 485096 271046
rect 485044 270982 485096 270988
rect 485056 266898 485084 270982
rect 486620 270774 486648 278052
rect 486792 274644 486844 274650
rect 486792 274586 486844 274592
rect 486608 270768 486660 270774
rect 486608 270710 486660 270716
rect 485044 266892 485096 266898
rect 485044 266834 485096 266840
rect 485044 266756 485096 266762
rect 485044 266698 485096 266704
rect 481732 266416 481784 266422
rect 481732 266358 481784 266364
rect 482836 266416 482888 266422
rect 482836 266358 482888 266364
rect 483388 266416 483440 266422
rect 483388 266358 483440 266364
rect 484216 266416 484268 266422
rect 484216 266358 484268 266364
rect 479996 264302 480102 264330
rect 480930 264302 481404 264330
rect 481744 264316 481772 266358
rect 482560 266076 482612 266082
rect 482560 266018 482612 266024
rect 482572 264316 482600 266018
rect 483400 264316 483428 266358
rect 484216 266212 484268 266218
rect 484216 266154 484268 266160
rect 484228 264316 484256 266154
rect 485056 264316 485084 266698
rect 486804 266422 486832 274586
rect 486976 270768 487028 270774
rect 486976 270710 487028 270716
rect 485872 266416 485924 266422
rect 485872 266358 485924 266364
rect 486792 266416 486844 266422
rect 486792 266358 486844 266364
rect 485884 264316 485912 266358
rect 486988 264330 487016 270710
rect 487816 270638 487844 278052
rect 488552 278038 489026 278066
rect 487988 277228 488040 277234
rect 487988 277170 488040 277176
rect 487804 270632 487856 270638
rect 487804 270574 487856 270580
rect 487160 266348 487212 266354
rect 487160 266290 487212 266296
rect 487172 266082 487200 266290
rect 487160 266076 487212 266082
rect 487160 266018 487212 266024
rect 488000 264330 488028 277170
rect 488356 274508 488408 274514
rect 488356 274450 488408 274456
rect 486726 264302 487016 264330
rect 487554 264302 488028 264330
rect 488368 264316 488396 274450
rect 488552 268938 488580 278038
rect 490208 270910 490236 278052
rect 490564 275868 490616 275874
rect 490564 275810 490616 275816
rect 490196 270904 490248 270910
rect 490196 270846 490248 270852
rect 489644 270632 489696 270638
rect 489644 270574 489696 270580
rect 488540 268932 488592 268938
rect 488540 268874 488592 268880
rect 489656 264330 489684 270574
rect 490576 267714 490604 275810
rect 491404 275194 491432 278052
rect 491680 278038 492614 278066
rect 491392 275188 491444 275194
rect 491392 275130 491444 275136
rect 491680 269074 491708 278038
rect 493704 271590 493732 278052
rect 494072 278038 494914 278066
rect 495452 278038 496110 278066
rect 493692 271584 493744 271590
rect 493692 271526 493744 271532
rect 492588 270904 492640 270910
rect 492588 270846 492640 270852
rect 491668 269068 491720 269074
rect 491668 269010 491720 269016
rect 490840 267980 490892 267986
rect 490840 267922 490892 267928
rect 490564 267708 490616 267714
rect 490564 267650 490616 267656
rect 490012 266756 490064 266762
rect 490012 266698 490064 266704
rect 489210 264302 489684 264330
rect 490024 264316 490052 266698
rect 490852 264316 490880 267922
rect 492600 266490 492628 270846
rect 493324 268252 493376 268258
rect 493324 268194 493376 268200
rect 491668 266484 491720 266490
rect 491668 266426 491720 266432
rect 492588 266484 492640 266490
rect 492588 266426 492640 266432
rect 491680 264316 491708 266426
rect 492496 266076 492548 266082
rect 492496 266018 492548 266024
rect 492508 264316 492536 266018
rect 493336 264316 493364 268194
rect 494072 268122 494100 278038
rect 494704 271856 494756 271862
rect 494704 271798 494756 271804
rect 494716 271046 494744 271798
rect 494704 271040 494756 271046
rect 494704 270982 494756 270988
rect 495072 271040 495124 271046
rect 495072 270982 495124 270988
rect 494060 268116 494112 268122
rect 494060 268058 494112 268064
rect 495084 266490 495112 270982
rect 495256 269544 495308 269550
rect 495256 269486 495308 269492
rect 494152 266484 494204 266490
rect 494152 266426 494204 266432
rect 495072 266484 495124 266490
rect 495072 266426 495124 266432
rect 494164 264316 494192 266426
rect 495268 264330 495296 269486
rect 495452 268802 495480 278038
rect 497292 271590 497320 278052
rect 497924 277092 497976 277098
rect 497924 277034 497976 277040
rect 497280 271584 497332 271590
rect 497280 271526 497332 271532
rect 496544 271448 496596 271454
rect 496544 271390 496596 271396
rect 495808 269068 495860 269074
rect 495808 269010 495860 269016
rect 495440 268796 495492 268802
rect 495440 268738 495492 268744
rect 495006 264302 495296 264330
rect 495820 264316 495848 269010
rect 496556 264330 496584 271390
rect 497936 264330 497964 277034
rect 498488 275738 498516 278052
rect 499684 277394 499712 278052
rect 499592 277366 499712 277394
rect 500696 278038 500894 278066
rect 501432 278038 501998 278066
rect 498476 275732 498528 275738
rect 498476 275674 498528 275680
rect 498844 275732 498896 275738
rect 498844 275674 498896 275680
rect 498292 268932 498344 268938
rect 498292 268874 498344 268880
rect 496556 264302 496662 264330
rect 497490 264302 497964 264330
rect 498304 264316 498332 268874
rect 498856 267578 498884 275674
rect 499304 271720 499356 271726
rect 499304 271662 499356 271668
rect 498844 267572 498896 267578
rect 498844 267514 498896 267520
rect 499316 264330 499344 271662
rect 499592 268666 499620 277366
rect 500696 271318 500724 278038
rect 501052 272808 501104 272814
rect 501052 272750 501104 272756
rect 501064 272406 501092 272750
rect 500868 272400 500920 272406
rect 500868 272342 500920 272348
rect 501052 272400 501104 272406
rect 501052 272342 501104 272348
rect 500880 272241 500908 272342
rect 500866 272232 500922 272241
rect 500866 272167 500922 272176
rect 501432 271862 501460 278038
rect 503180 273222 503208 278052
rect 504008 278038 504390 278066
rect 503444 275052 503496 275058
rect 503444 274994 503496 275000
rect 503168 273216 503220 273222
rect 503168 273158 503220 273164
rect 501602 271960 501658 271969
rect 501602 271895 501658 271904
rect 501420 271856 501472 271862
rect 501420 271798 501472 271804
rect 500684 271312 500736 271318
rect 500684 271254 500736 271260
rect 500776 268796 500828 268802
rect 500776 268738 500828 268744
rect 499580 268660 499632 268666
rect 499580 268602 499632 268608
rect 499948 266892 500000 266898
rect 499948 266834 500000 266840
rect 499146 264302 499344 264330
rect 499960 264316 499988 266834
rect 500788 264316 500816 268738
rect 501616 266626 501644 271895
rect 501972 271584 502024 271590
rect 501972 271526 502024 271532
rect 501604 266620 501656 266626
rect 501604 266562 501656 266568
rect 501984 264330 502012 271526
rect 503260 268660 503312 268666
rect 503260 268602 503312 268608
rect 502432 266484 502484 266490
rect 502432 266426 502484 266432
rect 501630 264302 502012 264330
rect 502444 264316 502472 266426
rect 503272 264316 503300 268602
rect 503456 266490 503484 274994
rect 504008 271182 504036 278038
rect 505572 275874 505600 278052
rect 506492 278038 506782 278066
rect 505560 275868 505612 275874
rect 505560 275810 505612 275816
rect 506204 274372 506256 274378
rect 506204 274314 506256 274320
rect 504180 273216 504232 273222
rect 504180 273158 504232 273164
rect 504192 272270 504220 273158
rect 504364 272808 504416 272814
rect 504364 272750 504416 272756
rect 504180 272264 504232 272270
rect 504180 272206 504232 272212
rect 504376 271998 504404 272750
rect 504548 272264 504600 272270
rect 504546 272232 504548 272241
rect 504600 272232 504602 272241
rect 504546 272167 504602 272176
rect 504364 271992 504416 271998
rect 504548 271992 504600 271998
rect 504364 271934 504416 271940
rect 504546 271960 504548 271969
rect 504600 271960 504602 271969
rect 504546 271895 504602 271904
rect 504364 271856 504416 271862
rect 504364 271798 504416 271804
rect 504376 271454 504404 271798
rect 504364 271448 504416 271454
rect 504364 271390 504416 271396
rect 505008 271448 505060 271454
rect 505008 271390 505060 271396
rect 503996 271176 504048 271182
rect 503996 271118 504048 271124
rect 504824 266620 504876 266626
rect 504824 266562 504876 266568
rect 503444 266484 503496 266490
rect 503444 266426 503496 266432
rect 504088 266484 504140 266490
rect 504088 266426 504140 266432
rect 504100 264316 504128 266426
rect 504836 264330 504864 266562
rect 505020 266490 505048 271390
rect 505008 266484 505060 266490
rect 505008 266426 505060 266432
rect 506216 264330 506244 274314
rect 506492 268530 506520 278038
rect 507492 275188 507544 275194
rect 507492 275130 507544 275136
rect 506480 268524 506532 268530
rect 506480 268466 506532 268472
rect 507504 267734 507532 275130
rect 507964 272270 507992 278052
rect 509068 276010 509096 278052
rect 509712 278038 510278 278066
rect 509056 276004 509108 276010
rect 509056 275946 509108 275952
rect 509712 272406 509740 278038
rect 511460 273222 511488 278052
rect 511632 276956 511684 276962
rect 511632 276898 511684 276904
rect 511448 273216 511500 273222
rect 511448 273158 511500 273164
rect 509700 272400 509752 272406
rect 509700 272342 509752 272348
rect 507952 272264 508004 272270
rect 507952 272206 508004 272212
rect 509700 272264 509752 272270
rect 509700 272206 509752 272212
rect 507676 271312 507728 271318
rect 507676 271254 507728 271260
rect 507412 267706 507532 267734
rect 506572 266484 506624 266490
rect 506572 266426 506624 266432
rect 504836 264302 504942 264330
rect 505770 264302 506244 264330
rect 506584 264316 506612 266426
rect 507412 264316 507440 267706
rect 507688 266490 507716 271254
rect 509238 269920 509294 269929
rect 509238 269855 509294 269864
rect 509252 269686 509280 269855
rect 509240 269680 509292 269686
rect 509240 269622 509292 269628
rect 509146 269512 509202 269521
rect 509146 269447 509202 269456
rect 508228 268524 508280 268530
rect 508228 268466 508280 268472
rect 507860 266892 507912 266898
rect 507860 266834 507912 266840
rect 507872 266490 507900 266834
rect 507676 266484 507728 266490
rect 507676 266426 507728 266432
rect 507860 266484 507912 266490
rect 507860 266426 507912 266432
rect 508240 264316 508268 268466
rect 509160 267734 509188 269447
rect 509068 267706 509188 267734
rect 509068 264316 509096 267706
rect 509712 266762 509740 272206
rect 509884 269544 509936 269550
rect 509882 269512 509884 269521
rect 509936 269512 509938 269521
rect 509882 269447 509938 269456
rect 511644 267734 511672 276898
rect 512656 275738 512684 278052
rect 513196 276004 513248 276010
rect 513196 275946 513248 275952
rect 512644 275732 512696 275738
rect 512644 275674 512696 275680
rect 511816 274236 511868 274242
rect 511816 274178 511868 274184
rect 509884 267708 509936 267714
rect 509884 267650 509936 267656
rect 511552 267706 511672 267734
rect 509700 266756 509752 266762
rect 509700 266698 509752 266704
rect 509896 264316 509924 267650
rect 510712 266756 510764 266762
rect 510712 266698 510764 266704
rect 510724 264316 510752 266698
rect 511552 264316 511580 267706
rect 511828 266762 511856 274178
rect 513208 266762 513236 275946
rect 513852 274106 513880 278052
rect 514484 276820 514536 276826
rect 514484 276762 514536 276768
rect 513840 274100 513892 274106
rect 513840 274042 513892 274048
rect 514208 272808 514260 272814
rect 514208 272750 514260 272756
rect 514220 272270 514248 272750
rect 514208 272264 514260 272270
rect 514208 272206 514260 272212
rect 511816 266756 511868 266762
rect 511816 266698 511868 266704
rect 512368 266756 512420 266762
rect 512368 266698 512420 266704
rect 513196 266756 513248 266762
rect 513196 266698 513248 266704
rect 512380 264316 512408 266698
rect 513196 265940 513248 265946
rect 513196 265882 513248 265888
rect 513208 264316 513236 265882
rect 514496 264330 514524 276762
rect 515048 273086 515076 278052
rect 516244 275602 516272 278052
rect 516520 278038 517362 278066
rect 516232 275596 516284 275602
rect 516232 275538 516284 275544
rect 515036 273080 515088 273086
rect 515036 273022 515088 273028
rect 515404 273080 515456 273086
rect 515404 273022 515456 273028
rect 514852 267572 514904 267578
rect 514852 267514 514904 267520
rect 514050 264302 514524 264330
rect 514864 264316 514892 267514
rect 515416 267170 515444 273022
rect 516520 269929 516548 278038
rect 516784 275596 516836 275602
rect 516784 275538 516836 275544
rect 516506 269920 516562 269929
rect 516506 269855 516562 269864
rect 516796 267442 516824 275538
rect 518544 273222 518572 278052
rect 518716 276684 518768 276690
rect 518716 276626 518768 276632
rect 518532 273216 518584 273222
rect 518532 273158 518584 273164
rect 517428 272400 517480 272406
rect 517428 272342 517480 272348
rect 516784 267436 516836 267442
rect 516784 267378 516836 267384
rect 515404 267164 515456 267170
rect 515404 267106 515456 267112
rect 517244 267164 517296 267170
rect 517244 267106 517296 267112
rect 516508 266756 516560 266762
rect 516508 266698 516560 266704
rect 515680 265804 515732 265810
rect 515680 265746 515732 265752
rect 515692 264316 515720 265746
rect 516520 264316 516548 266698
rect 517256 264330 517284 267106
rect 517440 266762 517468 272342
rect 518728 267734 518756 276626
rect 519740 273222 519768 278052
rect 520292 278038 520950 278066
rect 519728 273216 519780 273222
rect 519728 273158 519780 273164
rect 520096 272264 520148 272270
rect 520096 272206 520148 272212
rect 518544 267706 518756 267734
rect 517428 266756 517480 266762
rect 517428 266698 517480 266704
rect 518544 264330 518572 267706
rect 519820 267436 519872 267442
rect 519820 267378 519872 267384
rect 518992 266756 519044 266762
rect 518992 266698 519044 266704
rect 517256 264302 517362 264330
rect 518190 264302 518572 264330
rect 519004 264316 519032 266698
rect 519832 264316 519860 267378
rect 520108 266762 520136 272206
rect 520292 270502 520320 278038
rect 521476 273216 521528 273222
rect 521476 273158 521528 273164
rect 520280 270496 520332 270502
rect 520280 270438 520332 270444
rect 520096 266756 520148 266762
rect 520096 266698 520148 266704
rect 520648 265668 520700 265674
rect 520648 265610 520700 265616
rect 520660 264316 520688 265610
rect 521488 264316 521516 273158
rect 522132 272678 522160 278052
rect 522764 275868 522816 275874
rect 522764 275810 522816 275816
rect 522120 272672 522172 272678
rect 522120 272614 522172 272620
rect 522776 264330 522804 275810
rect 523328 274786 523356 278052
rect 524432 278038 524538 278066
rect 523316 274780 523368 274786
rect 523316 274722 523368 274728
rect 523684 274780 523736 274786
rect 523684 274722 523736 274728
rect 523132 270496 523184 270502
rect 523132 270438 523184 270444
rect 522330 264302 522804 264330
rect 523144 264316 523172 270438
rect 523696 267306 523724 274722
rect 524052 271176 524104 271182
rect 524052 271118 524104 271124
rect 524064 267734 524092 271118
rect 524432 270366 524460 278038
rect 525628 272950 525656 278052
rect 526824 275602 526852 278052
rect 527192 278038 528034 278066
rect 528572 278038 529230 278066
rect 526812 275596 526864 275602
rect 526812 275538 526864 275544
rect 526812 273080 526864 273086
rect 526812 273022 526864 273028
rect 525616 272944 525668 272950
rect 525616 272886 525668 272892
rect 524420 270360 524472 270366
rect 524420 270302 524472 270308
rect 525616 270360 525668 270366
rect 525616 270302 525668 270308
rect 523972 267706 524092 267734
rect 523684 267300 523736 267306
rect 523684 267242 523736 267248
rect 523972 264316 524000 267706
rect 524788 267300 524840 267306
rect 524788 267242 524840 267248
rect 524800 264316 524828 267242
rect 525628 264316 525656 270302
rect 526824 264330 526852 273022
rect 527192 270230 527220 278038
rect 528192 275732 528244 275738
rect 528192 275674 528244 275680
rect 527180 270224 527232 270230
rect 527180 270166 527232 270172
rect 527180 268116 527232 268122
rect 527180 268058 527232 268064
rect 527192 267170 527220 268058
rect 527180 267164 527232 267170
rect 527180 267106 527232 267112
rect 528204 266762 528232 275674
rect 528376 270224 528428 270230
rect 528376 270166 528428 270172
rect 527272 266756 527324 266762
rect 527272 266698 527324 266704
rect 528192 266756 528244 266762
rect 528192 266698 528244 266704
rect 526470 264302 526852 264330
rect 527284 264316 527312 266698
rect 528388 264330 528416 270166
rect 528572 268394 528600 278038
rect 530412 275466 530440 278052
rect 531332 278038 531622 278066
rect 530400 275460 530452 275466
rect 530400 275402 530452 275408
rect 529848 272672 529900 272678
rect 529848 272614 529900 272620
rect 528560 268388 528612 268394
rect 528560 268330 528612 268336
rect 529664 267164 529716 267170
rect 529664 267106 529716 267112
rect 528928 266756 528980 266762
rect 528928 266698 528980 266704
rect 528126 264302 528416 264330
rect 528940 264316 528968 266698
rect 529676 264330 529704 267106
rect 529860 266762 529888 272614
rect 530398 270192 530454 270201
rect 531332 270178 531360 278038
rect 532332 275596 532384 275602
rect 532332 275538 532384 275544
rect 530398 270127 530454 270136
rect 530780 270150 531360 270178
rect 530412 269822 530440 270127
rect 530780 270094 530808 270150
rect 530768 270088 530820 270094
rect 530768 270030 530820 270036
rect 530952 270088 531004 270094
rect 530952 270030 531004 270036
rect 530400 269816 530452 269822
rect 530400 269758 530452 269764
rect 529848 266756 529900 266762
rect 529848 266698 529900 266704
rect 530964 264330 530992 270030
rect 532344 267734 532372 275538
rect 532516 272944 532568 272950
rect 532516 272886 532568 272892
rect 532252 267706 532372 267734
rect 531412 266756 531464 266762
rect 531412 266698 531464 266704
rect 529676 264302 529782 264330
rect 530610 264302 530992 264330
rect 531424 264316 531452 266698
rect 532252 264316 532280 267706
rect 532528 266762 532556 272886
rect 532712 272542 532740 278052
rect 533908 274786 533936 278052
rect 534092 278038 535118 278066
rect 535748 278038 536314 278066
rect 533896 274780 533948 274786
rect 533896 274722 533948 274728
rect 533712 272672 533764 272678
rect 533712 272614 533764 272620
rect 532700 272536 532752 272542
rect 532700 272478 532752 272484
rect 532884 270496 532936 270502
rect 532884 270438 532936 270444
rect 532896 269686 532924 270438
rect 533528 270360 533580 270366
rect 533172 270308 533528 270314
rect 533172 270302 533580 270308
rect 533172 270286 533568 270302
rect 533172 270094 533200 270286
rect 533160 270088 533212 270094
rect 533160 270030 533212 270036
rect 532884 269680 532936 269686
rect 532884 269622 532936 269628
rect 532516 266756 532568 266762
rect 532516 266698 532568 266704
rect 533068 266756 533120 266762
rect 533068 266698 533120 266704
rect 533080 264316 533108 266698
rect 533724 264330 533752 272614
rect 534092 270201 534120 278038
rect 534724 274780 534776 274786
rect 534724 274722 534776 274728
rect 534078 270192 534134 270201
rect 534078 270127 534134 270136
rect 533988 269952 534040 269958
rect 533988 269894 534040 269900
rect 534000 266762 534028 269894
rect 534736 267034 534764 274722
rect 534724 267028 534776 267034
rect 534724 266970 534776 266976
rect 534724 266892 534776 266898
rect 534724 266834 534776 266840
rect 533988 266756 534040 266762
rect 533988 266698 534040 266704
rect 533724 264302 533922 264330
rect 534736 264316 534764 266834
rect 535552 266756 535604 266762
rect 535552 266698 535604 266704
rect 535564 264316 535592 266698
rect 535748 265130 535776 278038
rect 537496 275330 537524 278052
rect 538508 278038 538706 278066
rect 537668 275460 537720 275466
rect 537668 275402 537720 275408
rect 537484 275324 537536 275330
rect 537484 275266 537536 275272
rect 536748 274100 536800 274106
rect 536748 274042 536800 274048
rect 536378 272912 536434 272921
rect 536378 272847 536434 272856
rect 536392 272542 536420 272847
rect 536380 272536 536432 272542
rect 536380 272478 536432 272484
rect 536564 272536 536616 272542
rect 536564 272478 536616 272484
rect 535736 265124 535788 265130
rect 535736 265066 535788 265072
rect 536576 264330 536604 272478
rect 536760 266762 536788 274042
rect 536748 266756 536800 266762
rect 536748 266698 536800 266704
rect 537680 264330 537708 275402
rect 537944 272944 537996 272950
rect 538128 272944 538180 272950
rect 537944 272886 537996 272892
rect 538126 272912 538128 272921
rect 538180 272912 538182 272921
rect 537956 272649 537984 272886
rect 538126 272847 538182 272856
rect 537942 272640 537998 272649
rect 537942 272575 537998 272584
rect 538128 272536 538180 272542
rect 538180 272484 538260 272490
rect 538128 272478 538260 272484
rect 538140 272462 538260 272478
rect 538232 272377 538260 272462
rect 538218 272368 538274 272377
rect 538218 272303 538274 272312
rect 538508 270178 538536 278038
rect 539888 277394 539916 278052
rect 539888 277366 540008 277394
rect 539322 274000 539378 274009
rect 539322 273935 539378 273944
rect 538680 272672 538732 272678
rect 538678 272640 538680 272649
rect 538732 272640 538734 272649
rect 538678 272575 538734 272584
rect 538140 270150 538536 270178
rect 538140 270094 538168 270150
rect 538128 270088 538180 270094
rect 538128 270030 538180 270036
rect 538312 270088 538364 270094
rect 538312 270030 538364 270036
rect 537852 269952 537904 269958
rect 537850 269920 537852 269929
rect 538036 269952 538088 269958
rect 537904 269920 537906 269929
rect 538324 269929 538352 270030
rect 538036 269894 538088 269900
rect 538310 269920 538366 269929
rect 537850 269855 537906 269864
rect 536406 264302 536604 264330
rect 537234 264302 537708 264330
rect 538048 264316 538076 269894
rect 538310 269855 538366 269864
rect 538588 269816 538640 269822
rect 538588 269758 538640 269764
rect 538772 269816 538824 269822
rect 538772 269758 538824 269764
rect 538600 269414 538628 269758
rect 538588 269408 538640 269414
rect 538588 269350 538640 269356
rect 538220 269272 538272 269278
rect 538784 269226 538812 269758
rect 538272 269220 538812 269226
rect 538220 269214 538812 269220
rect 538232 269198 538812 269214
rect 539336 264330 539364 273935
rect 539692 267028 539744 267034
rect 539692 266970 539744 266976
rect 538890 264302 539364 264330
rect 539704 264316 539732 266970
rect 539980 265266 540008 277366
rect 540992 274786 541020 278052
rect 541176 278038 542202 278066
rect 540980 274780 541032 274786
rect 540980 274722 541032 274728
rect 541176 269362 541204 278038
rect 543384 276282 543412 278052
rect 543372 276276 543424 276282
rect 543372 276218 543424 276224
rect 542268 275324 542320 275330
rect 542268 275266 542320 275272
rect 540624 269334 541204 269362
rect 540624 269278 540652 269334
rect 540612 269272 540664 269278
rect 540612 269214 540664 269220
rect 540796 269272 540848 269278
rect 540796 269214 540848 269220
rect 539968 265260 540020 265266
rect 539968 265202 540020 265208
rect 540808 264330 540836 269214
rect 541348 268388 541400 268394
rect 541348 268330 541400 268336
rect 540546 264302 540836 264330
rect 541360 264316 541388 268330
rect 542280 267734 542308 275266
rect 544580 274922 544608 278052
rect 544568 274916 544620 274922
rect 544568 274858 544620 274864
rect 545776 273970 545804 278052
rect 546512 278038 546986 278066
rect 547892 278038 548090 278066
rect 545946 274000 546002 274009
rect 545764 273964 545816 273970
rect 545946 273935 545948 273944
rect 545764 273906 545816 273912
rect 546000 273935 546002 273944
rect 545948 273906 546000 273912
rect 543188 269952 543240 269958
rect 543188 269894 543240 269900
rect 542820 269816 542872 269822
rect 542820 269758 542872 269764
rect 542832 269090 542860 269758
rect 543200 269278 543228 269894
rect 543188 269272 543240 269278
rect 543188 269214 543240 269220
rect 546512 269210 546540 278038
rect 547694 272368 547750 272377
rect 547694 272303 547750 272312
rect 547708 272134 547736 272303
rect 547512 272128 547564 272134
rect 547510 272096 547512 272105
rect 547696 272128 547748 272134
rect 547564 272096 547566 272105
rect 547892 272105 547920 278038
rect 549272 273562 549300 278052
rect 550468 276418 550496 278052
rect 550652 278038 551678 278066
rect 550456 276412 550508 276418
rect 550456 276354 550508 276360
rect 549260 273556 549312 273562
rect 549260 273498 549312 273504
rect 549904 273556 549956 273562
rect 549904 273498 549956 273504
rect 547696 272070 547748 272076
rect 547878 272096 547934 272105
rect 547510 272031 547566 272040
rect 547878 272031 547934 272040
rect 543372 269204 543424 269210
rect 543372 269146 543424 269152
rect 546500 269204 546552 269210
rect 546500 269146 546552 269152
rect 543384 269090 543412 269146
rect 542832 269062 543412 269090
rect 542188 267706 542308 267734
rect 542188 264316 542216 267706
rect 543004 266756 543056 266762
rect 543004 266698 543056 266704
rect 543016 264316 543044 266698
rect 549916 266490 549944 273498
rect 549904 266484 549956 266490
rect 549904 266426 549956 266432
rect 550652 265402 550680 278038
rect 552860 273426 552888 278052
rect 553412 278038 554070 278066
rect 552848 273420 552900 273426
rect 552848 273362 552900 273368
rect 553412 265538 553440 278038
rect 555252 277370 555280 278052
rect 555240 277364 555292 277370
rect 555240 277306 555292 277312
rect 556356 273834 556384 278052
rect 557552 276554 557580 278052
rect 557736 278038 558762 278066
rect 557540 276548 557592 276554
rect 557540 276490 557592 276496
rect 556344 273828 556396 273834
rect 556344 273770 556396 273776
rect 556804 273828 556856 273834
rect 556804 273770 556856 273776
rect 556816 266626 556844 273770
rect 556804 266620 556856 266626
rect 556804 266562 556856 266568
rect 557736 266354 557764 278038
rect 559944 273698 559972 278052
rect 560680 278038 561154 278066
rect 561968 278038 562350 278066
rect 559932 273692 559984 273698
rect 559932 273634 559984 273640
rect 557724 266348 557776 266354
rect 557724 266290 557776 266296
rect 560680 266218 560708 278038
rect 561968 271998 561996 278038
rect 563440 274650 563468 278052
rect 563428 274644 563480 274650
rect 563428 274586 563480 274592
rect 562140 272808 562192 272814
rect 562140 272750 562192 272756
rect 562324 272808 562376 272814
rect 562324 272750 562376 272756
rect 562152 271998 562180 272750
rect 562336 272134 562364 272750
rect 562324 272128 562376 272134
rect 562324 272070 562376 272076
rect 561956 271992 562008 271998
rect 561956 271934 562008 271940
rect 562140 271992 562192 271998
rect 562140 271934 562192 271940
rect 564636 270774 564664 278052
rect 565832 277234 565860 278052
rect 565820 277228 565872 277234
rect 565820 277170 565872 277176
rect 567028 274514 567056 278052
rect 567016 274508 567068 274514
rect 567016 274450 567068 274456
rect 564624 270768 564676 270774
rect 564624 270710 564676 270716
rect 567844 270768 567896 270774
rect 567844 270710 567896 270716
rect 567856 267714 567884 270710
rect 568224 270638 568252 278052
rect 569420 271998 569448 278052
rect 570064 278038 570630 278066
rect 569408 271992 569460 271998
rect 569408 271934 569460 271940
rect 568212 270632 568264 270638
rect 568212 270574 568264 270580
rect 570064 267986 570092 278038
rect 571720 270910 571748 278052
rect 572732 278038 572930 278066
rect 571708 270904 571760 270910
rect 571708 270846 571760 270852
rect 570052 267980 570104 267986
rect 570052 267922 570104 267928
rect 567844 267708 567896 267714
rect 567844 267650 567896 267656
rect 560668 266212 560720 266218
rect 560668 266154 560720 266160
rect 572732 266082 572760 278038
rect 574112 268258 574140 278052
rect 575308 271046 575336 278052
rect 575492 278038 576518 278066
rect 576872 278038 577714 278066
rect 578528 278038 578910 278066
rect 575296 271040 575348 271046
rect 575296 270982 575348 270988
rect 575492 269414 575520 278038
rect 575480 269408 575532 269414
rect 575480 269350 575532 269356
rect 576872 269074 576900 278038
rect 578528 271862 578556 278038
rect 580000 277098 580028 278052
rect 581012 278038 581210 278066
rect 579988 277092 580040 277098
rect 579988 277034 580040 277040
rect 578516 271856 578568 271862
rect 578516 271798 578568 271804
rect 578884 271856 578936 271862
rect 578884 271798 578936 271804
rect 576860 269068 576912 269074
rect 576860 269010 576912 269016
rect 574100 268252 574152 268258
rect 574100 268194 574152 268200
rect 578896 267578 578924 271798
rect 581012 268938 581040 278038
rect 582392 271726 582420 278052
rect 583588 273562 583616 278052
rect 583772 278038 584798 278066
rect 583576 273556 583628 273562
rect 583576 273498 583628 273504
rect 582380 271720 582432 271726
rect 582380 271662 582432 271668
rect 583024 271720 583076 271726
rect 583024 271662 583076 271668
rect 581000 268932 581052 268938
rect 581000 268874 581052 268880
rect 578884 267572 578936 267578
rect 578884 267514 578936 267520
rect 583036 267442 583064 271662
rect 583772 268802 583800 278038
rect 585980 271590 586008 278052
rect 587084 275058 587112 278052
rect 587912 278038 588294 278066
rect 587072 275052 587124 275058
rect 587072 274994 587124 275000
rect 585968 271584 586020 271590
rect 585968 271526 586020 271532
rect 583760 268796 583812 268802
rect 583760 268738 583812 268744
rect 587912 268666 587940 278038
rect 589476 271454 589504 278052
rect 590672 273834 590700 278052
rect 591868 274378 591896 278052
rect 591856 274372 591908 274378
rect 591856 274314 591908 274320
rect 590660 273828 590712 273834
rect 590660 273770 590712 273776
rect 589464 271448 589516 271454
rect 589464 271390 589516 271396
rect 589924 271448 589976 271454
rect 589924 271390 589976 271396
rect 587900 268660 587952 268666
rect 587900 268602 587952 268608
rect 583024 267436 583076 267442
rect 583024 267378 583076 267384
rect 589936 266898 589964 271390
rect 593064 271318 593092 278052
rect 594260 275194 594288 278052
rect 594812 278038 595378 278066
rect 596192 278038 596574 278066
rect 594248 275188 594300 275194
rect 594248 275130 594300 275136
rect 593052 271312 593104 271318
rect 593052 271254 593104 271260
rect 594812 268530 594840 278038
rect 596192 269550 596220 278038
rect 597756 270774 597784 278052
rect 598952 274242 598980 278052
rect 600148 276962 600176 278052
rect 600136 276956 600188 276962
rect 600136 276898 600188 276904
rect 601344 276010 601372 278052
rect 601712 278038 602462 278066
rect 601332 276004 601384 276010
rect 601332 275946 601384 275952
rect 598940 274236 598992 274242
rect 598940 274178 598992 274184
rect 601148 272808 601200 272814
rect 601148 272750 601200 272756
rect 601160 272406 601188 272750
rect 600964 272400 601016 272406
rect 600964 272342 601016 272348
rect 601148 272400 601200 272406
rect 601148 272342 601200 272348
rect 600976 272134 601004 272342
rect 600964 272128 601016 272134
rect 600964 272070 601016 272076
rect 598204 271312 598256 271318
rect 598204 271254 598256 271260
rect 597744 270768 597796 270774
rect 597744 270710 597796 270716
rect 596180 269544 596232 269550
rect 596180 269486 596232 269492
rect 594800 268524 594852 268530
rect 594800 268466 594852 268472
rect 589924 266892 589976 266898
rect 589924 266834 589976 266840
rect 598216 266762 598244 271254
rect 598204 266756 598256 266762
rect 598204 266698 598256 266704
rect 572720 266076 572772 266082
rect 572720 266018 572772 266024
rect 601712 265946 601740 278038
rect 603644 276826 603672 278052
rect 603632 276820 603684 276826
rect 603632 276762 603684 276768
rect 604840 271862 604868 278052
rect 605852 278038 606050 278066
rect 604828 271856 604880 271862
rect 604828 271798 604880 271804
rect 601700 265940 601752 265946
rect 601700 265882 601752 265888
rect 605852 265810 605880 278038
rect 607232 272134 607260 278052
rect 607416 278038 608442 278066
rect 607220 272128 607272 272134
rect 607220 272070 607272 272076
rect 607416 268122 607444 278038
rect 609624 276690 609652 278052
rect 609612 276684 609664 276690
rect 609612 276626 609664 276632
rect 610728 272270 610756 278052
rect 610716 272264 610768 272270
rect 610716 272206 610768 272212
rect 611924 271726 611952 278052
rect 612752 278038 613134 278066
rect 611912 271720 611964 271726
rect 611912 271662 611964 271668
rect 612004 271584 612056 271590
rect 612004 271526 612056 271532
rect 607404 268116 607456 268122
rect 607404 268058 607456 268064
rect 612016 267306 612044 271526
rect 612004 267300 612056 267306
rect 612004 267242 612056 267248
rect 605840 265804 605892 265810
rect 605840 265746 605892 265752
rect 612752 265674 612780 278038
rect 614316 273222 614344 278052
rect 615512 275874 615540 278052
rect 616248 278038 616722 278066
rect 617352 278038 617826 278066
rect 615500 275868 615552 275874
rect 615500 275810 615552 275816
rect 614304 273216 614356 273222
rect 614304 273158 614356 273164
rect 616248 269686 616276 278038
rect 617352 271182 617380 278038
rect 619008 271590 619036 278052
rect 619652 278038 620218 278066
rect 618996 271584 619048 271590
rect 618996 271526 619048 271532
rect 617340 271176 617392 271182
rect 617340 271118 617392 271124
rect 617524 271176 617576 271182
rect 617524 271118 617576 271124
rect 616236 269680 616288 269686
rect 616236 269622 616288 269628
rect 617536 267170 617564 271118
rect 619652 270502 619680 278038
rect 621400 273086 621428 278052
rect 622596 275738 622624 278052
rect 623806 278038 624004 278066
rect 622584 275732 622636 275738
rect 622584 275674 622636 275680
rect 621388 273080 621440 273086
rect 621388 273022 621440 273028
rect 619640 270496 619692 270502
rect 619640 270438 619692 270444
rect 623976 270230 624004 278038
rect 624988 272950 625016 278052
rect 624976 272944 625028 272950
rect 624976 272886 625028 272892
rect 626092 271182 626120 278052
rect 626552 278038 627302 278066
rect 626080 271176 626132 271182
rect 626080 271118 626132 271124
rect 626552 270366 626580 278038
rect 628484 272678 628512 278052
rect 629680 275602 629708 278052
rect 629956 277778 629984 278122
rect 629944 277772 629996 277778
rect 629944 277714 629996 277720
rect 630140 277642 630168 278122
rect 630692 278038 630890 278066
rect 630128 277636 630180 277642
rect 630128 277578 630180 277584
rect 629668 275596 629720 275602
rect 629668 275538 629720 275544
rect 628472 272672 628524 272678
rect 628472 272614 628524 272620
rect 626540 270360 626592 270366
rect 626540 270302 626592 270308
rect 623964 270224 624016 270230
rect 623964 270166 624016 270172
rect 630692 270094 630720 278038
rect 632072 272542 632100 278052
rect 632060 272536 632112 272542
rect 632060 272478 632112 272484
rect 633268 271454 633296 278052
rect 634372 274106 634400 278052
rect 635096 278044 635148 278050
rect 635096 277986 635148 277992
rect 634360 274100 634412 274106
rect 634360 274042 634412 274048
rect 634084 272672 634136 272678
rect 634084 272614 634136 272620
rect 633256 271448 633308 271454
rect 633256 271390 633308 271396
rect 630680 270088 630732 270094
rect 630680 270030 630732 270036
rect 617524 267164 617576 267170
rect 617524 267106 617576 267112
rect 634096 267034 634124 272614
rect 634084 267028 634136 267034
rect 634084 266970 634136 266976
rect 612740 265668 612792 265674
rect 612740 265610 612792 265616
rect 553400 265532 553452 265538
rect 553400 265474 553452 265480
rect 550640 265396 550692 265402
rect 550640 265338 550692 265344
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 563704 259480 563756 259486
rect 563704 259422 563756 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 560944 256760 560996 256766
rect 560944 256702 560996 256708
rect 554502 255640 554558 255649
rect 554502 255575 554504 255584
rect 554556 255575 554558 255584
rect 558184 255604 558236 255610
rect 554504 255546 554556 255552
rect 558184 255546 558236 255552
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 554134 251288 554190 251297
rect 554134 251223 554136 251232
rect 554188 251223 554190 251232
rect 556804 251252 556856 251258
rect 554136 251194 554188 251200
rect 556804 251194 556856 251200
rect 554042 249112 554098 249121
rect 554042 249047 554098 249056
rect 553858 246936 553914 246945
rect 553858 246871 553914 246880
rect 553872 245682 553900 246871
rect 553860 245676 553912 245682
rect 553860 245618 553912 245624
rect 553490 244760 553546 244769
rect 553490 244695 553546 244704
rect 553504 244322 553532 244695
rect 553492 244316 553544 244322
rect 553492 244258 553544 244264
rect 553674 242584 553730 242593
rect 553674 242519 553730 242528
rect 553688 241534 553716 242519
rect 553676 241528 553728 241534
rect 553676 241470 553728 241476
rect 553768 236836 553820 236842
rect 553768 236778 553820 236784
rect 553780 236065 553808 236778
rect 553766 236056 553822 236065
rect 553766 235991 553822 236000
rect 135168 231464 135220 231470
rect 135168 231406 135220 231412
rect 137652 231464 137704 231470
rect 137652 231406 137704 231412
rect 92388 231192 92440 231198
rect 92388 231134 92440 231140
rect 82084 230036 82136 230042
rect 82084 229978 82136 229984
rect 86224 230036 86276 230042
rect 86224 229978 86276 229984
rect 68284 229764 68336 229770
rect 68284 229706 68336 229712
rect 67548 228676 67600 228682
rect 67548 228618 67600 228624
rect 64788 227724 64840 227730
rect 64788 227666 64840 227672
rect 63316 227180 63368 227186
rect 63316 227122 63368 227128
rect 63130 224496 63186 224505
rect 63130 224431 63186 224440
rect 62946 223544 63002 223553
rect 62946 223479 63002 223488
rect 62764 222896 62816 222902
rect 62764 222838 62816 222844
rect 62304 219020 62356 219026
rect 62304 218962 62356 218968
rect 61384 218204 61436 218210
rect 61384 218146 61436 218152
rect 61476 218068 61528 218074
rect 61476 218010 61528 218016
rect 58130 217110 58204 217138
rect 58958 217110 59032 217138
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 58130 216988 58158 217110
rect 58958 216988 58986 217110
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61488 217138 61516 218010
rect 62316 217138 62344 218962
rect 62776 218074 62804 222838
rect 63328 219434 63356 227122
rect 63144 219406 63356 219434
rect 62764 218068 62816 218074
rect 62764 218010 62816 218016
rect 63144 217274 63172 219406
rect 64604 219156 64656 219162
rect 64604 219098 64656 219104
rect 63960 218068 64012 218074
rect 63960 218010 64012 218016
rect 61442 217110 61516 217138
rect 62270 217110 62344 217138
rect 63098 217246 63172 217274
rect 61442 216988 61470 217110
rect 62270 216988 62298 217110
rect 63098 216988 63126 217246
rect 63972 217138 64000 218010
rect 64616 217274 64644 219098
rect 64800 218074 64828 227666
rect 66168 226024 66220 226030
rect 66168 225966 66220 225972
rect 66180 218074 66208 225966
rect 66904 223168 66956 223174
rect 66904 223110 66956 223116
rect 66916 219162 66944 223110
rect 66904 219156 66956 219162
rect 66904 219098 66956 219104
rect 67560 218210 67588 228618
rect 66444 218204 66496 218210
rect 66444 218146 66496 218152
rect 67548 218204 67600 218210
rect 67548 218146 67600 218152
rect 68100 218204 68152 218210
rect 68100 218146 68152 218152
rect 64788 218068 64840 218074
rect 64788 218010 64840 218016
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 64616 217246 64782 217274
rect 63926 217110 64000 217138
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217138 66484 218146
rect 67272 218068 67324 218074
rect 67272 218010 67324 218016
rect 67284 217138 67312 218010
rect 68112 217138 68140 218146
rect 68296 218074 68324 229706
rect 76564 225752 76616 225758
rect 76564 225694 76616 225700
rect 72424 225616 72476 225622
rect 72424 225558 72476 225564
rect 68928 224120 68980 224126
rect 68928 224062 68980 224068
rect 68284 218068 68336 218074
rect 68284 218010 68336 218016
rect 68940 217274 68968 224062
rect 69572 223304 69624 223310
rect 69572 223246 69624 223252
rect 69584 218210 69612 223246
rect 71412 223032 71464 223038
rect 71412 222974 71464 222980
rect 69756 220516 69808 220522
rect 69756 220458 69808 220464
rect 69572 218204 69624 218210
rect 69572 218146 69624 218152
rect 69768 217274 69796 220458
rect 70584 219428 70636 219434
rect 70584 219370 70636 219376
rect 65582 217110 65656 217138
rect 66410 217110 66484 217138
rect 67238 217110 67312 217138
rect 68066 217110 68140 217138
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217110
rect 67238 216988 67266 217110
rect 68066 216988 68094 217110
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 219370
rect 71424 217274 71452 222974
rect 72436 219026 72464 225558
rect 73712 224392 73764 224398
rect 73712 224334 73764 224340
rect 73068 220380 73120 220386
rect 73068 220322 73120 220328
rect 72424 219020 72476 219026
rect 72424 218962 72476 218968
rect 72240 218068 72292 218074
rect 72240 218010 72292 218016
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 218010
rect 73080 217274 73108 220322
rect 73724 218074 73752 224334
rect 75828 223440 75880 223446
rect 75828 223382 75880 223388
rect 73896 221604 73948 221610
rect 73896 221546 73948 221552
rect 73712 218068 73764 218074
rect 73712 218010 73764 218016
rect 73908 217274 73936 221546
rect 75552 218204 75604 218210
rect 75552 218146 75604 218152
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72206 217110 72280 217138
rect 73034 217246 73108 217274
rect 73862 217246 73936 217274
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73862 216988 73890 217246
rect 74736 217138 74764 218010
rect 75564 217138 75592 218146
rect 75840 218074 75868 223382
rect 76380 220108 76432 220114
rect 76380 220050 76432 220056
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220050
rect 76576 218210 76604 225694
rect 79968 224528 80020 224534
rect 79968 224470 80020 224476
rect 78588 222760 78640 222766
rect 78588 222702 78640 222708
rect 77208 219020 77260 219026
rect 77208 218962 77260 218968
rect 76564 218204 76616 218210
rect 76564 218146 76616 218152
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218962
rect 78600 218074 78628 222702
rect 79692 220244 79744 220250
rect 79692 220186 79744 220192
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217274 79732 220186
rect 79980 218074 80008 224470
rect 81348 223576 81400 223582
rect 81348 223518 81400 223524
rect 80520 221740 80572 221746
rect 80520 221682 80572 221688
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217274 80560 221682
rect 81360 217274 81388 223518
rect 82096 221610 82124 229978
rect 83464 225888 83516 225894
rect 83464 225830 83516 225836
rect 82084 221604 82136 221610
rect 82084 221546 82136 221552
rect 83004 220924 83056 220930
rect 83004 220866 83056 220872
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217246 79732 217274
rect 80486 217246 80560 217274
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217246
rect 80486 216988 80514 217246
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220866
rect 83476 218074 83504 225830
rect 85488 224664 85540 224670
rect 85488 224606 85540 224612
rect 85304 222352 85356 222358
rect 85304 222294 85356 222300
rect 83832 219156 83884 219162
rect 83832 219098 83884 219104
rect 83464 218068 83516 218074
rect 83464 218010 83516 218016
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 219098
rect 85316 218074 85344 222294
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 85304 218068 85356 218074
rect 85304 218010 85356 218016
rect 84672 217138 84700 218010
rect 85500 217274 85528 224606
rect 86236 221746 86264 229978
rect 88248 227860 88300 227866
rect 88248 227802 88300 227808
rect 87972 222488 88024 222494
rect 87972 222430 88024 222436
rect 86224 221740 86276 221746
rect 86224 221682 86276 221688
rect 86316 221604 86368 221610
rect 86316 221546 86368 221552
rect 86328 217274 86356 221546
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 85454 217246 85528 217274
rect 86282 217246 86356 217274
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86282 216988 86310 217246
rect 87156 217138 87184 218010
rect 87984 217274 88012 222430
rect 88260 218074 88288 227802
rect 89628 227316 89680 227322
rect 89628 227258 89680 227264
rect 88984 224392 89036 224398
rect 88984 224334 89036 224340
rect 89444 224392 89496 224398
rect 89444 224334 89496 224340
rect 88996 224126 89024 224334
rect 88984 224120 89036 224126
rect 88984 224062 89036 224068
rect 89456 218074 89484 224334
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227258
rect 91284 221740 91336 221746
rect 91284 221682 91336 221688
rect 91296 217274 91324 221682
rect 92400 219434 92428 231134
rect 128268 231056 128320 231062
rect 128268 230998 128320 231004
rect 118608 230920 118660 230926
rect 118608 230862 118660 230868
rect 94504 230784 94556 230790
rect 94504 230726 94556 230732
rect 93584 228812 93636 228818
rect 93584 228754 93636 228760
rect 92124 219406 92428 219434
rect 92124 217274 92152 219406
rect 93596 218074 93624 228754
rect 94516 219434 94544 230726
rect 104808 230648 104860 230654
rect 104808 230590 104860 230596
rect 95240 230172 95292 230178
rect 95240 230114 95292 230120
rect 95252 227866 95280 230114
rect 102140 229492 102192 229498
rect 102140 229434 102192 229440
rect 100668 228948 100720 228954
rect 100668 228890 100720 228896
rect 95240 227860 95292 227866
rect 95240 227802 95292 227808
rect 96436 227452 96488 227458
rect 96436 227394 96488 227400
rect 96252 224936 96304 224942
rect 96252 224878 96304 224884
rect 94688 222012 94740 222018
rect 94688 221954 94740 221960
rect 94700 219434 94728 221954
rect 94424 219406 94544 219434
rect 94608 219406 94728 219434
rect 94424 219298 94452 219406
rect 93768 219292 93820 219298
rect 93768 219234 93820 219240
rect 94412 219292 94464 219298
rect 94412 219234 94464 219240
rect 92940 218068 92992 218074
rect 92940 218010 92992 218016
rect 93584 218068 93636 218074
rect 93584 218010 93636 218016
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 90410 217252 90462 217258
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90410 217194 90462 217200
rect 91250 217246 91324 217274
rect 92078 217246 92152 217274
rect 90422 216988 90450 217194
rect 91250 216988 91278 217246
rect 92078 216988 92106 217246
rect 92952 217138 92980 218010
rect 93780 217138 93808 219234
rect 94608 217274 94636 219406
rect 96264 218074 96292 224878
rect 95424 218068 95476 218074
rect 95424 218010 95476 218016
rect 96252 218068 96304 218074
rect 96252 218010 96304 218016
rect 92906 217110 92980 217138
rect 93734 217110 93808 217138
rect 94562 217246 94636 217274
rect 92906 216988 92934 217110
rect 93734 216988 93762 217110
rect 94562 216988 94590 217246
rect 95436 217138 95464 218010
rect 96448 217274 96476 227394
rect 99288 222624 99340 222630
rect 99288 222566 99340 222572
rect 97908 222148 97960 222154
rect 97908 222090 97960 222096
rect 97080 218204 97132 218210
rect 97080 218146 97132 218152
rect 95390 217110 95464 217138
rect 96218 217246 96476 217274
rect 95390 216988 95418 217110
rect 96218 216988 96246 217246
rect 97092 217138 97120 218146
rect 97920 217274 97948 222090
rect 99300 218074 99328 222566
rect 100392 218340 100444 218346
rect 100392 218282 100444 218288
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97046 217110 97120 217138
rect 97874 217246 97948 217274
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218282
rect 100680 218074 100708 228890
rect 102152 227594 102180 229434
rect 102140 227588 102192 227594
rect 102140 227530 102192 227536
rect 103428 227588 103480 227594
rect 103428 227530 103480 227536
rect 102048 224800 102100 224806
rect 102048 224742 102100 224748
rect 101220 220652 101272 220658
rect 101220 220594 101272 220600
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101232 217274 101260 220594
rect 102060 217274 102088 224742
rect 103440 218142 103468 227530
rect 104348 222148 104400 222154
rect 104348 222090 104400 222096
rect 104360 221882 104388 222090
rect 104348 221876 104400 221882
rect 104348 221818 104400 221824
rect 104532 221332 104584 221338
rect 104532 221274 104584 221280
rect 102876 218136 102928 218142
rect 102876 218078 102928 218084
rect 103428 218136 103480 218142
rect 103428 218078 103480 218084
rect 103704 218136 103756 218142
rect 103704 218078 103756 218084
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217246 101260 217274
rect 102014 217246 102088 217274
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217246
rect 102014 216988 102042 217246
rect 102888 217138 102916 218078
rect 103716 217138 103744 218078
rect 104544 217274 104572 221274
rect 104820 218142 104848 230590
rect 110328 229356 110380 229362
rect 110328 229298 110380 229304
rect 106188 229084 106240 229090
rect 106188 229026 106240 229032
rect 105912 223984 105964 223990
rect 105912 223926 105964 223932
rect 105924 219434 105952 223926
rect 105924 219406 106044 219434
rect 106016 218142 106044 219406
rect 104808 218136 104860 218142
rect 104808 218078 104860 218084
rect 105360 218136 105412 218142
rect 105360 218078 105412 218084
rect 106004 218136 106056 218142
rect 106004 218078 106056 218084
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218078
rect 106200 217274 106228 229026
rect 110340 227730 110368 229298
rect 112996 228268 113048 228274
rect 112996 228210 113048 228216
rect 110328 227724 110380 227730
rect 110328 227666 110380 227672
rect 110512 227724 110564 227730
rect 110512 227666 110564 227672
rect 110524 227610 110552 227666
rect 110340 227582 110552 227610
rect 110144 225480 110196 225486
rect 110144 225422 110196 225428
rect 108672 223848 108724 223854
rect 108672 223790 108724 223796
rect 106372 222148 106424 222154
rect 106372 222090 106424 222096
rect 106384 221338 106412 222090
rect 106372 221332 106424 221338
rect 106372 221274 106424 221280
rect 107844 219972 107896 219978
rect 107844 219914 107896 219920
rect 107016 218272 107068 218278
rect 107016 218214 107068 218220
rect 107028 217274 107056 218214
rect 107856 217274 107884 219914
rect 108684 217274 108712 223790
rect 110156 219434 110184 225422
rect 110340 219434 110368 227582
rect 112812 223712 112864 223718
rect 112812 223654 112864 223660
rect 111156 221332 111208 221338
rect 111156 221274 111208 221280
rect 109500 219428 109552 219434
rect 110156 219406 110276 219434
rect 110340 219428 110472 219434
rect 110340 219406 110420 219428
rect 109500 219370 109552 219376
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 106982 217246 107056 217274
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 106982 216988 107010 217246
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 219370
rect 110248 217274 110276 219406
rect 110420 219370 110472 219376
rect 111168 217274 111196 221274
rect 112824 218142 112852 223654
rect 111984 218136 112036 218142
rect 111984 218078 112036 218084
rect 112812 218136 112864 218142
rect 112812 218078 112864 218084
rect 110248 217246 110322 217274
rect 109466 217110 109540 217138
rect 109466 216988 109494 217110
rect 110294 216988 110322 217246
rect 111122 217246 111196 217274
rect 111122 216988 111150 217246
rect 111996 217138 112024 218078
rect 113008 217274 113036 228210
rect 117228 226908 117280 226914
rect 117228 226850 117280 226856
rect 114284 220788 114336 220794
rect 114284 220730 114336 220736
rect 114296 219978 114324 220730
rect 114284 219972 114336 219978
rect 114284 219914 114336 219920
rect 114468 219972 114520 219978
rect 114468 219914 114520 219920
rect 113640 218612 113692 218618
rect 113640 218554 113692 218560
rect 111950 217110 112024 217138
rect 112778 217246 113036 217274
rect 111950 216988 111978 217110
rect 112778 216988 112806 217246
rect 113652 217138 113680 218554
rect 114480 217274 114508 219914
rect 117240 218346 117268 226850
rect 118422 222320 118478 222329
rect 118422 222255 118478 222264
rect 118436 219434 118464 222255
rect 118620 219434 118648 230862
rect 126888 230308 126940 230314
rect 126888 230250 126940 230256
rect 123484 229220 123536 229226
rect 123484 229162 123536 229168
rect 119988 228132 120040 228138
rect 119988 228074 120040 228080
rect 117780 219428 117832 219434
rect 118436 219406 118556 219434
rect 118620 219428 118752 219434
rect 118620 219406 118700 219428
rect 117780 219370 117832 219376
rect 116124 218340 116176 218346
rect 116124 218282 116176 218288
rect 117228 218340 117280 218346
rect 117228 218282 117280 218288
rect 115296 217456 115348 217462
rect 115296 217398 115348 217404
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115308 217138 115336 217398
rect 116136 217138 116164 218282
rect 116952 217592 117004 217598
rect 116952 217534 117004 217540
rect 116964 217138 116992 217534
rect 117792 217138 117820 219370
rect 118528 217274 118556 219406
rect 118700 219370 118752 219376
rect 120000 218346 120028 228074
rect 122748 226772 122800 226778
rect 122748 226714 122800 226720
rect 122564 226296 122616 226302
rect 122564 226238 122616 226244
rect 121092 219836 121144 219842
rect 121092 219778 121144 219784
rect 120264 219428 120316 219434
rect 120264 219370 120316 219376
rect 119436 218340 119488 218346
rect 119436 218282 119488 218288
rect 119988 218340 120040 218346
rect 119988 218282 120040 218288
rect 118528 217246 118602 217274
rect 115262 217110 115336 217138
rect 116090 217110 116164 217138
rect 116918 217110 116992 217138
rect 117746 217110 117820 217138
rect 115262 216988 115290 217110
rect 116090 216988 116118 217110
rect 116918 216988 116946 217110
rect 117746 216988 117774 217110
rect 118574 216988 118602 217246
rect 119448 217138 119476 218282
rect 120276 217138 120304 219370
rect 121104 217274 121132 219778
rect 122576 218346 122604 226238
rect 121920 218340 121972 218346
rect 121920 218282 121972 218288
rect 122564 218340 122616 218346
rect 122564 218282 122616 218288
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 218282
rect 122760 217274 122788 226714
rect 123496 219570 123524 229162
rect 126704 227996 126756 228002
rect 126704 227938 126756 227944
rect 125232 225344 125284 225350
rect 125232 225286 125284 225292
rect 124404 221060 124456 221066
rect 124404 221002 124456 221008
rect 123484 219564 123536 219570
rect 123484 219506 123536 219512
rect 123576 219428 123628 219434
rect 123576 219370 123628 219376
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123588 217138 123616 219370
rect 124416 217274 124444 221002
rect 125244 217274 125272 225286
rect 126716 218346 126744 227938
rect 126060 218340 126112 218346
rect 126060 218282 126112 218288
rect 126704 218340 126756 218346
rect 126704 218282 126756 218288
rect 123542 217110 123616 217138
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 123542 216988 123570 217110
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126072 217138 126100 218282
rect 126900 217274 126928 230250
rect 127624 226160 127676 226166
rect 127624 226102 127676 226108
rect 127636 225486 127664 226102
rect 127624 225480 127676 225486
rect 127624 225422 127676 225428
rect 127624 219972 127676 219978
rect 127624 219914 127676 219920
rect 127636 219706 127664 219914
rect 127624 219700 127676 219706
rect 127624 219642 127676 219648
rect 128280 218346 128308 230998
rect 133788 230444 133840 230450
rect 133788 230386 133840 230392
rect 133512 227860 133564 227866
rect 133512 227802 133564 227808
rect 129556 226636 129608 226642
rect 129556 226578 129608 226584
rect 129372 225344 129424 225350
rect 129372 225286 129424 225292
rect 129384 218346 129412 225286
rect 127716 218340 127768 218346
rect 127716 218282 127768 218288
rect 128268 218340 128320 218346
rect 128268 218282 128320 218288
rect 128544 218340 128596 218346
rect 128544 218282 128596 218288
rect 129372 218340 129424 218346
rect 129372 218282 129424 218288
rect 126026 217110 126100 217138
rect 126854 217246 126928 217274
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 218282
rect 128556 217138 128584 218282
rect 129568 217274 129596 226578
rect 132408 225072 132460 225078
rect 132408 225014 132460 225020
rect 131028 219700 131080 219706
rect 131028 219642 131080 219648
rect 129832 219428 129884 219434
rect 129832 219370 129884 219376
rect 130200 219428 130252 219434
rect 130200 219370 130252 219376
rect 129844 218346 129872 219370
rect 129832 218340 129884 218346
rect 129832 218282 129884 218288
rect 127682 217110 127756 217138
rect 128510 217110 128584 217138
rect 129338 217246 129596 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217110
rect 129338 216988 129366 217246
rect 130212 217138 130240 219370
rect 131040 217274 131068 219642
rect 132420 219434 132448 225014
rect 131856 219428 131908 219434
rect 131856 219370 131908 219376
rect 132408 219428 132460 219434
rect 132408 219370 132460 219376
rect 130166 217110 130240 217138
rect 130994 217246 131068 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217246
rect 131868 217138 131896 219370
rect 132498 218376 132554 218385
rect 133524 218346 133552 227802
rect 133800 219434 133828 230386
rect 135180 229094 135208 231406
rect 137664 230518 137692 231406
rect 137652 230512 137704 230518
rect 137652 230454 137704 230460
rect 137468 230444 137520 230450
rect 137468 230386 137520 230392
rect 137480 230042 137508 230386
rect 137284 230036 137336 230042
rect 137284 229978 137336 229984
rect 137468 230036 137520 230042
rect 137468 229978 137520 229984
rect 137296 229634 137324 229978
rect 137284 229628 137336 229634
rect 137284 229570 137336 229576
rect 133708 219406 133828 219434
rect 134352 229066 135208 229094
rect 140042 229120 140098 229129
rect 132498 218311 132500 218320
rect 132552 218311 132554 218320
rect 132684 218340 132736 218346
rect 132500 218282 132552 218288
rect 132684 218282 132736 218288
rect 133512 218340 133564 218346
rect 133512 218282 133564 218288
rect 132696 217138 132724 218282
rect 133708 217274 133736 219406
rect 134352 217274 134380 229066
rect 140042 229055 140098 229064
rect 137376 228540 137428 228546
rect 137376 228482 137428 228488
rect 137388 228426 137416 228482
rect 136824 228404 136876 228410
rect 136824 228346 136876 228352
rect 137204 228398 137416 228426
rect 139308 228404 139360 228410
rect 136638 227896 136694 227905
rect 136836 227866 136864 228346
rect 137204 228274 137232 228398
rect 139308 228346 139360 228352
rect 137192 228268 137244 228274
rect 137192 228210 137244 228216
rect 136638 227831 136640 227840
rect 136692 227831 136694 227840
rect 136824 227860 136876 227866
rect 136640 227802 136692 227808
rect 136824 227802 136876 227808
rect 136548 226500 136600 226506
rect 136548 226442 136600 226448
rect 135076 225208 135128 225214
rect 135076 225150 135128 225156
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133736 217274
rect 134306 217246 134380 217274
rect 135088 217274 135116 225150
rect 136560 218346 136588 226442
rect 136730 223952 136786 223961
rect 136730 223887 136786 223896
rect 136744 218385 136772 223887
rect 138480 221196 138532 221202
rect 138480 221138 138532 221144
rect 136916 220516 136968 220522
rect 136916 220458 136968 220464
rect 137100 220516 137152 220522
rect 137100 220458 137152 220464
rect 136928 219570 136956 220458
rect 137112 219842 137140 220458
rect 137100 219836 137152 219842
rect 137100 219778 137152 219784
rect 136916 219564 136968 219570
rect 136916 219506 136968 219512
rect 137652 219564 137704 219570
rect 137652 219506 137704 219512
rect 136730 218376 136786 218385
rect 135996 218340 136048 218346
rect 135996 218282 136048 218288
rect 136548 218340 136600 218346
rect 136730 218311 136786 218320
rect 136916 218340 136968 218346
rect 136548 218282 136600 218288
rect 136916 218282 136968 218288
rect 135088 217246 135162 217274
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134306 216988 134334 217246
rect 135134 216988 135162 217246
rect 136008 217138 136036 218282
rect 136928 217274 136956 218282
rect 137664 217274 137692 219506
rect 138492 217274 138520 221138
rect 139320 217274 139348 228346
rect 140056 219434 140084 229055
rect 141160 227866 141188 231676
rect 141344 231662 141818 231690
rect 141148 227860 141200 227866
rect 141148 227802 141200 227808
rect 141344 225060 141372 231662
rect 141514 227896 141570 227905
rect 141514 227831 141516 227840
rect 141568 227831 141570 227840
rect 141516 227802 141568 227808
rect 142448 227050 142476 231676
rect 143092 228274 143120 231676
rect 143552 231662 143750 231690
rect 144012 231662 144394 231690
rect 143552 229129 143580 231662
rect 143538 229120 143594 229129
rect 143538 229055 143594 229064
rect 143080 228268 143132 228274
rect 143080 228210 143132 228216
rect 143448 228268 143500 228274
rect 143448 228210 143500 228216
rect 142436 227044 142488 227050
rect 142436 226986 142488 226992
rect 143264 227044 143316 227050
rect 143264 226986 143316 226992
rect 141606 226536 141662 226545
rect 141606 226471 141608 226480
rect 141660 226471 141662 226480
rect 142250 226536 142306 226545
rect 142250 226471 142252 226480
rect 141608 226442 141660 226448
rect 142304 226471 142306 226480
rect 142252 226442 142304 226448
rect 141792 226432 141844 226438
rect 141792 226374 141844 226380
rect 142114 226432 142166 226438
rect 142166 226380 142292 226386
rect 142114 226374 142292 226380
rect 140792 225032 141372 225060
rect 140792 221474 140820 225032
rect 140780 221468 140832 221474
rect 140780 221410 140832 221416
rect 140964 221468 141016 221474
rect 140964 221410 141016 221416
rect 139964 219406 140084 219434
rect 139964 218890 139992 219406
rect 139952 218884 140004 218890
rect 139952 218826 140004 218832
rect 140136 218884 140188 218890
rect 140136 218826 140188 218832
rect 140148 218498 140176 218826
rect 139964 218470 140176 218498
rect 139964 218346 139992 218470
rect 139952 218340 140004 218346
rect 139952 218282 140004 218288
rect 140136 218340 140188 218346
rect 140136 218282 140188 218288
rect 135962 217110 136036 217138
rect 136790 217246 136956 217274
rect 137618 217246 137692 217274
rect 138446 217246 138520 217274
rect 139274 217246 139348 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217246
rect 137618 216988 137646 217246
rect 138446 216988 138474 217246
rect 139274 216988 139302 217246
rect 140148 217138 140176 218282
rect 140976 217274 141004 221410
rect 141804 217274 141832 226374
rect 142126 226358 142292 226374
rect 142264 226166 142292 226358
rect 142114 226160 142166 226166
rect 142114 226102 142166 226108
rect 142252 226160 142304 226166
rect 142252 226102 142304 226108
rect 142126 225978 142154 226102
rect 142620 226024 142672 226030
rect 142618 225992 142620 226001
rect 142804 226024 142856 226030
rect 142672 225992 142674 226001
rect 142126 225950 142292 225978
rect 142264 225622 142292 225950
rect 142804 225966 142856 225972
rect 142618 225927 142674 225936
rect 142816 225706 142844 225966
rect 142448 225678 142844 225706
rect 142114 225616 142166 225622
rect 142114 225558 142166 225564
rect 142252 225616 142304 225622
rect 142252 225558 142304 225564
rect 142126 225434 142154 225558
rect 142448 225434 142476 225678
rect 142126 225406 142476 225434
rect 142126 224182 142476 224210
rect 142126 224126 142154 224182
rect 142114 224120 142166 224126
rect 142114 224062 142166 224068
rect 142252 224120 142304 224126
rect 142252 224062 142304 224068
rect 142264 223961 142292 224062
rect 142448 223961 142476 224182
rect 142250 223952 142306 223961
rect 142250 223887 142306 223896
rect 142434 223952 142490 223961
rect 142434 223887 142490 223896
rect 142114 223304 142166 223310
rect 142166 223272 142214 223281
rect 142114 223246 142158 223252
rect 142126 223230 142158 223246
rect 142158 223207 142214 223216
rect 142436 223168 142488 223174
rect 142436 223110 142488 223116
rect 141976 222896 142028 222902
rect 141974 222864 141976 222873
rect 142160 222896 142212 222902
rect 142028 222864 142030 222873
rect 142448 222873 142476 223110
rect 142160 222838 142212 222844
rect 142434 222864 142490 222873
rect 141974 222799 142030 222808
rect 142172 222714 142200 222838
rect 142434 222799 142490 222808
rect 141988 222686 142200 222714
rect 141988 222329 142016 222686
rect 141974 222320 142030 222329
rect 141974 222255 142030 222264
rect 142112 220960 142168 220969
rect 142112 220895 142114 220904
rect 142166 220895 142168 220904
rect 142252 220924 142304 220930
rect 142114 220866 142166 220872
rect 142252 220866 142304 220872
rect 142264 220504 142292 220866
rect 142126 220476 142292 220504
rect 142126 220386 142154 220476
rect 142114 220380 142166 220386
rect 142114 220322 142166 220328
rect 142252 220380 142304 220386
rect 142252 220322 142304 220328
rect 142264 219722 142292 220322
rect 142126 219706 142292 219722
rect 142114 219700 142292 219706
rect 142166 219694 142292 219700
rect 142114 219642 142166 219648
rect 142434 218512 142490 218521
rect 143276 218482 143304 226986
rect 142434 218447 142436 218456
rect 142488 218447 142490 218456
rect 142620 218476 142672 218482
rect 142436 218418 142488 218424
rect 142620 218418 142672 218424
rect 143264 218476 143316 218482
rect 143264 218418 143316 218424
rect 140102 217110 140176 217138
rect 140930 217246 141004 217274
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217246
rect 141758 216988 141786 217246
rect 142632 217138 142660 218418
rect 143460 217274 143488 228210
rect 144012 223174 144040 231662
rect 144642 230480 144698 230489
rect 144642 230415 144698 230424
rect 144458 229800 144514 229809
rect 144458 229735 144460 229744
rect 144512 229735 144514 229744
rect 144460 229706 144512 229712
rect 144000 223168 144052 223174
rect 144000 223110 144052 223116
rect 144656 220386 144684 230415
rect 144828 229764 144880 229770
rect 144828 229706 144880 229712
rect 144840 227186 144868 229706
rect 144828 227180 144880 227186
rect 144828 227122 144880 227128
rect 144644 220380 144696 220386
rect 144644 220322 144696 220328
rect 144276 219564 144328 219570
rect 144276 219506 144328 219512
rect 144288 217274 144316 219506
rect 145024 218754 145052 231676
rect 145668 229498 145696 231676
rect 146312 229770 146340 231676
rect 146680 231662 146970 231690
rect 146300 229764 146352 229770
rect 146300 229706 146352 229712
rect 145656 229492 145708 229498
rect 145656 229434 145708 229440
rect 146024 229424 146076 229430
rect 145838 229392 145894 229401
rect 146024 229366 146076 229372
rect 145838 229327 145840 229336
rect 145892 229327 145894 229336
rect 145840 229298 145892 229304
rect 146036 228274 146064 229366
rect 146208 228676 146260 228682
rect 146208 228618 146260 228624
rect 146220 228274 146248 228618
rect 146024 228268 146076 228274
rect 146024 228210 146076 228216
rect 146208 228268 146260 228274
rect 146208 228210 146260 228216
rect 146114 228032 146170 228041
rect 146114 227967 146170 227976
rect 145930 223000 145986 223009
rect 145930 222935 145986 222944
rect 145012 218748 145064 218754
rect 145012 218690 145064 218696
rect 145944 218482 145972 222935
rect 145104 218476 145156 218482
rect 145104 218418 145156 218424
rect 145932 218476 145984 218482
rect 145932 218418 145984 218424
rect 142586 217110 142660 217138
rect 143414 217246 143488 217274
rect 144242 217246 144316 217274
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144242 216988 144270 217246
rect 145116 217138 145144 218418
rect 146128 217274 146156 227967
rect 146680 223310 146708 231662
rect 147128 228540 147180 228546
rect 147128 228482 147180 228488
rect 147140 228041 147168 228482
rect 147126 228032 147182 228041
rect 147126 227967 147182 227976
rect 147600 226030 147628 231676
rect 147968 231662 148258 231690
rect 147968 229401 147996 231662
rect 148138 229800 148194 229809
rect 148138 229735 148194 229744
rect 148152 229634 148180 229735
rect 148140 229628 148192 229634
rect 148140 229570 148192 229576
rect 147954 229392 148010 229401
rect 147954 229327 148010 229336
rect 148138 229256 148194 229265
rect 148138 229191 148140 229200
rect 148192 229191 148194 229200
rect 148324 229220 148376 229226
rect 148140 229162 148192 229168
rect 148324 229162 148376 229168
rect 147588 226024 147640 226030
rect 147588 225966 147640 225972
rect 147772 226024 147824 226030
rect 147772 225966 147824 225972
rect 147784 225706 147812 225966
rect 147692 225678 147812 225706
rect 147692 225622 147720 225678
rect 147680 225616 147732 225622
rect 147680 225558 147732 225564
rect 146668 223304 146720 223310
rect 146668 223246 146720 223252
rect 146944 223304 146996 223310
rect 146944 223246 146996 223252
rect 146576 223168 146628 223174
rect 146576 223110 146628 223116
rect 146588 218521 146616 223110
rect 146956 223038 146984 223246
rect 146944 223032 146996 223038
rect 147128 223032 147180 223038
rect 146944 222974 146996 222980
rect 147126 223000 147128 223009
rect 147180 223000 147182 223009
rect 147126 222935 147182 222944
rect 148336 220930 148364 229162
rect 148888 228274 148916 231676
rect 148876 228268 148928 228274
rect 148876 228210 148928 228216
rect 148874 225448 148930 225457
rect 148874 225383 148930 225392
rect 148506 220960 148562 220969
rect 148324 220924 148376 220930
rect 148506 220895 148508 220904
rect 148324 220866 148376 220872
rect 148560 220895 148562 220904
rect 148508 220866 148560 220872
rect 146760 220788 146812 220794
rect 146760 220730 146812 220736
rect 146944 220788 146996 220794
rect 146944 220730 146996 220736
rect 146772 220386 146800 220730
rect 146956 220522 146984 220730
rect 146944 220516 146996 220522
rect 146944 220458 146996 220464
rect 147588 220516 147640 220522
rect 147588 220458 147640 220464
rect 146760 220380 146812 220386
rect 146760 220322 146812 220328
rect 146760 219428 146812 219434
rect 146760 219370 146812 219376
rect 146944 219428 146996 219434
rect 146944 219370 146996 219376
rect 146772 218906 146800 219370
rect 146956 219026 146984 219370
rect 146944 219020 146996 219026
rect 146944 218962 146996 218968
rect 147128 219020 147180 219026
rect 147128 218962 147180 218968
rect 147140 218906 147168 218962
rect 146772 218878 147168 218906
rect 146760 218748 146812 218754
rect 146760 218690 146812 218696
rect 146574 218512 146630 218521
rect 146574 218447 146630 218456
rect 145070 217110 145144 217138
rect 145898 217246 146156 217274
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146772 217138 146800 218690
rect 147600 217274 147628 220458
rect 148888 218482 148916 225383
rect 149532 223281 149560 231676
rect 149808 231662 150190 231690
rect 149808 226001 149836 231662
rect 150820 229634 150848 231676
rect 151096 231662 151478 231690
rect 151096 230489 151124 231662
rect 151082 230480 151138 230489
rect 151082 230415 151138 230424
rect 151452 229900 151504 229906
rect 151452 229842 151504 229848
rect 151636 229900 151688 229906
rect 151636 229842 151688 229848
rect 150808 229628 150860 229634
rect 150808 229570 150860 229576
rect 150992 229628 151044 229634
rect 150992 229570 151044 229576
rect 150346 229528 150402 229537
rect 150346 229463 150402 229472
rect 150072 227180 150124 227186
rect 150072 227122 150124 227128
rect 149794 225992 149850 226001
rect 149794 225927 149850 225936
rect 149518 223272 149574 223281
rect 149518 223207 149574 223216
rect 150084 218482 150112 227122
rect 150360 219434 150388 229463
rect 151004 229265 151032 229570
rect 151464 229362 151492 229842
rect 151452 229356 151504 229362
rect 151452 229298 151504 229304
rect 150990 229256 151046 229265
rect 150990 229191 151046 229200
rect 151648 227338 151676 229842
rect 151188 227310 151676 227338
rect 151188 220930 151216 227310
rect 151450 226264 151506 226273
rect 151450 226199 151506 226208
rect 151176 220924 151228 220930
rect 151176 220866 151228 220872
rect 150714 220552 150770 220561
rect 150714 220487 150716 220496
rect 150768 220487 150770 220496
rect 150900 220516 150952 220522
rect 150716 220458 150768 220464
rect 150900 220458 150952 220464
rect 150268 219406 150388 219434
rect 148416 218476 148468 218482
rect 148416 218418 148468 218424
rect 148876 218476 148928 218482
rect 148876 218418 148928 218424
rect 149244 218476 149296 218482
rect 149244 218418 149296 218424
rect 150072 218476 150124 218482
rect 150072 218418 150124 218424
rect 146726 217110 146800 217138
rect 147554 217246 147628 217274
rect 146726 216988 146754 217110
rect 147554 216988 147582 217246
rect 148428 217138 148456 218418
rect 149256 217138 149284 218418
rect 150268 217274 150296 219406
rect 150912 217274 150940 220458
rect 151464 219434 151492 226199
rect 151634 224496 151690 224505
rect 151634 224431 151690 224440
rect 151648 224262 151676 224431
rect 151636 224256 151688 224262
rect 151636 224198 151688 224204
rect 151774 224256 151826 224262
rect 151774 224198 151826 224204
rect 151786 224074 151814 224198
rect 151648 224046 151814 224074
rect 151648 223961 151676 224046
rect 151634 223952 151690 223961
rect 151634 223887 151690 223896
rect 152108 223310 152136 231676
rect 152384 231662 152766 231690
rect 152384 224505 152412 231662
rect 153396 229634 153424 231676
rect 153384 229628 153436 229634
rect 153384 229570 153436 229576
rect 154040 229226 154068 231676
rect 154698 231662 154988 231690
rect 154396 229628 154448 229634
rect 154396 229570 154448 229576
rect 154028 229220 154080 229226
rect 154028 229162 154080 229168
rect 154212 229220 154264 229226
rect 154212 229162 154264 229168
rect 153016 228404 153068 228410
rect 153016 228346 153068 228352
rect 152370 224496 152426 224505
rect 152370 224431 152426 224440
rect 152096 223304 152148 223310
rect 152096 223246 152148 223252
rect 151910 220552 151966 220561
rect 151910 220487 151912 220496
rect 151964 220487 151966 220496
rect 151912 220458 151964 220464
rect 151648 220386 151952 220402
rect 151636 220380 151952 220386
rect 151688 220374 151952 220380
rect 151636 220322 151688 220328
rect 151924 220250 151952 220374
rect 151728 220244 151780 220250
rect 151728 220186 151780 220192
rect 151912 220244 151964 220250
rect 151912 220186 151964 220192
rect 151740 220130 151768 220186
rect 152186 220144 152242 220153
rect 151740 220102 151860 220130
rect 151832 219881 151860 220102
rect 152186 220079 152188 220088
rect 152240 220079 152242 220088
rect 152372 220108 152424 220114
rect 152188 220050 152240 220056
rect 152372 220050 152424 220056
rect 151818 219872 151874 219881
rect 151818 219807 151874 219816
rect 152384 219434 152412 220050
rect 153028 219434 153056 228346
rect 154224 227202 154252 229162
rect 153856 227174 154252 227202
rect 153200 223576 153252 223582
rect 153200 223518 153252 223524
rect 153212 223310 153240 223518
rect 153200 223304 153252 223310
rect 153200 223246 153252 223252
rect 153856 220114 153884 227174
rect 154408 224954 154436 229570
rect 154040 224926 154436 224954
rect 154040 220250 154068 224926
rect 154960 223582 154988 231662
rect 155132 231464 155184 231470
rect 155132 231406 155184 231412
rect 154948 223576 155000 223582
rect 154948 223518 155000 223524
rect 154212 223440 154264 223446
rect 154212 223382 154264 223388
rect 154028 220244 154080 220250
rect 154028 220186 154080 220192
rect 153844 220108 153896 220114
rect 153844 220050 153896 220056
rect 151464 219406 151676 219434
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150296 217274
rect 150866 217246 150940 217274
rect 151648 217274 151676 219406
rect 152372 219428 152424 219434
rect 152372 219370 152424 219376
rect 152556 219428 152608 219434
rect 153028 219406 153148 219434
rect 152556 219370 152608 219376
rect 152568 218362 152596 219370
rect 152384 218334 152596 218362
rect 152384 218210 152412 218334
rect 152372 218204 152424 218210
rect 152372 218146 152424 218152
rect 153120 218142 153148 219406
rect 153384 218476 153436 218482
rect 153384 218418 153436 218424
rect 152556 218136 152608 218142
rect 152556 218078 152608 218084
rect 153108 218136 153160 218142
rect 153108 218078 153160 218084
rect 151648 217246 151722 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150866 216988 150894 217246
rect 151694 216988 151722 217246
rect 152568 217138 152596 218078
rect 153396 217138 153424 218418
rect 154224 217274 154252 223382
rect 155144 222766 155172 231406
rect 155328 224262 155356 231676
rect 155972 229362 156000 231676
rect 156156 231662 156630 231690
rect 156984 231662 157274 231690
rect 157918 231662 158208 231690
rect 155960 229356 156012 229362
rect 155960 229298 156012 229304
rect 155590 227080 155646 227089
rect 155590 227015 155646 227024
rect 155316 224256 155368 224262
rect 155316 224198 155368 224204
rect 155604 223122 155632 227015
rect 155776 223576 155828 223582
rect 155776 223518 155828 223524
rect 155788 223310 155816 223518
rect 155776 223304 155828 223310
rect 155776 223246 155828 223252
rect 155604 223094 155908 223122
rect 155132 222760 155184 222766
rect 155132 222702 155184 222708
rect 155684 222760 155736 222766
rect 155684 222702 155736 222708
rect 154396 220176 154448 220182
rect 154394 220144 154396 220153
rect 154448 220144 154450 220153
rect 154394 220079 154450 220088
rect 155696 218142 155724 222702
rect 155040 218136 155092 218142
rect 155040 218078 155092 218084
rect 155684 218136 155736 218142
rect 155684 218078 155736 218084
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217246 154252 217274
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217246
rect 155052 217138 155080 218078
rect 155880 217274 155908 223094
rect 156156 220182 156184 231662
rect 156420 231600 156472 231606
rect 156420 231542 156472 231548
rect 156432 225894 156460 231542
rect 156984 231470 157012 231662
rect 156972 231464 157024 231470
rect 156972 231406 157024 231412
rect 157248 231464 157300 231470
rect 157248 231406 157300 231412
rect 156786 230072 156842 230081
rect 156786 230007 156788 230016
rect 156840 230007 156842 230016
rect 156788 229978 156840 229984
rect 157260 229906 157288 231406
rect 157614 230208 157670 230217
rect 157614 230143 157616 230152
rect 157668 230143 157670 230152
rect 157800 230172 157852 230178
rect 157616 230114 157668 230120
rect 157800 230114 157852 230120
rect 157430 230072 157486 230081
rect 157430 230007 157432 230016
rect 157484 230007 157486 230016
rect 157432 229978 157484 229984
rect 157248 229900 157300 229906
rect 157248 229842 157300 229848
rect 156786 229800 156842 229809
rect 156786 229735 156788 229744
rect 156840 229735 156842 229744
rect 156788 229706 156840 229712
rect 157812 229362 157840 230114
rect 157982 229664 158038 229673
rect 157982 229599 157984 229608
rect 158036 229599 158038 229608
rect 157984 229570 158036 229576
rect 157800 229356 157852 229362
rect 157800 229298 157852 229304
rect 157984 229356 158036 229362
rect 157984 229298 158036 229304
rect 157338 227488 157394 227497
rect 157338 227423 157394 227432
rect 157352 227338 157380 227423
rect 157306 227322 157380 227338
rect 157294 227316 157380 227322
rect 157346 227310 157380 227316
rect 157524 227316 157576 227322
rect 157294 227258 157346 227264
rect 157524 227258 157576 227264
rect 157536 227089 157564 227258
rect 157522 227080 157578 227089
rect 157522 227015 157578 227024
rect 157154 226264 157210 226273
rect 157154 226199 157210 226208
rect 157168 226012 157196 226199
rect 157340 226024 157392 226030
rect 157168 225984 157340 226012
rect 157340 225966 157392 225972
rect 156420 225888 156472 225894
rect 156420 225830 156472 225836
rect 156602 225856 156658 225865
rect 156602 225791 156658 225800
rect 156616 225690 156644 225791
rect 156604 225684 156656 225690
rect 156604 225626 156656 225632
rect 157340 225616 157392 225622
rect 157168 225564 157340 225570
rect 157168 225558 157392 225564
rect 157168 225542 157380 225558
rect 157168 225457 157196 225542
rect 157154 225448 157210 225457
rect 157154 225383 157210 225392
rect 157248 224256 157300 224262
rect 157248 224198 157300 224204
rect 156788 223440 156840 223446
rect 156788 223382 156840 223388
rect 156420 223304 156472 223310
rect 156420 223246 156472 223252
rect 156432 222358 156460 223246
rect 156800 222902 156828 223382
rect 156604 222896 156656 222902
rect 156604 222838 156656 222844
rect 156788 222896 156840 222902
rect 156788 222838 156840 222844
rect 156420 222352 156472 222358
rect 156420 222294 156472 222300
rect 156616 222290 156644 222838
rect 156604 222284 156656 222290
rect 156604 222226 156656 222232
rect 156328 220244 156380 220250
rect 156328 220186 156380 220192
rect 156144 220176 156196 220182
rect 156144 220118 156196 220124
rect 156340 219881 156368 220186
rect 156326 219872 156382 219881
rect 156326 219807 156382 219816
rect 156236 219428 156288 219434
rect 156236 219370 156288 219376
rect 156420 219428 156472 219434
rect 156420 219370 156472 219376
rect 156248 218872 156276 219370
rect 156432 219026 156460 219370
rect 156420 219020 156472 219026
rect 156420 218962 156472 218968
rect 156788 218884 156840 218890
rect 156248 218844 156788 218872
rect 156788 218826 156840 218832
rect 157260 218142 157288 224198
rect 157432 222148 157484 222154
rect 157432 222090 157484 222096
rect 157444 221649 157472 222090
rect 157614 222048 157670 222057
rect 157614 221983 157616 221992
rect 157668 221983 157670 221992
rect 157616 221954 157668 221960
rect 157430 221640 157486 221649
rect 157430 221575 157486 221584
rect 157524 220108 157576 220114
rect 157524 220050 157576 220056
rect 156696 218136 156748 218142
rect 156696 218078 156748 218084
rect 157248 218136 157300 218142
rect 157248 218078 157300 218084
rect 155006 217110 155080 217138
rect 155834 217246 155908 217274
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156708 217138 156736 218078
rect 157536 217138 157564 220050
rect 157996 219162 158024 229298
rect 158180 225865 158208 231662
rect 158548 230178 158576 231676
rect 158916 231662 159206 231690
rect 158536 230172 158588 230178
rect 158536 230114 158588 230120
rect 158166 225856 158222 225865
rect 158166 225791 158222 225800
rect 158720 223440 158772 223446
rect 158720 223382 158772 223388
rect 158350 222048 158406 222057
rect 158350 221983 158352 221992
rect 158404 221983 158406 221992
rect 158352 221954 158404 221960
rect 158168 221876 158220 221882
rect 158168 221818 158220 221824
rect 158180 221649 158208 221818
rect 158166 221640 158222 221649
rect 158166 221575 158222 221584
rect 158352 220924 158404 220930
rect 158352 220866 158404 220872
rect 157984 219156 158036 219162
rect 157984 219098 158036 219104
rect 158364 217138 158392 220866
rect 158732 218890 158760 223382
rect 158916 220250 158944 231662
rect 159362 228848 159418 228857
rect 159362 228783 159364 228792
rect 159416 228783 159418 228792
rect 159364 228754 159416 228760
rect 159836 223582 159864 231676
rect 160006 228440 160062 228449
rect 160006 228375 160062 228384
rect 159824 223576 159876 223582
rect 159824 223518 159876 223524
rect 158904 220244 158956 220250
rect 158904 220186 158956 220192
rect 160020 219434 160048 228375
rect 160480 224534 160508 231676
rect 160756 231662 161138 231690
rect 160756 229634 160784 231662
rect 161768 231470 161796 231676
rect 161952 231662 162426 231690
rect 162688 231662 163070 231690
rect 161756 231464 161808 231470
rect 161756 231406 161808 231412
rect 160744 229628 160796 229634
rect 160744 229570 160796 229576
rect 160928 229628 160980 229634
rect 160928 229570 160980 229576
rect 160468 224528 160520 224534
rect 160468 224470 160520 224476
rect 160940 224262 160968 229570
rect 161664 224528 161716 224534
rect 161664 224470 161716 224476
rect 160928 224256 160980 224262
rect 160928 224198 160980 224204
rect 160836 221604 160888 221610
rect 160836 221546 160888 221552
rect 160650 220960 160706 220969
rect 160848 220930 160876 221546
rect 161018 221232 161074 221241
rect 161018 221167 161074 221176
rect 160650 220895 160652 220904
rect 160704 220895 160706 220904
rect 160836 220924 160888 220930
rect 160652 220866 160704 220872
rect 160836 220866 160888 220872
rect 158996 219428 159048 219434
rect 158996 219370 159048 219376
rect 159180 219428 159232 219434
rect 159180 219370 159232 219376
rect 160008 219428 160060 219434
rect 160008 219370 160060 219376
rect 159008 218890 159036 219370
rect 158720 218884 158772 218890
rect 158720 218826 158772 218832
rect 158996 218884 159048 218890
rect 158996 218826 159048 218832
rect 159192 217138 159220 219370
rect 160008 218204 160060 218210
rect 160008 218146 160060 218152
rect 160020 217138 160048 218146
rect 161032 217274 161060 221167
rect 156662 217110 156736 217138
rect 157490 217110 157564 217138
rect 158318 217110 158392 217138
rect 159146 217110 159220 217138
rect 159974 217110 160048 217138
rect 160802 217246 161060 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217110
rect 158318 216988 158346 217110
rect 159146 216988 159174 217110
rect 159974 216988 160002 217110
rect 160802 216988 160830 217246
rect 161676 217138 161704 224470
rect 161952 223310 161980 231662
rect 162688 231606 162716 231662
rect 162676 231600 162728 231606
rect 162676 231542 162728 231548
rect 162306 230208 162362 230217
rect 162306 230143 162362 230152
rect 162492 230172 162544 230178
rect 162320 229906 162348 230143
rect 162492 230114 162544 230120
rect 162308 229900 162360 229906
rect 162308 229842 162360 229848
rect 162124 229764 162176 229770
rect 162124 229706 162176 229712
rect 162136 229226 162164 229706
rect 162504 229401 162532 230114
rect 162490 229392 162546 229401
rect 163700 229362 163728 231676
rect 163964 229764 164016 229770
rect 163964 229706 164016 229712
rect 162490 229327 162546 229336
rect 163688 229356 163740 229362
rect 163688 229298 163740 229304
rect 162124 229220 162176 229226
rect 162124 229162 162176 229168
rect 162490 228848 162546 228857
rect 162490 228783 162546 228792
rect 162676 228812 162728 228818
rect 162504 228682 162532 228783
rect 162676 228754 162728 228760
rect 162308 228676 162360 228682
rect 162308 228618 162360 228624
rect 162492 228676 162544 228682
rect 162492 228618 162544 228624
rect 162320 228562 162348 228618
rect 162688 228562 162716 228754
rect 162320 228534 162716 228562
rect 161940 223304 161992 223310
rect 161940 223246 161992 223252
rect 162492 223304 162544 223310
rect 162492 223246 162544 223252
rect 161952 223094 162348 223122
rect 161952 222766 161980 223094
rect 162320 223038 162348 223094
rect 162124 223032 162176 223038
rect 162124 222974 162176 222980
rect 162308 223032 162360 223038
rect 162308 222974 162360 222980
rect 162136 222766 162164 222974
rect 161940 222760 161992 222766
rect 161940 222702 161992 222708
rect 162124 222760 162176 222766
rect 162124 222702 162176 222708
rect 162124 221604 162176 221610
rect 162124 221546 162176 221552
rect 162136 221202 162164 221546
rect 162306 221232 162362 221241
rect 162124 221196 162176 221202
rect 162306 221167 162308 221176
rect 162124 221138 162176 221144
rect 162360 221167 162362 221176
rect 162308 221138 162360 221144
rect 162504 219586 162532 223246
rect 162228 219558 162532 219586
rect 162228 218618 162256 219558
rect 163976 219434 164004 229706
rect 164344 220930 164372 231676
rect 164988 222494 165016 231676
rect 165632 224670 165660 231676
rect 166276 229906 166304 231676
rect 166552 231662 166934 231690
rect 167196 231662 167578 231690
rect 167840 231662 168222 231690
rect 168576 231662 168866 231690
rect 169128 231662 169510 231690
rect 169772 231662 170154 231690
rect 166264 229900 166316 229906
rect 166264 229842 166316 229848
rect 166552 227497 166580 231662
rect 166816 229356 166868 229362
rect 166816 229298 166868 229304
rect 166828 228682 166856 229298
rect 166816 228676 166868 228682
rect 166816 228618 166868 228624
rect 166954 228676 167006 228682
rect 166954 228618 167006 228624
rect 166966 228562 166994 228618
rect 166828 228534 166994 228562
rect 166828 228449 166856 228534
rect 166814 228440 166870 228449
rect 166814 228375 166870 228384
rect 166538 227488 166594 227497
rect 166538 227423 166594 227432
rect 165620 224664 165672 224670
rect 165620 224606 165672 224612
rect 165160 224256 165212 224262
rect 165160 224198 165212 224204
rect 164976 222488 165028 222494
rect 164976 222430 165028 222436
rect 164514 220960 164570 220969
rect 164332 220924 164384 220930
rect 164514 220895 164516 220904
rect 164332 220866 164384 220872
rect 164568 220895 164570 220904
rect 164516 220866 164568 220872
rect 164148 220244 164200 220250
rect 164148 220186 164200 220192
rect 162400 219428 162452 219434
rect 162400 219370 162452 219376
rect 163320 219428 163372 219434
rect 163320 219370 163372 219376
rect 163964 219428 164016 219434
rect 163964 219370 164016 219376
rect 162412 219162 162440 219370
rect 162400 219156 162452 219162
rect 162400 219098 162452 219104
rect 162676 219020 162728 219026
rect 162676 218962 162728 218968
rect 162216 218612 162268 218618
rect 162216 218554 162268 218560
rect 162492 218612 162544 218618
rect 162492 218554 162544 218560
rect 162504 217138 162532 218554
rect 162688 218210 162716 218962
rect 162676 218204 162728 218210
rect 162676 218146 162728 218152
rect 163332 217138 163360 219370
rect 164160 217138 164188 220186
rect 165172 217274 165200 224198
rect 165620 223576 165672 223582
rect 165620 223518 165672 223524
rect 165632 219162 165660 223518
rect 166814 222048 166870 222057
rect 166814 221983 166816 221992
rect 166868 221983 166870 221992
rect 166998 222048 167054 222057
rect 166998 221983 167000 221992
rect 166816 221954 166868 221960
rect 167052 221983 167054 221992
rect 167000 221954 167052 221960
rect 167196 221746 167224 231662
rect 167840 224398 167868 231662
rect 167828 224392 167880 224398
rect 167828 224334 167880 224340
rect 168288 224392 168340 224398
rect 168288 224334 168340 224340
rect 167184 221740 167236 221746
rect 167184 221682 167236 221688
rect 167460 221740 167512 221746
rect 167460 221682 167512 221688
rect 165620 219156 165672 219162
rect 165620 219098 165672 219104
rect 165804 219156 165856 219162
rect 165804 219098 165856 219104
rect 161630 217110 161704 217138
rect 162458 217110 162532 217138
rect 163286 217110 163360 217138
rect 164114 217110 164188 217138
rect 164942 217246 165200 217274
rect 161630 216988 161658 217110
rect 162458 216988 162486 217110
rect 163286 216988 163314 217110
rect 164114 216988 164142 217110
rect 164942 216988 164970 217246
rect 165816 217138 165844 219098
rect 166632 218204 166684 218210
rect 166632 218146 166684 218152
rect 166644 217138 166672 218146
rect 167472 217138 167500 221682
rect 168300 217138 168328 224334
rect 168576 217326 168604 231662
rect 169128 229362 169156 231662
rect 169116 229356 169168 229362
rect 169116 229298 169168 229304
rect 169574 227216 169630 227225
rect 169574 227151 169630 227160
rect 169588 219298 169616 227151
rect 169772 222018 169800 231662
rect 170784 231198 170812 231676
rect 170772 231192 170824 231198
rect 170772 231134 170824 231140
rect 171428 230790 171456 231676
rect 171704 231662 172086 231690
rect 171416 230784 171468 230790
rect 171416 230726 171468 230732
rect 170956 229356 171008 229362
rect 170956 229298 171008 229304
rect 170770 227488 170826 227497
rect 170770 227423 170772 227432
rect 170824 227423 170826 227432
rect 170772 227394 170824 227400
rect 169760 222012 169812 222018
rect 169760 221954 169812 221960
rect 170968 219298 170996 229298
rect 171704 227497 171732 231662
rect 171690 227488 171746 227497
rect 171094 227452 171146 227458
rect 171690 227423 171746 227432
rect 171094 227394 171146 227400
rect 171106 227225 171134 227394
rect 171092 227216 171148 227225
rect 171092 227151 171148 227160
rect 171968 223576 172020 223582
rect 171968 223518 172020 223524
rect 171600 223168 171652 223174
rect 171600 223110 171652 223116
rect 171784 223168 171836 223174
rect 171784 223110 171836 223116
rect 171612 222630 171640 223110
rect 171796 222766 171824 223110
rect 171980 222766 172008 223518
rect 171784 222760 171836 222766
rect 171784 222702 171836 222708
rect 171968 222760 172020 222766
rect 171968 222702 172020 222708
rect 171600 222624 171652 222630
rect 171600 222566 171652 222572
rect 172242 222456 172298 222465
rect 172242 222391 172298 222400
rect 171784 222012 171836 222018
rect 171784 221954 171836 221960
rect 171416 221740 171468 221746
rect 171416 221682 171468 221688
rect 171600 221740 171652 221746
rect 171600 221682 171652 221688
rect 171428 221377 171456 221682
rect 171414 221368 171470 221377
rect 171414 221303 171470 221312
rect 169116 219292 169168 219298
rect 169116 219234 169168 219240
rect 169576 219292 169628 219298
rect 169576 219234 169628 219240
rect 169944 219292 169996 219298
rect 169944 219234 169996 219240
rect 170956 219292 171008 219298
rect 170956 219234 171008 219240
rect 171416 219292 171468 219298
rect 171416 219234 171468 219240
rect 168564 217320 168616 217326
rect 168564 217262 168616 217268
rect 169128 217138 169156 219234
rect 169956 217138 169984 219234
rect 171428 218890 171456 219234
rect 171416 218884 171468 218890
rect 171416 218826 171468 218832
rect 170588 218340 170640 218346
rect 170588 218282 170640 218288
rect 170772 218340 170824 218346
rect 170772 218282 170824 218288
rect 170600 218074 170628 218282
rect 170588 218068 170640 218074
rect 170588 218010 170640 218016
rect 170784 217138 170812 218282
rect 171612 217138 171640 221682
rect 171796 221338 171824 221954
rect 171966 221368 172022 221377
rect 171784 221332 171836 221338
rect 171966 221303 171968 221312
rect 171784 221274 171836 221280
rect 172020 221303 172022 221312
rect 171968 221274 172020 221280
rect 172256 219298 172284 222391
rect 172716 222154 172744 231676
rect 172992 231662 173374 231690
rect 174018 231662 174216 231690
rect 172992 224942 173020 231662
rect 173900 229764 173952 229770
rect 173900 229706 173952 229712
rect 173912 229226 173940 229706
rect 173900 229220 173952 229226
rect 173900 229162 173952 229168
rect 173162 228848 173218 228857
rect 173162 228783 173218 228792
rect 172980 224936 173032 224942
rect 172980 224878 173032 224884
rect 172704 222148 172756 222154
rect 172704 222090 172756 222096
rect 173176 219298 173204 228783
rect 174188 224954 174216 231662
rect 174648 228954 174676 231676
rect 175306 231662 175596 231690
rect 175568 229094 175596 231662
rect 175752 231662 175950 231690
rect 175752 229094 175780 231662
rect 175924 229764 175976 229770
rect 175924 229706 175976 229712
rect 176384 229764 176436 229770
rect 176384 229706 176436 229712
rect 175936 229226 175964 229706
rect 175924 229220 175976 229226
rect 175924 229162 175976 229168
rect 175384 229066 175596 229094
rect 175660 229066 175780 229094
rect 174636 228948 174688 228954
rect 174636 228890 174688 228896
rect 175186 227624 175242 227633
rect 175186 227559 175188 227568
rect 175240 227559 175242 227568
rect 175188 227530 175240 227536
rect 175384 224954 175412 229066
rect 174188 224926 174308 224954
rect 175384 224926 175504 224954
rect 174084 222148 174136 222154
rect 174084 222090 174136 222096
rect 172244 219292 172296 219298
rect 172244 219234 172296 219240
rect 172428 219292 172480 219298
rect 172428 219234 172480 219240
rect 173164 219292 173216 219298
rect 173164 219234 173216 219240
rect 171784 218884 171836 218890
rect 171784 218826 171836 218832
rect 171796 218618 171824 218826
rect 171784 218612 171836 218618
rect 171784 218554 171836 218560
rect 171968 218612 172020 218618
rect 171968 218554 172020 218560
rect 171980 218074 172008 218554
rect 171968 218068 172020 218074
rect 171968 218010 172020 218016
rect 172440 217138 172468 219234
rect 173256 218068 173308 218074
rect 173256 218010 173308 218016
rect 173268 217138 173296 218010
rect 174096 217138 174124 222090
rect 174280 217938 174308 224926
rect 174912 224664 174964 224670
rect 174912 224606 174964 224612
rect 174268 217932 174320 217938
rect 174268 217874 174320 217880
rect 174924 217138 174952 224606
rect 175280 223576 175332 223582
rect 175280 223518 175332 223524
rect 175292 222630 175320 223518
rect 175280 222624 175332 222630
rect 175280 222566 175332 222572
rect 175476 220658 175504 224926
rect 175660 222494 175688 229066
rect 176106 228848 176162 228857
rect 176106 228783 176108 228792
rect 176160 228783 176162 228792
rect 176108 228754 176160 228760
rect 175924 227520 175976 227526
rect 175924 227462 175976 227468
rect 175936 227361 175964 227462
rect 175922 227352 175978 227361
rect 175922 227287 175978 227296
rect 176016 222556 176068 222562
rect 176016 222498 176068 222504
rect 175648 222488 175700 222494
rect 175648 222430 175700 222436
rect 175830 222456 175886 222465
rect 175830 222391 175832 222400
rect 175884 222391 175886 222400
rect 175832 222362 175884 222368
rect 175464 220652 175516 220658
rect 175464 220594 175516 220600
rect 175740 219292 175792 219298
rect 175740 219234 175792 219240
rect 175752 217138 175780 219234
rect 176028 218618 176056 222498
rect 176016 218612 176068 218618
rect 176016 218554 176068 218560
rect 176396 217274 176424 229706
rect 176580 223582 176608 231676
rect 177224 227633 177252 231676
rect 177408 231662 177882 231690
rect 177210 227624 177266 227633
rect 177210 227559 177266 227568
rect 176750 227352 176806 227361
rect 176750 227287 176752 227296
rect 176804 227287 176806 227296
rect 176752 227258 176804 227264
rect 176568 223576 176620 223582
rect 176568 223518 176620 223524
rect 177408 221921 177436 231662
rect 178512 224942 178540 231676
rect 179156 230654 179184 231676
rect 179144 230648 179196 230654
rect 179144 230590 179196 230596
rect 179800 229090 179828 231676
rect 180444 229226 180472 231676
rect 180432 229220 180484 229226
rect 180432 229162 180484 229168
rect 179788 229084 179840 229090
rect 179788 229026 179840 229032
rect 180064 229084 180116 229090
rect 180064 229026 180116 229032
rect 178500 224936 178552 224942
rect 178500 224878 178552 224884
rect 178684 224936 178736 224942
rect 178684 224878 178736 224884
rect 178040 224800 178092 224806
rect 178040 224742 178092 224748
rect 176566 221912 176622 221921
rect 176566 221847 176568 221856
rect 176620 221847 176622 221856
rect 177394 221912 177450 221921
rect 177394 221847 177450 221856
rect 176568 221818 176620 221824
rect 176566 220688 176622 220697
rect 176566 220623 176622 220632
rect 177396 220652 177448 220658
rect 176580 218346 176608 220623
rect 177396 220594 177448 220600
rect 176568 218340 176620 218346
rect 176568 218282 176620 218288
rect 177408 217274 177436 220594
rect 178052 219434 178080 224742
rect 178696 224670 178724 224878
rect 178684 224664 178736 224670
rect 178684 224606 178736 224612
rect 179328 224664 179380 224670
rect 179328 224606 179380 224612
rect 178040 219428 178092 219434
rect 178040 219370 178092 219376
rect 178224 219428 178276 219434
rect 178224 219370 178276 219376
rect 178236 218226 178264 219370
rect 179052 218340 179104 218346
rect 179052 218282 179104 218288
rect 178052 218198 178264 218226
rect 178052 218074 178080 218198
rect 178040 218068 178092 218074
rect 178040 218010 178092 218016
rect 178224 218068 178276 218074
rect 178224 218010 178276 218016
rect 176396 217246 176562 217274
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 168254 217110 168328 217138
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217110 170812 217138
rect 171566 217110 171640 217138
rect 172394 217110 172468 217138
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217110 174952 217138
rect 175706 217110 175780 217138
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217110
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217110
rect 171566 216988 171594 217110
rect 172394 216988 172422 217110
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217110
rect 175706 216988 175734 217110
rect 176534 216988 176562 217246
rect 177362 217246 177436 217274
rect 177362 216988 177390 217246
rect 178236 217138 178264 218010
rect 179064 217138 179092 218282
rect 179340 218074 179368 224606
rect 180076 219162 180104 229026
rect 181088 223990 181116 231676
rect 181536 227588 181588 227594
rect 181536 227530 181588 227536
rect 181076 223984 181128 223990
rect 181076 223926 181128 223932
rect 181260 222148 181312 222154
rect 181260 222090 181312 222096
rect 181272 221882 181300 222090
rect 181548 222034 181576 227530
rect 181732 223446 181760 231676
rect 182376 227730 182404 231676
rect 182652 231662 183034 231690
rect 183678 231662 183876 231690
rect 182364 227724 182416 227730
rect 182364 227666 182416 227672
rect 181720 223440 181772 223446
rect 181720 223382 181772 223388
rect 182652 222154 182680 231662
rect 183376 229220 183428 229226
rect 183376 229162 183428 229168
rect 182640 222148 182692 222154
rect 182640 222090 182692 222096
rect 181456 222006 181576 222034
rect 181260 221876 181312 221882
rect 181260 221818 181312 221824
rect 180798 220960 180854 220969
rect 180798 220895 180854 220904
rect 180812 220810 180840 220895
rect 180766 220794 180840 220810
rect 180754 220788 180840 220794
rect 180806 220782 180840 220788
rect 180904 220794 181300 220810
rect 180904 220788 181312 220794
rect 180904 220782 181260 220788
rect 180754 220730 180806 220736
rect 180904 220674 180932 220782
rect 181260 220730 181312 220736
rect 180812 220658 180932 220674
rect 180800 220652 180932 220658
rect 180852 220646 180932 220652
rect 181074 220688 181130 220697
rect 181074 220623 181076 220632
rect 180800 220594 180852 220600
rect 181128 220623 181130 220632
rect 181076 220594 181128 220600
rect 181456 219434 181484 222006
rect 181628 221876 181680 221882
rect 181628 221818 181680 221824
rect 181640 219434 181668 221818
rect 183388 219434 183416 229162
rect 183652 225888 183704 225894
rect 183652 225830 183704 225836
rect 180708 219428 180760 219434
rect 180708 219370 180760 219376
rect 181364 219406 181484 219434
rect 181548 219406 181668 219434
rect 183204 219406 183416 219434
rect 183664 219434 183692 225830
rect 183848 223854 183876 231662
rect 184112 227588 184164 227594
rect 184112 227530 184164 227536
rect 184124 226914 184152 227530
rect 184112 226908 184164 226914
rect 184112 226850 184164 226856
rect 184308 225758 184336 231676
rect 184952 228970 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 186608 231662 186898 231690
rect 185136 229094 185164 231662
rect 185584 230172 185636 230178
rect 185584 230114 185636 230120
rect 185398 229936 185454 229945
rect 185398 229871 185454 229880
rect 185412 229770 185440 229871
rect 185596 229770 185624 230114
rect 185400 229764 185452 229770
rect 185400 229706 185452 229712
rect 185584 229764 185636 229770
rect 185584 229706 185636 229712
rect 184860 228954 184980 228970
rect 184848 228948 184980 228954
rect 184900 228942 184980 228948
rect 185044 229066 185164 229094
rect 185872 229094 185900 231662
rect 186044 230172 186096 230178
rect 186044 230114 186096 230120
rect 186056 229945 186084 230114
rect 186042 229936 186098 229945
rect 186042 229871 186098 229880
rect 185584 229084 185636 229090
rect 184848 228890 184900 228896
rect 184296 225752 184348 225758
rect 184296 225694 184348 225700
rect 183836 223848 183888 223854
rect 183836 223790 183888 223796
rect 184848 223712 184900 223718
rect 184848 223654 184900 223660
rect 184664 223440 184716 223446
rect 184664 223382 184716 223388
rect 183664 219406 183784 219434
rect 180064 219156 180116 219162
rect 180064 219098 180116 219104
rect 179512 218884 179564 218890
rect 179512 218826 179564 218832
rect 179524 218074 179552 218826
rect 179880 218612 179932 218618
rect 179880 218554 179932 218560
rect 179328 218068 179380 218074
rect 179328 218010 179380 218016
rect 179512 218068 179564 218074
rect 179512 218010 179564 218016
rect 179892 217138 179920 218554
rect 180720 217138 180748 219370
rect 181364 218074 181392 219406
rect 181352 218068 181404 218074
rect 181352 218010 181404 218016
rect 181548 217274 181576 219406
rect 182364 218884 182416 218890
rect 182364 218826 182416 218832
rect 178190 217110 178264 217138
rect 179018 217110 179092 217138
rect 179846 217110 179920 217138
rect 180674 217110 180748 217138
rect 181502 217246 181576 217274
rect 178190 216988 178218 217110
rect 179018 216988 179046 217110
rect 179846 216988 179874 217110
rect 180674 216988 180702 217110
rect 181502 216988 181530 217246
rect 182376 217138 182404 218826
rect 183204 217274 183232 219406
rect 183756 218754 183784 219406
rect 183744 218748 183796 218754
rect 183744 218690 183796 218696
rect 184676 218074 184704 223382
rect 184020 218068 184072 218074
rect 184020 218010 184072 218016
rect 184664 218068 184716 218074
rect 184664 218010 184716 218016
rect 182330 217110 182404 217138
rect 183158 217246 183232 217274
rect 182330 216988 182358 217110
rect 183158 216988 183186 217246
rect 184032 217138 184060 218010
rect 184860 217274 184888 223654
rect 185044 220969 185072 229066
rect 185872 229066 185992 229094
rect 185584 229026 185636 229032
rect 185216 228948 185268 228954
rect 185216 228890 185268 228896
rect 185228 228138 185256 228890
rect 185596 228682 185624 229026
rect 185400 228676 185452 228682
rect 185400 228618 185452 228624
rect 185584 228676 185636 228682
rect 185584 228618 185636 228624
rect 185412 228138 185440 228618
rect 185216 228132 185268 228138
rect 185216 228074 185268 228080
rect 185400 228132 185452 228138
rect 185400 228074 185452 228080
rect 185228 227854 185624 227882
rect 185228 227730 185256 227854
rect 185216 227724 185268 227730
rect 185216 227666 185268 227672
rect 185400 227724 185452 227730
rect 185400 227666 185452 227672
rect 185412 226778 185440 227666
rect 185596 227610 185624 227854
rect 185596 227582 185808 227610
rect 185780 227458 185808 227582
rect 185584 227452 185636 227458
rect 185584 227394 185636 227400
rect 185768 227452 185820 227458
rect 185768 227394 185820 227400
rect 185596 226914 185624 227394
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 185400 226772 185452 226778
rect 185400 226714 185452 226720
rect 185412 224998 185808 225026
rect 185412 224670 185440 224998
rect 185780 224942 185808 224998
rect 185584 224936 185636 224942
rect 185584 224878 185636 224884
rect 185768 224936 185820 224942
rect 185768 224878 185820 224884
rect 185596 224670 185624 224878
rect 185400 224664 185452 224670
rect 185400 224606 185452 224612
rect 185584 224664 185636 224670
rect 185584 224606 185636 224612
rect 185964 223854 185992 229066
rect 186136 226772 186188 226778
rect 186136 226714 186188 226720
rect 185952 223848 186004 223854
rect 185952 223790 186004 223796
rect 185400 223304 185452 223310
rect 185400 223246 185452 223252
rect 185412 222766 185440 223246
rect 185584 223168 185636 223174
rect 185584 223110 185636 223116
rect 185596 222766 185624 223110
rect 185400 222760 185452 222766
rect 185400 222702 185452 222708
rect 185584 222760 185636 222766
rect 185584 222702 185636 222708
rect 185030 220960 185086 220969
rect 185030 220895 185086 220904
rect 185858 220824 185914 220833
rect 185858 220759 185914 220768
rect 185872 219434 185900 220759
rect 185860 219428 185912 219434
rect 185860 219370 185912 219376
rect 186148 218074 186176 226714
rect 186608 223582 186636 231662
rect 187528 227594 187556 231676
rect 188172 230926 188200 231676
rect 188448 231662 188830 231690
rect 189092 231662 189474 231690
rect 188160 230920 188212 230926
rect 188160 230862 188212 230868
rect 187516 227588 187568 227594
rect 187516 227530 187568 227536
rect 186964 223848 187016 223854
rect 186964 223790 187016 223796
rect 186596 223576 186648 223582
rect 186596 223518 186648 223524
rect 186504 219428 186556 219434
rect 186504 219370 186556 219376
rect 185676 218068 185728 218074
rect 185676 218010 185728 218016
rect 186136 218068 186188 218074
rect 186136 218010 186188 218016
rect 183986 217110 184060 217138
rect 184814 217246 184888 217274
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185688 217138 185716 218010
rect 186516 217138 186544 219370
rect 186976 218482 187004 223790
rect 187332 223576 187384 223582
rect 187332 223518 187384 223524
rect 186964 218476 187016 218482
rect 186964 218418 187016 218424
rect 187344 217274 187372 223518
rect 188448 219434 188476 231662
rect 189092 229094 189120 231662
rect 189092 229066 189212 229094
rect 188896 223304 188948 223310
rect 188896 223246 188948 223252
rect 187988 219406 188476 219434
rect 187988 217462 188016 219406
rect 188712 218476 188764 218482
rect 188712 218418 188764 218424
rect 188160 218068 188212 218074
rect 188160 218010 188212 218016
rect 187976 217456 188028 217462
rect 187976 217398 188028 217404
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217246 187372 217274
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217246
rect 188172 217138 188200 218010
rect 188724 217274 188752 218418
rect 188908 218074 188936 223246
rect 188896 218068 188948 218074
rect 188896 218010 188948 218016
rect 189184 217598 189212 229066
rect 189724 229084 189776 229090
rect 189724 229026 189776 229032
rect 189736 218890 189764 229026
rect 190104 228954 190132 231676
rect 190656 231662 190762 231690
rect 191024 231662 191406 231690
rect 190092 228948 190144 228954
rect 190092 228890 190144 228896
rect 189908 227588 189960 227594
rect 189908 227530 189960 227536
rect 189920 219162 189948 227530
rect 190412 220824 190468 220833
rect 190276 220788 190328 220794
rect 190412 220759 190414 220768
rect 190276 220730 190328 220736
rect 190466 220759 190468 220768
rect 190414 220730 190466 220736
rect 190288 220130 190316 220730
rect 190288 220102 190454 220130
rect 190274 220008 190330 220017
rect 190426 219978 190454 220102
rect 190656 220017 190684 231662
rect 191024 222222 191052 231662
rect 192036 223174 192064 231676
rect 192484 229084 192536 229090
rect 192484 229026 192536 229032
rect 192496 227866 192524 229026
rect 192484 227860 192536 227866
rect 192484 227802 192536 227808
rect 192680 227730 192708 231676
rect 193324 230194 193352 231676
rect 193324 230166 193444 230194
rect 193034 228984 193090 228993
rect 193034 228919 193090 228928
rect 192668 227724 192720 227730
rect 192668 227666 192720 227672
rect 192024 223168 192076 223174
rect 192024 223110 192076 223116
rect 191012 222216 191064 222222
rect 191012 222158 191064 222164
rect 191472 222148 191524 222154
rect 191472 222090 191524 222096
rect 190642 220008 190698 220017
rect 190274 219943 190276 219952
rect 190328 219943 190330 219952
rect 190414 219972 190466 219978
rect 190276 219914 190328 219920
rect 190642 219943 190698 219952
rect 190414 219914 190466 219920
rect 189908 219156 189960 219162
rect 189908 219098 189960 219104
rect 190644 219156 190696 219162
rect 190644 219098 190696 219104
rect 189724 218884 189776 218890
rect 189724 218826 189776 218832
rect 189816 218068 189868 218074
rect 189816 218010 189868 218016
rect 189172 217592 189224 217598
rect 189172 217534 189224 217540
rect 188724 217246 188982 217274
rect 188126 217110 188200 217138
rect 188126 216988 188154 217110
rect 188954 216988 188982 217246
rect 189828 217138 189856 218010
rect 190656 217138 190684 219098
rect 191484 217274 191512 222090
rect 192852 218884 192904 218890
rect 192852 218826 192904 218832
rect 192116 218748 192168 218754
rect 192116 218690 192168 218696
rect 192128 218074 192156 218690
rect 192116 218068 192168 218074
rect 192116 218010 192168 218016
rect 192300 218068 192352 218074
rect 192300 218010 192352 218016
rect 189782 217110 189856 217138
rect 190610 217110 190684 217138
rect 191438 217246 191512 217274
rect 189782 216988 189810 217110
rect 190610 216988 190638 217110
rect 191438 216988 191466 217246
rect 192312 217138 192340 218010
rect 192864 217274 192892 218826
rect 193048 218074 193076 228919
rect 193416 221066 193444 230166
rect 193968 226302 193996 231676
rect 194416 230648 194468 230654
rect 194416 230590 194468 230596
rect 194428 230314 194456 230590
rect 194416 230308 194468 230314
rect 194416 230250 194468 230256
rect 193956 226296 194008 226302
rect 193956 226238 194008 226244
rect 194140 226296 194192 226302
rect 194140 226238 194192 226244
rect 193404 221060 193456 221066
rect 193404 221002 193456 221008
rect 194152 219434 194180 226238
rect 194612 224126 194640 231676
rect 194876 230308 194928 230314
rect 194876 230250 194928 230256
rect 194888 229770 194916 230250
rect 195060 230036 195112 230042
rect 195060 229978 195112 229984
rect 195072 229770 195100 229978
rect 194876 229764 194928 229770
rect 194876 229706 194928 229712
rect 195060 229764 195112 229770
rect 195060 229706 195112 229712
rect 195256 229094 195284 231676
rect 195900 231062 195928 231676
rect 196176 231662 196558 231690
rect 196912 231662 197202 231690
rect 197372 231662 197846 231690
rect 198016 231662 198490 231690
rect 195888 231056 195940 231062
rect 195888 230998 195940 231004
rect 195428 230308 195480 230314
rect 195428 230250 195480 230256
rect 195612 230308 195664 230314
rect 195612 230250 195664 230256
rect 195440 230042 195468 230250
rect 195428 230036 195480 230042
rect 195428 229978 195480 229984
rect 195072 229066 195284 229094
rect 195072 227866 195100 229066
rect 195426 228984 195482 228993
rect 195244 228948 195296 228954
rect 195426 228919 195428 228928
rect 195244 228890 195296 228896
rect 195480 228919 195482 228928
rect 195428 228890 195480 228896
rect 195256 228138 195284 228890
rect 195244 228132 195296 228138
rect 195244 228074 195296 228080
rect 195060 227860 195112 227866
rect 195060 227802 195112 227808
rect 195244 227724 195296 227730
rect 195244 227666 195296 227672
rect 195256 226778 195284 227666
rect 195244 226772 195296 226778
rect 195244 226714 195296 226720
rect 195244 224936 195296 224942
rect 195244 224878 195296 224884
rect 195428 224936 195480 224942
rect 195428 224878 195480 224884
rect 195256 224126 195284 224878
rect 194600 224120 194652 224126
rect 194600 224062 194652 224068
rect 195244 224120 195296 224126
rect 195244 224062 195296 224068
rect 195440 223718 195468 224878
rect 195428 223712 195480 223718
rect 195428 223654 195480 223660
rect 194324 223168 194376 223174
rect 194324 223110 194376 223116
rect 194336 222358 194364 223110
rect 194324 222352 194376 222358
rect 194324 222294 194376 222300
rect 194508 222352 194560 222358
rect 194508 222294 194560 222300
rect 193784 219406 194180 219434
rect 193784 218482 193812 219406
rect 193772 218476 193824 218482
rect 193772 218418 193824 218424
rect 194520 218074 194548 222294
rect 195624 219434 195652 230250
rect 196176 225486 196204 231662
rect 196912 230654 196940 231662
rect 196900 230648 196952 230654
rect 196900 230590 196952 230596
rect 197372 226642 197400 231662
rect 198016 229094 198044 231662
rect 197648 229066 198044 229094
rect 197360 226636 197412 226642
rect 197360 226578 197412 226584
rect 196164 225480 196216 225486
rect 196164 225422 196216 225428
rect 196348 225480 196400 225486
rect 196348 225422 196400 225428
rect 195888 223712 195940 223718
rect 195888 223654 195940 223660
rect 195256 219406 195652 219434
rect 195256 218754 195284 219406
rect 195244 218748 195296 218754
rect 195244 218690 195296 218696
rect 195612 218476 195664 218482
rect 195612 218418 195664 218424
rect 193036 218068 193088 218074
rect 193036 218010 193088 218016
rect 193956 218068 194008 218074
rect 193956 218010 194008 218016
rect 194508 218068 194560 218074
rect 194508 218010 194560 218016
rect 194784 218068 194836 218074
rect 194784 218010 194836 218016
rect 192864 217246 193122 217274
rect 192266 217110 192340 217138
rect 192266 216988 192294 217110
rect 193094 216988 193122 217246
rect 193968 217138 193996 218010
rect 194796 217138 194824 218010
rect 195624 217138 195652 218418
rect 195900 218074 195928 223654
rect 196360 219434 196388 225422
rect 197176 222624 197228 222630
rect 197176 222566 197228 222572
rect 196268 219406 196388 219434
rect 196268 218346 196296 219406
rect 196256 218340 196308 218346
rect 196256 218282 196308 218288
rect 195888 218068 195940 218074
rect 195888 218010 195940 218016
rect 196440 218068 196492 218074
rect 196440 218010 196492 218016
rect 196452 217138 196480 218010
rect 197188 217274 197216 222566
rect 197648 219842 197676 229066
rect 198004 225888 198056 225894
rect 198004 225830 198056 225836
rect 197636 219836 197688 219842
rect 197636 219778 197688 219784
rect 197820 219836 197872 219842
rect 197820 219778 197872 219784
rect 197832 219162 197860 219778
rect 197820 219156 197872 219162
rect 197820 219098 197872 219104
rect 198016 218482 198044 225830
rect 199120 225350 199148 231676
rect 199108 225344 199160 225350
rect 199108 225286 199160 225292
rect 199764 223174 199792 231676
rect 200408 229090 200436 231676
rect 201052 230518 201080 231676
rect 201040 230512 201092 230518
rect 201040 230454 201092 230460
rect 200396 229084 200448 229090
rect 200396 229026 200448 229032
rect 201408 229084 201460 229090
rect 201408 229026 201460 229032
rect 200396 228540 200448 228546
rect 200396 228482 200448 228488
rect 200408 228002 200436 228482
rect 200396 227996 200448 228002
rect 200396 227938 200448 227944
rect 200028 226772 200080 226778
rect 200028 226714 200080 226720
rect 199752 223168 199804 223174
rect 199752 223110 199804 223116
rect 200040 218890 200068 226714
rect 201224 223984 201276 223990
rect 201224 223926 201276 223932
rect 201236 219434 201264 223926
rect 201236 219406 201356 219434
rect 198924 218884 198976 218890
rect 198924 218826 198976 218832
rect 200028 218884 200080 218890
rect 200028 218826 200080 218832
rect 200212 218884 200264 218890
rect 200212 218826 200264 218832
rect 198004 218476 198056 218482
rect 198004 218418 198056 218424
rect 198280 218476 198332 218482
rect 198280 218418 198332 218424
rect 198096 218340 198148 218346
rect 198096 218282 198148 218288
rect 197188 217246 197262 217274
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217110 195652 217138
rect 196406 217110 196480 217138
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217110
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198108 217138 198136 218282
rect 198292 218074 198320 218418
rect 198280 218068 198332 218074
rect 198280 218010 198332 218016
rect 198936 217138 198964 218826
rect 200224 218770 200252 218826
rect 199764 218742 200252 218770
rect 199764 217274 199792 218742
rect 200580 218204 200632 218210
rect 200580 218146 200632 218152
rect 198062 217110 198136 217138
rect 198890 217110 198964 217138
rect 199718 217246 199792 217274
rect 198062 216988 198090 217110
rect 198890 216988 198918 217110
rect 199718 216988 199746 217246
rect 200592 217138 200620 218146
rect 201328 217274 201356 219406
rect 201420 218226 201448 229026
rect 201696 225078 201724 231676
rect 202340 229770 202368 231676
rect 202328 229764 202380 229770
rect 202328 229706 202380 229712
rect 202984 226506 203012 231676
rect 203168 231662 203642 231690
rect 202972 226500 203024 226506
rect 202972 226442 203024 226448
rect 201684 225072 201736 225078
rect 201684 225014 201736 225020
rect 202696 225072 202748 225078
rect 202696 225014 202748 225020
rect 202512 221604 202564 221610
rect 202512 221546 202564 221552
rect 202524 221066 202552 221546
rect 202512 221060 202564 221066
rect 202512 221002 202564 221008
rect 201420 218210 201540 218226
rect 202708 218210 202736 225014
rect 203168 219706 203196 231662
rect 204076 227044 204128 227050
rect 204076 226986 204128 226992
rect 204088 226642 204116 226986
rect 204076 226636 204128 226642
rect 204076 226578 204128 226584
rect 203524 226500 203576 226506
rect 203524 226442 203576 226448
rect 203156 219700 203208 219706
rect 203156 219642 203208 219648
rect 203536 219026 203564 226442
rect 204272 225214 204300 231676
rect 204640 231662 204930 231690
rect 204640 229094 204668 231662
rect 204904 230308 204956 230314
rect 204904 230250 204956 230256
rect 204916 229770 204944 230250
rect 204904 229764 204956 229770
rect 204904 229706 204956 229712
rect 204548 229066 204668 229094
rect 204260 225208 204312 225214
rect 204260 225150 204312 225156
rect 204548 224806 204576 229066
rect 204904 228540 204956 228546
rect 204904 228482 204956 228488
rect 204916 227866 204944 228482
rect 205560 228274 205588 231676
rect 205744 231662 206218 231690
rect 206388 231662 206862 231690
rect 205548 228268 205600 228274
rect 205548 228210 205600 228216
rect 204904 227860 204956 227866
rect 204904 227802 204956 227808
rect 205456 227860 205508 227866
rect 205456 227802 205508 227808
rect 205088 227588 205140 227594
rect 205088 227530 205140 227536
rect 205272 227588 205324 227594
rect 205272 227530 205324 227536
rect 205100 226914 205128 227530
rect 205088 226908 205140 226914
rect 205088 226850 205140 226856
rect 205284 226778 205312 227530
rect 205272 226772 205324 226778
rect 205272 226714 205324 226720
rect 205088 225888 205140 225894
rect 205088 225830 205140 225836
rect 204720 225752 204772 225758
rect 204720 225694 204772 225700
rect 204732 225486 204760 225694
rect 204720 225480 204772 225486
rect 204720 225422 204772 225428
rect 205100 225350 205128 225830
rect 205088 225344 205140 225350
rect 205088 225286 205140 225292
rect 204536 224800 204588 224806
rect 204536 224742 204588 224748
rect 204720 224800 204772 224806
rect 204720 224742 204772 224748
rect 204732 224210 204760 224742
rect 204640 224182 204760 224210
rect 204640 224126 204668 224182
rect 204628 224120 204680 224126
rect 204628 224062 204680 224068
rect 205088 223984 205140 223990
rect 205088 223926 205140 223932
rect 205100 223718 205128 223926
rect 205088 223712 205140 223718
rect 205088 223654 205140 223660
rect 204260 223168 204312 223174
rect 204260 223110 204312 223116
rect 204272 222766 204300 223110
rect 204260 222760 204312 222766
rect 204260 222702 204312 222708
rect 204444 222760 204496 222766
rect 204444 222702 204496 222708
rect 204456 222358 204484 222702
rect 204444 222352 204496 222358
rect 204444 222294 204496 222300
rect 204168 221332 204220 221338
rect 204168 221274 204220 221280
rect 203892 219564 203944 219570
rect 203892 219506 203944 219512
rect 203524 219020 203576 219026
rect 203524 218962 203576 218968
rect 201420 218204 201552 218210
rect 201420 218198 201500 218204
rect 201500 218146 201552 218152
rect 202236 218204 202288 218210
rect 202236 218146 202288 218152
rect 202696 218204 202748 218210
rect 202696 218146 202748 218152
rect 203064 218204 203116 218210
rect 203064 218146 203116 218152
rect 201328 217246 201402 217274
rect 200546 217110 200620 217138
rect 200546 216988 200574 217110
rect 201374 216988 201402 217246
rect 202248 217138 202276 218146
rect 203076 217138 203104 218146
rect 203904 217274 203932 219506
rect 204180 218346 204208 221274
rect 204168 218340 204220 218346
rect 204168 218282 204220 218288
rect 204720 218340 204772 218346
rect 204720 218282 204772 218288
rect 202202 217110 202276 217138
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 202202 216988 202230 217110
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218282
rect 205468 217274 205496 227802
rect 205744 221610 205772 231662
rect 205916 228268 205968 228274
rect 205916 228210 205968 228216
rect 205928 227866 205956 228210
rect 205916 227860 205968 227866
rect 205916 227802 205968 227808
rect 205732 221604 205784 221610
rect 205732 221546 205784 221552
rect 206388 221066 206416 231662
rect 206560 230308 206612 230314
rect 206560 230250 206612 230256
rect 206376 221060 206428 221066
rect 206376 221002 206428 221008
rect 206572 219434 206600 230250
rect 207492 222494 207520 231676
rect 208136 226642 208164 231676
rect 208596 231662 208794 231690
rect 208124 226636 208176 226642
rect 208124 226578 208176 226584
rect 208124 225344 208176 225350
rect 208124 225286 208176 225292
rect 207480 222488 207532 222494
rect 207480 222430 207532 222436
rect 207664 222488 207716 222494
rect 207664 222430 207716 222436
rect 206296 219406 206600 219434
rect 206296 218210 206324 219406
rect 206468 219020 206520 219026
rect 206468 218962 206520 218968
rect 206284 218204 206336 218210
rect 206284 218146 206336 218152
rect 206480 217274 206508 218962
rect 207676 218346 207704 222430
rect 207664 218340 207716 218346
rect 207664 218282 207716 218288
rect 208136 218210 208164 225286
rect 208400 221604 208452 221610
rect 208400 221546 208452 221552
rect 208412 219434 208440 221546
rect 208596 219706 208624 231662
rect 209424 226166 209452 231676
rect 210068 229498 210096 231676
rect 210056 229492 210108 229498
rect 210056 229434 210108 229440
rect 210712 228002 210740 231676
rect 210700 227996 210752 228002
rect 210700 227938 210752 227944
rect 210332 227860 210384 227866
rect 210332 227802 210384 227808
rect 209412 226160 209464 226166
rect 209412 226102 209464 226108
rect 209688 226160 209740 226166
rect 209688 226102 209740 226108
rect 208584 219700 208636 219706
rect 208584 219642 208636 219648
rect 208320 219406 208440 219434
rect 207204 218204 207256 218210
rect 207204 218146 207256 218152
rect 208124 218204 208176 218210
rect 208124 218146 208176 218152
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206342 217246 206508 217274
rect 206342 216988 206370 217246
rect 207216 217138 207244 218146
rect 208320 217274 208348 219406
rect 209700 219162 209728 226102
rect 208860 219156 208912 219162
rect 208860 219098 208912 219104
rect 209688 219156 209740 219162
rect 209688 219098 209740 219104
rect 207170 217110 207244 217138
rect 207998 217246 208348 217274
rect 207170 216988 207198 217110
rect 207998 216988 208026 217246
rect 208872 217138 208900 219098
rect 210344 218618 210372 227802
rect 211356 220522 211384 231676
rect 212000 223174 212028 231676
rect 212552 231662 212658 231690
rect 212172 226636 212224 226642
rect 212172 226578 212224 226584
rect 211988 223168 212040 223174
rect 211988 223110 212040 223116
rect 211804 222352 211856 222358
rect 211804 222294 211856 222300
rect 211344 220516 211396 220522
rect 211344 220458 211396 220464
rect 210516 219700 210568 219706
rect 210516 219642 210568 219648
rect 210332 218612 210384 218618
rect 210332 218554 210384 218560
rect 209688 218340 209740 218346
rect 209688 218282 209740 218288
rect 209700 217138 209728 218282
rect 210528 217274 210556 219642
rect 211344 218204 211396 218210
rect 211344 218146 211396 218152
rect 208826 217110 208900 217138
rect 209654 217110 209728 217138
rect 210482 217246 210556 217274
rect 208826 216988 208854 217110
rect 209654 216988 209682 217110
rect 210482 216988 210510 217246
rect 211356 217138 211384 218146
rect 211816 218074 211844 222294
rect 211804 218068 211856 218074
rect 211804 218010 211856 218016
rect 212184 217274 212212 226578
rect 212552 225486 212580 231662
rect 213092 230444 213144 230450
rect 213092 230386 213144 230392
rect 212540 225480 212592 225486
rect 212540 225422 212592 225428
rect 213104 219434 213132 230386
rect 213288 227186 213316 231676
rect 213946 231662 214144 231690
rect 213276 227180 213328 227186
rect 213276 227122 213328 227128
rect 213828 226500 213880 226506
rect 213828 226442 213880 226448
rect 213644 220380 213696 220386
rect 213644 220322 213696 220328
rect 213656 219978 213684 220322
rect 213644 219972 213696 219978
rect 213644 219914 213696 219920
rect 212828 219406 213132 219434
rect 212828 218346 212856 219406
rect 212816 218340 212868 218346
rect 212816 218282 212868 218288
rect 213000 218340 213052 218346
rect 213000 218282 213052 218288
rect 211310 217110 211384 217138
rect 212138 217246 212212 217274
rect 211310 216988 211338 217110
rect 212138 216988 212166 217246
rect 213012 217138 213040 218282
rect 213840 217274 213868 226442
rect 214116 220522 214144 231662
rect 214380 227180 214432 227186
rect 214380 227122 214432 227128
rect 214392 226914 214420 227122
rect 214380 226908 214432 226914
rect 214380 226850 214432 226856
rect 214576 225622 214604 231676
rect 215220 230042 215248 231676
rect 215208 230036 215260 230042
rect 215208 229978 215260 229984
rect 215864 228410 215892 231676
rect 216232 231662 216522 231690
rect 215852 228404 215904 228410
rect 215852 228346 215904 228352
rect 214760 227854 215156 227882
rect 214760 227730 214788 227854
rect 214748 227724 214800 227730
rect 214748 227666 214800 227672
rect 214932 227724 214984 227730
rect 214932 227666 214984 227672
rect 214944 226642 214972 227666
rect 215128 227050 215156 227854
rect 215116 227044 215168 227050
rect 215116 226986 215168 226992
rect 214932 226636 214984 226642
rect 214932 226578 214984 226584
rect 214564 225616 214616 225622
rect 214564 225558 214616 225564
rect 215208 225616 215260 225622
rect 215208 225558 215260 225564
rect 214104 220516 214156 220522
rect 214104 220458 214156 220464
rect 214288 220516 214340 220522
rect 214288 220458 214340 220464
rect 214300 220114 214328 220458
rect 214288 220108 214340 220114
rect 214288 220050 214340 220056
rect 214748 219972 214800 219978
rect 214748 219914 214800 219920
rect 214760 219570 214788 219914
rect 214748 219564 214800 219570
rect 214748 219506 214800 219512
rect 215220 218074 215248 225558
rect 216232 223174 216260 231662
rect 216496 228404 216548 228410
rect 216496 228346 216548 228352
rect 215392 223168 215444 223174
rect 215392 223110 215444 223116
rect 216220 223168 216272 223174
rect 216220 223110 216272 223116
rect 215404 222902 215432 223110
rect 215392 222896 215444 222902
rect 215392 222838 215444 222844
rect 215944 222896 215996 222902
rect 215944 222838 215996 222844
rect 215956 219298 215984 222838
rect 215944 219292 215996 219298
rect 215944 219234 215996 219240
rect 216312 218340 216364 218346
rect 216312 218282 216364 218288
rect 214656 218068 214708 218074
rect 214656 218010 214708 218016
rect 215208 218068 215260 218074
rect 215208 218010 215260 218016
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214668 217138 214696 218010
rect 215496 217138 215524 218010
rect 216324 217138 216352 218282
rect 216508 218074 216536 228346
rect 217152 226030 217180 231676
rect 217140 226024 217192 226030
rect 217140 225966 217192 225972
rect 217796 223854 217824 231676
rect 218440 226914 218468 231676
rect 218716 231662 219098 231690
rect 218428 226908 218480 226914
rect 218428 226850 218480 226856
rect 217784 223848 217836 223854
rect 217784 223790 217836 223796
rect 218716 220522 218744 231662
rect 219348 226636 219400 226642
rect 219348 226578 219400 226584
rect 218704 220516 218756 220522
rect 218704 220458 218756 220464
rect 217140 219700 217192 219706
rect 217140 219642 217192 219648
rect 216496 218068 216548 218074
rect 216496 218010 216548 218016
rect 217152 217274 217180 219642
rect 219360 219162 219388 226578
rect 219728 223038 219756 231676
rect 220372 229634 220400 231676
rect 220360 229628 220412 229634
rect 220360 229570 220412 229576
rect 220084 229492 220136 229498
rect 220084 229434 220136 229440
rect 219716 223032 219768 223038
rect 219716 222974 219768 222980
rect 219808 221060 219860 221066
rect 219808 221002 219860 221008
rect 219624 219292 219676 219298
rect 219624 219234 219676 219240
rect 218796 219156 218848 219162
rect 218796 219098 218848 219104
rect 219348 219156 219400 219162
rect 219348 219098 219400 219104
rect 217968 218204 218020 218210
rect 217968 218146 218020 218152
rect 214622 217110 214696 217138
rect 215450 217110 215524 217138
rect 216278 217110 216352 217138
rect 217106 217246 217180 217274
rect 214622 216988 214650 217110
rect 215450 216988 215478 217110
rect 216278 216988 216306 217110
rect 217106 216988 217134 217246
rect 217980 217138 218008 218146
rect 218808 217138 218836 219098
rect 219636 217138 219664 219234
rect 219820 218074 219848 221002
rect 220096 218618 220124 229434
rect 221016 228546 221044 231676
rect 221292 231662 221674 231690
rect 221004 228540 221056 228546
rect 221004 228482 221056 228488
rect 221292 221202 221320 231662
rect 221830 226808 221886 226817
rect 221830 226743 221886 226752
rect 221280 221196 221332 221202
rect 221280 221138 221332 221144
rect 220452 219564 220504 219570
rect 220452 219506 220504 219512
rect 220084 218612 220136 218618
rect 220084 218554 220136 218560
rect 219808 218068 219860 218074
rect 219808 218010 219860 218016
rect 220464 217274 220492 219506
rect 221844 218074 221872 226743
rect 222016 226024 222068 226030
rect 222016 225966 222068 225972
rect 221280 218068 221332 218074
rect 221280 218010 221332 218016
rect 221832 218068 221884 218074
rect 221832 218010 221884 218016
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218010
rect 222028 217274 222056 225966
rect 222304 220930 222332 231676
rect 222476 227316 222528 227322
rect 222476 227258 222528 227264
rect 222488 226914 222516 227258
rect 222476 226908 222528 226914
rect 222476 226850 222528 226856
rect 222948 226778 222976 231676
rect 223592 227458 223620 231676
rect 223776 231662 224250 231690
rect 223776 229094 223804 231662
rect 223776 229066 223896 229094
rect 223580 227452 223632 227458
rect 223580 227394 223632 227400
rect 223118 226808 223174 226817
rect 222936 226772 222988 226778
rect 223118 226743 223120 226752
rect 222936 226714 222988 226720
rect 223172 226743 223174 226752
rect 223120 226714 223172 226720
rect 222752 221196 222804 221202
rect 222752 221138 222804 221144
rect 222292 220924 222344 220930
rect 222292 220866 222344 220872
rect 222764 218210 222792 221138
rect 223672 220516 223724 220522
rect 223672 220458 223724 220464
rect 223684 219706 223712 220458
rect 223868 220250 223896 229066
rect 224684 228404 224736 228410
rect 224684 228346 224736 228352
rect 224224 227452 224276 227458
rect 224224 227394 224276 227400
rect 224040 227180 224092 227186
rect 224040 227122 224092 227128
rect 224052 226506 224080 227122
rect 224236 227050 224264 227394
rect 224224 227044 224276 227050
rect 224224 226986 224276 226992
rect 224040 226500 224092 226506
rect 224040 226442 224092 226448
rect 224696 223938 224724 228346
rect 224880 224534 224908 231676
rect 225524 229906 225552 231676
rect 225512 229900 225564 229906
rect 225512 229842 225564 229848
rect 225696 229900 225748 229906
rect 225696 229842 225748 229848
rect 224868 224528 224920 224534
rect 224868 224470 224920 224476
rect 224696 223910 224816 223938
rect 224592 223848 224644 223854
rect 224592 223790 224644 223796
rect 224224 220652 224276 220658
rect 224224 220594 224276 220600
rect 223856 220244 223908 220250
rect 223856 220186 223908 220192
rect 223672 219700 223724 219706
rect 223672 219642 223724 219648
rect 224236 219570 224264 220594
rect 224408 220380 224460 220386
rect 224408 220322 224460 220328
rect 224420 219706 224448 220322
rect 224408 219700 224460 219706
rect 224408 219642 224460 219648
rect 224224 219564 224276 219570
rect 224224 219506 224276 219512
rect 224408 219428 224460 219434
rect 224408 219370 224460 219376
rect 224224 219156 224276 219162
rect 224224 219098 224276 219104
rect 224236 218482 224264 219098
rect 224420 218482 224448 219370
rect 224224 218476 224276 218482
rect 224224 218418 224276 218424
rect 224408 218476 224460 218482
rect 224408 218418 224460 218424
rect 222752 218204 222804 218210
rect 222752 218146 222804 218152
rect 222936 218204 222988 218210
rect 222936 218146 222988 218152
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218146
rect 224604 218074 224632 223790
rect 223764 218068 223816 218074
rect 223764 218010 223816 218016
rect 224592 218068 224644 218074
rect 224592 218010 224644 218016
rect 223776 217138 223804 218010
rect 224788 217274 224816 223910
rect 225708 219434 225736 229842
rect 226168 228682 226196 231676
rect 226536 231662 226826 231690
rect 226156 228676 226208 228682
rect 226156 228618 226208 228624
rect 226340 228676 226392 228682
rect 226340 228618 226392 228624
rect 226352 228562 226380 228618
rect 225616 219406 225736 219434
rect 226168 228534 226380 228562
rect 225616 218210 225644 219406
rect 225972 218612 226024 218618
rect 225972 218554 226024 218560
rect 225604 218204 225656 218210
rect 225604 218146 225656 218152
rect 225420 218068 225472 218074
rect 225420 218010 225472 218016
rect 222902 217110 222976 217138
rect 223730 217110 223804 217138
rect 224558 217246 224816 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217110
rect 224558 216988 224586 217246
rect 225432 217138 225460 218010
rect 225984 217274 226012 218554
rect 226168 218074 226196 228534
rect 226536 221474 226564 231662
rect 227456 224262 227484 231676
rect 227444 224256 227496 224262
rect 227444 224198 227496 224204
rect 228100 222358 228128 231676
rect 228744 226914 228772 231676
rect 229296 231662 229402 231690
rect 228732 226908 228784 226914
rect 228732 226850 228784 226856
rect 228732 224528 228784 224534
rect 228732 224470 228784 224476
rect 228088 222352 228140 222358
rect 228088 222294 228140 222300
rect 226524 221468 226576 221474
rect 226524 221410 226576 221416
rect 227904 221468 227956 221474
rect 227904 221410 227956 221416
rect 227076 219700 227128 219706
rect 227076 219642 227128 219648
rect 226156 218068 226208 218074
rect 226156 218010 226208 218016
rect 227088 217274 227116 219642
rect 227916 217274 227944 221410
rect 228744 217274 228772 224470
rect 229296 219570 229324 231662
rect 230032 224398 230060 231676
rect 230480 230036 230532 230042
rect 230480 229978 230532 229984
rect 230020 224392 230072 224398
rect 230020 224334 230072 224340
rect 230492 223666 230520 229978
rect 230676 229362 230704 231676
rect 230664 229356 230716 229362
rect 230664 229298 230716 229304
rect 231320 228818 231348 231676
rect 231872 231662 231978 231690
rect 232240 231662 232622 231690
rect 231308 228812 231360 228818
rect 231308 228754 231360 228760
rect 231032 226772 231084 226778
rect 231032 226714 231084 226720
rect 230400 223638 230520 223666
rect 230204 223032 230256 223038
rect 230204 222974 230256 222980
rect 229284 219564 229336 219570
rect 229284 219506 229336 219512
rect 230216 219434 230244 222974
rect 230400 219434 230428 223638
rect 229560 219428 229612 219434
rect 230216 219406 230336 219434
rect 230400 219428 230532 219434
rect 230400 219406 230480 219428
rect 229560 219370 229612 219376
rect 225984 217246 226242 217274
rect 225386 217110 225460 217138
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227042 217246 227116 217274
rect 227870 217246 227944 217274
rect 228698 217246 228772 217274
rect 227042 216988 227070 217246
rect 227870 216988 227898 217246
rect 228698 216988 228726 217246
rect 229572 217138 229600 219370
rect 230308 217274 230336 219406
rect 230480 219370 230532 219376
rect 231044 218482 231072 226714
rect 231676 224256 231728 224262
rect 231676 224198 231728 224204
rect 231032 218476 231084 218482
rect 231032 218418 231084 218424
rect 231688 218074 231716 224198
rect 231872 222018 231900 231662
rect 231860 222012 231912 222018
rect 231860 221954 231912 221960
rect 232240 221746 232268 231662
rect 233252 229094 233280 231676
rect 233252 229066 233372 229094
rect 233148 224392 233200 224398
rect 233148 224334 233200 224340
rect 232228 221740 232280 221746
rect 232228 221682 232280 221688
rect 232872 218340 232924 218346
rect 232872 218282 232924 218288
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 230308 217246 230382 217274
rect 229526 217110 229600 217138
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217274 232912 218282
rect 233160 218074 233188 224334
rect 233344 222902 233372 229066
rect 233896 227322 233924 231676
rect 234172 231662 234554 231690
rect 233884 227316 233936 227322
rect 233884 227258 233936 227264
rect 233332 222896 233384 222902
rect 233332 222838 233384 222844
rect 233700 222012 233752 222018
rect 233700 221954 233752 221960
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233712 217274 233740 221954
rect 234172 220250 234200 231662
rect 235184 224670 235212 231676
rect 235828 230178 235856 231676
rect 235816 230172 235868 230178
rect 235816 230114 235868 230120
rect 235816 227316 235868 227322
rect 235816 227258 235868 227264
rect 235172 224664 235224 224670
rect 235172 224606 235224 224612
rect 234528 222896 234580 222902
rect 234528 222838 234580 222844
rect 234160 220244 234212 220250
rect 234160 220186 234212 220192
rect 234540 217274 234568 222838
rect 235828 218074 235856 227258
rect 236472 225894 236500 231676
rect 236656 231662 237130 231690
rect 236460 225888 236512 225894
rect 236460 225830 236512 225836
rect 236656 220794 236684 231662
rect 237288 225888 237340 225894
rect 237288 225830 237340 225836
rect 236644 220788 236696 220794
rect 236644 220730 236696 220736
rect 237012 220244 237064 220250
rect 237012 220186 237064 220192
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235816 218068 235868 218074
rect 235816 218010 235868 218016
rect 236184 218068 236236 218074
rect 236184 218010 236236 218016
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217246 232912 217274
rect 233666 217246 233740 217274
rect 234494 217246 234568 217274
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217246
rect 233666 216988 233694 217246
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217138 236224 218010
rect 237024 217274 237052 220186
rect 237300 218074 237328 225830
rect 237760 224806 237788 231676
rect 238404 228002 238432 231676
rect 239048 228138 239076 231676
rect 239036 228132 239088 228138
rect 239036 228074 239088 228080
rect 238392 227996 238444 228002
rect 238392 227938 238444 227944
rect 238668 227996 238720 228002
rect 238668 227938 238720 227944
rect 237748 224800 237800 224806
rect 237748 224742 237800 224748
rect 238024 223712 238076 223718
rect 238024 223654 238076 223660
rect 237840 219428 237892 219434
rect 237840 219370 237892 219376
rect 237288 218068 237340 218074
rect 237288 218010 237340 218016
rect 235322 217110 235396 217138
rect 236150 217110 236224 217138
rect 236978 217246 237052 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217110
rect 236978 216988 237006 217246
rect 237852 217138 237880 219370
rect 238036 218482 238064 223654
rect 238024 218476 238076 218482
rect 238024 218418 238076 218424
rect 238680 217274 238708 227938
rect 239692 223446 239720 231676
rect 240152 231662 240350 231690
rect 239680 223440 239732 223446
rect 239680 223382 239732 223388
rect 240152 221882 240180 231662
rect 240324 230172 240376 230178
rect 240324 230114 240376 230120
rect 240336 225894 240364 230114
rect 240980 229226 241008 231676
rect 240968 229220 241020 229226
rect 240968 229162 241020 229168
rect 241624 227458 241652 231676
rect 241612 227452 241664 227458
rect 241612 227394 241664 227400
rect 240324 225888 240376 225894
rect 240324 225830 240376 225836
rect 241152 225344 241204 225350
rect 241152 225286 241204 225292
rect 240140 221876 240192 221882
rect 240140 221818 240192 221824
rect 239312 221740 239364 221746
rect 239312 221682 239364 221688
rect 239324 219434 239352 221682
rect 239312 219428 239364 219434
rect 239312 219370 239364 219376
rect 239496 219428 239548 219434
rect 239496 219370 239548 219376
rect 237806 217110 237880 217138
rect 238634 217246 238708 217274
rect 237806 216988 237834 217110
rect 238634 216988 238662 217246
rect 239508 217138 239536 219370
rect 240324 218068 240376 218074
rect 240324 218010 240376 218016
rect 240336 217138 240364 218010
rect 241164 217274 241192 225286
rect 242268 223582 242296 231676
rect 242716 225208 242768 225214
rect 242716 225150 242768 225156
rect 242256 223576 242308 223582
rect 242256 223518 242308 223524
rect 241336 223168 241388 223174
rect 241336 223110 241388 223116
rect 241348 218074 241376 223110
rect 242728 220946 242756 225150
rect 242912 224942 242940 231676
rect 243280 231662 243570 231690
rect 243280 226778 243308 231662
rect 243268 226772 243320 226778
rect 243268 226714 243320 226720
rect 243452 226704 243504 226710
rect 243452 226646 243504 226652
rect 242900 224936 242952 224942
rect 242900 224878 242952 224884
rect 242728 220918 242848 220946
rect 242624 220788 242676 220794
rect 242624 220730 242676 220736
rect 242636 219434 242664 220730
rect 242820 219434 242848 220918
rect 241796 219428 241848 219434
rect 241796 219370 241848 219376
rect 241980 219428 242032 219434
rect 242636 219406 242756 219434
rect 242820 219428 242952 219434
rect 242820 219406 242900 219428
rect 241980 219370 242032 219376
rect 241808 218890 241836 219370
rect 241612 218884 241664 218890
rect 241612 218826 241664 218832
rect 241796 218884 241848 218890
rect 241796 218826 241848 218832
rect 241624 218346 241652 218826
rect 241612 218340 241664 218346
rect 241612 218282 241664 218288
rect 241336 218068 241388 218074
rect 241336 218010 241388 218016
rect 239462 217110 239536 217138
rect 240290 217110 240364 217138
rect 241118 217246 241192 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217110
rect 241118 216988 241146 217246
rect 241992 217138 242020 219370
rect 242728 217274 242756 219406
rect 242900 219370 242952 219376
rect 243464 218754 243492 226646
rect 244200 226302 244228 231676
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 244476 229094 244504 231662
rect 244384 229066 244504 229094
rect 244188 226296 244240 226302
rect 244188 226238 244240 226244
rect 244096 223440 244148 223446
rect 244096 223382 244148 223388
rect 243452 218748 243504 218754
rect 243452 218690 243504 218696
rect 244108 218074 244136 223382
rect 244384 220266 244412 229066
rect 245120 223310 245148 231662
rect 246132 229770 246160 231676
rect 246120 229764 246172 229770
rect 246120 229706 246172 229712
rect 246488 229764 246540 229770
rect 246488 229706 246540 229712
rect 246304 228812 246356 228818
rect 246304 228754 246356 228760
rect 245292 224800 245344 224806
rect 245292 224742 245344 224748
rect 245108 223304 245160 223310
rect 245108 223246 245160 223252
rect 244292 220238 244412 220266
rect 244292 220114 244320 220238
rect 244280 220108 244332 220114
rect 244280 220050 244332 220056
rect 244464 220108 244516 220114
rect 244464 220050 244516 220056
rect 243636 218068 243688 218074
rect 243636 218010 243688 218016
rect 244096 218068 244148 218074
rect 244096 218010 244148 218016
rect 242728 217246 242802 217274
rect 241946 217110 242020 217138
rect 241946 216988 241974 217110
rect 242774 216988 242802 217246
rect 243648 217138 243676 218010
rect 244476 217274 244504 220050
rect 244924 219428 244976 219434
rect 244924 219370 244976 219376
rect 244936 218890 244964 219370
rect 244924 218884 244976 218890
rect 244924 218826 244976 218832
rect 245304 217274 245332 224742
rect 246316 218346 246344 228754
rect 246500 220794 246528 229706
rect 246776 228954 246804 231676
rect 246764 228948 246816 228954
rect 246764 228890 246816 228896
rect 246856 223304 246908 223310
rect 246856 223246 246908 223252
rect 246488 220788 246540 220794
rect 246488 220730 246540 220736
rect 246304 218340 246356 218346
rect 246304 218282 246356 218288
rect 246120 218204 246172 218210
rect 246120 218146 246172 218152
rect 243602 217110 243676 217138
rect 244430 217246 244504 217274
rect 245258 217246 245332 217274
rect 243602 216988 243630 217110
rect 244430 216988 244458 217246
rect 245258 216988 245286 217246
rect 246132 217138 246160 218146
rect 246868 217274 246896 223246
rect 247420 222766 247448 231676
rect 247604 231662 248078 231690
rect 247408 222760 247460 222766
rect 247408 222702 247460 222708
rect 247604 222154 247632 231662
rect 248236 228812 248288 228818
rect 248236 228754 248288 228760
rect 247592 222148 247644 222154
rect 247592 222090 247644 222096
rect 248248 218074 248276 228754
rect 248708 226710 248736 231676
rect 248696 226704 248748 226710
rect 248696 226646 248748 226652
rect 249352 225758 249380 231676
rect 249616 226772 249668 226778
rect 249616 226714 249668 226720
rect 249340 225752 249392 225758
rect 249340 225694 249392 225700
rect 249432 218884 249484 218890
rect 249432 218826 249484 218832
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248236 218068 248288 218074
rect 248236 218010 248288 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 246868 217246 246942 217274
rect 246086 217110 246160 217138
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217138 249472 218826
rect 249628 218074 249656 226714
rect 249996 222630 250024 231676
rect 250640 223990 250668 231676
rect 251284 229634 251312 231676
rect 251272 229628 251324 229634
rect 251272 229570 251324 229576
rect 251732 229628 251784 229634
rect 251732 229570 251784 229576
rect 251088 224664 251140 224670
rect 251088 224606 251140 224612
rect 250628 223984 250680 223990
rect 250628 223926 250680 223932
rect 250904 223576 250956 223582
rect 250904 223518 250956 223524
rect 249984 222624 250036 222630
rect 249984 222566 250036 222572
rect 250916 218074 250944 223518
rect 249616 218068 249668 218074
rect 249616 218010 249668 218016
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250904 218068 250956 218074
rect 250904 218010 250956 218016
rect 250272 217138 250300 218010
rect 251100 217274 251128 224606
rect 251744 218890 251772 229570
rect 251928 227594 251956 231676
rect 252572 229090 252600 231676
rect 252756 231662 253230 231690
rect 252560 229084 252612 229090
rect 252560 229026 252612 229032
rect 251916 227588 251968 227594
rect 251916 227530 251968 227536
rect 252468 225888 252520 225894
rect 252468 225830 252520 225836
rect 251732 218884 251784 218890
rect 251732 218826 251784 218832
rect 251732 218748 251784 218754
rect 251732 218690 251784 218696
rect 251744 218210 251772 218690
rect 251732 218204 251784 218210
rect 251732 218146 251784 218152
rect 252480 218074 252508 225830
rect 252756 221338 252784 231662
rect 253860 228954 253888 231676
rect 253848 228948 253900 228954
rect 253848 228890 253900 228896
rect 254504 225078 254532 231676
rect 254780 231662 255162 231690
rect 254492 225072 254544 225078
rect 254492 225014 254544 225020
rect 252744 221332 252796 221338
rect 252744 221274 252796 221280
rect 253848 220856 253900 220862
rect 253848 220798 253900 220804
rect 253572 220652 253624 220658
rect 253572 220594 253624 220600
rect 253204 219156 253256 219162
rect 253204 219098 253256 219104
rect 252744 218884 252796 218890
rect 252744 218826 252796 218832
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217110 249472 217138
rect 250226 217110 250300 217138
rect 251054 217246 251128 217274
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217110
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218826
rect 253216 218346 253244 219098
rect 253204 218340 253256 218346
rect 253204 218282 253256 218288
rect 253584 217274 253612 220594
rect 253860 219026 253888 220798
rect 254780 219978 254808 231662
rect 255228 228948 255280 228954
rect 255228 228890 255280 228896
rect 255044 225752 255096 225758
rect 255044 225694 255096 225700
rect 254768 219972 254820 219978
rect 254768 219914 254820 219920
rect 253848 219020 253900 219026
rect 253848 218962 253900 218968
rect 255056 218074 255084 225694
rect 254400 218068 254452 218074
rect 254400 218010 254452 218016
rect 255044 218068 255096 218074
rect 255044 218010 255096 218016
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254412 217138 254440 218010
rect 255240 217274 255268 228890
rect 255792 224126 255820 231676
rect 256436 230314 256464 231676
rect 256424 230308 256476 230314
rect 256424 230250 256476 230256
rect 256608 230308 256660 230314
rect 256608 230250 256660 230256
rect 255780 224120 255832 224126
rect 255780 224062 255832 224068
rect 256620 219434 256648 230250
rect 257080 228274 257108 231676
rect 257528 229084 257580 229090
rect 257528 229026 257580 229032
rect 257068 228268 257120 228274
rect 257068 228210 257120 228216
rect 256528 219406 256648 219434
rect 256528 218074 256556 219406
rect 257540 218074 257568 229026
rect 257724 225486 257752 231676
rect 257896 227452 257948 227458
rect 257896 227394 257948 227400
rect 257712 225480 257764 225486
rect 257712 225422 257764 225428
rect 257908 219434 257936 227394
rect 258368 222494 258396 231676
rect 258644 231662 259026 231690
rect 258356 222488 258408 222494
rect 258356 222430 258408 222436
rect 258080 222148 258132 222154
rect 258080 222090 258132 222096
rect 257724 219406 257936 219434
rect 256056 218068 256108 218074
rect 256056 218010 256108 218016
rect 256516 218068 256568 218074
rect 256516 218010 256568 218016
rect 256884 218068 256936 218074
rect 256884 218010 256936 218016
rect 257528 218068 257580 218074
rect 257528 218010 257580 218016
rect 254366 217110 254440 217138
rect 255194 217246 255268 217274
rect 254366 216988 254394 217110
rect 255194 216988 255222 217246
rect 256068 217138 256096 218010
rect 256896 217138 256924 218010
rect 257724 217274 257752 219406
rect 258092 218346 258120 222090
rect 258644 220862 258672 231662
rect 259276 227588 259328 227594
rect 259276 227530 259328 227536
rect 258632 220856 258684 220862
rect 258632 220798 258684 220804
rect 259092 219020 259144 219026
rect 259092 218962 259144 218968
rect 258080 218340 258132 218346
rect 258080 218282 258132 218288
rect 258540 218068 258592 218074
rect 258540 218010 258592 218016
rect 256022 217110 256096 217138
rect 256850 217110 256924 217138
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217110
rect 257678 216988 257706 217246
rect 258552 217138 258580 218010
rect 259104 217274 259132 218962
rect 259288 218074 259316 227530
rect 259656 226166 259684 231676
rect 259932 231662 260314 231690
rect 260852 231662 260958 231690
rect 259644 226160 259696 226166
rect 259644 226102 259696 226108
rect 259932 219842 259960 231662
rect 260852 221610 260880 231662
rect 261588 230450 261616 231676
rect 261576 230444 261628 230450
rect 261576 230386 261628 230392
rect 262232 227730 262260 231676
rect 262220 227724 262272 227730
rect 262220 227666 262272 227672
rect 262876 227186 262904 231676
rect 263060 231662 263534 231690
rect 263704 231662 264178 231690
rect 262864 227180 262916 227186
rect 262864 227122 262916 227128
rect 261852 226160 261904 226166
rect 261852 226102 261904 226108
rect 260840 221604 260892 221610
rect 260840 221546 260892 221552
rect 261024 221604 261076 221610
rect 261024 221546 261076 221552
rect 260196 220788 260248 220794
rect 260196 220730 260248 220736
rect 259920 219836 259972 219842
rect 259920 219778 259972 219784
rect 259276 218068 259328 218074
rect 259276 218010 259328 218016
rect 260208 217274 260236 220730
rect 261036 217274 261064 221546
rect 261864 217274 261892 226102
rect 263060 221066 263088 231662
rect 263508 227180 263560 227186
rect 263508 227122 263560 227128
rect 263324 221876 263376 221882
rect 263324 221818 263376 221824
rect 263048 221060 263100 221066
rect 263048 221002 263100 221008
rect 263336 219434 263364 221818
rect 263336 219406 263456 219434
rect 262680 218068 262732 218074
rect 262680 218010 262732 218016
rect 259104 217246 259362 217274
rect 258506 217110 258580 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217246
rect 260162 217246 260236 217274
rect 260990 217246 261064 217274
rect 261818 217246 261892 217274
rect 260162 216988 260190 217246
rect 260990 216988 261018 217246
rect 261818 216988 261846 217246
rect 262692 217138 262720 218010
rect 263428 217274 263456 219406
rect 263520 218090 263548 227122
rect 263704 222154 263732 231662
rect 264808 228546 264836 231676
rect 265176 231662 265466 231690
rect 264796 228540 264848 228546
rect 264796 228482 264848 228488
rect 264152 226568 264204 226574
rect 264152 226510 264204 226516
rect 263692 222148 263744 222154
rect 263692 222090 263744 222096
rect 264164 219298 264192 226510
rect 264796 222760 264848 222766
rect 264796 222702 264848 222708
rect 264152 219292 264204 219298
rect 264152 219234 264204 219240
rect 263520 218074 263640 218090
rect 264808 218074 264836 222702
rect 265176 220522 265204 231662
rect 266096 225622 266124 231676
rect 266084 225616 266136 225622
rect 266084 225558 266136 225564
rect 266176 224120 266228 224126
rect 266176 224062 266228 224068
rect 265164 220516 265216 220522
rect 265164 220458 265216 220464
rect 265992 219156 266044 219162
rect 265992 219098 266044 219104
rect 263520 218068 263652 218074
rect 263520 218062 263600 218068
rect 263600 218010 263652 218016
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 263428 217246 263502 217274
rect 262646 217110 262720 217138
rect 262646 216988 262674 217110
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217138 266032 219098
rect 266188 218074 266216 224062
rect 266740 223718 266768 231676
rect 267384 226914 267412 231676
rect 267936 231662 268042 231690
rect 268304 231662 268686 231690
rect 267372 226908 267424 226914
rect 267372 226850 267424 226856
rect 267004 226296 267056 226302
rect 267004 226238 267056 226244
rect 266728 223712 266780 223718
rect 266728 223654 266780 223660
rect 266820 221332 266872 221338
rect 266820 221274 266872 221280
rect 266176 218068 266228 218074
rect 266176 218010 266228 218016
rect 266832 217274 266860 221274
rect 267016 218618 267044 226238
rect 267648 220516 267700 220522
rect 267648 220458 267700 220464
rect 267004 218612 267056 218618
rect 267004 218554 267056 218560
rect 267660 217274 267688 220458
rect 267936 220386 267964 231662
rect 268304 221202 268332 231662
rect 268936 228268 268988 228274
rect 268936 228210 268988 228216
rect 268292 221196 268344 221202
rect 268292 221138 268344 221144
rect 267924 220380 267976 220386
rect 267924 220322 267976 220328
rect 268948 218074 268976 228210
rect 269316 226574 269344 231676
rect 269304 226568 269356 226574
rect 269304 226510 269356 226516
rect 269960 226030 269988 231676
rect 269948 226024 270000 226030
rect 269948 225966 270000 225972
rect 270040 225616 270092 225622
rect 270040 225558 270092 225564
rect 270052 218074 270080 225558
rect 270604 223854 270632 231676
rect 271248 227050 271276 231676
rect 271892 229906 271920 231676
rect 271880 229900 271932 229906
rect 271880 229842 271932 229848
rect 272536 228682 272564 231676
rect 272720 231662 273194 231690
rect 272524 228676 272576 228682
rect 272524 228618 272576 228624
rect 272524 228540 272576 228546
rect 272524 228482 272576 228488
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 271144 226432 271196 226438
rect 271144 226374 271196 226380
rect 270592 223848 270644 223854
rect 270592 223790 270644 223796
rect 270224 222148 270276 222154
rect 270224 222090 270276 222096
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 268936 218068 268988 218074
rect 268936 218010 268988 218016
rect 269304 218068 269356 218074
rect 269304 218010 269356 218016
rect 270040 218068 270092 218074
rect 270040 218010 270092 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217110 266032 217138
rect 266786 217246 266860 217274
rect 267614 217246 267688 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217110
rect 266786 216988 266814 217246
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218010
rect 270236 217274 270264 222090
rect 271156 218482 271184 226374
rect 271144 218476 271196 218482
rect 271144 218418 271196 218424
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 270098 217246 270264 217274
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272340 219428 272392 219434
rect 272340 219370 272392 219376
rect 272352 218618 272380 219370
rect 272340 218612 272392 218618
rect 272340 218554 272392 218560
rect 272536 218074 272564 228482
rect 272720 219706 272748 231662
rect 273824 228410 273852 231676
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274468 226302 274496 231676
rect 275112 229094 275140 231676
rect 274928 229066 275140 229094
rect 275480 231662 275770 231690
rect 276124 231662 276414 231690
rect 274456 226296 274508 226302
rect 274456 226238 274508 226244
rect 274272 224936 274324 224942
rect 274272 224878 274324 224884
rect 273444 220380 273496 220386
rect 273444 220322 273496 220328
rect 272708 219700 272760 219706
rect 272708 219642 272760 219648
rect 272708 219428 272760 219434
rect 272708 219370 272760 219376
rect 272524 218068 272576 218074
rect 272524 218010 272576 218016
rect 272720 217274 272748 219370
rect 273456 217274 273484 220322
rect 274284 217274 274312 224878
rect 274928 224534 274956 229066
rect 274916 224528 274968 224534
rect 274916 224470 274968 224476
rect 275100 224528 275152 224534
rect 275100 224470 275152 224476
rect 275112 217274 275140 224470
rect 275480 223038 275508 231662
rect 275652 229900 275704 229906
rect 275652 229842 275704 229848
rect 275664 229094 275692 229842
rect 275664 229066 275876 229094
rect 275468 223032 275520 223038
rect 275468 222974 275520 222980
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 272582 217246 272748 217274
rect 273410 217246 273484 217274
rect 274238 217246 274312 217274
rect 275066 217246 275140 217274
rect 275848 217274 275876 229066
rect 276124 221474 276152 231662
rect 277044 230042 277072 231676
rect 277032 230036 277084 230042
rect 277032 229978 277084 229984
rect 277216 230036 277268 230042
rect 277216 229978 277268 229984
rect 277032 227724 277084 227730
rect 277032 227666 277084 227672
rect 276112 221468 276164 221474
rect 276112 221410 276164 221416
rect 277044 219434 277072 227666
rect 277228 227186 277256 229978
rect 277216 227180 277268 227186
rect 277216 227122 277268 227128
rect 277688 224398 277716 231676
rect 277964 231662 278346 231690
rect 277676 224392 277728 224398
rect 277676 224334 277728 224340
rect 277964 222018 277992 231662
rect 278412 226024 278464 226030
rect 278412 225966 278464 225972
rect 277952 222012 278004 222018
rect 277952 221954 278004 221960
rect 277044 219406 277256 219434
rect 277228 218074 277256 219406
rect 276756 218068 276808 218074
rect 276756 218010 276808 218016
rect 277216 218068 277268 218074
rect 277216 218010 277268 218016
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272582 216988 272610 217246
rect 273410 216988 273438 217246
rect 274238 216988 274266 217246
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276768 217138 276796 218010
rect 277596 217138 277624 218010
rect 278424 217274 278452 225966
rect 278976 224262 279004 231676
rect 279620 226438 279648 231676
rect 280264 227322 280292 231676
rect 280448 231662 280922 231690
rect 280252 227316 280304 227322
rect 280252 227258 280304 227264
rect 279608 226432 279660 226438
rect 279608 226374 279660 226380
rect 278964 224256 279016 224262
rect 278964 224198 279016 224204
rect 279424 223916 279476 223922
rect 279424 223858 279476 223864
rect 278596 223032 278648 223038
rect 278596 222974 278648 222980
rect 278608 218074 278636 222974
rect 279436 218618 279464 223858
rect 280068 222012 280120 222018
rect 280068 221954 280120 221960
rect 279424 218612 279476 218618
rect 279424 218554 279476 218560
rect 279240 218476 279292 218482
rect 279240 218418 279292 218424
rect 278596 218068 278648 218074
rect 278596 218010 278648 218016
rect 276722 217110 276796 217138
rect 277550 217110 277624 217138
rect 278378 217246 278452 217274
rect 276722 216988 276750 217110
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218418
rect 280080 217274 280108 221954
rect 280448 220250 280476 231662
rect 281356 227180 281408 227186
rect 281356 227122 281408 227128
rect 280436 220244 280488 220250
rect 280436 220186 280488 220192
rect 281368 219434 281396 227122
rect 281552 222902 281580 231676
rect 282196 230178 282224 231676
rect 282184 230172 282236 230178
rect 282184 230114 282236 230120
rect 282644 230172 282696 230178
rect 282644 230114 282696 230120
rect 282656 225622 282684 230114
rect 282840 228002 282868 231676
rect 282828 227996 282880 228002
rect 282828 227938 282880 227944
rect 282644 225616 282696 225622
rect 282644 225558 282696 225564
rect 283484 223174 283512 231676
rect 283668 231662 284142 231690
rect 283472 223168 283524 223174
rect 283472 223110 283524 223116
rect 281540 222896 281592 222902
rect 281540 222838 281592 222844
rect 282460 222896 282512 222902
rect 282460 222838 282512 222844
rect 281368 219406 281488 219434
rect 281460 218074 281488 219406
rect 282472 218074 282500 222838
rect 283668 221746 283696 231662
rect 284116 225616 284168 225622
rect 284116 225558 284168 225564
rect 283656 221740 283708 221746
rect 283656 221682 283708 221688
rect 282644 220924 282696 220930
rect 282644 220866 282696 220872
rect 280896 218068 280948 218074
rect 280896 218010 280948 218016
rect 281448 218068 281500 218074
rect 281448 218010 281500 218016
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 282460 218068 282512 218074
rect 282460 218010 282512 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280908 217138 280936 218010
rect 281736 217138 281764 218010
rect 282656 217274 282684 220866
rect 283380 220244 283432 220250
rect 283380 220186 283432 220192
rect 283392 217274 283420 220186
rect 280862 217110 280936 217138
rect 281690 217110 281764 217138
rect 282518 217246 282684 217274
rect 283346 217246 283420 217274
rect 284128 217274 284156 225558
rect 284772 223922 284800 231676
rect 285048 231662 285430 231690
rect 285048 225214 285076 231662
rect 285496 228404 285548 228410
rect 285496 228346 285548 228352
rect 285036 225208 285088 225214
rect 285036 225150 285088 225156
rect 284760 223916 284812 223922
rect 284760 223858 284812 223864
rect 285508 218074 285536 228346
rect 286060 223446 286088 231676
rect 286324 226296 286376 226302
rect 286324 226238 286376 226244
rect 286048 223440 286100 223446
rect 286048 223382 286100 223388
rect 285864 219428 285916 219434
rect 285864 219370 285916 219376
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 280862 216988 280890 217110
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283346 216988 283374 217246
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 219370
rect 286336 218754 286364 226238
rect 286704 225350 286732 231676
rect 287348 229770 287376 231676
rect 287336 229764 287388 229770
rect 287336 229706 287388 229712
rect 287704 229764 287756 229770
rect 287704 229706 287756 229712
rect 286692 225344 286744 225350
rect 286692 225286 286744 225292
rect 286692 224392 286744 224398
rect 286692 224334 286744 224340
rect 286324 218748 286376 218754
rect 286324 218690 286376 218696
rect 286704 217274 286732 224334
rect 287716 220930 287744 229706
rect 287992 224806 288020 231676
rect 287980 224800 288032 224806
rect 287980 224742 288032 224748
rect 288636 223310 288664 231676
rect 288820 231662 289294 231690
rect 288624 223304 288676 223310
rect 288624 223246 288676 223252
rect 288256 223168 288308 223174
rect 288256 223110 288308 223116
rect 287888 222352 287940 222358
rect 287888 222294 287940 222300
rect 287704 220924 287756 220930
rect 287704 220866 287756 220872
rect 287900 218890 287928 222294
rect 287888 218884 287940 218890
rect 287888 218826 287940 218832
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288268 217274 288296 223110
rect 288820 222194 288848 231662
rect 289924 226302 289952 231676
rect 290568 226778 290596 231676
rect 290556 226772 290608 226778
rect 290556 226714 290608 226720
rect 289912 226296 289964 226302
rect 289912 226238 289964 226244
rect 291016 226296 291068 226302
rect 291016 226238 291068 226244
rect 290832 224256 290884 224262
rect 290832 224198 290884 224204
rect 289728 223304 289780 223310
rect 289728 223246 289780 223252
rect 288544 222166 288848 222194
rect 288544 220114 288572 222166
rect 288532 220108 288584 220114
rect 288532 220050 288584 220056
rect 288716 220108 288768 220114
rect 288716 220050 288768 220056
rect 288728 218074 288756 220050
rect 289740 218074 289768 223246
rect 288716 218068 288768 218074
rect 288716 218010 288768 218016
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289728 218068 289780 218074
rect 289728 218010 289780 218016
rect 290004 218068 290056 218074
rect 290004 218010 290056 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217138 290044 218010
rect 290844 217274 290872 224198
rect 291028 219434 291056 226238
rect 291212 223582 291240 231676
rect 291856 228818 291884 231676
rect 292500 229634 292528 231676
rect 292488 229628 292540 229634
rect 292488 229570 292540 229576
rect 291844 228812 291896 228818
rect 291844 228754 291896 228760
rect 291660 228676 291712 228682
rect 291660 228618 291712 228624
rect 291200 223576 291252 223582
rect 291200 223518 291252 223524
rect 291028 219406 291148 219434
rect 291120 218074 291148 219406
rect 291672 219026 291700 228618
rect 293144 225894 293172 231676
rect 293328 231662 293802 231690
rect 293132 225888 293184 225894
rect 293132 225830 293184 225836
rect 292488 221468 292540 221474
rect 292488 221410 292540 221416
rect 291660 219020 291712 219026
rect 291660 218962 291712 218968
rect 291660 218884 291712 218890
rect 291660 218826 291712 218832
rect 291108 218068 291160 218074
rect 291108 218010 291160 218016
rect 289142 217110 289216 217138
rect 289970 217110 290044 217138
rect 290798 217246 290872 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217110
rect 290798 216988 290826 217246
rect 291672 217138 291700 218826
rect 292500 217274 292528 221410
rect 293328 220658 293356 231662
rect 293776 226908 293828 226914
rect 293776 226850 293828 226856
rect 293316 220652 293368 220658
rect 293316 220594 293368 220600
rect 293788 218074 293816 226850
rect 294432 224670 294460 231676
rect 294420 224664 294472 224670
rect 294420 224606 294472 224612
rect 295076 222358 295104 231676
rect 295720 228954 295748 231676
rect 296364 229090 296392 231676
rect 296352 229084 296404 229090
rect 296352 229026 296404 229032
rect 295708 228948 295760 228954
rect 295708 228890 295760 228896
rect 296628 228676 296680 228682
rect 296628 228618 296680 228624
rect 296444 225888 296496 225894
rect 296444 225830 296496 225836
rect 295064 222352 295116 222358
rect 295064 222294 295116 222300
rect 294972 219972 295024 219978
rect 294972 219914 295024 219920
rect 294144 218476 294196 218482
rect 294144 218418 294196 218424
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 291626 217110 291700 217138
rect 292454 217246 292528 217274
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 218418
rect 294984 217274 295012 219914
rect 296456 219434 296484 225830
rect 296456 219406 296576 219434
rect 295800 219156 295852 219162
rect 295800 219098 295852 219104
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 219098
rect 296548 217274 296576 219406
rect 296640 219178 296668 228618
rect 297008 225758 297036 231676
rect 297652 230314 297680 231676
rect 297640 230308 297692 230314
rect 297640 230250 297692 230256
rect 297824 230308 297876 230314
rect 297824 230250 297876 230256
rect 297836 229094 297864 230250
rect 297744 229066 297864 229094
rect 296996 225752 297048 225758
rect 296996 225694 297048 225700
rect 297272 225072 297324 225078
rect 297272 225014 297324 225020
rect 296640 219162 296760 219178
rect 296640 219156 296772 219162
rect 296640 219150 296720 219156
rect 296720 219098 296772 219104
rect 297284 219026 297312 225014
rect 297744 223310 297772 229066
rect 298296 227594 298324 231676
rect 298572 231662 298954 231690
rect 298284 227588 298336 227594
rect 298284 227530 298336 227536
rect 297916 223576 297968 223582
rect 297916 223518 297968 223524
rect 297732 223304 297784 223310
rect 297732 223246 297784 223252
rect 297272 219020 297324 219026
rect 297272 218962 297324 218968
rect 297928 218074 297956 223518
rect 298572 220794 298600 231662
rect 299584 227458 299612 231676
rect 300228 228818 300256 231676
rect 300216 228812 300268 228818
rect 300216 228754 300268 228760
rect 300676 228812 300728 228818
rect 300676 228754 300728 228760
rect 299572 227452 299624 227458
rect 299572 227394 299624 227400
rect 299296 224664 299348 224670
rect 299296 224606 299348 224612
rect 299112 223304 299164 223310
rect 299112 223246 299164 223252
rect 298560 220788 298612 220794
rect 298560 220730 298612 220736
rect 299124 218074 299152 223246
rect 297456 218068 297508 218074
rect 297456 218010 297508 218016
rect 297916 218068 297968 218074
rect 297916 218010 297968 218016
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 299112 218068 299164 218074
rect 299112 218010 299164 218016
rect 296548 217246 296622 217274
rect 295766 217110 295840 217138
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218010
rect 298296 217138 298324 218010
rect 299308 217274 299336 224606
rect 300492 218884 300544 218890
rect 300492 218826 300544 218832
rect 299940 218068 299992 218074
rect 299940 218010 299992 218016
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217246 299336 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217246
rect 299952 217138 299980 218010
rect 300504 217274 300532 218826
rect 300688 218074 300716 228754
rect 300872 226166 300900 231676
rect 301240 231662 301530 231690
rect 301792 231662 302174 231690
rect 300860 226160 300912 226166
rect 300860 226102 300912 226108
rect 301240 221882 301268 231662
rect 301504 227588 301556 227594
rect 301504 227530 301556 227536
rect 301516 227050 301544 227530
rect 301504 227044 301556 227050
rect 301504 226986 301556 226992
rect 301228 221876 301280 221882
rect 301228 221818 301280 221824
rect 301792 221610 301820 231662
rect 302804 230042 302832 231676
rect 302792 230036 302844 230042
rect 302792 229978 302844 229984
rect 303252 230036 303304 230042
rect 303252 229978 303304 229984
rect 302148 228948 302200 228954
rect 302148 228890 302200 228896
rect 301964 221876 302016 221882
rect 301964 221818 302016 221824
rect 301780 221604 301832 221610
rect 301780 221546 301832 221552
rect 301976 219298 302004 221818
rect 301964 219292 302016 219298
rect 301964 219234 302016 219240
rect 302160 218074 302188 228890
rect 303264 223582 303292 229978
rect 303448 224126 303476 231676
rect 303816 231662 304106 231690
rect 304368 231662 304750 231690
rect 303436 224120 303488 224126
rect 303436 224062 303488 224068
rect 303252 223576 303304 223582
rect 303252 223518 303304 223524
rect 303252 221740 303304 221746
rect 303252 221682 303304 221688
rect 302424 220652 302476 220658
rect 302424 220594 302476 220600
rect 300676 218068 300728 218074
rect 300676 218010 300728 218016
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 300504 217246 300762 217274
rect 299906 217110 299980 217138
rect 299906 216988 299934 217110
rect 300734 216988 300762 217246
rect 301608 217138 301636 218010
rect 302436 217274 302464 220594
rect 303264 217274 303292 221682
rect 303816 221338 303844 231662
rect 304368 222766 304396 231662
rect 304908 227452 304960 227458
rect 304908 227394 304960 227400
rect 304724 223440 304776 223446
rect 304724 223382 304776 223388
rect 304356 222760 304408 222766
rect 304356 222702 304408 222708
rect 303804 221332 303856 221338
rect 303804 221274 303856 221280
rect 304736 218074 304764 223382
rect 304080 218068 304132 218074
rect 304080 218010 304132 218016
rect 304724 218068 304776 218074
rect 304724 218010 304776 218016
rect 301562 217110 301636 217138
rect 302390 217246 302464 217274
rect 303218 217246 303292 217274
rect 301562 216988 301590 217110
rect 302390 216988 302418 217246
rect 303218 216988 303246 217246
rect 304092 217138 304120 218010
rect 304920 217274 304948 227394
rect 305380 225078 305408 231676
rect 305552 229084 305604 229090
rect 305552 229026 305604 229032
rect 305368 225072 305420 225078
rect 305368 225014 305420 225020
rect 305564 218618 305592 229026
rect 306024 228274 306052 231676
rect 306392 231662 306682 231690
rect 306852 231662 307326 231690
rect 306012 228268 306064 228274
rect 306012 228210 306064 228216
rect 306196 227316 306248 227322
rect 306196 227258 306248 227264
rect 305552 218612 305604 218618
rect 305552 218554 305604 218560
rect 306208 218074 306236 227258
rect 306392 222154 306420 231662
rect 306380 222148 306432 222154
rect 306380 222090 306432 222096
rect 306852 220522 306880 231662
rect 307956 230178 307984 231676
rect 307944 230172 307996 230178
rect 307944 230114 307996 230120
rect 308128 230172 308180 230178
rect 308128 230114 308180 230120
rect 307668 223576 307720 223582
rect 307668 223518 307720 223524
rect 306840 220516 306892 220522
rect 306840 220458 306892 220464
rect 307392 219020 307444 219026
rect 307392 218962 307444 218968
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306196 218068 306248 218074
rect 306196 218010 306248 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217274 307432 218962
rect 307680 218074 307708 223518
rect 308140 223446 308168 230114
rect 308600 227594 308628 231676
rect 308588 227588 308640 227594
rect 308588 227530 308640 227536
rect 309048 226160 309100 226166
rect 309048 226102 309100 226108
rect 308128 223440 308180 223446
rect 308128 223382 308180 223388
rect 308864 221604 308916 221610
rect 308864 221546 308916 221552
rect 308876 219434 308904 221546
rect 309060 219434 309088 226102
rect 309244 220386 309272 231676
rect 309888 228546 309916 231676
rect 310546 231662 310744 231690
rect 310716 229094 310744 231662
rect 310716 229066 310928 229094
rect 309876 228540 309928 228546
rect 309876 228482 309928 228488
rect 310428 227044 310480 227050
rect 310428 226986 310480 226992
rect 309232 220380 309284 220386
rect 309232 220322 309284 220328
rect 308220 219428 308272 219434
rect 308876 219406 308996 219434
rect 309060 219428 309192 219434
rect 309060 219406 309140 219428
rect 308220 219370 308272 219376
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217246 307432 217274
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217246
rect 308232 217138 308260 219370
rect 308968 217274 308996 219406
rect 309140 219370 309192 219376
rect 310440 218074 310468 226986
rect 310704 222148 310756 222154
rect 310704 222090 310756 222096
rect 309876 218068 309928 218074
rect 309876 218010 309928 218016
rect 310428 218068 310480 218074
rect 310428 218010 310480 218016
rect 308968 217246 309042 217274
rect 308186 217110 308260 217138
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309888 217138 309916 218010
rect 310716 217274 310744 222090
rect 310900 221882 310928 229066
rect 311176 224534 311204 231676
rect 311820 227730 311848 231676
rect 311992 230444 312044 230450
rect 311992 230386 312044 230392
rect 312004 229906 312032 230386
rect 311992 229900 312044 229906
rect 311992 229842 312044 229848
rect 311808 227724 311860 227730
rect 311808 227666 311860 227672
rect 312464 224942 312492 231676
rect 313108 230450 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230444 313148 230450
rect 313096 230386 313148 230392
rect 312636 229900 312688 229906
rect 312636 229842 312688 229848
rect 312452 224936 312504 224942
rect 312452 224878 312504 224884
rect 311164 224528 311216 224534
rect 311164 224470 311216 224476
rect 311532 224528 311584 224534
rect 311532 224470 311584 224476
rect 310888 221876 310940 221882
rect 310888 221818 310940 221824
rect 311544 217274 311572 224470
rect 312648 222154 312676 229842
rect 313292 226030 313320 231662
rect 313936 229094 313964 231662
rect 313752 229066 313964 229094
rect 313280 226024 313332 226030
rect 313280 225966 313332 225972
rect 312912 223440 312964 223446
rect 312912 223382 312964 223388
rect 312636 222148 312688 222154
rect 312636 222090 312688 222096
rect 312924 218074 312952 223382
rect 313752 222018 313780 229066
rect 313924 228540 313976 228546
rect 313924 228482 313976 228488
rect 313740 222012 313792 222018
rect 313740 221954 313792 221960
rect 313188 221876 313240 221882
rect 313188 221818 313240 221824
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 312912 218068 312964 218074
rect 312912 218010 312964 218016
rect 309842 217110 309916 217138
rect 310670 217246 310744 217274
rect 311498 217246 311572 217274
rect 309842 216988 309870 217110
rect 310670 216988 310698 217246
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313200 217274 313228 221818
rect 313936 219298 313964 228482
rect 315040 223038 315068 231676
rect 315684 229090 315712 231676
rect 315672 229084 315724 229090
rect 315672 229026 315724 229032
rect 315672 225752 315724 225758
rect 315672 225694 315724 225700
rect 315028 223032 315080 223038
rect 315028 222974 315080 222980
rect 314844 220380 314896 220386
rect 314844 220322 314896 220328
rect 313924 219292 313976 219298
rect 313924 219234 313976 219240
rect 314016 219156 314068 219162
rect 314016 219098 314068 219104
rect 312326 217110 312400 217138
rect 313154 217246 313228 217274
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 219098
rect 314856 217274 314884 220322
rect 315684 217274 315712 225694
rect 316328 222902 316356 231676
rect 316512 231662 316986 231690
rect 316316 222896 316368 222902
rect 316316 222838 316368 222844
rect 316512 221218 316540 231662
rect 317616 227186 317644 231676
rect 318260 229770 318288 231676
rect 318248 229764 318300 229770
rect 318248 229706 318300 229712
rect 318064 229628 318116 229634
rect 318064 229570 318116 229576
rect 317604 227180 317656 227186
rect 317604 227122 317656 227128
rect 316684 223032 316736 223038
rect 316684 222974 316736 222980
rect 316328 221190 316540 221218
rect 316328 220250 316356 221190
rect 316316 220244 316368 220250
rect 316316 220186 316368 220192
rect 316500 220244 316552 220250
rect 316500 220186 316552 220192
rect 316512 217274 316540 220186
rect 316696 218482 316724 222974
rect 318076 219434 318104 229570
rect 318904 228410 318932 231676
rect 318892 228404 318944 228410
rect 318892 228346 318944 228352
rect 319548 224398 319576 231676
rect 320192 225622 320220 231676
rect 320836 228546 320864 231676
rect 321112 231662 321494 231690
rect 320824 228540 320876 228546
rect 320824 228482 320876 228488
rect 320180 225616 320232 225622
rect 320180 225558 320232 225564
rect 319996 224800 320048 224806
rect 319996 224742 320048 224748
rect 319536 224392 319588 224398
rect 319536 224334 319588 224340
rect 319812 224392 319864 224398
rect 319812 224334 319864 224340
rect 318248 222012 318300 222018
rect 318248 221954 318300 221960
rect 318260 219434 318288 221954
rect 317984 219406 318104 219434
rect 318168 219406 318288 219434
rect 316684 218476 316736 218482
rect 316684 218418 316736 218424
rect 317984 218074 318012 219406
rect 317328 218068 317380 218074
rect 317328 218010 317380 218016
rect 317972 218068 318024 218074
rect 317972 218010 318024 218016
rect 313982 217110 314056 217138
rect 314810 217246 314884 217274
rect 315638 217246 315712 217274
rect 316466 217246 316540 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217246
rect 315638 216988 315666 217246
rect 316466 216988 316494 217246
rect 317340 217138 317368 218010
rect 318168 217274 318196 219406
rect 319824 218074 319852 224334
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 319812 218068 319864 218074
rect 319812 218010 319864 218016
rect 317294 217110 317368 217138
rect 318122 217246 318196 217274
rect 317294 216988 317322 217110
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 320008 217274 320036 224742
rect 321112 223174 321140 231662
rect 322124 226302 322152 231676
rect 322400 231662 322782 231690
rect 322112 226296 322164 226302
rect 322112 226238 322164 226244
rect 321376 225616 321428 225622
rect 321376 225558 321428 225564
rect 321100 223168 321152 223174
rect 321100 223110 321152 223116
rect 320640 219292 320692 219298
rect 320640 219234 320692 219240
rect 318950 217110 319024 217138
rect 319778 217246 320036 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 219234
rect 321388 217274 321416 225558
rect 321560 220788 321612 220794
rect 321560 220730 321612 220736
rect 321572 218754 321600 220730
rect 322400 220114 322428 231662
rect 323412 230314 323440 231676
rect 323688 231662 324070 231690
rect 324516 231662 324714 231690
rect 324976 231662 325358 231690
rect 325896 231662 326002 231690
rect 326264 231662 326646 231690
rect 323400 230308 323452 230314
rect 323400 230250 323452 230256
rect 322848 227180 322900 227186
rect 322848 227122 322900 227128
rect 322388 220108 322440 220114
rect 322388 220050 322440 220056
rect 321560 218748 321612 218754
rect 321560 218690 321612 218696
rect 322860 218074 322888 227122
rect 323688 224262 323716 231662
rect 323676 224256 323728 224262
rect 323676 224198 323728 224204
rect 323952 224256 324004 224262
rect 323952 224198 324004 224204
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 323124 218068 323176 218074
rect 323124 218010 323176 218016
rect 321388 217246 321462 217274
rect 320606 217110 320680 217138
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217138 323164 218010
rect 323964 217274 323992 224198
rect 324136 222896 324188 222902
rect 324136 222838 324188 222844
rect 324148 218074 324176 222838
rect 324516 220794 324544 231662
rect 324976 226914 325004 231662
rect 325424 228540 325476 228546
rect 325424 228482 325476 228488
rect 324964 226908 325016 226914
rect 324964 226850 325016 226856
rect 324504 220788 324556 220794
rect 324504 220730 324556 220736
rect 325436 218074 325464 228482
rect 325608 220108 325660 220114
rect 325608 220050 325660 220056
rect 324136 218068 324188 218074
rect 324136 218010 324188 218016
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 325424 218068 325476 218074
rect 325424 218010 325476 218016
rect 322262 217110 322336 217138
rect 323090 217110 323164 217138
rect 323918 217246 323992 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217110
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325620 217274 325648 220050
rect 325896 219978 325924 231662
rect 326264 221474 326292 231662
rect 326896 229084 326948 229090
rect 326896 229026 326948 229032
rect 326252 221468 326304 221474
rect 326252 221410 326304 221416
rect 325884 219972 325936 219978
rect 325884 219914 325936 219920
rect 326908 218074 326936 229026
rect 327276 223038 327304 231676
rect 327552 231662 327934 231690
rect 327552 225894 327580 231662
rect 327540 225888 327592 225894
rect 327540 225830 327592 225836
rect 327724 225004 327776 225010
rect 327724 224946 327776 224952
rect 327264 223032 327316 223038
rect 327264 222974 327316 222980
rect 327736 218890 327764 224946
rect 328564 223310 328592 231676
rect 329208 228682 329236 231676
rect 329852 230042 329880 231676
rect 329840 230036 329892 230042
rect 329840 229978 329892 229984
rect 330496 228818 330524 231676
rect 330944 230036 330996 230042
rect 330944 229978 330996 229984
rect 330956 229094 330984 229978
rect 330956 229066 331076 229094
rect 330484 228812 330536 228818
rect 330484 228754 330536 228760
rect 329196 228676 329248 228682
rect 329196 228618 329248 228624
rect 330484 228404 330536 228410
rect 330484 228346 330536 228352
rect 329748 226024 329800 226030
rect 329748 225966 329800 225972
rect 328552 223304 328604 223310
rect 328552 223246 328604 223252
rect 328092 223032 328144 223038
rect 328092 222974 328144 222980
rect 327724 218884 327776 218890
rect 327724 218826 327776 218832
rect 327264 218748 327316 218754
rect 327264 218690 327316 218696
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 324746 217110 324820 217138
rect 325574 217246 325648 217274
rect 324746 216988 324774 217110
rect 325574 216988 325602 217246
rect 326448 217138 326476 218010
rect 327276 217138 327304 218690
rect 328104 217274 328132 222974
rect 328920 218204 328972 218210
rect 328920 218146 328972 218152
rect 326402 217110 326476 217138
rect 327230 217110 327304 217138
rect 328058 217246 328132 217274
rect 326402 216988 326430 217110
rect 327230 216988 327258 217110
rect 328058 216988 328086 217246
rect 328932 217138 328960 218146
rect 329760 217274 329788 225966
rect 330496 218210 330524 228346
rect 330484 218204 330536 218210
rect 330484 218146 330536 218152
rect 331048 218074 331076 229066
rect 331140 228970 331168 231676
rect 331140 228954 331260 228970
rect 331140 228948 331272 228954
rect 331140 228942 331220 228948
rect 331220 228890 331272 228896
rect 331784 224670 331812 231676
rect 332060 231662 332442 231690
rect 332796 231662 333086 231690
rect 332060 225010 332088 231662
rect 332232 225888 332284 225894
rect 332232 225830 332284 225836
rect 332048 225004 332100 225010
rect 332048 224946 332100 224952
rect 331772 224664 331824 224670
rect 331772 224606 331824 224612
rect 331404 222148 331456 222154
rect 331404 222090 331456 222096
rect 330576 218068 330628 218074
rect 330576 218010 330628 218016
rect 331036 218068 331088 218074
rect 331036 218010 331088 218016
rect 328886 217110 328960 217138
rect 329714 217246 329788 217274
rect 328886 216988 328914 217110
rect 329714 216988 329742 217246
rect 330588 217138 330616 218010
rect 331416 217274 331444 222090
rect 332244 217274 332272 225830
rect 332796 221746 332824 231662
rect 333716 227458 333744 231676
rect 334084 231662 334374 231690
rect 333704 227452 333756 227458
rect 333704 227394 333756 227400
rect 333888 227452 333940 227458
rect 333888 227394 333940 227400
rect 332784 221740 332836 221746
rect 332784 221682 332836 221688
rect 332692 219564 332744 219570
rect 332692 219506 332744 219512
rect 332704 219026 332732 219506
rect 333704 219428 333756 219434
rect 333704 219370 333756 219376
rect 332692 219020 332744 219026
rect 332692 218962 332744 218968
rect 333060 218068 333112 218074
rect 333060 218010 333112 218016
rect 330542 217110 330616 217138
rect 331370 217246 331444 217274
rect 332198 217246 332272 217274
rect 330542 216988 330570 217110
rect 331370 216988 331398 217246
rect 332198 216988 332226 217246
rect 333072 217138 333100 218010
rect 333716 217274 333744 219370
rect 333900 218074 333928 227394
rect 334084 220658 334112 231662
rect 335004 230178 335032 231676
rect 334992 230172 335044 230178
rect 334992 230114 335044 230120
rect 335176 230172 335228 230178
rect 335176 230114 335228 230120
rect 335188 229094 335216 230114
rect 335004 229066 335216 229094
rect 335004 224262 335032 229066
rect 335176 224664 335228 224670
rect 335176 224606 335228 224612
rect 334992 224256 335044 224262
rect 334992 224198 335044 224204
rect 334072 220652 334124 220658
rect 334072 220594 334124 220600
rect 335188 218074 335216 224606
rect 335648 223582 335676 231676
rect 336292 226166 336320 231676
rect 336464 228676 336516 228682
rect 336464 228618 336516 228624
rect 336280 226160 336332 226166
rect 336280 226102 336332 226108
rect 335636 223576 335688 223582
rect 335636 223518 335688 223524
rect 336004 223372 336056 223378
rect 336004 223314 336056 223320
rect 336016 219162 336044 223314
rect 336476 219434 336504 228618
rect 336936 227322 336964 231676
rect 337212 231662 337594 231690
rect 336924 227316 336976 227322
rect 336924 227258 336976 227264
rect 337212 219570 337240 231662
rect 338224 227050 338252 231676
rect 338212 227044 338264 227050
rect 338212 226986 338264 226992
rect 338672 227044 338724 227050
rect 338672 226986 338724 226992
rect 338028 220516 338080 220522
rect 338028 220458 338080 220464
rect 337200 219564 337252 219570
rect 337200 219506 337252 219512
rect 336384 219406 336504 219434
rect 336004 219156 336056 219162
rect 336004 219098 336056 219104
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335176 218068 335228 218074
rect 335176 218010 335228 218016
rect 335544 218068 335596 218074
rect 335544 218010 335596 218016
rect 333716 217246 333882 217274
rect 333026 217110 333100 217138
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218010
rect 336384 217274 336412 219406
rect 337200 219020 337252 219026
rect 337200 218962 337252 218968
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336412 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218962
rect 338040 217274 338068 220458
rect 338684 218074 338712 226986
rect 338868 224534 338896 231676
rect 339526 231662 339724 231690
rect 338856 224528 338908 224534
rect 338856 224470 338908 224476
rect 339408 224256 339460 224262
rect 339408 224198 339460 224204
rect 339420 218074 339448 224198
rect 339696 221610 339724 231662
rect 340156 229906 340184 231676
rect 340432 231662 340814 231690
rect 341076 231662 341458 231690
rect 340144 229900 340196 229906
rect 340144 229842 340196 229848
rect 340432 221882 340460 231662
rect 340696 227316 340748 227322
rect 340696 227258 340748 227264
rect 340420 221876 340472 221882
rect 340420 221818 340472 221824
rect 339684 221604 339736 221610
rect 339684 221546 339736 221552
rect 340512 218884 340564 218890
rect 340512 218826 340564 218832
rect 338672 218068 338724 218074
rect 338672 218010 338724 218016
rect 338856 218068 338908 218074
rect 338856 218010 338908 218016
rect 339408 218068 339460 218074
rect 339408 218010 339460 218016
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337166 217110 337240 217138
rect 337994 217246 338068 217274
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338868 217138 338896 218010
rect 339696 217138 339724 218010
rect 340524 217138 340552 218826
rect 340708 218074 340736 227258
rect 341076 220386 341104 231662
rect 342088 223514 342116 231676
rect 342272 231662 342746 231690
rect 342916 231662 343390 231690
rect 343836 231662 344034 231690
rect 342076 223508 342128 223514
rect 342076 223450 342128 223456
rect 342272 223378 342300 231662
rect 342916 229094 342944 231662
rect 342640 229066 342944 229094
rect 342260 223372 342312 223378
rect 342260 223314 342312 223320
rect 341340 221604 341392 221610
rect 341340 221546 341392 221552
rect 341064 220380 341116 220386
rect 341064 220322 341116 220328
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341352 217274 341380 221546
rect 342168 221468 342220 221474
rect 342168 221410 342220 221416
rect 342180 217274 342208 221410
rect 342640 220250 342668 229066
rect 342812 223440 342864 223446
rect 342812 223382 342864 223388
rect 342628 220244 342680 220250
rect 342628 220186 342680 220192
rect 342824 219298 342852 223382
rect 343836 222018 343864 231662
rect 344664 225758 344692 231676
rect 345308 229770 345336 231676
rect 345664 229900 345716 229906
rect 345664 229842 345716 229848
rect 345296 229764 345348 229770
rect 345296 229706 345348 229712
rect 344652 225752 344704 225758
rect 344652 225694 344704 225700
rect 344652 223168 344704 223174
rect 344652 223110 344704 223116
rect 343824 222012 343876 222018
rect 343824 221954 343876 221960
rect 342996 220380 343048 220386
rect 342996 220322 343048 220328
rect 342812 219292 342864 219298
rect 342812 219234 342864 219240
rect 343008 217274 343036 220322
rect 343824 219156 343876 219162
rect 343824 219098 343876 219104
rect 338822 217110 338896 217138
rect 339650 217110 339724 217138
rect 340478 217110 340552 217138
rect 341306 217246 341380 217274
rect 342134 217246 342208 217274
rect 342962 217246 343036 217274
rect 338822 216988 338850 217110
rect 339650 216988 339678 217110
rect 340478 216988 340506 217110
rect 341306 216988 341334 217246
rect 342134 216988 342162 217246
rect 342962 216988 342990 217246
rect 343836 217138 343864 219098
rect 344664 217274 344692 223110
rect 345676 219026 345704 229842
rect 345952 224806 345980 231676
rect 346596 225622 346624 231676
rect 346584 225616 346636 225622
rect 346584 225558 346636 225564
rect 347044 225616 347096 225622
rect 347044 225558 347096 225564
rect 345940 224800 345992 224806
rect 345940 224742 345992 224748
rect 346216 224528 346268 224534
rect 346216 224470 346268 224476
rect 345664 219020 345716 219026
rect 345664 218962 345716 218968
rect 345480 218068 345532 218074
rect 345480 218010 345532 218016
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345492 217138 345520 218010
rect 346228 217274 346256 224470
rect 347056 218074 347084 225558
rect 347240 224398 347268 231676
rect 347228 224392 347280 224398
rect 347228 224334 347280 224340
rect 347884 223446 347912 231676
rect 347872 223440 347924 223446
rect 347872 223382 347924 223388
rect 347228 223304 347280 223310
rect 347228 223246 347280 223252
rect 347240 219434 347268 223246
rect 348528 222902 348556 231676
rect 349172 228546 349200 231676
rect 349160 228540 349212 228546
rect 349160 228482 349212 228488
rect 349816 227186 349844 231676
rect 350460 230178 350488 231676
rect 350448 230172 350500 230178
rect 350448 230114 350500 230120
rect 351104 229090 351132 231676
rect 351472 231662 351762 231690
rect 352116 231662 352406 231690
rect 351092 229084 351144 229090
rect 351092 229026 351144 229032
rect 350448 228540 350500 228546
rect 350448 228482 350500 228488
rect 349804 227180 349856 227186
rect 349804 227122 349856 227128
rect 350264 226364 350316 226370
rect 350264 226306 350316 226312
rect 348516 222896 348568 222902
rect 348516 222838 348568 222844
rect 349068 222896 349120 222902
rect 349068 222838 349120 222844
rect 348792 220244 348844 220250
rect 348792 220186 348844 220192
rect 347228 219428 347280 219434
rect 347228 219370 347280 219376
rect 347228 219020 347280 219026
rect 347228 218962 347280 218968
rect 347044 218068 347096 218074
rect 347044 218010 347096 218016
rect 347240 217274 347268 218962
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 346228 217246 346302 217274
rect 345446 217110 345520 217138
rect 345446 216988 345474 217110
rect 346274 216988 346302 217246
rect 347102 217246 347268 217274
rect 347102 216988 347130 217246
rect 347976 217138 348004 218010
rect 348804 217274 348832 220186
rect 349080 218074 349108 222838
rect 350276 219434 350304 226306
rect 350460 219434 350488 228482
rect 351092 226500 351144 226506
rect 351092 226442 351144 226448
rect 349620 219428 349672 219434
rect 350276 219406 350396 219434
rect 350460 219428 350592 219434
rect 350460 219406 350540 219428
rect 349620 219370 349672 219376
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 347930 217110 348004 217138
rect 348758 217246 348832 217274
rect 347930 216988 347958 217110
rect 348758 216988 348786 217246
rect 349632 217138 349660 219370
rect 350368 217274 350396 219406
rect 350540 219370 350592 219376
rect 351104 218754 351132 226442
rect 351472 223038 351500 231662
rect 351736 229764 351788 229770
rect 351736 229706 351788 229712
rect 351748 226370 351776 229706
rect 351736 226364 351788 226370
rect 351736 226306 351788 226312
rect 351460 223032 351512 223038
rect 351460 222974 351512 222980
rect 351276 221876 351328 221882
rect 351276 221818 351328 221824
rect 351092 218748 351144 218754
rect 351092 218690 351144 218696
rect 351288 217274 351316 221818
rect 352116 220114 352144 231662
rect 353036 226506 353064 231676
rect 353024 226500 353076 226506
rect 353024 226442 353076 226448
rect 353680 226030 353708 231676
rect 353864 231662 354338 231690
rect 353668 226024 353720 226030
rect 353668 225966 353720 225972
rect 352932 225752 352984 225758
rect 352932 225694 352984 225700
rect 352104 220108 352156 220114
rect 352104 220050 352156 220056
rect 352104 219428 352156 219434
rect 352104 219370 352156 219376
rect 350368 217246 350442 217274
rect 349586 217110 349660 217138
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351316 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 219370
rect 352944 217274 352972 225694
rect 353864 223122 353892 231662
rect 354968 228410 354996 231676
rect 355612 230042 355640 231676
rect 355600 230036 355652 230042
rect 355600 229978 355652 229984
rect 354956 228404 355008 228410
rect 354956 228346 355008 228352
rect 355324 228404 355376 228410
rect 355324 228346 355376 228352
rect 354588 226024 354640 226030
rect 354588 225966 354640 225972
rect 353772 223094 353892 223122
rect 353772 222154 353800 223094
rect 353944 223032 353996 223038
rect 353944 222974 353996 222980
rect 353760 222148 353812 222154
rect 353760 222090 353812 222096
rect 353956 219162 353984 222974
rect 353944 219156 353996 219162
rect 353944 219098 353996 219104
rect 353760 218748 353812 218754
rect 353760 218690 353812 218696
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218690
rect 354600 217274 354628 225966
rect 355336 219434 355364 228346
rect 356256 227458 356284 231676
rect 356244 227452 356296 227458
rect 356244 227394 356296 227400
rect 355876 227180 355928 227186
rect 355876 227122 355928 227128
rect 355324 219428 355376 219434
rect 355324 219370 355376 219376
rect 355888 218074 355916 227122
rect 356900 224670 356928 231676
rect 357072 227452 357124 227458
rect 357072 227394 357124 227400
rect 356888 224664 356940 224670
rect 356888 224606 356940 224612
rect 357084 222034 357112 227394
rect 357544 225894 357572 231676
rect 357912 231662 358202 231690
rect 357532 225888 357584 225894
rect 357532 225830 357584 225836
rect 357912 223310 357940 231662
rect 358832 228682 358860 231676
rect 359016 231662 359490 231690
rect 358820 228676 358872 228682
rect 358820 228618 358872 228624
rect 358084 224256 358136 224262
rect 358084 224198 358136 224204
rect 357900 223304 357952 223310
rect 357900 223246 357952 223252
rect 356992 222006 357112 222034
rect 356992 218074 357020 222006
rect 357164 221740 357216 221746
rect 357164 221682 357216 221688
rect 355416 218068 355468 218074
rect 355416 218010 355468 218016
rect 355876 218068 355928 218074
rect 355876 218010 355928 218016
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 356980 218068 357032 218074
rect 356980 218010 357032 218016
rect 353726 217110 353800 217138
rect 354554 217246 354628 217274
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355428 217138 355456 218010
rect 356256 217138 356284 218010
rect 357176 217274 357204 221682
rect 357900 220652 357952 220658
rect 357900 220594 357952 220600
rect 357912 217274 357940 220594
rect 358096 218890 358124 224198
rect 359016 220522 359044 231662
rect 359924 228676 359976 228682
rect 359924 228618 359976 228624
rect 359004 220516 359056 220522
rect 359004 220458 359056 220464
rect 358820 220108 358872 220114
rect 358820 220050 358872 220056
rect 358832 219434 358860 220050
rect 358740 219406 358860 219434
rect 359936 219434 359964 228618
rect 360120 227050 360148 231676
rect 360764 229906 360792 231676
rect 360752 229900 360804 229906
rect 360752 229842 360804 229848
rect 361212 229900 361264 229906
rect 361212 229842 361264 229848
rect 361224 229094 361252 229842
rect 361040 229066 361252 229094
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359936 219406 360148 219434
rect 358084 218884 358136 218890
rect 358084 218826 358136 218832
rect 358740 217274 358768 219406
rect 360120 218074 360148 219406
rect 361040 218074 361068 229066
rect 361408 227322 361436 231676
rect 361776 231662 362066 231690
rect 362328 231662 362710 231690
rect 361396 227316 361448 227322
rect 361396 227258 361448 227264
rect 361212 224392 361264 224398
rect 361212 224334 361264 224340
rect 359556 218068 359608 218074
rect 359556 218010 359608 218016
rect 360108 218068 360160 218074
rect 360108 218010 360160 218016
rect 360384 218068 360436 218074
rect 360384 218010 360436 218016
rect 361028 218068 361080 218074
rect 361028 218010 361080 218016
rect 355382 217110 355456 217138
rect 356210 217110 356284 217138
rect 357038 217246 357204 217274
rect 357866 217246 357940 217274
rect 358694 217246 358768 217274
rect 355382 216988 355410 217110
rect 356210 216988 356238 217110
rect 357038 216988 357066 217246
rect 357866 216988 357894 217246
rect 358694 216988 358722 217246
rect 359568 217138 359596 218010
rect 360396 217138 360424 218010
rect 361224 217274 361252 224334
rect 361776 221610 361804 231662
rect 362328 224126 362356 231662
rect 362776 227044 362828 227050
rect 362776 226986 362828 226992
rect 362316 224120 362368 224126
rect 362316 224062 362368 224068
rect 361764 221604 361816 221610
rect 361764 221546 361816 221552
rect 362040 219428 362092 219434
rect 362040 219370 362092 219376
rect 359522 217110 359596 217138
rect 360350 217110 360424 217138
rect 361178 217246 361252 217274
rect 359522 216988 359550 217110
rect 360350 216988 360378 217110
rect 361178 216988 361206 217246
rect 362052 217138 362080 219370
rect 362788 217274 362816 226986
rect 363340 224262 363368 231676
rect 363524 231662 363998 231690
rect 363524 229094 363552 231662
rect 363432 229066 363552 229094
rect 363432 224346 363460 229066
rect 363604 224664 363656 224670
rect 363604 224606 363656 224612
rect 363432 224318 363552 224346
rect 363328 224256 363380 224262
rect 363328 224198 363380 224204
rect 363524 220402 363552 224318
rect 363432 220386 363552 220402
rect 363420 220380 363552 220386
rect 363472 220374 363552 220380
rect 363420 220322 363472 220328
rect 363616 219026 363644 224606
rect 364628 223174 364656 231676
rect 364812 231662 365286 231690
rect 364616 223168 364668 223174
rect 364616 223110 364668 223116
rect 364812 221474 364840 231662
rect 365536 223168 365588 223174
rect 365536 223110 365588 223116
rect 364800 221468 364852 221474
rect 364800 221410 364852 221416
rect 363604 219020 363656 219026
rect 363604 218962 363656 218968
rect 363696 218884 363748 218890
rect 363696 218826 363748 218832
rect 362788 217246 362862 217274
rect 362006 217110 362080 217138
rect 362006 216988 362034 217110
rect 362834 216988 362862 217246
rect 363708 217138 363736 218826
rect 365352 218204 365404 218210
rect 365352 218146 365404 218152
rect 364524 218068 364576 218074
rect 364524 218010 364576 218016
rect 364536 217138 364564 218010
rect 365364 217138 365392 218146
rect 365548 218074 365576 223110
rect 365916 223038 365944 231676
rect 366560 224534 366588 231676
rect 366548 224528 366600 224534
rect 366548 224470 366600 224476
rect 366732 224256 366784 224262
rect 366732 224198 366784 224204
rect 365904 223032 365956 223038
rect 365904 222974 365956 222980
rect 366744 218074 366772 224198
rect 366916 223032 366968 223038
rect 366916 222974 366968 222980
rect 365536 218068 365588 218074
rect 365536 218010 365588 218016
rect 366180 218068 366232 218074
rect 366180 218010 366232 218016
rect 366732 218068 366784 218074
rect 366732 218010 366784 218016
rect 366192 217138 366220 218010
rect 366928 217274 366956 222974
rect 367204 222902 367232 231676
rect 367848 225622 367876 231676
rect 367836 225616 367888 225622
rect 367836 225558 367888 225564
rect 368492 224670 368520 231676
rect 369136 228546 369164 231676
rect 369320 231662 369794 231690
rect 369964 231662 370438 231690
rect 369124 228540 369176 228546
rect 369124 228482 369176 228488
rect 369124 225004 369176 225010
rect 369124 224946 369176 224952
rect 368480 224664 368532 224670
rect 368480 224606 368532 224612
rect 367192 222896 367244 222902
rect 367192 222838 367244 222844
rect 368388 222896 368440 222902
rect 368388 222838 368440 222844
rect 367652 222012 367704 222018
rect 367652 221954 367704 221960
rect 367664 219434 367692 221954
rect 367652 219428 367704 219434
rect 367652 219370 367704 219376
rect 368400 218074 368428 222838
rect 368664 219020 368716 219026
rect 368664 218962 368716 218968
rect 367836 218068 367888 218074
rect 367836 218010 367888 218016
rect 368388 218068 368440 218074
rect 368388 218010 368440 218016
rect 366928 217246 367002 217274
rect 363662 217110 363736 217138
rect 364490 217110 364564 217138
rect 365318 217110 365392 217138
rect 366146 217110 366220 217138
rect 363662 216988 363690 217110
rect 364490 216988 364518 217110
rect 365318 216988 365346 217110
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367848 217138 367876 218010
rect 368676 217138 368704 218962
rect 369136 218754 369164 224946
rect 369320 221882 369348 231662
rect 369308 221876 369360 221882
rect 369308 221818 369360 221824
rect 369492 221604 369544 221610
rect 369492 221546 369544 221552
rect 369124 218748 369176 218754
rect 369124 218690 369176 218696
rect 369504 217274 369532 221546
rect 369964 220250 369992 231662
rect 371068 229770 371096 231676
rect 371056 229764 371108 229770
rect 371056 229706 371108 229712
rect 371712 229094 371740 231676
rect 371620 229066 371740 229094
rect 371056 228540 371108 228546
rect 371056 228482 371108 228488
rect 369952 220244 370004 220250
rect 369952 220186 370004 220192
rect 370504 220244 370556 220250
rect 370504 220186 370556 220192
rect 370516 218890 370544 220186
rect 370504 218884 370556 218890
rect 370504 218826 370556 218832
rect 370320 218748 370372 218754
rect 370320 218690 370372 218696
rect 370332 217274 370360 218690
rect 367802 217110 367876 217138
rect 368630 217110 368704 217138
rect 369458 217246 369532 217274
rect 370286 217246 370360 217274
rect 371068 217274 371096 228482
rect 371620 225758 371648 229066
rect 372356 226030 372384 231676
rect 373000 228410 373028 231676
rect 372988 228404 373040 228410
rect 372988 228346 373040 228352
rect 373448 228404 373500 228410
rect 373448 228346 373500 228352
rect 372344 226024 372396 226030
rect 372344 225966 372396 225972
rect 371608 225752 371660 225758
rect 371608 225694 371660 225700
rect 371792 225752 371844 225758
rect 371792 225694 371844 225700
rect 371804 218210 371832 225694
rect 372528 225616 372580 225622
rect 372528 225558 372580 225564
rect 371792 218204 371844 218210
rect 371792 218146 371844 218152
rect 372540 218074 372568 225558
rect 373460 218074 373488 228346
rect 373644 225010 373672 231676
rect 374288 227458 374316 231676
rect 374472 231662 374946 231690
rect 374276 227452 374328 227458
rect 374276 227394 374328 227400
rect 373816 225888 373868 225894
rect 373816 225830 373868 225836
rect 373632 225004 373684 225010
rect 373632 224946 373684 224952
rect 373828 219434 373856 225830
rect 374472 220658 374500 231662
rect 374644 230444 374696 230450
rect 374644 230386 374696 230392
rect 374656 221746 374684 230386
rect 375576 227186 375604 231676
rect 376220 230450 376248 231676
rect 376208 230444 376260 230450
rect 376208 230386 376260 230392
rect 376024 228812 376076 228818
rect 376024 228754 376076 228760
rect 375564 227180 375616 227186
rect 375564 227122 375616 227128
rect 374644 221740 374696 221746
rect 374644 221682 374696 221688
rect 375288 221468 375340 221474
rect 375288 221410 375340 221416
rect 374460 220652 374512 220658
rect 374460 220594 374512 220600
rect 373644 219406 373856 219434
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 373448 218068 373500 218074
rect 373448 218010 373500 218016
rect 371068 217246 371142 217274
rect 367802 216988 367830 217110
rect 368630 216988 368658 217110
rect 369458 216988 369486 217246
rect 370286 216988 370314 217246
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373644 217274 373672 219406
rect 374460 218204 374512 218210
rect 374460 218146 374512 218152
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217246 373672 217274
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217246
rect 374472 217138 374500 218146
rect 375300 217274 375328 221410
rect 376036 218210 376064 228754
rect 376864 228682 376892 231676
rect 376852 228676 376904 228682
rect 376852 228618 376904 228624
rect 376668 227180 376720 227186
rect 376668 227122 376720 227128
rect 376024 218204 376076 218210
rect 376024 218146 376076 218152
rect 376680 218074 376708 227122
rect 377508 224398 377536 231676
rect 378166 231662 378364 231690
rect 377680 229764 377732 229770
rect 377680 229706 377732 229712
rect 377692 225894 377720 229706
rect 377680 225888 377732 225894
rect 377680 225830 377732 225836
rect 377864 225888 377916 225894
rect 377864 225830 377916 225836
rect 377496 224392 377548 224398
rect 377496 224334 377548 224340
rect 377404 224120 377456 224126
rect 377404 224062 377456 224068
rect 377416 219026 377444 224062
rect 377876 219434 377904 225830
rect 378336 220114 378364 231662
rect 378796 229906 378824 231676
rect 378784 229900 378836 229906
rect 378784 229842 378836 229848
rect 379440 227050 379468 231676
rect 379624 231662 380098 231690
rect 380268 231662 380742 231690
rect 381096 231662 381386 231690
rect 381648 231662 382030 231690
rect 382384 231662 382674 231690
rect 382844 231662 383318 231690
rect 379428 227044 379480 227050
rect 379428 226986 379480 226992
rect 379244 224392 379296 224398
rect 379244 224334 379296 224340
rect 378324 220108 378376 220114
rect 378324 220050 378376 220056
rect 377784 219406 377904 219434
rect 377404 219020 377456 219026
rect 377404 218962 377456 218968
rect 376944 218884 376996 218890
rect 376944 218826 376996 218832
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376668 218068 376720 218074
rect 376668 218010 376720 218016
rect 374426 217110 374500 217138
rect 375254 217246 375328 217274
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217138 376984 218826
rect 377784 217274 377812 219406
rect 379256 218074 379284 224334
rect 379624 223174 379652 231662
rect 379612 223168 379664 223174
rect 379612 223110 379664 223116
rect 380072 223168 380124 223174
rect 380072 223110 380124 223116
rect 379428 220108 379480 220114
rect 379428 220050 379480 220056
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 379244 218068 379296 218074
rect 379244 218010 379296 218016
rect 376082 217110 376156 217138
rect 376910 217110 376984 217138
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217110
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379440 217274 379468 220050
rect 380084 218754 380112 223110
rect 380268 222018 380296 231662
rect 380256 222012 380308 222018
rect 380256 221954 380308 221960
rect 381096 220250 381124 231662
rect 381648 224262 381676 231662
rect 382096 227316 382148 227322
rect 382096 227258 382148 227264
rect 381636 224256 381688 224262
rect 381636 224198 381688 224204
rect 381084 220244 381136 220250
rect 381084 220186 381136 220192
rect 380256 219428 380308 219434
rect 380256 219370 380308 219376
rect 380072 218748 380124 218754
rect 380072 218690 380124 218696
rect 378566 217110 378640 217138
rect 379394 217246 379468 217274
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 219370
rect 381912 218204 381964 218210
rect 381912 218146 381964 218152
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381096 217138 381124 218010
rect 381924 217138 381952 218146
rect 382108 218074 382136 227258
rect 382384 222902 382412 231662
rect 382844 229094 382872 231662
rect 383948 229094 383976 231676
rect 384132 231662 384606 231690
rect 384132 229094 384160 231662
rect 382752 229066 382872 229094
rect 383856 229066 383976 229094
rect 384040 229066 384160 229094
rect 382752 225758 382780 229066
rect 382740 225752 382792 225758
rect 382740 225694 382792 225700
rect 382924 225752 382976 225758
rect 382924 225694 382976 225700
rect 382372 222896 382424 222902
rect 382372 222838 382424 222844
rect 382740 218884 382792 218890
rect 382740 218826 382792 218832
rect 382096 218068 382148 218074
rect 382096 218010 382148 218016
rect 382752 217138 382780 218826
rect 382936 218210 382964 225694
rect 383856 223038 383884 229066
rect 383844 223032 383896 223038
rect 383844 222974 383896 222980
rect 383476 222896 383528 222902
rect 383476 222838 383528 222844
rect 383488 218890 383516 222838
rect 384040 221610 384068 229066
rect 385236 228546 385264 231676
rect 385224 228540 385276 228546
rect 385224 228482 385276 228488
rect 385880 224126 385908 231676
rect 386052 228540 386104 228546
rect 386052 228482 386104 228488
rect 385868 224120 385920 224126
rect 385868 224062 385920 224068
rect 384212 223032 384264 223038
rect 384212 222974 384264 222980
rect 384028 221604 384080 221610
rect 384028 221546 384080 221552
rect 384224 219434 384252 222974
rect 384396 221604 384448 221610
rect 384396 221546 384448 221552
rect 384212 219428 384264 219434
rect 384212 219370 384264 219376
rect 383476 218884 383528 218890
rect 383476 218826 383528 218832
rect 383568 218748 383620 218754
rect 383568 218690 383620 218696
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 383580 217138 383608 218690
rect 384408 217274 384436 221546
rect 385224 220788 385276 220794
rect 385224 220730 385276 220736
rect 385236 217274 385264 220730
rect 386064 217274 386092 228482
rect 386524 223174 386552 231676
rect 387168 228410 387196 231676
rect 387432 230376 387484 230382
rect 387432 230318 387484 230324
rect 387156 228404 387208 228410
rect 387156 228346 387208 228352
rect 387444 225622 387472 230318
rect 387812 228818 387840 231676
rect 388456 230382 388484 231676
rect 388444 230376 388496 230382
rect 388444 230318 388496 230324
rect 389100 229770 389128 231676
rect 389088 229764 389140 229770
rect 389088 229706 389140 229712
rect 388628 229628 388680 229634
rect 388628 229570 388680 229576
rect 388640 229094 388668 229570
rect 388640 229066 388760 229094
rect 387800 228812 387852 228818
rect 387800 228754 387852 228760
rect 388536 226364 388588 226370
rect 388536 226306 388588 226312
rect 387432 225616 387484 225622
rect 387432 225558 387484 225564
rect 387708 224528 387760 224534
rect 387708 224470 387760 224476
rect 386512 223168 386564 223174
rect 386512 223110 386564 223116
rect 386880 219020 386932 219026
rect 386880 218962 386932 218968
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217110 381952 217138
rect 382706 217110 382780 217138
rect 383534 217110 383608 217138
rect 384362 217246 384436 217274
rect 385190 217246 385264 217274
rect 386018 217246 386092 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217110
rect 382706 216988 382734 217110
rect 383534 216988 383562 217110
rect 384362 216988 384390 217246
rect 385190 216988 385218 217246
rect 386018 216988 386046 217246
rect 386892 217138 386920 218962
rect 387720 217274 387748 224470
rect 388548 218890 388576 226306
rect 388732 220794 388760 229066
rect 389744 227186 389772 231676
rect 390008 228404 390060 228410
rect 390008 228346 390060 228352
rect 389732 227180 389784 227186
rect 389732 227122 389784 227128
rect 388720 220788 388772 220794
rect 388720 220730 388772 220736
rect 388720 220244 388772 220250
rect 388720 220186 388772 220192
rect 388536 218884 388588 218890
rect 388536 218826 388588 218832
rect 388732 217274 388760 220186
rect 390020 218074 390048 228346
rect 390388 225894 390416 231676
rect 390756 231662 391046 231690
rect 390376 225888 390428 225894
rect 390376 225830 390428 225836
rect 390192 225616 390244 225622
rect 390192 225558 390244 225564
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 390008 218068 390060 218074
rect 390008 218010 390060 218016
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 388502 217246 388760 217274
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388502 216988 388530 217246
rect 389376 217138 389404 218010
rect 390204 217274 390232 225558
rect 390756 221474 390784 231662
rect 391676 226370 391704 231676
rect 392136 231662 392334 231690
rect 391848 227044 391900 227050
rect 391848 226986 391900 226992
rect 391664 226364 391716 226370
rect 391664 226306 391716 226312
rect 391020 221740 391072 221746
rect 391020 221682 391072 221688
rect 390744 221468 390796 221474
rect 390744 221410 390796 221416
rect 391032 217274 391060 221682
rect 391860 219434 391888 226986
rect 392136 220114 392164 231662
rect 392964 227322 392992 231676
rect 392952 227316 393004 227322
rect 392952 227258 393004 227264
rect 393136 227180 393188 227186
rect 393136 227122 393188 227128
rect 392124 220108 392176 220114
rect 392124 220050 392176 220056
rect 389330 217110 389404 217138
rect 390158 217246 390232 217274
rect 390986 217246 391060 217274
rect 391768 219406 391888 219434
rect 391768 217274 391796 219406
rect 393148 218074 393176 227122
rect 393608 224398 393636 231676
rect 393976 231662 394266 231690
rect 393596 224392 393648 224398
rect 393596 224334 393648 224340
rect 393976 223038 394004 231662
rect 394332 225888 394384 225894
rect 394332 225830 394384 225836
rect 393964 223032 394016 223038
rect 393964 222974 394016 222980
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393136 218068 393188 218074
rect 393136 218010 393188 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 391768 217246 391842 217274
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217274 394372 225830
rect 394516 224256 394568 224262
rect 394516 224198 394568 224204
rect 394528 218074 394556 224198
rect 394896 222902 394924 231676
rect 395172 231662 395554 231690
rect 394884 222896 394936 222902
rect 394884 222838 394936 222844
rect 395172 221610 395200 231662
rect 396184 225758 396212 231676
rect 396368 231662 396842 231690
rect 396172 225752 396224 225758
rect 396172 225694 396224 225700
rect 395804 222896 395856 222902
rect 395804 222838 395856 222844
rect 395160 221604 395212 221610
rect 395160 221546 395212 221552
rect 395816 218074 395844 222838
rect 395988 220108 396040 220114
rect 395988 220050 396040 220056
rect 394516 218068 394568 218074
rect 394516 218010 394568 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395804 218068 395856 218074
rect 395804 218010 395856 218016
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217246 394372 217274
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217246
rect 395172 217138 395200 218010
rect 396000 217274 396028 220050
rect 396368 219434 396396 231662
rect 397472 228546 397500 231676
rect 397840 231662 398130 231690
rect 397460 228540 397512 228546
rect 397460 228482 397512 228488
rect 397840 224534 397868 231662
rect 398104 230376 398156 230382
rect 398104 230318 398156 230324
rect 397828 224528 397880 224534
rect 397828 224470 397880 224476
rect 396816 221468 396868 221474
rect 396816 221410 396868 221416
rect 396276 219406 396396 219434
rect 396276 218754 396304 219406
rect 396264 218748 396316 218754
rect 396264 218690 396316 218696
rect 396828 217274 396856 221410
rect 398116 219026 398144 230318
rect 398760 229634 398788 231676
rect 399404 230382 399432 231676
rect 399392 230376 399444 230382
rect 399392 230318 399444 230324
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 398748 229628 398800 229634
rect 398748 229570 398800 229576
rect 399864 219434 399892 229706
rect 400048 228410 400076 231676
rect 400416 231662 400706 231690
rect 400968 231662 401350 231690
rect 400036 228404 400088 228410
rect 400036 228346 400088 228352
rect 400128 228132 400180 228138
rect 400128 228074 400180 228080
rect 400140 219434 400168 228074
rect 400416 221746 400444 231662
rect 400404 221740 400456 221746
rect 400404 221682 400456 221688
rect 400588 221604 400640 221610
rect 400588 221546 400640 221552
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 398104 219020 398156 219026
rect 398104 218962 398156 218968
rect 398472 218612 398524 218618
rect 398472 218554 398524 218560
rect 397644 218068 397696 218074
rect 397644 218010 397696 218016
rect 395126 217110 395200 217138
rect 395954 217246 396028 217274
rect 396782 217246 396856 217274
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396782 216988 396810 217246
rect 397656 217138 397684 218010
rect 398484 217138 398512 218554
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 400600 218074 400628 221546
rect 400968 220250 400996 231662
rect 401980 225622 402008 231676
rect 402624 227322 402652 231676
rect 402796 228404 402848 228410
rect 402796 228346 402848 228352
rect 402612 227316 402664 227322
rect 402612 227258 402664 227264
rect 402244 227180 402296 227186
rect 402244 227122 402296 227128
rect 401968 225616 402020 225622
rect 401968 225558 402020 225564
rect 400956 220244 401008 220250
rect 400956 220186 401008 220192
rect 401784 218204 401836 218210
rect 401784 218146 401836 218152
rect 400588 218068 400640 218074
rect 400588 218010 400640 218016
rect 400956 218068 401008 218074
rect 400956 218010 401008 218016
rect 400048 217246 400122 217274
rect 397610 217110 397684 217138
rect 398438 217110 398512 217138
rect 399266 217110 399340 217138
rect 397610 216988 397638 217110
rect 398438 216988 398466 217110
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218010
rect 401796 217138 401824 218146
rect 402256 218074 402284 227122
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218068 402296 218074
rect 402244 218010 402296 218016
rect 402624 217138 402652 218826
rect 402808 218210 402836 228346
rect 403268 225894 403296 231676
rect 403544 231662 403926 231690
rect 403544 227050 403572 231662
rect 403532 227044 403584 227050
rect 403532 226986 403584 226992
rect 403992 226500 404044 226506
rect 403992 226442 404044 226448
rect 403256 225888 403308 225894
rect 403256 225830 403308 225836
rect 402796 218204 402848 218210
rect 402796 218146 402848 218152
rect 404004 218074 404032 226442
rect 404176 225004 404228 225010
rect 404176 224946 404228 224952
rect 403440 218068 403492 218074
rect 403440 218010 403492 218016
rect 403992 218068 404044 218074
rect 403992 218010 404044 218016
rect 403452 217138 403480 218010
rect 404188 217274 404216 224946
rect 404556 224262 404584 231676
rect 404740 231662 405214 231690
rect 404544 224256 404596 224262
rect 404544 224198 404596 224204
rect 404740 220114 404768 231662
rect 405556 224256 405608 224262
rect 405556 224198 405608 224204
rect 404728 220108 404780 220114
rect 404728 220050 404780 220056
rect 405568 218074 405596 224198
rect 405844 221610 405872 231676
rect 406488 222902 406516 231676
rect 407146 231662 407344 231690
rect 406752 223576 406804 223582
rect 406752 223518 406804 223524
rect 406476 222896 406528 222902
rect 406476 222838 406528 222844
rect 405832 221604 405884 221610
rect 405832 221546 405884 221552
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405096 218068 405148 218074
rect 405096 218010 405148 218016
rect 405556 218068 405608 218074
rect 405556 218010 405608 218016
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405108 217138 405136 218010
rect 405936 217274 405964 219438
rect 406764 217274 406792 223518
rect 407316 221474 407344 231662
rect 407776 228546 407804 231676
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 408420 227186 408448 231676
rect 408696 231662 409078 231690
rect 408408 227180 408460 227186
rect 408408 227122 408460 227128
rect 408696 226370 408724 231662
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228540 409840 228546
rect 409788 228482 409840 228488
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 407764 226364 407816 226370
rect 407764 226306 407816 226312
rect 408684 226364 408736 226370
rect 408684 226306 408736 226312
rect 407304 221468 407356 221474
rect 407304 221410 407356 221416
rect 407776 218618 407804 226306
rect 408408 221468 408460 221474
rect 408408 221410 408460 221416
rect 407764 218612 407816 218618
rect 407764 218554 407816 218560
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 405062 217110 405136 217138
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217110
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 221410
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228482
rect 410352 227798 410380 231676
rect 410720 231662 411010 231690
rect 410720 229094 410748 231662
rect 410892 229900 410944 229906
rect 410892 229842 410944 229848
rect 410904 229094 410932 229842
rect 410628 229066 410748 229094
rect 410812 229066 410932 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410628 225010 410656 229066
rect 410616 225004 410668 225010
rect 410616 224946 410668 224952
rect 410812 219434 410840 229066
rect 411640 228410 411668 231676
rect 411628 228404 411680 228410
rect 411628 228346 411680 228352
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 410984 225616 411036 225622
rect 410984 225558 411036 225564
rect 410996 219434 411024 225558
rect 410720 219406 410840 219434
rect 410904 219406 411024 219434
rect 410720 218074 410748 219406
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 219406
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412284 226506 412312 231676
rect 412744 231662 412942 231690
rect 412548 227044 412600 227050
rect 412548 226986 412600 226992
rect 412272 226500 412324 226506
rect 412272 226442 412324 226448
rect 412560 218890 412588 226986
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229356 413888 229362
rect 413836 229298 413888 229304
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412548 218884 412600 218890
rect 412548 218826 412600 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229298
rect 414216 224262 414244 231676
rect 414204 224256 414256 224262
rect 414204 224198 414256 224204
rect 414860 223582 414888 231676
rect 415504 228546 415532 231676
rect 415492 228540 415544 228546
rect 415492 228482 415544 228488
rect 415032 228064 415084 228070
rect 415032 228006 415084 228012
rect 414848 223576 414900 223582
rect 414848 223518 414900 223524
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 228006
rect 416148 225622 416176 231676
rect 416792 229094 416820 231676
rect 417436 229906 417464 231676
rect 417712 231662 418094 231690
rect 418356 231662 418738 231690
rect 417424 229900 417476 229906
rect 417424 229842 417476 229848
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416688 227928 416740 227934
rect 416688 227870 416740 227876
rect 416136 225616 416188 225622
rect 416136 225558 416188 225564
rect 416504 225004 416556 225010
rect 416504 224946 416556 224952
rect 416516 219434 416544 224946
rect 416700 219434 416728 227870
rect 416884 221474 416912 229066
rect 417160 229066 417740 229094
rect 416872 221468 416924 221474
rect 416872 221410 416924 221416
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418356 224954 418384 231662
rect 419368 227050 419396 231676
rect 420012 229362 420040 231676
rect 420000 229356 420052 229362
rect 420000 229298 420052 229304
rect 420656 227934 420684 231676
rect 421024 231662 421314 231690
rect 420644 227928 420696 227934
rect 420644 227870 420696 227876
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 419356 227044 419408 227050
rect 419356 226986 419408 226992
rect 418172 224926 418384 224954
rect 418172 220794 418200 224926
rect 418344 220856 418396 220862
rect 418344 220798 418396 220804
rect 418160 220788 418212 220794
rect 418160 220730 418212 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 418356 217274 418384 220798
rect 420656 219434 420684 227734
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420656 219406 420776 219434
rect 419172 219292 419224 219298
rect 419172 219234 419224 219240
rect 419184 217274 419212 219234
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 417482 217110 417556 217138
rect 418310 217246 418384 217274
rect 419138 217246 419212 217274
rect 417482 216988 417510 217110
rect 418310 216988 418338 217246
rect 419138 216988 419166 217246
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 228070 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 421932 228064 421984 228070
rect 421932 228006 421984 228012
rect 422220 225010 422248 229066
rect 422208 225004 422260 225010
rect 422208 224946 422260 224952
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423496 229152 423548 229158
rect 423496 229094 423548 229100
rect 423508 219434 423536 229094
rect 423876 227798 423904 231676
rect 424060 231662 424534 231690
rect 423864 227792 423916 227798
rect 423864 227734 423916 227740
rect 424060 220862 424088 231662
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 222148 425020 222154
rect 424968 222090 425020 222096
rect 424048 220856 424100 220862
rect 424048 220798 424100 220804
rect 422680 219406 422892 219434
rect 423324 219406 423536 219434
rect 422680 219298 422708 219406
rect 422668 219292 422720 219298
rect 422668 219234 422720 219240
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 419966 217110 420040 217138
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 219406
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 222090
rect 425440 218210 425468 231662
rect 426452 224330 426480 231676
rect 426820 231662 427110 231690
rect 426440 224324 426492 224330
rect 426440 224266 426492 224272
rect 426820 220114 426848 231662
rect 427740 229158 427768 231676
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 428384 229094 428412 231676
rect 428752 231662 429042 231690
rect 429304 231662 429686 231690
rect 429948 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 428384 229066 428504 229094
rect 426992 224324 427044 224330
rect 426992 224266 427044 224272
rect 426808 220108 426860 220114
rect 426808 220050 426860 220056
rect 426624 218476 426676 218482
rect 426624 218418 426676 218424
rect 425796 218340 425848 218346
rect 425796 218282 425848 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218282
rect 426636 217138 426664 218418
rect 427004 218074 427032 224266
rect 427912 224256 427964 224262
rect 427912 224198 427964 224204
rect 427924 218074 427952 224198
rect 428476 218346 428504 229066
rect 428752 224262 428780 231662
rect 428740 224256 428792 224262
rect 428740 224198 428792 224204
rect 429304 222154 429332 231662
rect 429292 222148 429344 222154
rect 429292 222090 429344 222096
rect 429948 219434 429976 231662
rect 430120 220244 430172 220250
rect 430120 220186 430172 220192
rect 429580 219406 429976 219434
rect 429580 218482 429608 219406
rect 429936 218748 429988 218754
rect 429936 218690 429988 218696
rect 429568 218476 429620 218482
rect 429568 218418 429620 218424
rect 428464 218340 428516 218346
rect 428464 218282 428516 218288
rect 428280 218204 428332 218210
rect 428280 218146 428332 218152
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 427912 218068 427964 218074
rect 427912 218010 427964 218016
rect 427464 217138 427492 218010
rect 428292 217138 428320 218146
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217138 429148 218010
rect 429948 217138 429976 218690
rect 430132 218210 430160 220186
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 220250 432092 231662
rect 432052 220244 432104 220250
rect 432052 220186 432104 220192
rect 431960 220108 432012 220114
rect 431960 220050 432012 220056
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 430120 218204 430172 218210
rect 430120 218146 430172 218152
rect 430592 218074 430620 219406
rect 430580 218068 430632 218074
rect 430580 218010 430632 218016
rect 430776 217274 430804 219406
rect 431972 218090 432000 220050
rect 432708 218754 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432696 218748 432748 218754
rect 432696 218690 432748 218696
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217110 428320 217138
rect 429074 217110 429148 217138
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217110
rect 429074 216988 429102 217110
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220114 434852 231676
rect 435192 231662 435482 231690
rect 436126 231662 436324 231690
rect 434812 220108 434864 220114
rect 434812 220050 434864 220056
rect 435192 219434 435220 231662
rect 434732 219406 435220 219434
rect 434732 218210 434760 219406
rect 434720 218204 434772 218210
rect 434720 218146 434772 218152
rect 434904 218204 434956 218210
rect 434904 218146 434956 218152
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218146
rect 436296 218074 436324 231662
rect 436572 231662 436770 231690
rect 437032 231662 437414 231690
rect 437584 231662 438058 231690
rect 436572 229094 436600 231662
rect 436572 229066 436692 229094
rect 435732 218068 435784 218074
rect 435732 218010 435784 218016
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436468 218068 436520 218074
rect 436468 218010 436520 218016
rect 435744 217138 435772 218010
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436480 217138 436508 218010
rect 436664 217546 436692 229066
rect 437032 219434 437060 231662
rect 437584 219434 437612 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 219434 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 219434 439360 230318
rect 436848 219406 437060 219434
rect 437492 219406 437612 219434
rect 438872 219406 438992 219434
rect 439056 219406 439360 219434
rect 436848 218210 436876 219406
rect 436836 218204 436888 218210
rect 436836 218146 436888 218152
rect 437492 218074 437520 219406
rect 438872 218074 438900 219406
rect 437480 218068 437532 218074
rect 437480 218010 437532 218016
rect 438216 218068 438268 218074
rect 438216 218010 438268 218016
rect 438860 218068 438912 218074
rect 438860 218010 438912 218016
rect 436664 217518 437336 217546
rect 437308 217274 437336 217518
rect 437308 217246 437382 217274
rect 436480 217110 436554 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217246
rect 438228 217138 438256 218010
rect 439056 217274 439084 219406
rect 440344 218074 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 218068 439924 218074
rect 439872 218010 439924 218016
rect 440332 218068 440384 218074
rect 440332 218010 440384 218016
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 218010
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 219434 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 219406 441752 219434
rect 441632 218090 441660 219406
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441540 218062 441660 218090
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441540 217138 441568 218062
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 229362 443868 231676
rect 444484 230178 444512 231676
rect 444668 231662 445142 231690
rect 444472 230172 444524 230178
rect 444472 230114 444524 230120
rect 443828 229356 443880 229362
rect 443828 229298 443880 229304
rect 444668 229094 444696 231662
rect 444840 229356 444892 229362
rect 444840 229298 444892 229304
rect 444852 229094 444880 229298
rect 445772 229094 445800 231676
rect 446416 229430 446444 231676
rect 446404 229424 446456 229430
rect 446404 229366 446456 229372
rect 443472 229066 443960 229094
rect 444668 229066 444788 229094
rect 444852 229066 445616 229094
rect 445772 229066 446444 229094
rect 443932 217274 443960 229066
rect 444760 217274 444788 229066
rect 445588 217274 445616 229066
rect 446416 217274 446444 229066
rect 447060 227934 447088 231676
rect 447520 231662 447718 231690
rect 447048 227928 447100 227934
rect 447048 227870 447100 227876
rect 447520 224262 447548 231662
rect 447692 230172 447744 230178
rect 447692 230114 447744 230120
rect 447508 224256 447560 224262
rect 447508 224198 447560 224204
rect 447704 219434 447732 230114
rect 448348 229094 448376 231676
rect 448992 229566 449020 231676
rect 449636 229906 449664 231676
rect 449624 229900 449676 229906
rect 449624 229842 449676 229848
rect 448980 229560 449032 229566
rect 448980 229502 449032 229508
rect 448980 229424 449032 229430
rect 448980 229366 449032 229372
rect 448348 229066 448652 229094
rect 448060 224256 448112 224262
rect 448060 224198 448112 224204
rect 447336 219406 447732 219434
rect 447336 217274 447364 219406
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444760 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 441494 217110 441568 217138
rect 441494 216988 441522 217110
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447290 217246 447364 217274
rect 448072 217274 448100 224198
rect 448072 217246 448146 217274
rect 448624 217258 448652 229066
rect 448992 217274 449020 229366
rect 450280 229294 450308 231676
rect 450544 229900 450596 229906
rect 450544 229842 450596 229848
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 229842
rect 450924 229158 450952 231676
rect 451568 230450 451596 231676
rect 452226 231662 452608 231690
rect 451556 230444 451608 230450
rect 451556 230386 451608 230392
rect 451924 229560 451976 229566
rect 451924 229502 451976 229508
rect 451740 229288 451792 229294
rect 451740 229230 451792 229236
rect 450912 229152 450964 229158
rect 450912 229094 450964 229100
rect 450556 229066 450768 229094
rect 450544 227928 450596 227934
rect 450544 227870 450596 227876
rect 447290 216988 447318 217246
rect 448118 216988 448146 217246
rect 448612 217252 448664 217258
rect 448612 217194 448664 217200
rect 448946 217246 449020 217274
rect 450556 217274 450584 227870
rect 450740 218346 450768 229066
rect 451752 219434 451780 229230
rect 451936 229094 451964 229502
rect 451936 229066 452240 229094
rect 451476 219406 451780 219434
rect 450728 218340 450780 218346
rect 450728 218282 450780 218288
rect 451476 217274 451504 219406
rect 449762 217252 449814 217258
rect 448946 216988 448974 217246
rect 450556 217246 450630 217274
rect 449762 217194 449814 217200
rect 449774 216988 449802 217194
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 229066
rect 452580 222154 452608 231662
rect 452856 230246 452884 231676
rect 453304 230444 453356 230450
rect 453304 230386 453356 230392
rect 452844 230240 452896 230246
rect 452844 230182 452896 230188
rect 452752 229152 452804 229158
rect 452752 229094 452804 229100
rect 452764 229066 453068 229094
rect 452568 222148 452620 222154
rect 452568 222090 452620 222096
rect 453040 217274 453068 229066
rect 453316 218074 453344 230386
rect 453500 229974 453528 231676
rect 454144 230110 454172 231676
rect 454316 230240 454368 230246
rect 454316 230182 454368 230188
rect 454132 230104 454184 230110
rect 454132 230046 454184 230052
rect 453488 229968 453540 229974
rect 453488 229910 453540 229916
rect 454328 229094 454356 230182
rect 454788 229094 454816 231676
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455328 230104 455380 230110
rect 455328 230046 455380 230052
rect 454328 229066 454724 229094
rect 454788 229066 454908 229094
rect 453856 218340 453908 218346
rect 453856 218282 453908 218288
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 218282
rect 454696 217274 454724 229066
rect 454880 223582 454908 229066
rect 454868 223576 454920 223582
rect 454868 223518 454920 223524
rect 455340 220794 455368 230046
rect 455788 229968 455840 229974
rect 455788 229910 455840 229916
rect 455604 222148 455656 222154
rect 455604 222090 455656 222096
rect 455328 220788 455380 220794
rect 455328 220730 455380 220736
rect 455616 218074 455644 222090
rect 455800 219434 455828 229910
rect 456076 224534 456104 231676
rect 456064 224528 456116 224534
rect 456064 224470 456116 224476
rect 456720 220930 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 220924 456760 220930
rect 456708 220866 456760 220872
rect 457180 219434 457208 230318
rect 457364 229770 457392 231676
rect 457352 229764 457404 229770
rect 457352 229706 457404 229712
rect 458008 229094 458036 231676
rect 458008 229066 458128 229094
rect 455800 219406 456380 219434
rect 457180 219406 458036 219434
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455604 218068 455656 218074
rect 455604 218010 455656 218016
rect 455432 217274 455460 218010
rect 456352 217274 456380 219406
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 454696 217246 454770 217274
rect 455432 217246 455598 217274
rect 456352 217246 456426 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455570 216988 455598 217246
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458100 218498 458128 229066
rect 458652 226302 458680 231676
rect 459310 231662 459508 231690
rect 458640 226296 458692 226302
rect 458640 226238 458692 226244
rect 458824 220788 458876 220794
rect 458824 220730 458876 220736
rect 458100 218470 458220 218498
rect 458192 218414 458220 218470
rect 458180 218408 458232 218414
rect 458180 218350 458232 218356
rect 458836 217274 458864 220730
rect 459480 220250 459508 231662
rect 459744 224528 459796 224534
rect 459744 224470 459796 224476
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459756 217274 459784 224470
rect 459940 222902 459968 231676
rect 460584 224942 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224936 460624 224942
rect 460572 224878 460624 224884
rect 460480 223576 460532 223582
rect 460480 223518 460532 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 217246 459784 217274
rect 460492 217274 460520 223518
rect 461308 218340 461360 218346
rect 461308 218282 461360 218288
rect 460492 217246 460566 217274
rect 459710 216988 459738 217246
rect 460538 216988 460566 217246
rect 461320 217138 461348 218282
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224806 462544 231676
rect 462964 226296 463016 226302
rect 462964 226238 463016 226244
rect 462504 224800 462556 224806
rect 462504 224742 462556 224748
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 220856 462188 220862
rect 462136 220798 462188 220804
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 220798
rect 462976 217274 463004 226238
rect 463160 225418 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 229764 463936 229770
rect 463884 229706 463936 229712
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 224936 463200 224942
rect 463148 224878 463200 224884
rect 463160 218074 463188 224878
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 229706
rect 465000 219638 465028 231662
rect 465460 229770 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 229764 465500 229770
rect 465448 229706 465500 229712
rect 465736 220794 465764 230318
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220930 466132 231662
rect 467024 229906 467052 231676
rect 467012 229900 467064 229906
rect 467012 229842 467064 229848
rect 467472 229764 467524 229770
rect 467472 229706 467524 229712
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220924 466144 220930
rect 466092 220866 466144 220872
rect 465724 220788 465776 220794
rect 465724 220730 465776 220736
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 461320 217110 461394 217138
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229706
rect 467668 225622 467696 231676
rect 468312 230246 468340 231676
rect 468300 230240 468352 230246
rect 468300 230182 468352 230188
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 468956 221474 468984 231676
rect 469128 230240 469180 230246
rect 469128 230182 469180 230188
rect 468944 221468 468996 221474
rect 468944 221410 468996 221416
rect 469140 220522 469168 230182
rect 469600 229770 469628 231676
rect 469588 229764 469640 229770
rect 469588 229706 469640 229712
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224800 469364 224806
rect 469312 224742 469364 224748
rect 469128 220516 469180 220522
rect 469128 220458 469180 220464
rect 468772 217246 468846 217274
rect 469324 217258 469352 224742
rect 469588 220788 469640 220794
rect 469588 220730 469640 220736
rect 469600 217274 469628 220730
rect 469876 218618 469904 227598
rect 470244 224262 470272 231676
rect 470888 230382 470916 231676
rect 470876 230376 470928 230382
rect 470876 230318 470928 230324
rect 471532 227798 471560 231676
rect 471888 230376 471940 230382
rect 471888 230318 471940 230324
rect 471520 227792 471572 227798
rect 471520 227734 471572 227740
rect 470232 224256 470284 224262
rect 470232 224198 470284 224204
rect 471900 222154 471928 230318
rect 472176 229362 472204 231676
rect 472834 231662 473216 231690
rect 472164 229356 472216 229362
rect 472164 229298 472216 229304
rect 472992 229356 473044 229362
rect 472992 229298 473044 229304
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 471428 220924 471480 220930
rect 471428 220866 471480 220872
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 471440 218074 471468 220866
rect 473004 220386 473032 229298
rect 472992 220380 473044 220386
rect 472992 220322 473044 220328
rect 473188 220250 473216 231662
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474004 229900 474056 229906
rect 474004 229842 474056 229848
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 473176 220244 473228 220250
rect 473176 220186 473228 220192
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471428 218068 471480 218074
rect 471428 218010 471480 218016
rect 472084 217274 472112 219574
rect 472900 218068 472952 218074
rect 472900 218010 472952 218016
rect 472084 217246 472158 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472912 217138 472940 218010
rect 473740 217274 473768 222838
rect 474016 220794 474044 229842
rect 474476 228410 474504 231662
rect 474464 228404 474516 228410
rect 474464 228346 474516 228352
rect 474752 226506 474780 231676
rect 475410 231662 475976 231690
rect 474740 226500 474792 226506
rect 474740 226442 474792 226448
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 474004 220788 474056 220794
rect 474004 220730 474056 220736
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474556 220516 474608 220522
rect 474556 220458 474608 220464
rect 474568 217274 474596 220458
rect 475396 217274 475424 220730
rect 475580 218618 475608 223518
rect 475948 221746 475976 231662
rect 476040 230466 476068 231676
rect 476040 230450 476160 230466
rect 476040 230444 476172 230450
rect 476040 230438 476120 230444
rect 476120 230386 476172 230392
rect 476684 229906 476712 231676
rect 476672 229900 476724 229906
rect 476672 229842 476724 229848
rect 476764 229764 476816 229770
rect 476764 229706 476816 229712
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475936 221740 475988 221746
rect 475936 221682 475988 221688
rect 476212 221468 476264 221474
rect 476212 221410 476264 221416
rect 475568 218612 475620 218618
rect 475568 218554 475620 218560
rect 476224 217274 476252 221410
rect 476592 217274 476620 225558
rect 476776 220794 476804 229706
rect 477328 225622 477356 231676
rect 477986 231662 478368 231690
rect 478630 231662 478828 231690
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478340 220114 478368 231662
rect 478604 230444 478656 230450
rect 478604 230386 478656 230392
rect 478616 227186 478644 230386
rect 478800 229094 478828 231662
rect 479260 229770 479288 231676
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 478800 229066 478920 229094
rect 478892 228818 478920 229066
rect 478880 228812 478932 228818
rect 478880 228754 478932 228760
rect 479524 227792 479576 227798
rect 479524 227734 479576 227740
rect 478604 227180 478656 227186
rect 478604 227122 478656 227128
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478328 220108 478380 220114
rect 478328 220050 478380 220056
rect 478708 217274 478736 220730
rect 479536 217274 479564 227734
rect 479904 222902 479932 231676
rect 480548 224398 480576 231676
rect 480824 231662 481206 231690
rect 480536 224392 480588 224398
rect 480536 224334 480588 224340
rect 480444 224256 480496 224262
rect 480444 224198 480496 224204
rect 479892 222896 479944 222902
rect 479892 222838 479944 222844
rect 480456 217274 480484 224198
rect 480824 221610 480852 231662
rect 481836 229906 481864 231676
rect 482494 231662 482968 231690
rect 481640 229900 481692 229906
rect 481640 229842 481692 229848
rect 481824 229900 481876 229906
rect 481824 229842 481876 229848
rect 481652 226370 481680 229842
rect 482744 226500 482796 226506
rect 482744 226442 482796 226448
rect 481640 226364 481692 226370
rect 481640 226306 481692 226312
rect 482756 222222 482784 226442
rect 482744 222216 482796 222222
rect 482744 222158 482796 222164
rect 480812 221604 480864 221610
rect 480812 221546 480864 221552
rect 481180 220380 481232 220386
rect 481180 220322 481232 220328
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480410 217246 480484 217274
rect 481192 217274 481220 220322
rect 482008 220244 482060 220250
rect 482008 220186 482060 220192
rect 482020 217274 482048 220186
rect 482756 218754 482784 222158
rect 482940 220250 482968 231662
rect 483124 223310 483152 231676
rect 483768 225894 483796 231676
rect 484412 230042 484440 231676
rect 484400 230036 484452 230042
rect 484400 229978 484452 229984
rect 485056 228546 485084 231676
rect 485700 228682 485728 231676
rect 486358 231662 486648 231690
rect 485688 228676 485740 228682
rect 485688 228618 485740 228624
rect 485044 228540 485096 228546
rect 485044 228482 485096 228488
rect 484492 228404 484544 228410
rect 484492 228346 484544 228352
rect 483756 225888 483808 225894
rect 483756 225830 483808 225836
rect 483112 223304 483164 223310
rect 483112 223246 483164 223252
rect 484504 222358 484532 228346
rect 486620 224262 486648 231662
rect 486792 227180 486844 227186
rect 486792 227122 486844 227128
rect 486804 224954 486832 227122
rect 486988 227050 487016 231676
rect 487632 230246 487660 231676
rect 488290 231662 488488 231690
rect 488460 230330 488488 231662
rect 488460 230302 488672 230330
rect 487620 230240 487672 230246
rect 487620 230182 487672 230188
rect 488448 230240 488500 230246
rect 488448 230182 488500 230188
rect 486976 227044 487028 227050
rect 486976 226986 487028 226992
rect 487804 226364 487856 226370
rect 487804 226306 487856 226312
rect 486804 224926 487016 224954
rect 486608 224256 486660 224262
rect 486608 224198 486660 224204
rect 484492 222352 484544 222358
rect 484492 222294 484544 222300
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 482928 220244 482980 220250
rect 482928 220186 482980 220192
rect 482744 218748 482796 218754
rect 482744 218690 482796 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 480410 216988 480438 217246
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483768 217274 483796 221410
rect 483722 217246 483796 217274
rect 484504 217274 484532 222294
rect 486148 221740 486200 221746
rect 486148 221682 486200 221688
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 484504 217246 484578 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485332 217138 485360 218690
rect 486160 217138 486188 221682
rect 486988 220289 487016 224926
rect 486974 220280 487030 220289
rect 486974 220215 487030 220224
rect 486988 217274 487016 220215
rect 487816 218113 487844 226306
rect 488460 220522 488488 230182
rect 488644 223174 488672 230302
rect 488920 225758 488948 231676
rect 489564 227186 489592 231676
rect 489920 229764 489972 229770
rect 489920 229706 489972 229712
rect 489552 227180 489604 227186
rect 489552 227122 489604 227128
rect 488908 225752 488960 225758
rect 488908 225694 488960 225700
rect 488816 225616 488868 225622
rect 488816 225558 488868 225564
rect 488632 223168 488684 223174
rect 488632 223110 488684 223116
rect 488448 220516 488500 220522
rect 488448 220458 488500 220464
rect 487802 218104 487858 218113
rect 487802 218039 487858 218048
rect 487816 217274 487844 218039
rect 488828 217274 488856 225558
rect 489932 222358 489960 229706
rect 490208 228410 490236 231676
rect 490866 231662 491248 231690
rect 491220 229094 491248 231662
rect 491496 230110 491524 231676
rect 491484 230104 491536 230110
rect 491484 230046 491536 230052
rect 492140 229770 492168 231676
rect 492798 231662 493088 231690
rect 492496 230104 492548 230110
rect 492496 230046 492548 230052
rect 492128 229764 492180 229770
rect 492128 229706 492180 229712
rect 491220 229066 491340 229094
rect 490380 228812 490432 228818
rect 490380 228754 490432 228760
rect 490196 228404 490248 228410
rect 490196 228346 490248 228352
rect 489920 222352 489972 222358
rect 489920 222294 489972 222300
rect 489460 220108 489512 220114
rect 489460 220050 489512 220056
rect 486988 217246 487062 217274
rect 487816 217246 487890 217274
rect 485332 217110 485406 217138
rect 486160 217110 486234 217138
rect 485378 216988 485406 217110
rect 486206 216988 486234 217110
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488690 217246 488856 217274
rect 488690 216988 488718 217246
rect 488828 217161 488856 217246
rect 488814 217152 488870 217161
rect 489472 217138 489500 220050
rect 490392 218074 490420 228754
rect 491312 224534 491340 229066
rect 491300 224528 491352 224534
rect 491300 224470 491352 224476
rect 491944 222896 491996 222902
rect 491944 222838 491996 222844
rect 491116 222352 491168 222358
rect 491116 222294 491168 222300
rect 490380 218068 490432 218074
rect 490380 218010 490432 218016
rect 490392 217274 490420 218010
rect 490346 217246 490420 217274
rect 489472 217110 489546 217138
rect 488814 217087 488870 217096
rect 489518 216988 489546 217110
rect 490346 216988 490374 217246
rect 491128 217138 491156 222294
rect 491956 218210 491984 222838
rect 492508 220114 492536 230046
rect 492772 224392 492824 224398
rect 492772 224334 492824 224340
rect 492496 220108 492548 220114
rect 492496 220050 492548 220056
rect 491944 218204 491996 218210
rect 491944 218146 491996 218152
rect 491956 217138 491984 218146
rect 492784 217138 492812 224334
rect 493060 223038 493088 231662
rect 493428 230382 493456 231676
rect 493416 230376 493468 230382
rect 493416 230318 493468 230324
rect 493692 229900 493744 229906
rect 493692 229842 493744 229848
rect 493704 225010 493732 229842
rect 494072 225622 494100 231676
rect 494716 227322 494744 231676
rect 495164 230240 495216 230246
rect 495164 230182 495216 230188
rect 494704 227316 494756 227322
rect 494704 227258 494756 227264
rect 494060 225616 494112 225622
rect 494060 225558 494112 225564
rect 495176 225010 495204 230182
rect 495360 229294 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 229288 495400 229294
rect 495348 229230 495400 229236
rect 496188 229094 496216 231662
rect 497292 230382 497320 231676
rect 497476 231662 497950 231690
rect 496360 230376 496412 230382
rect 496360 230318 496412 230324
rect 497280 230376 497332 230382
rect 497280 230318 497332 230324
rect 496372 229094 496400 230318
rect 496188 229066 496308 229094
rect 496372 229066 496492 229094
rect 493692 225004 493744 225010
rect 493692 224946 493744 224952
rect 494704 225004 494756 225010
rect 494704 224946 494756 224952
rect 495164 225004 495216 225010
rect 495164 224946 495216 224952
rect 493048 223032 493100 223038
rect 493048 222974 493100 222980
rect 492956 221604 493008 221610
rect 492956 221546 493008 221552
rect 492968 219745 492996 221546
rect 492954 219736 493010 219745
rect 492954 219671 493010 219680
rect 493690 219736 493746 219745
rect 493690 219671 493746 219680
rect 493704 217138 493732 219671
rect 494716 218385 494744 224946
rect 495176 222086 495204 224946
rect 496084 223304 496136 223310
rect 496084 223246 496136 223252
rect 495164 222080 495216 222086
rect 495164 222022 495216 222028
rect 495256 220244 495308 220250
rect 495256 220186 495308 220192
rect 494702 218376 494758 218385
rect 494532 218334 494702 218362
rect 494532 217274 494560 218334
rect 494702 218311 494758 218320
rect 495268 217274 495296 220186
rect 491128 217110 491202 217138
rect 491956 217110 492030 217138
rect 492784 217110 492858 217138
rect 491174 216988 491202 217110
rect 492002 216988 492030 217110
rect 492830 216988 492858 217110
rect 493658 217110 493732 217138
rect 494486 217246 494560 217274
rect 495176 217246 495342 217274
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 495176 217161 495204 217246
rect 495162 217152 495218 217161
rect 495162 217087 495218 217096
rect 495314 216988 495342 217246
rect 496096 217138 496124 223246
rect 496280 221746 496308 229066
rect 496268 221740 496320 221746
rect 496268 221682 496320 221688
rect 496464 220386 496492 229066
rect 497280 225888 497332 225894
rect 497280 225830 497332 225836
rect 497292 224954 497320 225830
rect 497016 224926 497320 224954
rect 496452 220380 496504 220386
rect 496452 220322 496504 220328
rect 497016 218346 497044 224926
rect 497476 221610 497504 231662
rect 498108 230376 498160 230382
rect 498108 230318 498160 230324
rect 498120 226030 498148 230318
rect 498580 228682 498608 231676
rect 498292 228676 498344 228682
rect 498292 228618 498344 228624
rect 498568 228676 498620 228682
rect 498568 228618 498620 228624
rect 498108 226024 498160 226030
rect 498108 225966 498160 225972
rect 497740 222080 497792 222086
rect 497740 222022 497792 222028
rect 497464 221604 497516 221610
rect 497464 221546 497516 221552
rect 497004 218340 497056 218346
rect 497004 218282 497056 218288
rect 497016 217274 497044 218282
rect 496970 217246 497044 217274
rect 496096 217110 496170 217138
rect 496142 216988 496170 217110
rect 496970 216988 496998 217246
rect 497752 217138 497780 222022
rect 498304 217258 498332 228618
rect 498660 228540 498712 228546
rect 498660 228482 498712 228488
rect 498672 217274 498700 228482
rect 499224 224398 499252 231676
rect 499868 228818 499896 231676
rect 500526 231662 500816 231690
rect 500224 229288 500276 229294
rect 500224 229230 500276 229236
rect 499856 228812 499908 228818
rect 499856 228754 499908 228760
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 500040 224256 500092 224262
rect 500040 224198 500092 224204
rect 500052 218482 500080 224198
rect 500236 220658 500264 229230
rect 500788 222902 500816 231662
rect 500960 227044 501012 227050
rect 500960 226986 501012 226992
rect 500972 224954 501000 226986
rect 501156 225894 501184 231676
rect 501340 231662 501814 231690
rect 501144 225888 501196 225894
rect 501144 225830 501196 225836
rect 500972 224926 501184 224954
rect 500776 222896 500828 222902
rect 500776 222838 500828 222844
rect 500224 220652 500276 220658
rect 500224 220594 500276 220600
rect 501156 219502 501184 224926
rect 501340 220250 501368 231662
rect 502444 228546 502472 231676
rect 503102 231662 503392 231690
rect 502432 228540 502484 228546
rect 502432 228482 502484 228488
rect 503364 223310 503392 231662
rect 503732 229158 503760 231676
rect 503720 229152 503772 229158
rect 503720 229094 503772 229100
rect 504180 227180 504232 227186
rect 504180 227122 504232 227128
rect 503628 225752 503680 225758
rect 503628 225694 503680 225700
rect 503352 223304 503404 223310
rect 503352 223246 503404 223252
rect 502708 223168 502760 223174
rect 502708 223110 502760 223116
rect 501880 220516 501932 220522
rect 501880 220458 501932 220464
rect 501328 220244 501380 220250
rect 501328 220186 501380 220192
rect 501144 219496 501196 219502
rect 501144 219438 501196 219444
rect 500040 218476 500092 218482
rect 500040 218418 500092 218424
rect 498292 217252 498344 217258
rect 498292 217194 498344 217200
rect 498626 217246 498700 217274
rect 500052 217274 500080 218418
rect 500960 218204 501012 218210
rect 500960 218146 501012 218152
rect 500972 217297 501000 218146
rect 500958 217288 501014 217297
rect 499442 217252 499494 217258
rect 497752 217110 497826 217138
rect 498626 217122 498654 217246
rect 500052 217246 500310 217274
rect 499442 217194 499494 217200
rect 497798 216988 497826 217110
rect 498614 217116 498666 217122
rect 498614 217058 498666 217064
rect 498626 216988 498654 217058
rect 499454 216988 499482 217194
rect 500282 216988 500310 217246
rect 501156 217274 501184 219438
rect 500958 217223 501014 217232
rect 501110 217246 501184 217274
rect 501110 216988 501138 217246
rect 501892 217138 501920 220458
rect 502720 218618 502748 223110
rect 503640 219638 503668 225694
rect 504192 224954 504220 227122
rect 504376 224954 504404 231676
rect 505020 227050 505048 231676
rect 505664 229430 505692 231676
rect 506216 231662 506322 231690
rect 505652 229424 505704 229430
rect 505652 229366 505704 229372
rect 505192 228404 505244 228410
rect 505192 228346 505244 228352
rect 505008 227044 505060 227050
rect 505008 226986 505060 226992
rect 504192 224926 504312 224954
rect 504376 224926 504496 224954
rect 503628 219632 503680 219638
rect 503628 219574 503680 219580
rect 502708 218612 502760 218618
rect 502708 218554 502760 218560
rect 502720 217138 502748 218554
rect 503640 217274 503668 219574
rect 503594 217246 503668 217274
rect 504284 217274 504312 224926
rect 504468 224262 504496 224926
rect 504456 224256 504508 224262
rect 504456 224198 504508 224204
rect 505204 223650 505232 228346
rect 506216 227186 506244 231662
rect 506388 229900 506440 229906
rect 506388 229842 506440 229848
rect 506400 228954 506428 229842
rect 506388 228948 506440 228954
rect 506388 228890 506440 228896
rect 506204 227180 506256 227186
rect 506204 227122 506256 227128
rect 506952 224806 506980 231676
rect 507596 229906 507624 231676
rect 507584 229900 507636 229906
rect 507584 229842 507636 229848
rect 507124 229764 507176 229770
rect 507124 229706 507176 229712
rect 506940 224800 506992 224806
rect 506940 224742 506992 224748
rect 506020 224528 506072 224534
rect 506020 224470 506072 224476
rect 505192 223644 505244 223650
rect 505192 223586 505244 223592
rect 505204 217274 505232 223586
rect 506032 217274 506060 224470
rect 506848 220108 506900 220114
rect 506848 220050 506900 220056
rect 506860 217274 506888 220050
rect 507136 218210 507164 229706
rect 508240 223174 508268 231676
rect 508884 225758 508912 231676
rect 509528 229702 509556 231676
rect 509516 229696 509568 229702
rect 509516 229638 509568 229644
rect 509884 229152 509936 229158
rect 509884 229094 509936 229100
rect 508872 225752 508924 225758
rect 508872 225694 508924 225700
rect 509516 225616 509568 225622
rect 509516 225558 509568 225564
rect 509528 223786 509556 225558
rect 509516 223780 509568 223786
rect 509516 223722 509568 223728
rect 508228 223168 508280 223174
rect 508228 223110 508280 223116
rect 508596 223032 508648 223038
rect 508596 222974 508648 222980
rect 507124 218204 507176 218210
rect 507124 218146 507176 218152
rect 507676 218204 507728 218210
rect 507676 218146 507728 218152
rect 504284 217246 504450 217274
rect 505204 217246 505278 217274
rect 506032 217246 506106 217274
rect 506860 217246 506934 217274
rect 501892 217110 501966 217138
rect 502720 217110 502794 217138
rect 501938 216988 501966 217110
rect 502766 216988 502794 217110
rect 503594 216988 503622 217246
rect 504422 216988 504450 217246
rect 505250 216988 505278 217246
rect 506078 217190 506106 217246
rect 506066 217184 506118 217190
rect 506066 217126 506118 217132
rect 506078 216988 506106 217126
rect 506906 216988 506934 217246
rect 507688 217138 507716 218146
rect 508608 217326 508636 222974
rect 509896 221882 509924 229094
rect 510172 225622 510200 231676
rect 510816 230382 510844 231676
rect 510804 230376 510856 230382
rect 510804 230318 510856 230324
rect 511460 230246 511488 231676
rect 511908 230376 511960 230382
rect 511908 230318 511960 230324
rect 511448 230240 511500 230246
rect 511448 230182 511500 230188
rect 510620 229424 510672 229430
rect 510620 229366 510672 229372
rect 510632 227322 510660 229366
rect 511920 229094 511948 230318
rect 511828 229066 511948 229094
rect 510620 227316 510672 227322
rect 510620 227258 510672 227264
rect 510988 226908 511040 226914
rect 510988 226850 511040 226856
rect 510160 225616 510212 225622
rect 510160 225558 510212 225564
rect 510160 223780 510212 223786
rect 510160 223722 510212 223728
rect 509884 221876 509936 221882
rect 509884 221818 509936 221824
rect 509332 220380 509384 220386
rect 509332 220322 509384 220328
rect 508596 217320 508648 217326
rect 508596 217262 508648 217268
rect 509344 217274 509372 220322
rect 510172 217274 510200 223722
rect 511000 217569 511028 226850
rect 511828 220794 511856 229066
rect 512104 228410 512132 231676
rect 512762 231662 513144 231690
rect 512736 228948 512788 228954
rect 512736 228890 512788 228896
rect 512092 228404 512144 228410
rect 512092 228346 512144 228352
rect 511816 220788 511868 220794
rect 511816 220730 511868 220736
rect 511816 220652 511868 220658
rect 511816 220594 511868 220600
rect 510986 217560 511042 217569
rect 510986 217495 511042 217504
rect 508608 217138 508636 217262
rect 509344 217246 509418 217274
rect 510172 217246 510246 217274
rect 507688 217110 507762 217138
rect 507734 216988 507762 217110
rect 508562 217110 508636 217138
rect 508562 216988 508590 217110
rect 509390 216988 509418 217246
rect 510218 216988 510246 217246
rect 511000 217138 511028 217495
rect 511828 217274 511856 220594
rect 512748 218890 512776 228890
rect 513116 220114 513144 231662
rect 513392 229294 513420 231676
rect 513380 229288 513432 229294
rect 513380 229230 513432 229236
rect 514036 227458 514064 231676
rect 514024 227452 514076 227458
rect 514024 227394 514076 227400
rect 514300 226024 514352 226030
rect 514300 225966 514352 225972
rect 513564 221740 513616 221746
rect 513564 221682 513616 221688
rect 513576 220969 513604 221682
rect 513562 220960 513618 220969
rect 513562 220895 513618 220904
rect 513104 220108 513156 220114
rect 513104 220050 513156 220056
rect 512736 218884 512788 218890
rect 512736 218826 512788 218832
rect 512748 217274 512776 218826
rect 513576 217274 513604 220895
rect 513840 218748 513892 218754
rect 513840 218690 513892 218696
rect 513852 218210 513880 218690
rect 514024 218612 514076 218618
rect 514024 218554 514076 218560
rect 514036 218210 514064 218554
rect 513840 218204 513892 218210
rect 513840 218146 513892 218152
rect 514024 218204 514076 218210
rect 514024 218146 514076 218152
rect 511828 217246 511902 217274
rect 511000 217110 511074 217138
rect 511046 216988 511074 217110
rect 511874 216988 511902 217246
rect 512702 217246 512776 217274
rect 513530 217246 513604 217274
rect 514312 217274 514340 225966
rect 514680 223310 514708 231676
rect 515324 229158 515352 231676
rect 515496 229696 515548 229702
rect 515496 229638 515548 229644
rect 515312 229152 515364 229158
rect 515312 229094 515364 229100
rect 514668 223304 514720 223310
rect 514668 223246 514720 223252
rect 515508 222086 515536 229638
rect 515772 228676 515824 228682
rect 515772 228618 515824 228624
rect 515496 222080 515548 222086
rect 515496 222022 515548 222028
rect 515128 221604 515180 221610
rect 515128 221546 515180 221552
rect 515140 220017 515168 221546
rect 515784 221241 515812 228618
rect 515968 224534 515996 231676
rect 516612 226030 516640 231676
rect 517256 230042 517284 231676
rect 517520 230240 517572 230246
rect 517520 230182 517572 230188
rect 517244 230036 517296 230042
rect 517244 229978 517296 229984
rect 516784 229900 516836 229906
rect 516784 229842 516836 229848
rect 516796 229094 516824 229842
rect 516796 229066 517008 229094
rect 516600 226024 516652 226030
rect 516600 225966 516652 225972
rect 515956 224528 516008 224534
rect 515956 224470 516008 224476
rect 516784 224392 516836 224398
rect 516784 224334 516836 224340
rect 515770 221232 515826 221241
rect 515770 221167 515826 221176
rect 515126 220008 515182 220017
rect 515126 219943 515182 219952
rect 515140 217274 515168 219943
rect 515784 219434 515812 221167
rect 515784 219406 516088 219434
rect 516060 217274 516088 219406
rect 514312 217246 514386 217274
rect 515140 217246 515214 217274
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515186 216988 515214 217246
rect 516014 217246 516088 217274
rect 516796 217274 516824 224334
rect 516980 220386 517008 229066
rect 517532 223446 517560 230182
rect 517900 228682 517928 231676
rect 518544 228818 518572 231676
rect 519188 229906 519216 231676
rect 519176 229900 519228 229906
rect 519176 229842 519228 229848
rect 519084 229288 519136 229294
rect 519084 229230 519136 229236
rect 518164 228812 518216 228818
rect 518164 228754 518216 228760
rect 518532 228812 518584 228818
rect 518532 228754 518584 228760
rect 517888 228676 517940 228682
rect 517888 228618 517940 228624
rect 517520 223440 517572 223446
rect 517520 223382 517572 223388
rect 517520 222896 517572 222902
rect 517520 222838 517572 222844
rect 517532 220862 517560 222838
rect 517520 220856 517572 220862
rect 517520 220798 517572 220804
rect 516968 220380 517020 220386
rect 516968 220322 517020 220328
rect 518176 218754 518204 228754
rect 519096 224126 519124 229230
rect 519268 225888 519320 225894
rect 519268 225830 519320 225836
rect 519084 224120 519136 224126
rect 519084 224062 519136 224068
rect 518532 220856 518584 220862
rect 518532 220798 518584 220804
rect 517704 218748 517756 218754
rect 517704 218690 517756 218696
rect 518164 218748 518216 218754
rect 518164 218690 518216 218696
rect 517716 217274 517744 218690
rect 518544 217274 518572 220798
rect 516796 217246 516870 217274
rect 516014 216988 516042 217246
rect 516842 216988 516870 217246
rect 517670 217246 517744 217274
rect 518498 217246 518572 217274
rect 519280 217274 519308 225830
rect 519832 222902 519860 231676
rect 520476 224670 520504 231676
rect 521120 230382 521148 231676
rect 521108 230376 521160 230382
rect 521108 230318 521160 230324
rect 520924 229152 520976 229158
rect 520924 229094 520976 229100
rect 520464 224664 520516 224670
rect 520464 224606 520516 224612
rect 519820 222896 519872 222902
rect 519820 222838 519872 222844
rect 520936 220658 520964 229094
rect 521108 228540 521160 228546
rect 521108 228482 521160 228488
rect 521120 220998 521148 228482
rect 521764 225894 521792 231676
rect 522422 231662 522896 231690
rect 521752 225888 521804 225894
rect 521752 225830 521804 225836
rect 521752 223168 521804 223174
rect 521752 223110 521804 223116
rect 521108 220992 521160 220998
rect 521108 220934 521160 220940
rect 520924 220652 520976 220658
rect 520924 220594 520976 220600
rect 520188 220244 520240 220250
rect 520188 220186 520240 220192
rect 520200 219473 520228 220186
rect 520186 219464 520242 219473
rect 521120 219434 521148 220934
rect 520186 219399 520242 219408
rect 521028 219406 521148 219434
rect 520004 218748 520056 218754
rect 520004 218690 520056 218696
rect 520016 217569 520044 218690
rect 520002 217560 520058 217569
rect 520002 217495 520058 217504
rect 520200 217274 520228 219399
rect 521028 217274 521056 219406
rect 519280 217246 519354 217274
rect 517670 216988 517698 217246
rect 518498 216988 518526 217246
rect 519326 216988 519354 217246
rect 520154 217246 520228 217274
rect 520982 217246 521056 217274
rect 521764 217274 521792 223110
rect 522580 221876 522632 221882
rect 522580 221818 522632 221824
rect 522592 221513 522620 221818
rect 522868 221610 522896 231662
rect 523052 229770 523080 231676
rect 523040 229764 523092 229770
rect 523040 229706 523092 229712
rect 523696 227050 523724 231676
rect 524248 231662 524354 231690
rect 523040 227044 523092 227050
rect 523040 226986 523092 226992
rect 523684 227044 523736 227050
rect 523684 226986 523736 226992
rect 522856 221604 522908 221610
rect 522856 221546 522908 221552
rect 522578 221504 522634 221513
rect 522578 221439 522634 221448
rect 522592 217274 522620 221439
rect 523052 217870 523080 226986
rect 523500 224256 523552 224262
rect 523500 224198 523552 224204
rect 523512 221134 523540 224198
rect 524248 221746 524276 231662
rect 524604 230036 524656 230042
rect 524604 229978 524656 229984
rect 524616 227594 524644 229978
rect 524984 229158 525012 231676
rect 524972 229152 525024 229158
rect 524972 229094 525024 229100
rect 524604 227588 524656 227594
rect 524604 227530 524656 227536
rect 524420 227316 524472 227322
rect 524420 227258 524472 227264
rect 524432 223922 524460 227258
rect 525628 224398 525656 231676
rect 526272 227322 526300 231676
rect 526444 230376 526496 230382
rect 526444 230318 526496 230324
rect 526456 228954 526484 230318
rect 526916 229634 526944 231676
rect 526904 229628 526956 229634
rect 526904 229570 526956 229576
rect 526444 228948 526496 228954
rect 526444 228890 526496 228896
rect 527560 228546 527588 231676
rect 528218 231662 528416 231690
rect 527548 228540 527600 228546
rect 527548 228482 527600 228488
rect 526260 227316 526312 227322
rect 526260 227258 526312 227264
rect 525984 227180 526036 227186
rect 525984 227122 526036 227128
rect 525616 224392 525668 224398
rect 525616 224334 525668 224340
rect 524420 223916 524472 223922
rect 524420 223858 524472 223864
rect 525064 223916 525116 223922
rect 525064 223858 525116 223864
rect 524236 221740 524288 221746
rect 524236 221682 524288 221688
rect 523500 221128 523552 221134
rect 523500 221070 523552 221076
rect 523040 217864 523092 217870
rect 523040 217806 523092 217812
rect 523512 217274 523540 221070
rect 524236 217864 524288 217870
rect 524236 217806 524288 217812
rect 521764 217246 521838 217274
rect 522592 217246 522666 217274
rect 520154 216988 520182 217246
rect 520982 216988 521010 217246
rect 521810 216988 521838 217246
rect 522638 216988 522666 217246
rect 523466 217246 523540 217274
rect 523466 216988 523494 217246
rect 524248 217138 524276 217806
rect 525076 217274 525104 223858
rect 525996 221338 526024 227122
rect 526720 224800 526772 224806
rect 526720 224742 526772 224748
rect 525984 221332 526036 221338
rect 525984 221274 526036 221280
rect 525996 217274 526024 221274
rect 525076 217246 525150 217274
rect 524248 217110 524322 217138
rect 524294 216988 524322 217110
rect 525122 216988 525150 217246
rect 525950 217246 526024 217274
rect 526732 217274 526760 224742
rect 527824 223032 527876 223038
rect 527824 222974 527876 222980
rect 527548 220380 527600 220386
rect 527548 220322 527600 220328
rect 527560 219774 527588 220322
rect 527548 219768 527600 219774
rect 527548 219710 527600 219716
rect 527560 217274 527588 219710
rect 527836 217462 527864 222974
rect 528388 220250 528416 231662
rect 528848 230042 528876 231676
rect 528836 230036 528888 230042
rect 528836 229978 528888 229984
rect 528560 229900 528612 229906
rect 528560 229842 528612 229848
rect 528572 226166 528600 229842
rect 528560 226160 528612 226166
rect 528560 226102 528612 226108
rect 529204 225752 529256 225758
rect 529204 225694 529256 225700
rect 528376 220244 528428 220250
rect 528376 220186 528428 220192
rect 527824 217456 527876 217462
rect 527824 217398 527876 217404
rect 528468 217456 528520 217462
rect 528468 217398 528520 217404
rect 526732 217246 526806 217274
rect 527560 217246 527634 217274
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527606 216988 527634 217246
rect 528480 217138 528508 217398
rect 529216 217274 529244 225694
rect 529492 223038 529520 231676
rect 530136 230382 530164 231676
rect 530124 230376 530176 230382
rect 530124 230318 530176 230324
rect 530780 230246 530808 231676
rect 531136 230376 531188 230382
rect 531136 230318 531188 230324
rect 530768 230240 530820 230246
rect 530768 230182 530820 230188
rect 529940 229152 529992 229158
rect 529940 229094 529992 229100
rect 529952 224806 529980 229094
rect 530952 225616 531004 225622
rect 530952 225558 531004 225564
rect 529940 224800 529992 224806
rect 529940 224742 529992 224748
rect 529480 223032 529532 223038
rect 529480 222974 529532 222980
rect 529848 222624 529900 222630
rect 529848 222566 529900 222572
rect 529860 222086 529888 222566
rect 529848 222080 529900 222086
rect 529848 222022 529900 222028
rect 529860 221354 529888 222022
rect 529860 221326 530072 221354
rect 530044 217274 530072 221326
rect 530964 217598 530992 225558
rect 531148 220386 531176 230318
rect 531424 225622 531452 231676
rect 531412 225616 531464 225622
rect 531412 225558 531464 225564
rect 531504 223440 531556 223446
rect 531504 223382 531556 223388
rect 531136 220380 531188 220386
rect 531136 220322 531188 220328
rect 530952 217592 531004 217598
rect 531516 217569 531544 223382
rect 532068 223174 532096 231676
rect 532712 230178 532740 231676
rect 532700 230172 532752 230178
rect 532700 230114 532752 230120
rect 532976 228404 533028 228410
rect 532976 228346 533028 228352
rect 532056 223168 532108 223174
rect 532056 223110 532108 223116
rect 531688 220516 531740 220522
rect 531688 220458 531740 220464
rect 530952 217534 531004 217540
rect 531502 217560 531558 217569
rect 529216 217246 529290 217274
rect 530044 217246 530118 217274
rect 528434 217110 528508 217138
rect 528434 216988 528462 217110
rect 529262 216988 529290 217246
rect 530090 216988 530118 217246
rect 530964 217138 530992 217534
rect 531502 217495 531558 217504
rect 531700 217274 531728 220458
rect 532988 219434 533016 228346
rect 533356 227186 533384 231676
rect 533528 230308 533580 230314
rect 533528 230250 533580 230256
rect 533540 230042 533568 230250
rect 533528 230036 533580 230042
rect 533528 229978 533580 229984
rect 533344 227180 533396 227186
rect 533344 227122 533396 227128
rect 534000 222086 534028 231676
rect 534644 230042 534672 231676
rect 534632 230036 534684 230042
rect 534632 229978 534684 229984
rect 534816 229764 534868 229770
rect 534816 229706 534868 229712
rect 534828 223446 534856 229706
rect 535288 224262 535316 231676
rect 535736 227452 535788 227458
rect 535736 227394 535788 227400
rect 535276 224256 535328 224262
rect 535276 224198 535328 224204
rect 535000 224120 535052 224126
rect 535000 224062 535052 224068
rect 534816 223440 534868 223446
rect 534816 223382 534868 223388
rect 533988 222080 534040 222086
rect 533988 222022 534040 222028
rect 533620 221604 533672 221610
rect 533620 221546 533672 221552
rect 533632 221490 533660 221546
rect 533172 221462 533660 221490
rect 533172 221338 533200 221462
rect 533160 221332 533212 221338
rect 533160 221274 533212 221280
rect 534172 220108 534224 220114
rect 534172 220050 534224 220056
rect 532988 219406 533476 219434
rect 533448 217734 533476 219406
rect 533436 217728 533488 217734
rect 533436 217670 533488 217676
rect 532514 217560 532570 217569
rect 532514 217495 532570 217504
rect 531700 217246 531774 217274
rect 530918 217110 530992 217138
rect 530918 216988 530946 217110
rect 531746 216988 531774 217246
rect 532528 217138 532556 217495
rect 533448 217138 533476 217670
rect 534184 217274 534212 220050
rect 535012 217274 535040 224062
rect 535460 223304 535512 223310
rect 535460 223246 535512 223252
rect 535472 217870 535500 223246
rect 535748 220522 535776 227394
rect 535932 225758 535960 231676
rect 536576 229906 536604 231676
rect 536564 229900 536616 229906
rect 536564 229842 536616 229848
rect 536104 229628 536156 229634
rect 536104 229570 536156 229576
rect 535920 225752 535972 225758
rect 535920 225694 535972 225700
rect 536116 221950 536144 229570
rect 537220 228410 537248 231676
rect 537878 231662 538168 231690
rect 537208 228404 537260 228410
rect 537208 228346 537260 228352
rect 536104 221944 536156 221950
rect 536104 221886 536156 221892
rect 537484 220652 537536 220658
rect 537484 220594 537536 220600
rect 535736 220516 535788 220522
rect 535736 220458 535788 220464
rect 535748 219434 535776 220458
rect 535748 219406 535960 219434
rect 535460 217864 535512 217870
rect 535460 217806 535512 217812
rect 535932 217274 535960 219406
rect 537496 219026 537524 220594
rect 538140 220114 538168 231662
rect 538312 230308 538364 230314
rect 538312 230250 538364 230256
rect 538324 227458 538352 230250
rect 538508 229770 538536 231676
rect 538784 231662 539166 231690
rect 538496 229764 538548 229770
rect 538496 229706 538548 229712
rect 538784 229094 538812 231662
rect 539600 230444 539652 230450
rect 539600 230386 539652 230392
rect 538508 229066 538812 229094
rect 538312 227452 538364 227458
rect 538312 227394 538364 227400
rect 538508 221354 538536 229066
rect 539612 228682 539640 230386
rect 547144 230172 547196 230178
rect 547144 230114 547196 230120
rect 544292 228948 544344 228954
rect 544292 228890 544344 228896
rect 541624 228812 541676 228818
rect 541624 228754 541676 228760
rect 539416 228676 539468 228682
rect 539416 228618 539468 228624
rect 539600 228676 539652 228682
rect 539600 228618 539652 228624
rect 539428 228274 539456 228618
rect 539416 228268 539468 228274
rect 539416 228210 539468 228216
rect 540796 228268 540848 228274
rect 540796 228210 540848 228216
rect 539968 227588 540020 227594
rect 539968 227530 540020 227536
rect 538680 226024 538732 226030
rect 538680 225966 538732 225972
rect 538324 221338 538536 221354
rect 538312 221332 538536 221338
rect 538364 221326 538536 221332
rect 538312 221274 538364 221280
rect 538496 221264 538548 221270
rect 538496 221206 538548 221212
rect 538508 220726 538536 221206
rect 538496 220720 538548 220726
rect 538496 220662 538548 220668
rect 538692 220538 538720 225966
rect 539980 224534 540008 227530
rect 538864 224528 538916 224534
rect 538864 224470 538916 224476
rect 539968 224528 540020 224534
rect 539968 224470 540020 224476
rect 538876 220726 538904 224470
rect 538864 220720 538916 220726
rect 538864 220662 538916 220668
rect 538324 220510 538720 220538
rect 538128 220108 538180 220114
rect 538128 220050 538180 220056
rect 538324 219434 538352 220510
rect 538876 219434 538904 220662
rect 538232 219406 538352 219434
rect 538416 219406 538904 219434
rect 537484 219020 537536 219026
rect 537484 218962 537536 218968
rect 536656 217864 536708 217870
rect 536656 217806 536708 217812
rect 534184 217246 534258 217274
rect 535012 217246 535086 217274
rect 532528 217110 532602 217138
rect 532574 216988 532602 217110
rect 533402 217110 533476 217138
rect 533402 216988 533430 217110
rect 534230 216988 534258 217246
rect 535058 216988 535086 217246
rect 535886 217246 535960 217274
rect 535886 216988 535914 217246
rect 536668 217138 536696 217806
rect 537496 217274 537524 218962
rect 538232 217598 538260 219406
rect 538220 217592 538272 217598
rect 538220 217534 538272 217540
rect 538416 217274 538444 219406
rect 539140 217592 539192 217598
rect 539140 217534 539192 217540
rect 537496 217246 537570 217274
rect 536668 217110 536742 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217246
rect 538370 217246 538444 217274
rect 538370 216988 538398 217246
rect 539152 217138 539180 217534
rect 539980 217274 540008 224470
rect 540808 219774 540836 228210
rect 540796 219768 540848 219774
rect 540796 219710 540848 219716
rect 540808 217274 540836 219710
rect 541636 217274 541664 228754
rect 542636 226160 542688 226166
rect 542636 226102 542688 226108
rect 542452 224528 542504 224534
rect 542450 224496 542452 224505
rect 542504 224496 542506 224505
rect 542450 224431 542506 224440
rect 542648 219434 542676 226102
rect 544304 224670 544332 228890
rect 545764 225888 545816 225894
rect 545764 225830 545816 225836
rect 544108 224664 544160 224670
rect 544108 224606 544160 224612
rect 544292 224664 544344 224670
rect 544292 224606 544344 224612
rect 545028 224664 545080 224670
rect 545028 224606 545080 224612
rect 542820 224528 542872 224534
rect 542820 224470 542872 224476
rect 543186 224496 543242 224505
rect 542832 223786 542860 224470
rect 543186 224431 543242 224440
rect 543200 224058 543228 224431
rect 543004 224052 543056 224058
rect 543004 223994 543056 224000
rect 543188 224052 543240 224058
rect 543188 223994 543240 224000
rect 543016 223786 543044 223994
rect 542820 223780 542872 223786
rect 542820 223722 542872 223728
rect 543004 223780 543056 223786
rect 543004 223722 543056 223728
rect 543372 222896 543424 222902
rect 543372 222838 543424 222844
rect 542648 219406 543044 219434
rect 543016 219162 543044 219406
rect 542544 219156 542596 219162
rect 542544 219098 542596 219104
rect 543004 219156 543056 219162
rect 543004 219098 543056 219104
rect 539980 217246 540054 217274
rect 540808 217246 540882 217274
rect 541636 217246 541710 217274
rect 539152 217110 539226 217138
rect 539198 216988 539226 217110
rect 540026 216988 540054 217246
rect 540854 216988 540882 217246
rect 541682 216988 541710 217246
rect 542556 217138 542584 219098
rect 543188 219020 543240 219026
rect 543188 218962 543240 218968
rect 543200 218618 543228 218962
rect 543188 218612 543240 218618
rect 543188 218554 543240 218560
rect 543384 217598 543412 222838
rect 543832 222760 543884 222766
rect 543832 222702 543884 222708
rect 543844 222034 543872 222702
rect 543706 222006 543872 222034
rect 543706 221950 543734 222006
rect 543694 221944 543746 221950
rect 543694 221886 543746 221892
rect 543372 217592 543424 217598
rect 543372 217534 543424 217540
rect 543384 217138 543412 217534
rect 542510 217110 542584 217138
rect 543338 217110 543412 217138
rect 544120 217138 544148 224606
rect 544292 221740 544344 221746
rect 544292 221682 544344 221688
rect 544304 220726 544332 221682
rect 544292 220720 544344 220726
rect 544292 220662 544344 220668
rect 545040 217138 545068 224606
rect 545776 221785 545804 225830
rect 547156 221950 547184 230114
rect 549260 230036 549312 230042
rect 549260 229978 549312 229984
rect 548708 227044 548760 227050
rect 548708 226986 548760 226992
rect 548720 224954 548748 226986
rect 548444 224926 548748 224954
rect 548064 224800 548116 224806
rect 548062 224768 548064 224777
rect 548248 224800 548300 224806
rect 548116 224768 548118 224777
rect 548248 224742 548300 224748
rect 548062 224703 548118 224712
rect 548260 224398 548288 224742
rect 548248 224392 548300 224398
rect 548248 224334 548300 224340
rect 547420 223440 547472 223446
rect 547420 223382 547472 223388
rect 547144 221944 547196 221950
rect 547144 221886 547196 221892
rect 546960 221876 547012 221882
rect 546960 221818 547012 221824
rect 545762 221776 545818 221785
rect 545762 221711 545818 221720
rect 545776 217274 545804 221711
rect 546972 221474 547000 221818
rect 546592 221468 546644 221474
rect 546592 221410 546644 221416
rect 546960 221468 547012 221474
rect 546960 221410 547012 221416
rect 545776 217246 545850 217274
rect 544120 217110 544194 217138
rect 542510 216988 542538 217110
rect 543338 216988 543366 217110
rect 544166 216988 544194 217110
rect 544994 217110 545068 217138
rect 544994 216988 545022 217110
rect 545822 216988 545850 217246
rect 546604 217138 546632 221410
rect 547432 218793 547460 223382
rect 548444 219722 548472 224926
rect 549272 224806 549300 229978
rect 553216 228540 553268 228546
rect 553216 228482 553268 228488
rect 551560 227316 551612 227322
rect 551560 227258 551612 227264
rect 549260 224800 549312 224806
rect 549260 224742 549312 224748
rect 549994 224768 550050 224777
rect 549994 224703 550050 224712
rect 550454 224768 550510 224777
rect 550510 224726 550818 224754
rect 550454 224703 550510 224712
rect 549258 221776 549314 221785
rect 549258 221711 549314 221720
rect 549272 221474 549300 221711
rect 549076 221468 549128 221474
rect 549076 221410 549128 221416
rect 549260 221468 549312 221474
rect 549260 221410 549312 221416
rect 548708 220244 548760 220250
rect 548708 220186 548760 220192
rect 548720 219910 548748 220186
rect 548708 219904 548760 219910
rect 548708 219846 548760 219852
rect 548892 219904 548944 219910
rect 548892 219846 548944 219852
rect 548904 219722 548932 219846
rect 548444 219694 548932 219722
rect 548248 219292 548300 219298
rect 548248 219234 548300 219240
rect 548260 218890 548288 219234
rect 548248 218884 548300 218890
rect 548248 218826 548300 218832
rect 547418 218784 547474 218793
rect 547418 218719 547474 218728
rect 547432 217138 547460 218719
rect 548444 217274 548472 219694
rect 548800 219156 548852 219162
rect 548800 219098 548852 219104
rect 548812 218890 548840 219098
rect 548800 218884 548852 218890
rect 548800 218826 548852 218832
rect 548614 218784 548670 218793
rect 548614 218719 548616 218728
rect 548668 218719 548670 218728
rect 548616 218690 548668 218696
rect 548306 217246 548472 217274
rect 546604 217110 546678 217138
rect 547432 217110 547506 217138
rect 546650 216988 546678 217110
rect 547478 216988 547506 217110
rect 548306 216988 548334 217246
rect 549088 217138 549116 221410
rect 550008 217138 550036 224703
rect 550790 224670 550818 224726
rect 550640 224664 550692 224670
rect 550640 224606 550692 224612
rect 550778 224664 550830 224670
rect 550778 224606 550830 224612
rect 550652 220658 550680 224606
rect 550640 220652 550692 220658
rect 550640 220594 550692 220600
rect 550652 217274 550680 220594
rect 551572 217274 551600 227258
rect 553228 224954 553256 228482
rect 553228 224926 553348 224954
rect 552388 222760 552440 222766
rect 552388 222702 552440 222708
rect 550652 217246 550818 217274
rect 551572 217246 551646 217274
rect 549088 217110 549162 217138
rect 549134 216988 549162 217110
rect 549962 217110 550036 217138
rect 549962 216988 549990 217110
rect 550790 216988 550818 217246
rect 551618 216988 551646 217246
rect 552400 217138 552428 222702
rect 553320 222329 553348 224926
rect 554056 222902 554084 249047
rect 555424 244316 555476 244322
rect 555424 244258 555476 244264
rect 554502 240408 554558 240417
rect 554502 240343 554558 240352
rect 554516 240174 554544 240343
rect 554504 240168 554556 240174
rect 554504 240110 554556 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 555436 227050 555464 244258
rect 556816 228546 556844 251194
rect 557172 228676 557224 228682
rect 557172 228618 557224 228624
rect 556804 228540 556856 228546
rect 556804 228482 556856 228488
rect 556068 227452 556120 227458
rect 556068 227394 556120 227400
rect 555424 227044 555476 227050
rect 555424 226986 555476 226992
rect 556080 224505 556108 227394
rect 554870 224496 554926 224505
rect 554870 224431 554926 224440
rect 556066 224496 556122 224505
rect 556066 224431 556122 224440
rect 554044 222896 554096 222902
rect 554044 222838 554096 222844
rect 553306 222320 553362 222329
rect 553306 222255 553362 222264
rect 553320 217274 553348 222255
rect 554228 220652 554280 220658
rect 554228 220594 554280 220600
rect 554240 220386 554268 220594
rect 554044 220380 554096 220386
rect 554044 220322 554096 220328
rect 554228 220380 554280 220386
rect 554228 220322 554280 220328
rect 553274 217246 553348 217274
rect 554056 217274 554084 220322
rect 554884 217274 554912 224431
rect 555700 223032 555752 223038
rect 555700 222974 555752 222980
rect 555712 220658 555740 222974
rect 556988 221944 557040 221950
rect 556986 221912 556988 221921
rect 557040 221912 557042 221921
rect 556986 221847 557042 221856
rect 555700 220652 555752 220658
rect 555700 220594 555752 220600
rect 555712 217274 555740 220594
rect 556528 220516 556580 220522
rect 556528 220458 556580 220464
rect 556540 217274 556568 220458
rect 557184 219434 557212 228618
rect 558196 225894 558224 255546
rect 559564 246356 559616 246362
rect 559564 246298 559616 246304
rect 559576 236842 559604 246298
rect 559564 236836 559616 236842
rect 559564 236778 559616 236784
rect 560956 230110 560984 256702
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 560944 230104 560996 230110
rect 560944 230046 560996 230052
rect 559564 229900 559616 229906
rect 559564 229842 559616 229848
rect 558184 225888 558236 225894
rect 558184 225830 558236 225836
rect 558276 225616 558328 225622
rect 558276 225558 558328 225564
rect 557632 225140 557684 225146
rect 557632 225082 557684 225088
rect 557644 224806 557672 225082
rect 557632 224800 557684 224806
rect 557632 224742 557684 224748
rect 557816 224800 557868 224806
rect 557816 224742 557868 224748
rect 557828 224210 557856 224742
rect 557998 224632 558054 224641
rect 557998 224567 558054 224576
rect 558012 224398 558040 224567
rect 558000 224392 558052 224398
rect 558000 224334 558052 224340
rect 557552 224194 557856 224210
rect 557540 224188 557856 224194
rect 557592 224182 557856 224188
rect 557540 224130 557592 224136
rect 557540 223032 557592 223038
rect 557540 222974 557592 222980
rect 557354 222320 557410 222329
rect 557354 222255 557410 222264
rect 557368 221882 557396 222255
rect 557552 221921 557580 222974
rect 557538 221912 557594 221921
rect 557356 221876 557408 221882
rect 557538 221847 557594 221856
rect 557356 221818 557408 221824
rect 558288 220522 558316 225558
rect 559012 223168 559064 223174
rect 559012 223110 559064 223116
rect 558276 220516 558328 220522
rect 558276 220458 558328 220464
rect 557184 219406 557396 219434
rect 557368 219298 557396 219406
rect 557356 219292 557408 219298
rect 557356 219234 557408 219240
rect 557368 217274 557396 219234
rect 558288 217274 558316 220458
rect 554056 217246 554130 217274
rect 554884 217246 554958 217274
rect 555712 217246 555786 217274
rect 556540 217246 556614 217274
rect 557368 217246 557442 217274
rect 552400 217110 552474 217138
rect 552446 216988 552474 217110
rect 553274 216988 553302 217246
rect 554102 216988 554130 217246
rect 554930 216988 554958 217246
rect 555758 216988 555786 217246
rect 556586 216988 556614 217246
rect 557414 216988 557442 217246
rect 558242 217246 558316 217274
rect 559024 217274 559052 223110
rect 559576 222086 559604 229842
rect 560944 227180 560996 227186
rect 560944 227122 560996 227128
rect 559840 223032 559892 223038
rect 559840 222974 559892 222980
rect 559380 222080 559432 222086
rect 559378 222048 559380 222057
rect 559564 222080 559616 222086
rect 559432 222048 559434 222057
rect 559564 222022 559616 222028
rect 559378 221983 559434 221992
rect 559852 217274 559880 222974
rect 560668 219292 560720 219298
rect 560668 219234 560720 219240
rect 560680 218890 560708 219234
rect 560484 218884 560536 218890
rect 560484 218826 560536 218832
rect 560668 218884 560720 218890
rect 560668 218826 560720 218832
rect 560298 218648 560354 218657
rect 560298 218583 560354 218592
rect 560312 218210 560340 218583
rect 560496 218210 560524 218826
rect 560300 218204 560352 218210
rect 560300 218146 560352 218152
rect 560484 218204 560536 218210
rect 560484 218146 560536 218152
rect 560956 217569 560984 227122
rect 561956 225140 562008 225146
rect 561956 225082 562008 225088
rect 561968 223310 561996 225082
rect 562336 224806 562364 252554
rect 563716 225010 563744 259422
rect 568120 230104 568172 230110
rect 568120 230046 568172 230052
rect 566832 229764 566884 229770
rect 566832 229706 566884 229712
rect 565636 228404 565688 228410
rect 565636 228346 565688 228352
rect 563980 225752 564032 225758
rect 563980 225694 564032 225700
rect 563704 225004 563756 225010
rect 563704 224946 563756 224952
rect 562140 224800 562192 224806
rect 562138 224768 562140 224777
rect 562324 224800 562376 224806
rect 562192 224768 562194 224777
rect 562324 224742 562376 224748
rect 563702 224768 563758 224777
rect 562138 224703 562194 224712
rect 563702 224703 563758 224712
rect 561956 223304 562008 223310
rect 561956 223246 562008 223252
rect 561494 222048 561550 222057
rect 561494 221983 561550 221992
rect 560758 217560 560814 217569
rect 560758 217495 560814 217504
rect 560942 217560 560998 217569
rect 560942 217495 560998 217504
rect 559024 217246 559098 217274
rect 559852 217246 559926 217274
rect 558242 216988 558270 217246
rect 559070 216988 559098 217246
rect 559898 216988 559926 217246
rect 560772 217138 560800 217495
rect 561508 217274 561536 221983
rect 561968 220674 561996 223246
rect 562324 223168 562376 223174
rect 562324 223110 562376 223116
rect 562336 222494 562364 223110
rect 562324 222488 562376 222494
rect 562324 222430 562376 222436
rect 562324 221944 562376 221950
rect 562324 221886 562376 221892
rect 562336 221762 562364 221886
rect 563716 221785 563744 224703
rect 563702 221776 563758 221785
rect 562336 221746 562732 221762
rect 562336 221740 562744 221746
rect 562336 221734 562692 221740
rect 563702 221711 563758 221720
rect 562692 221682 562744 221688
rect 561968 220646 562180 220674
rect 561770 220552 561826 220561
rect 561770 220487 561772 220496
rect 561824 220487 561826 220496
rect 561956 220516 562008 220522
rect 561772 220458 561824 220464
rect 561956 220458 562008 220464
rect 561968 220114 561996 220458
rect 561956 220108 562008 220114
rect 561956 220050 562008 220056
rect 562152 219434 562180 220646
rect 563150 220552 563206 220561
rect 563150 220487 563152 220496
rect 563204 220487 563206 220496
rect 563152 220458 563204 220464
rect 562324 220380 562376 220386
rect 562324 220322 562376 220328
rect 562336 220046 562364 220322
rect 562324 220040 562376 220046
rect 562324 219982 562376 219988
rect 562152 219406 562364 219434
rect 561680 219020 561732 219026
rect 561680 218962 561732 218968
rect 561692 218657 561720 218962
rect 561678 218648 561734 218657
rect 561678 218583 561734 218592
rect 562336 217274 562364 219406
rect 563012 219056 563068 219065
rect 563012 218991 563014 219000
rect 563066 218991 563068 219000
rect 563152 219020 563204 219026
rect 563014 218962 563066 218968
rect 563152 218962 563204 218968
rect 563164 218226 563192 218962
rect 563026 218210 563192 218226
rect 563014 218204 563192 218210
rect 563066 218198 563192 218204
rect 563014 218146 563066 218152
rect 563520 218000 563572 218006
rect 563072 217948 563520 217954
rect 563072 217942 563572 217948
rect 563072 217926 563560 217942
rect 563072 217682 563100 217926
rect 563026 217654 563100 217682
rect 563026 217326 563054 217654
rect 563150 217560 563206 217569
rect 563150 217495 563206 217504
rect 563164 217326 563192 217495
rect 563014 217320 563066 217326
rect 561508 217246 561582 217274
rect 562336 217246 562410 217274
rect 563014 217262 563066 217268
rect 563152 217320 563204 217326
rect 563152 217262 563204 217268
rect 560726 217110 560800 217138
rect 560726 216988 560754 217110
rect 561554 216988 561582 217246
rect 562382 216988 562410 217246
rect 563716 217138 563744 221711
rect 563992 217274 564020 225694
rect 564808 222080 564860 222086
rect 564808 222022 564860 222028
rect 564820 217841 564848 222022
rect 565648 220561 565676 228346
rect 566844 224618 566872 229706
rect 567016 225072 567068 225078
rect 567016 225014 567068 225020
rect 567028 224806 567056 225014
rect 567016 224800 567068 224806
rect 567016 224742 567068 224748
rect 567200 224800 567252 224806
rect 567200 224742 567252 224748
rect 567212 224618 567240 224742
rect 566844 224590 567240 224618
rect 565634 220552 565690 220561
rect 565634 220487 565690 220496
rect 564806 217832 564862 217841
rect 564806 217767 564862 217776
rect 563992 217246 564066 217274
rect 563210 217110 563744 217138
rect 563210 216988 563238 217110
rect 564038 216988 564066 217246
rect 564820 217138 564848 217767
rect 565648 217274 565676 220487
rect 566844 220386 566872 224590
rect 567844 223304 567896 223310
rect 567844 223246 567896 223252
rect 567856 222494 567884 223246
rect 567844 222488 567896 222494
rect 567844 222430 567896 222436
rect 566464 220380 566516 220386
rect 566464 220322 566516 220328
rect 566832 220380 566884 220386
rect 566832 220322 566884 220328
rect 567292 220380 567344 220386
rect 567292 220322 567344 220328
rect 565648 217246 565722 217274
rect 564820 217110 564894 217138
rect 564866 216988 564894 217110
rect 565694 216988 565722 217246
rect 566476 217138 566504 220322
rect 567304 217274 567332 220322
rect 567660 219020 567712 219026
rect 567660 218962 567712 218968
rect 567844 219020 567896 219026
rect 567844 218962 567896 218968
rect 567672 218793 567700 218962
rect 567658 218784 567714 218793
rect 567856 218754 567884 218962
rect 567658 218719 567714 218728
rect 567844 218748 567896 218754
rect 567844 218690 567896 218696
rect 568132 217274 568160 230046
rect 568592 220386 568620 260850
rect 570616 234598 570644 261462
rect 596824 245676 596876 245682
rect 596824 245618 596876 245624
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 570604 228540 570656 228546
rect 570604 228482 570656 228488
rect 569132 225072 569184 225078
rect 569132 225014 569184 225020
rect 569144 224954 569172 225014
rect 568856 224936 568908 224942
rect 569144 224926 569264 224954
rect 568856 224878 568908 224884
rect 568580 220380 568632 220386
rect 568580 220322 568632 220328
rect 568302 218784 568358 218793
rect 568302 218719 568304 218728
rect 568356 218719 568358 218728
rect 568304 218690 568356 218696
rect 568868 217274 568896 224878
rect 569236 224806 569264 224926
rect 569224 224800 569276 224806
rect 569224 224742 569276 224748
rect 569958 220552 570014 220561
rect 569958 220487 570014 220496
rect 569776 220380 569828 220386
rect 569776 220322 569828 220328
rect 567304 217246 567378 217274
rect 568132 217246 568206 217274
rect 568868 217246 569034 217274
rect 566476 217110 566550 217138
rect 566522 216988 566550 217110
rect 567350 216988 567378 217246
rect 568178 216988 568206 217246
rect 569006 216988 569034 217246
rect 569788 217138 569816 220322
rect 569972 220318 570000 220487
rect 569960 220312 570012 220318
rect 569960 220254 570012 220260
rect 570616 217274 570644 228482
rect 571340 225888 571392 225894
rect 571340 225830 571392 225836
rect 571352 224954 571380 225830
rect 571352 224926 571564 224954
rect 571340 224800 571392 224806
rect 571340 224742 571392 224748
rect 570616 217246 570690 217274
rect 569788 217110 569862 217138
rect 569834 216988 569862 217110
rect 570662 216988 570690 217246
rect 571352 217138 571380 224742
rect 571536 217274 571564 224926
rect 572444 224936 572496 224942
rect 572444 224878 572496 224884
rect 571708 224800 571760 224806
rect 571708 224742 571760 224748
rect 571720 224194 571748 224742
rect 572456 224194 572484 224878
rect 571708 224188 571760 224194
rect 571708 224130 571760 224136
rect 572444 224188 572496 224194
rect 572444 224130 572496 224136
rect 572626 221776 572682 221785
rect 572626 221711 572682 221720
rect 572640 220402 572668 221711
rect 572640 220386 572714 220402
rect 572640 220380 572726 220386
rect 572640 220374 572674 220380
rect 572674 220322 572726 220328
rect 572076 220176 572128 220182
rect 572076 220118 572128 220124
rect 572088 219450 572116 220118
rect 572088 219422 572714 219450
rect 572686 219366 572714 219422
rect 572536 219360 572588 219366
rect 572536 219302 572588 219308
rect 572674 219360 572726 219366
rect 572674 219302 572726 219308
rect 572548 219201 572576 219302
rect 572534 219192 572590 219201
rect 572534 219127 572590 219136
rect 574742 219192 574798 219201
rect 574742 219127 574798 219136
rect 574560 219020 574612 219026
rect 574560 218962 574612 218968
rect 572534 218920 572590 218929
rect 572534 218855 572590 218864
rect 571708 218748 571760 218754
rect 571708 218690 571760 218696
rect 571892 218748 571944 218754
rect 571892 218690 571944 218696
rect 571720 217682 571748 218690
rect 571904 217841 571932 218690
rect 572548 218226 572576 218855
rect 572548 218210 572714 218226
rect 572548 218204 572726 218210
rect 572548 218198 572674 218204
rect 572674 218146 572726 218152
rect 572168 218000 572220 218006
rect 572220 217948 572300 217954
rect 572168 217942 572300 217948
rect 572180 217926 572300 217942
rect 571890 217832 571946 217841
rect 571890 217767 571946 217776
rect 572074 217832 572130 217841
rect 572074 217767 572130 217776
rect 572088 217682 572116 217767
rect 571720 217654 572116 217682
rect 572272 217682 572300 217926
rect 574374 217832 574430 217841
rect 574374 217767 574430 217776
rect 572272 217654 572714 217682
rect 572534 217560 572590 217569
rect 572534 217495 572590 217504
rect 572548 217326 572576 217495
rect 572686 217326 572714 217654
rect 574190 217560 574246 217569
rect 574190 217495 574246 217504
rect 572536 217320 572588 217326
rect 571536 217246 572346 217274
rect 572536 217262 572588 217268
rect 572674 217320 572726 217326
rect 572674 217262 572726 217268
rect 571352 217110 571518 217138
rect 571490 216988 571518 217110
rect 572318 216988 572346 217246
rect 574204 217054 574232 217495
rect 574192 217048 574244 217054
rect 574192 216990 574244 216996
rect 53286 215112 53342 215121
rect 53286 215047 53342 215056
rect 574388 214742 574416 217767
rect 574376 214736 574428 214742
rect 574376 214678 574428 214684
rect 574572 214606 574600 218962
rect 574756 214878 574784 219127
rect 575478 216744 575534 216753
rect 575478 216679 575534 216688
rect 574744 214872 574796 214878
rect 574744 214814 574796 214820
rect 574560 214600 574612 214606
rect 574560 214542 574612 214548
rect 575492 213246 575520 216679
rect 575480 213240 575532 213246
rect 575480 213182 575532 213188
rect 51722 180840 51778 180849
rect 51722 180775 51778 180784
rect 577516 99142 577544 240110
rect 591486 224224 591542 224233
rect 591486 224159 591542 224168
rect 586980 223304 587032 223310
rect 586980 223246 587032 223252
rect 586992 222222 587020 223246
rect 587164 223168 587216 223174
rect 587164 223110 587216 223116
rect 587176 222222 587204 223110
rect 586980 222216 587032 222222
rect 586980 222158 587032 222164
rect 587164 222216 587216 222222
rect 587164 222158 587216 222164
rect 586980 219156 587032 219162
rect 586980 219098 587032 219104
rect 586992 218346 587020 219098
rect 587164 219020 587216 219026
rect 587164 218962 587216 218968
rect 587176 218346 587204 218962
rect 586980 218340 587032 218346
rect 586980 218282 587032 218288
rect 587164 218340 587216 218346
rect 587164 218282 587216 218288
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578514 211712 578570 211721
rect 578514 211647 578570 211656
rect 578528 211206 578556 211647
rect 578516 211200 578568 211206
rect 578516 211142 578568 211148
rect 578896 208350 578924 213959
rect 591304 212560 591356 212566
rect 591304 212502 591356 212508
rect 580908 211200 580960 211206
rect 580908 211142 580960 211148
rect 579528 209840 579580 209846
rect 579526 209808 579528 209817
rect 579580 209808 579582 209817
rect 579526 209743 579582 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 580920 206922 580948 211142
rect 582288 209840 582340 209846
rect 582288 209782 582340 209788
rect 581644 208616 581696 208622
rect 581644 208558 581696 208564
rect 580908 206916 580960 206922
rect 580908 206858 580960 206864
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 580264 171148 580316 171154
rect 580264 171090 580316 171096
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 580276 167346 580304 171090
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 578240 167340 578292 167346
rect 578240 167282 578292 167288
rect 580264 167340 580316 167346
rect 580264 167282 580316 167288
rect 578252 166977 578280 167282
rect 579988 167068 580040 167074
rect 579988 167010 580040 167016
rect 578238 166968 578294 166977
rect 578238 166903 578294 166912
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579344 165232 579396 165238
rect 579344 165174 579396 165180
rect 578240 163668 578292 163674
rect 578240 163610 578292 163616
rect 578252 159905 578280 163610
rect 579356 162761 579384 165174
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 580000 163674 580028 167010
rect 579988 163668 580040 163674
rect 579988 163610 580040 163616
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579342 162752 579398 162761
rect 578424 162716 578476 162722
rect 579342 162687 579398 162696
rect 578424 162658 578476 162664
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162658
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 580552 154698 580580 161434
rect 580724 160132 580776 160138
rect 580724 160074 580776 160080
rect 578332 154692 578384 154698
rect 578332 154634 578384 154640
rect 580540 154692 580592 154698
rect 580540 154634 580592 154640
rect 578344 154057 578372 154634
rect 578330 154048 578386 154057
rect 578330 153983 578386 153992
rect 580736 152794 580764 160074
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 580724 152788 580776 152794
rect 580724 152730 580776 152736
rect 578252 151745 578280 152730
rect 580264 151836 580316 151842
rect 580264 151778 580316 151784
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 148368 579580 148374
rect 579528 148310 579580 148316
rect 579540 147529 579568 148310
rect 579526 147520 579582 147529
rect 579526 147455 579582 147464
rect 578884 146328 578936 146334
rect 578884 146270 578936 146276
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 578896 136649 578924 146270
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580276 140758 580304 151778
rect 580448 140820 580500 140826
rect 580448 140762 580500 140768
rect 580264 140752 580316 140758
rect 580264 140694 580316 140700
rect 579528 138712 579580 138718
rect 579528 138654 579580 138660
rect 579068 137352 579120 137358
rect 579068 137294 579120 137300
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 579080 132297 579108 137294
rect 579540 134473 579568 138654
rect 580264 134564 580316 134570
rect 580264 134506 580316 134512
rect 579526 134464 579582 134473
rect 579526 134399 579582 134408
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578884 131164 578936 131170
rect 578884 131106 578936 131112
rect 578896 129713 578924 131106
rect 578882 129704 578938 129713
rect 578882 129639 578938 129648
rect 579528 129056 579580 129062
rect 579528 128998 579580 129004
rect 579540 127945 579568 128998
rect 579526 127936 579582 127945
rect 579526 127871 579582 127880
rect 579068 127016 579120 127022
rect 579068 126958 579120 126964
rect 578332 125656 578384 125662
rect 578332 125598 578384 125604
rect 578344 125361 578372 125598
rect 578330 125352 578386 125361
rect 578330 125287 578386 125296
rect 578424 123616 578476 123622
rect 578422 123584 578424 123593
rect 578476 123584 578478 123593
rect 578422 123519 578478 123528
rect 578884 122188 578936 122194
rect 578884 122130 578936 122136
rect 578896 121417 578924 122130
rect 578882 121408 578938 121417
rect 578882 121343 578938 121352
rect 578516 118448 578568 118454
rect 578514 118416 578516 118425
rect 578568 118416 578570 118425
rect 578514 118351 578570 118360
rect 578332 108724 578384 108730
rect 578332 108666 578384 108672
rect 578344 108361 578372 108666
rect 578330 108352 578386 108361
rect 578330 108287 578386 108296
rect 578884 107636 578936 107642
rect 578884 107578 578936 107584
rect 578608 99272 578660 99278
rect 578606 99240 578608 99249
rect 578660 99240 578662 99249
rect 578606 99175 578662 99184
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578332 97980 578384 97986
rect 578332 97922 578384 97928
rect 578344 97481 578372 97922
rect 578330 97472 578386 97481
rect 578330 97407 578386 97416
rect 578516 93492 578568 93498
rect 578516 93434 578568 93440
rect 578528 93129 578556 93434
rect 578514 93120 578570 93129
rect 578514 93055 578570 93064
rect 578896 80073 578924 107578
rect 579080 105913 579108 126958
rect 580276 118454 580304 134506
rect 580460 125662 580488 140762
rect 580448 125656 580500 125662
rect 580448 125598 580500 125604
rect 580448 124228 580500 124234
rect 580448 124170 580500 124176
rect 580264 118448 580316 118454
rect 580264 118390 580316 118396
rect 579528 116952 579580 116958
rect 579526 116920 579528 116929
rect 579580 116920 579582 116929
rect 579526 116855 579582 116864
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 579528 112872 579580 112878
rect 579528 112814 579580 112820
rect 579540 112577 579568 112814
rect 579526 112568 579582 112577
rect 579526 112503 579582 112512
rect 579344 110152 579396 110158
rect 579342 110120 579344 110129
rect 579396 110120 579398 110129
rect 579342 110055 579398 110064
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 580264 104916 580316 104922
rect 580264 104858 580316 104864
rect 579528 103488 579580 103494
rect 579528 103430 579580 103436
rect 579540 103329 579568 103430
rect 579526 103320 579582 103329
rect 579526 103255 579582 103264
rect 579528 101856 579580 101862
rect 579528 101798 579580 101804
rect 579540 101697 579568 101798
rect 579526 101688 579582 101697
rect 579526 101623 579582 101632
rect 579068 99408 579120 99414
rect 579068 99350 579120 99356
rect 579080 90953 579108 99350
rect 579528 95056 579580 95062
rect 579526 95024 579528 95033
rect 579580 95024 579582 95033
rect 579526 94959 579582 94968
rect 579344 91112 579396 91118
rect 579344 91054 579396 91060
rect 579066 90944 579122 90953
rect 579066 90879 579122 90888
rect 579356 86465 579384 91054
rect 579528 88120 579580 88126
rect 579526 88088 579528 88097
rect 579580 88088 579582 88097
rect 579526 88023 579582 88032
rect 579342 86456 579398 86465
rect 579342 86391 579398 86400
rect 579160 84176 579212 84182
rect 579160 84118 579212 84124
rect 579172 84017 579200 84118
rect 579158 84008 579214 84017
rect 579158 83943 579214 83952
rect 579068 82408 579120 82414
rect 579068 82350 579120 82356
rect 579080 82249 579108 82350
rect 579066 82240 579122 82249
rect 579066 82175 579122 82184
rect 579528 82136 579580 82142
rect 579528 82078 579580 82084
rect 578882 80064 578938 80073
rect 578882 79999 578938 80008
rect 579068 79348 579120 79354
rect 579068 79290 579120 79296
rect 578240 75880 578292 75886
rect 578240 75822 578292 75828
rect 578252 75585 578280 75822
rect 578238 75576 578294 75585
rect 578238 75511 578294 75520
rect 579080 73137 579108 79290
rect 579540 77897 579568 82078
rect 579526 77888 579582 77897
rect 579526 77823 579582 77832
rect 580276 75886 580304 104858
rect 580460 99278 580488 124170
rect 580632 122052 580684 122058
rect 580632 121994 580684 122000
rect 580644 108730 580672 121994
rect 581656 114510 581684 208558
rect 582300 205562 582328 209782
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 206916 589516 206922
rect 589464 206858 589516 206864
rect 589476 206417 589504 206858
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 582288 205556 582340 205562
rect 582288 205498 582340 205504
rect 589464 205556 589516 205562
rect 589464 205498 589516 205504
rect 589476 204785 589504 205498
rect 589462 204776 589518 204785
rect 589462 204711 589518 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589646 170504 589702 170513
rect 589646 170439 589702 170448
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 582380 168428 582432 168434
rect 582380 168370 582432 168376
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 582392 165238 582420 168370
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589660 166326 589688 170439
rect 589648 166320 589700 166326
rect 589648 166262 589700 166268
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 582380 165232 582432 165238
rect 582380 165174 582432 165180
rect 589476 164286 589504 165543
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 582484 162722 582512 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 582472 162716 582524 162722
rect 582472 162658 582524 162664
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158778 589504 159015
rect 585784 158772 585836 158778
rect 585784 158714 585836 158720
rect 589464 158772 589516 158778
rect 589464 158714 589516 158720
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 150618 585824 158714
rect 589278 157448 589334 157457
rect 587164 157412 587216 157418
rect 589278 157383 589280 157392
rect 587164 157354 587216 157360
rect 589332 157383 589334 157392
rect 589280 157354 589332 157360
rect 585784 150612 585836 150618
rect 585784 150554 585836 150560
rect 585140 149116 585192 149122
rect 585140 149058 585192 149064
rect 585152 146334 585180 149058
rect 587176 148374 587204 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 590014 150920 590070 150929
rect 590014 150855 590070 150864
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 587164 148368 587216 148374
rect 587164 148310 587216 148316
rect 588542 147656 588598 147665
rect 588542 147591 588598 147600
rect 585140 146328 585192 146334
rect 585140 146270 585192 146276
rect 584772 144968 584824 144974
rect 584772 144910 584824 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 139460 583076 139466
rect 583024 139402 583076 139408
rect 581828 131300 581880 131306
rect 581828 131242 581880 131248
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 110492 581696 110498
rect 581644 110434 581696 110440
rect 580632 108724 580684 108730
rect 580632 108666 580684 108672
rect 580448 99272 580500 99278
rect 580448 99214 580500 99220
rect 581656 84182 581684 110434
rect 581840 110158 581868 131242
rect 583036 123622 583064 139402
rect 584784 137358 584812 144910
rect 585968 143608 586020 143614
rect 585968 143550 586020 143556
rect 584772 137352 584824 137358
rect 584772 137294 584824 137300
rect 584588 136672 584640 136678
rect 584588 136614 584640 136620
rect 583208 129192 583260 129198
rect 583208 129134 583260 129140
rect 583024 123616 583076 123622
rect 583024 123558 583076 123564
rect 583220 116958 583248 129134
rect 584404 122868 584456 122874
rect 584404 122810 584456 122816
rect 583208 116952 583260 116958
rect 583208 116894 583260 116900
rect 583208 115252 583260 115258
rect 583208 115194 583260 115200
rect 583024 113212 583076 113218
rect 583024 113154 583076 113160
rect 581828 110152 581880 110158
rect 581828 110094 581880 110100
rect 581644 84176 581696 84182
rect 581644 84118 581696 84124
rect 583036 82414 583064 113154
rect 583220 95062 583248 115194
rect 584416 101862 584444 122810
rect 584600 122194 584628 136614
rect 585784 132524 585836 132530
rect 585784 132466 585836 132472
rect 584588 122188 584640 122194
rect 584588 122130 584640 122136
rect 585796 112878 585824 132466
rect 585980 131170 586008 143550
rect 587164 142452 587216 142458
rect 587164 142394 587216 142400
rect 585968 131164 586020 131170
rect 585968 131106 586020 131112
rect 587176 129062 587204 142394
rect 588556 138718 588584 147591
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589830 142760 589886 142769
rect 589830 142695 589886 142704
rect 589844 142458 589872 142695
rect 589832 142452 589884 142458
rect 589832 142394 589884 142400
rect 590028 142154 590056 150855
rect 589936 142126 590056 142154
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589936 139330 589964 142126
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 588544 138712 588596 138718
rect 588544 138654 588596 138660
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 134570 589504 136167
rect 590382 134600 590438 134609
rect 589464 134564 589516 134570
rect 590382 134535 590438 134544
rect 589464 134506 589516 134512
rect 589462 132968 589518 132977
rect 589462 132903 589518 132912
rect 589476 132530 589504 132903
rect 589464 132524 589516 132530
rect 589464 132466 589516 132472
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 588542 129704 588598 129713
rect 588542 129639 588598 129648
rect 587164 129056 587216 129062
rect 587164 128998 587216 129004
rect 587348 118720 587400 118726
rect 587348 118662 587400 118668
rect 586152 116000 586204 116006
rect 586152 115942 586204 115948
rect 585784 112872 585836 112878
rect 585784 112814 585836 112820
rect 585968 112464 586020 112470
rect 585968 112406 586020 112412
rect 584588 109064 584640 109070
rect 584588 109006 584640 109012
rect 584404 101856 584456 101862
rect 584404 101798 584456 101804
rect 584404 100156 584456 100162
rect 584404 100098 584456 100104
rect 583208 95056 583260 95062
rect 583208 94998 583260 95004
rect 583024 82408 583076 82414
rect 583024 82350 583076 82356
rect 581642 77888 581698 77897
rect 581642 77823 581698 77832
rect 580264 75880 580316 75886
rect 580264 75822 580316 75828
rect 579066 73128 579122 73137
rect 579066 73063 579122 73072
rect 578884 72480 578936 72486
rect 578884 72422 578936 72428
rect 577504 60036 577556 60042
rect 577504 59978 577556 59984
rect 576124 58676 576176 58682
rect 576124 58618 576176 58624
rect 574928 57248 574980 57254
rect 574928 57190 574980 57196
rect 574744 56024 574796 56030
rect 574744 55966 574796 55972
rect 574560 55888 574612 55894
rect 574560 55830 574612 55836
rect 574572 53990 574600 55830
rect 574756 54126 574784 55966
rect 574744 54120 574796 54126
rect 574744 54062 574796 54068
rect 574560 53984 574612 53990
rect 574560 53926 574612 53932
rect 574940 53854 574968 57190
rect 576136 55049 576164 58618
rect 576122 55040 576178 55049
rect 576122 54975 576178 54984
rect 577516 54233 577544 59978
rect 578896 54505 578924 72422
rect 579068 71392 579120 71398
rect 579068 71334 579120 71340
rect 579080 71233 579108 71334
rect 579066 71224 579122 71233
rect 579066 71159 579122 71168
rect 580264 68332 580316 68338
rect 580264 68274 580316 68280
rect 580276 54777 580304 68274
rect 580262 54768 580318 54777
rect 580262 54703 580318 54712
rect 578882 54496 578938 54505
rect 578882 54431 578938 54440
rect 581656 54262 581684 77823
rect 584416 71398 584444 100098
rect 584600 91118 584628 109006
rect 585980 93498 586008 112406
rect 586164 99414 586192 115942
rect 587164 106344 587216 106350
rect 587164 106286 587216 106292
rect 586152 99408 586204 99414
rect 586152 99350 586204 99356
rect 585968 93492 586020 93498
rect 585968 93434 586020 93440
rect 584588 91112 584640 91118
rect 584588 91054 584640 91060
rect 585140 89004 585192 89010
rect 585140 88946 585192 88952
rect 585152 88126 585180 88946
rect 585140 88120 585192 88126
rect 585140 88062 585192 88068
rect 587176 82142 587204 106286
rect 587360 97986 587388 118662
rect 588556 103494 588584 129639
rect 590396 129198 590424 134535
rect 590384 129192 590436 129198
rect 590384 129134 590436 129140
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 589922 126440 589978 126449
rect 589922 126375 589978 126384
rect 589462 124808 589518 124817
rect 589462 124743 589518 124752
rect 589476 124234 589504 124743
rect 589464 124228 589516 124234
rect 589464 124170 589516 124176
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589936 122058 589964 126375
rect 589924 122052 589976 122058
rect 589924 121994 589976 122000
rect 590014 121544 590070 121553
rect 590014 121479 590070 121488
rect 589646 119912 589702 119921
rect 589646 119847 589702 119856
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589660 115258 589688 119847
rect 590028 118726 590056 121479
rect 590016 118720 590068 118726
rect 590016 118662 590068 118668
rect 590106 118280 590162 118289
rect 590106 118215 590162 118224
rect 589648 115252 589700 115258
rect 589648 115194 589700 115200
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 590120 112470 590148 118215
rect 590290 115016 590346 115025
rect 590290 114951 590346 114960
rect 590108 112464 590160 112470
rect 590108 112406 590160 112412
rect 589462 111752 589518 111761
rect 589462 111687 589518 111696
rect 589476 110498 589504 111687
rect 589464 110492 589516 110498
rect 589464 110434 589516 110440
rect 589278 110120 589334 110129
rect 589278 110055 589334 110064
rect 589292 109070 589320 110055
rect 589280 109064 589332 109070
rect 589280 109006 589332 109012
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589830 106856 589886 106865
rect 589830 106791 589886 106800
rect 589844 106350 589872 106791
rect 589832 106344 589884 106350
rect 589832 106286 589884 106292
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 588726 103592 588782 103601
rect 588726 103527 588782 103536
rect 588544 103488 588596 103494
rect 588544 103430 588596 103436
rect 587348 97980 587400 97986
rect 587348 97922 587400 97928
rect 587164 82136 587216 82142
rect 587164 82078 587216 82084
rect 588740 79354 588768 103527
rect 590304 103514 590332 114951
rect 589936 103486 590332 103514
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100162 589504 101895
rect 589464 100156 589516 100162
rect 589464 100098 589516 100104
rect 589936 89010 589964 103486
rect 589924 89004 589976 89010
rect 589924 88946 589976 88952
rect 588728 79348 588780 79354
rect 588728 79290 588780 79296
rect 584404 71392 584456 71398
rect 584404 71334 584456 71340
rect 581644 54256 581696 54262
rect 577502 54224 577558 54233
rect 581644 54198 581696 54204
rect 577502 54159 577558 54168
rect 574928 53848 574980 53854
rect 574928 53790 574980 53796
rect 459834 53680 459890 53689
rect 459834 53615 459890 53624
rect 460754 53680 460810 53689
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 461674 53615 461730 53624
rect 462594 53680 462650 53689
rect 462594 53615 462650 53624
rect 464160 53644 464212 53650
rect 129004 53236 129056 53242
rect 129004 53178 129056 53184
rect 128820 51740 128872 51746
rect 128820 51682 128872 51688
rect 50528 49156 50580 49162
rect 50528 49098 50580 49104
rect 46204 49020 46256 49026
rect 46204 48962 46256 48968
rect 128832 44810 128860 51682
rect 129016 45354 129044 53178
rect 312360 53168 312412 53174
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 130384 53100 130436 53106
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 130384 53042 130436 53048
rect 129188 51876 129240 51882
rect 129188 51818 129240 51824
rect 129556 51876 129608 51882
rect 129556 51818 129608 51824
rect 129004 45348 129056 45354
rect 129004 45290 129056 45296
rect 128820 44804 128872 44810
rect 128820 44746 128872 44752
rect 129200 44538 129228 51818
rect 129372 49156 129424 49162
rect 129372 49098 129424 49104
rect 129384 44946 129412 49098
rect 129568 45082 129596 51818
rect 129556 45076 129608 45082
rect 129556 45018 129608 45024
rect 129372 44940 129424 44946
rect 129372 44882 129424 44888
rect 129188 44532 129240 44538
rect 129188 44474 129240 44480
rect 43628 44328 43680 44334
rect 130396 44305 130424 53042
rect 130568 52012 130620 52018
rect 130568 51954 130620 51960
rect 130580 45558 130608 51954
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459468 53100 459520 53106
rect 459468 53042 459520 53048
rect 459480 52578 459508 53042
rect 459848 52578 459876 53615
rect 460066 52828 460118 52834
rect 460066 52770 460118 52776
rect 459172 52550 459508 52578
rect 459632 52550 459876 52578
rect 460078 52564 460106 52770
rect 460768 52578 460796 53615
rect 461308 53372 461360 53378
rect 461308 53314 461360 53320
rect 461320 52578 461348 53314
rect 461688 52578 461716 53615
rect 462228 53508 462280 53514
rect 462228 53450 462280 53456
rect 462240 52578 462268 53450
rect 462608 52578 462636 53615
rect 464160 53586 464212 53592
rect 464344 53644 464396 53650
rect 464344 53586 464396 53592
rect 464528 53644 464580 53650
rect 464528 53586 464580 53592
rect 464896 53644 464948 53650
rect 464896 53586 464948 53592
rect 465908 53644 465960 53650
rect 465908 53586 465960 53592
rect 466092 53644 466144 53650
rect 466092 53586 466144 53592
rect 473728 53644 473780 53650
rect 473728 53586 473780 53592
rect 464172 53417 464200 53586
rect 464158 53408 464214 53417
rect 464158 53343 464214 53352
rect 464068 53236 464120 53242
rect 464068 53178 464120 53184
rect 463148 52964 463200 52970
rect 463148 52906 463200 52912
rect 463160 52578 463188 52906
rect 463608 52692 463660 52698
rect 463608 52634 463660 52640
rect 463620 52578 463648 52634
rect 464080 52578 464108 53178
rect 464356 52578 464384 53586
rect 464540 52698 464568 53586
rect 464710 53408 464766 53417
rect 464710 53343 464766 53352
rect 464528 52692 464580 52698
rect 464528 52634 464580 52640
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461932 52550 462268 52578
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463648 52578
rect 463772 52550 464108 52578
rect 464232 52550 464384 52578
rect 464724 52442 464752 53343
rect 464908 53106 464936 53586
rect 464896 53100 464948 53106
rect 464896 53042 464948 53048
rect 465448 52692 465500 52698
rect 465448 52634 465500 52640
rect 465460 52578 465488 52634
rect 465920 52578 465948 53586
rect 466104 52834 466132 53586
rect 471980 53576 472032 53582
rect 471794 53544 471850 53553
rect 471980 53518 472032 53524
rect 472808 53576 472860 53582
rect 472808 53518 472860 53524
rect 473542 53544 473598 53553
rect 471794 53479 471796 53488
rect 471848 53479 471850 53488
rect 471796 53450 471848 53456
rect 471992 53242 472020 53518
rect 471980 53236 472032 53242
rect 471980 53178 472032 53184
rect 466092 52828 466144 52834
rect 466092 52770 466144 52776
rect 472820 52698 472848 53518
rect 473542 53479 473544 53488
rect 473596 53479 473598 53488
rect 473544 53450 473596 53456
rect 473740 52970 473768 53586
rect 473728 52964 473780 52970
rect 473728 52906 473780 52912
rect 472808 52692 472860 52698
rect 472808 52634 472860 52640
rect 465152 52550 465488 52578
rect 465612 52550 465948 52578
rect 464692 52414 464752 52442
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458180 50516 458232 50522
rect 458180 50458 458232 50464
rect 130752 50380 130804 50386
rect 130752 50322 130804 50328
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 130568 45552 130620 45558
rect 130568 45494 130620 45500
rect 43628 44270 43680 44276
rect 130382 44296 130438 44305
rect 130382 44231 130438 44240
rect 43444 44192 43496 44198
rect 43444 44134 43496 44140
rect 130764 44062 130792 50322
rect 130936 49020 130988 49026
rect 130936 48962 130988 48968
rect 130948 45234 130976 48962
rect 458192 47025 458220 50458
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 458364 50380 458416 50386
rect 458364 50322 458416 50328
rect 522948 50380 523000 50386
rect 522948 50322 523000 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50322
rect 522960 47841 522988 50322
rect 522946 47832 523002 47841
rect 522946 47767 523002 47776
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461072 47682
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 462392 47654 462728 47682
rect 462852 47654 462912 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132592 45552 132644 45558
rect 132592 45494 132644 45500
rect 130948 45218 131436 45234
rect 130948 45212 131448 45218
rect 130948 45206 131396 45212
rect 131396 45154 131448 45160
rect 131580 44668 131632 44674
rect 131580 44610 131632 44616
rect 131592 44198 131620 44610
rect 132604 44422 132632 45494
rect 133144 45212 133196 45218
rect 133144 45154 133196 45160
rect 132592 44416 132644 44422
rect 132592 44358 132644 44364
rect 132408 44328 132460 44334
rect 132406 44296 132408 44305
rect 132460 44296 132462 44305
rect 132406 44231 132462 44240
rect 133156 44198 133184 45154
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 131580 44192 131632 44198
rect 131580 44134 131632 44140
rect 133144 44192 133196 44198
rect 133144 44134 133196 44140
rect 255870 44160 255926 44169
rect 255870 44095 255926 44104
rect 130752 44056 130804 44062
rect 130752 43998 130804 44004
rect 255884 42838 255912 44095
rect 361762 43888 361818 43897
rect 361762 43823 361818 43832
rect 440238 43888 440294 43897
rect 440238 43823 440240 43832
rect 187332 42832 187384 42838
rect 187332 42774 187384 42780
rect 255872 42832 255924 42838
rect 255872 42774 255924 42780
rect 187344 42092 187372 42774
rect 307300 42764 307352 42770
rect 307300 42706 307352 42712
rect 307312 42106 307340 42706
rect 310428 42628 310480 42634
rect 310428 42570 310480 42576
rect 310440 42106 310468 42570
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361776 42092 361804 43823
rect 440292 43823 440294 43832
rect 441066 43888 441122 43897
rect 441066 43823 441068 43832
rect 440240 43794 440292 43800
rect 441120 43823 441122 43832
rect 441068 43794 441120 43800
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 441068 42764 441120 42770
rect 441068 42706 441120 42712
rect 449164 42764 449216 42770
rect 449164 42706 449216 42712
rect 453580 42764 453632 42770
rect 453580 42706 453632 42712
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 415582 42392 415638 42401
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405188 42356 405240 42362
rect 415582 42327 415638 42336
rect 420736 42356 420788 42362
rect 405188 42298 405240 42304
rect 365074 41848 365130 41857
rect 364918 41806 365074 41834
rect 365074 41783 365130 41792
rect 404464 41478 404492 42298
rect 405200 42106 405228 42298
rect 415596 42106 415624 42327
rect 420736 42298 420788 42304
rect 426900 42356 426952 42362
rect 426900 42298 426952 42304
rect 405200 42078 405582 42106
rect 415426 42078 415624 42106
rect 416686 41848 416742 41857
rect 416622 41806 416686 41834
rect 419906 41848 419962 41857
rect 419750 41806 419906 41834
rect 416686 41783 416742 41792
rect 419906 41783 419962 41792
rect 420748 41478 420776 42298
rect 426912 41478 426940 42298
rect 427096 42022 427124 42570
rect 431236 42022 431264 42706
rect 441080 42022 441108 42706
rect 441252 42628 441304 42634
rect 441252 42570 441304 42576
rect 446404 42628 446456 42634
rect 446404 42570 446456 42576
rect 427084 42016 427136 42022
rect 427084 41958 427136 41964
rect 431224 42016 431276 42022
rect 431224 41958 431276 41964
rect 441068 42016 441120 42022
rect 441068 41958 441120 41964
rect 441264 41886 441292 42570
rect 446218 42256 446274 42265
rect 446218 42191 446274 42200
rect 441252 41880 441304 41886
rect 441252 41822 441304 41828
rect 446232 41585 446260 42191
rect 446416 42022 446444 42570
rect 446404 42016 446456 42022
rect 446404 41958 446456 41964
rect 449176 41886 449204 42706
rect 453592 41886 453620 42706
rect 454500 42492 454552 42498
rect 454500 42434 454552 42440
rect 454512 42022 454540 42434
rect 454500 42016 454552 42022
rect 454500 41958 454552 41964
rect 449164 41880 449216 41886
rect 449164 41822 449216 41828
rect 453580 41880 453632 41886
rect 453580 41822 453632 41828
rect 446218 41576 446274 41585
rect 446218 41511 446274 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44169 460152 47654
rect 460110 44160 460166 44169
rect 460110 44095 460166 44104
rect 460860 43489 460888 47654
rect 461044 44441 461072 47654
rect 461030 44432 461086 44441
rect 461030 44367 461086 44376
rect 460846 43480 460902 43489
rect 460846 43415 460902 43424
rect 461780 42945 461808 47654
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 461964 42265 461992 47654
rect 462700 43217 462728 47654
rect 462884 44441 462912 47654
rect 463068 47654 463312 47682
rect 463772 47654 463832 47682
rect 462870 44432 462926 44441
rect 462870 44367 462926 44376
rect 462686 43208 462742 43217
rect 462686 43143 462742 43152
rect 463068 42498 463096 47654
rect 463804 44441 463832 47654
rect 464218 47410 464246 47668
rect 464172 47382 464246 47410
rect 464356 47654 464692 47682
rect 463790 44432 463846 44441
rect 463790 44367 463846 44376
rect 463974 42936 464030 42945
rect 463974 42871 464030 42880
rect 463988 42514 464016 42871
rect 464172 42770 464200 47382
rect 464356 44169 464384 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 47025 465120 47382
rect 465078 47016 465134 47025
rect 465078 46951 465134 46960
rect 465276 46753 465304 47654
rect 545684 47297 545712 53094
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 553688 48113 553716 53094
rect 591316 51882 591344 212502
rect 591500 101697 591528 224159
rect 593972 223304 594024 223310
rect 593972 223246 594024 223252
rect 591684 219694 592034 219722
rect 591684 219366 591712 219694
rect 592006 219638 592034 219694
rect 591856 219632 591908 219638
rect 591856 219574 591908 219580
rect 591994 219632 592046 219638
rect 591994 219574 592046 219580
rect 591868 219366 591896 219574
rect 591672 219360 591724 219366
rect 591672 219302 591724 219308
rect 591856 219360 591908 219366
rect 591856 219302 591908 219308
rect 592684 212696 592736 212702
rect 592684 212638 592736 212644
rect 591486 101688 591542 101697
rect 591486 101623 591542 101632
rect 591304 51876 591356 51882
rect 591304 51818 591356 51824
rect 592696 51746 592724 212638
rect 593984 210202 594012 223246
rect 596836 221882 596864 245618
rect 629944 241528 629996 241534
rect 629944 241470 629996 241476
rect 629956 229094 629984 241470
rect 629956 229066 630076 229094
rect 616052 224800 616104 224806
rect 616052 224742 616104 224748
rect 614948 223644 615000 223650
rect 614948 223586 615000 223592
rect 600596 222012 600648 222018
rect 600596 221954 600648 221960
rect 600964 222012 601016 222018
rect 600964 221954 601016 221960
rect 606668 222012 606720 222018
rect 606668 221954 606720 221960
rect 596824 221876 596876 221882
rect 596824 221818 596876 221824
rect 600608 220998 600636 221954
rect 600976 221474 601004 221954
rect 601792 221604 601844 221610
rect 601792 221546 601844 221552
rect 600964 221468 601016 221474
rect 600964 221410 601016 221416
rect 600870 221232 600926 221241
rect 600870 221167 600926 221176
rect 600412 220992 600464 220998
rect 599490 220960 599546 220969
rect 600412 220934 600464 220940
rect 600596 220992 600648 220998
rect 600596 220934 600648 220940
rect 599490 220895 599546 220904
rect 598572 219904 598624 219910
rect 598572 219846 598624 219852
rect 598584 219502 598612 219846
rect 596180 219496 596232 219502
rect 596180 219438 596232 219444
rect 597744 219496 597796 219502
rect 597744 219438 597796 219444
rect 598572 219496 598624 219502
rect 598572 219438 598624 219444
rect 594800 219156 594852 219162
rect 594800 219098 594852 219104
rect 594812 216782 594840 219098
rect 595166 217288 595222 217297
rect 595166 217223 595222 217232
rect 594800 216776 594852 216782
rect 594800 216718 594852 216724
rect 594800 213240 594852 213246
rect 594800 213182 594852 213188
rect 594812 210202 594840 213182
rect 595180 210202 595208 217223
rect 595718 217016 595774 217025
rect 596192 217002 596220 219438
rect 596192 216974 596772 217002
rect 595718 216951 595774 216960
rect 595732 210202 595760 216951
rect 596364 216912 596416 216918
rect 596364 216854 596416 216860
rect 596376 210202 596404 216854
rect 596744 210202 596772 216974
rect 597756 210202 597784 219438
rect 598848 218612 598900 218618
rect 598848 218554 598900 218560
rect 598860 217326 598888 218554
rect 598480 217320 598532 217326
rect 598480 217262 598532 217268
rect 598848 217320 598900 217326
rect 598848 217262 598900 217268
rect 597928 217184 597980 217190
rect 597928 217126 597980 217132
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596744 210174 597172 210202
rect 597724 210174 597784 210202
rect 597940 210202 597968 217126
rect 598492 210202 598520 217262
rect 599030 215656 599086 215665
rect 599030 215591 599086 215600
rect 599044 210202 599072 215591
rect 599504 210202 599532 220895
rect 600424 213042 600452 220934
rect 600688 220856 600740 220862
rect 600688 220798 600740 220804
rect 600412 213036 600464 213042
rect 600412 212978 600464 212984
rect 600504 212900 600556 212906
rect 600504 212842 600556 212848
rect 600516 210202 600544 212842
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600484 210174 600544 210202
rect 600700 209930 600728 220798
rect 600884 212906 600912 221167
rect 601240 218476 601292 218482
rect 601240 218418 601292 218424
rect 601056 218340 601108 218346
rect 601056 218282 601108 218288
rect 601068 218074 601096 218282
rect 601252 218074 601280 218418
rect 601056 218068 601108 218074
rect 601056 218010 601108 218016
rect 601240 218068 601292 218074
rect 601240 218010 601292 218016
rect 601804 214470 601832 221546
rect 604828 221264 604880 221270
rect 604828 221206 604880 221212
rect 601976 221128 602028 221134
rect 601976 221070 602028 221076
rect 601792 214464 601844 214470
rect 601792 214406 601844 214412
rect 601240 213036 601292 213042
rect 601240 212978 601292 212984
rect 600872 212900 600924 212906
rect 600872 212842 600924 212848
rect 601252 210202 601280 212978
rect 601988 210202 602016 221070
rect 604644 220992 604696 220998
rect 604644 220934 604696 220940
rect 603080 218748 603132 218754
rect 603080 218690 603132 218696
rect 603092 217462 603120 218690
rect 604460 218612 604512 218618
rect 604460 218554 604512 218560
rect 604000 217864 604052 217870
rect 604000 217806 604052 217812
rect 603448 217728 603500 217734
rect 603448 217670 603500 217676
rect 603080 217456 603132 217462
rect 603080 217398 603132 217404
rect 603080 217184 603132 217190
rect 603080 217126 603132 217132
rect 602344 214464 602396 214470
rect 602344 214406 602396 214412
rect 602356 210202 602384 214406
rect 603092 210202 603120 217126
rect 603460 210202 603488 217670
rect 604012 210202 604040 217806
rect 604472 217734 604500 218554
rect 604460 217728 604512 217734
rect 604460 217670 604512 217676
rect 604656 214470 604684 220934
rect 604644 214464 604696 214470
rect 604644 214406 604696 214412
rect 604840 210202 604868 221206
rect 606024 219904 606076 219910
rect 606024 219846 606076 219852
rect 605104 214464 605156 214470
rect 605104 214406 605156 214412
rect 605116 210202 605144 214406
rect 606036 210202 606064 219846
rect 606208 217592 606260 217598
rect 606208 217534 606260 217540
rect 601252 210174 601588 210202
rect 601988 210174 602140 210202
rect 602356 210174 602692 210202
rect 603092 210174 603244 210202
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604840 210174 604900 210202
rect 605116 210174 605452 210202
rect 606004 210174 606064 210202
rect 606220 210202 606248 217534
rect 606680 210202 606708 221954
rect 608600 221740 608652 221746
rect 608600 221682 608652 221688
rect 607312 220040 607364 220046
rect 607312 219982 607364 219988
rect 607128 218340 607180 218346
rect 607128 218282 607180 218288
rect 607140 216918 607168 218282
rect 607128 216912 607180 216918
rect 607128 216854 607180 216860
rect 607324 214606 607352 219982
rect 607496 219496 607548 219502
rect 607496 219438 607548 219444
rect 607312 214600 607364 214606
rect 607312 214542 607364 214548
rect 607508 210202 607536 219438
rect 607864 214600 607916 214606
rect 607864 214542 607916 214548
rect 607876 210202 607904 214542
rect 608612 210202 608640 221682
rect 608876 220652 608928 220658
rect 608876 220594 608928 220600
rect 608888 210202 608916 220594
rect 609428 220516 609480 220522
rect 609428 220458 609480 220464
rect 609440 210202 609468 220458
rect 610532 220380 610584 220386
rect 610532 220322 610584 220328
rect 610072 217048 610124 217054
rect 610072 216990 610124 216996
rect 610084 210202 610112 216990
rect 610544 210202 610572 220322
rect 611634 220280 611690 220289
rect 611452 220244 611504 220250
rect 611634 220215 611690 220224
rect 611452 220186 611504 220192
rect 611464 210202 611492 220186
rect 611648 210202 611676 220215
rect 612738 219736 612794 219745
rect 612738 219671 612794 219680
rect 612280 216912 612332 216918
rect 612280 216854 612332 216860
rect 612292 210202 612320 216854
rect 612752 210202 612780 219671
rect 614120 218884 614172 218890
rect 614120 218826 614172 218832
rect 613568 218204 613620 218210
rect 613568 218146 613620 218152
rect 613384 216776 613436 216782
rect 613384 216718 613436 216724
rect 613396 210202 613424 216718
rect 613580 216714 613608 218146
rect 614132 217598 614160 218826
rect 614304 217728 614356 217734
rect 614304 217670 614356 217676
rect 614120 217592 614172 217598
rect 614120 217534 614172 217540
rect 613568 216708 613620 216714
rect 613568 216650 613620 216656
rect 614316 210202 614344 217670
rect 614488 216708 614540 216714
rect 614488 216650 614540 216656
rect 606220 210174 606556 210202
rect 606680 210174 607108 210202
rect 607508 210174 607660 210202
rect 607876 210174 608212 210202
rect 608612 210174 608764 210202
rect 608888 210174 609316 210202
rect 609440 210174 609868 210202
rect 610084 210174 610420 210202
rect 610544 210174 610972 210202
rect 611464 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612752 210174 613180 210202
rect 613396 210174 613732 210202
rect 614284 210174 614344 210202
rect 614500 210202 614528 216650
rect 614960 210202 614988 223586
rect 615684 218000 615736 218006
rect 615684 217942 615736 217948
rect 615696 210202 615724 217942
rect 616064 210202 616092 224742
rect 625252 224664 625304 224670
rect 625252 224606 625304 224612
rect 623780 224528 623832 224534
rect 623780 224470 623832 224476
rect 622676 224052 622728 224058
rect 622676 223994 622728 224000
rect 619640 223916 619692 223922
rect 619640 223858 619692 223864
rect 618258 221504 618314 221513
rect 618258 221439 618314 221448
rect 617154 220008 617210 220017
rect 617154 219943 617210 219952
rect 616880 214872 616932 214878
rect 616880 214814 616932 214820
rect 616892 210202 616920 214814
rect 617168 210202 617196 219943
rect 617798 215928 617854 215937
rect 617798 215863 617854 215872
rect 617812 210202 617840 215863
rect 618272 214606 618300 221439
rect 618442 219464 618498 219473
rect 618442 219399 618498 219408
rect 618260 214600 618312 214606
rect 618260 214542 618312 214548
rect 618456 210202 618484 219399
rect 618904 214600 618956 214606
rect 618904 214542 618956 214548
rect 618916 210202 618944 214542
rect 619652 210202 619680 223858
rect 621572 223780 621624 223786
rect 621572 223722 621624 223728
rect 619916 222624 619968 222630
rect 619916 222566 619968 222572
rect 619928 214606 619956 222566
rect 620100 219768 620152 219774
rect 620100 219710 620152 219716
rect 619916 214600 619968 214606
rect 619916 214542 619968 214548
rect 620112 210202 620140 219710
rect 621110 215384 621166 215393
rect 621110 215319 621166 215328
rect 620560 214600 620612 214606
rect 620560 214542 620612 214548
rect 620572 210202 620600 214542
rect 621124 210202 621152 215319
rect 621584 210202 621612 223722
rect 622400 217320 622452 217326
rect 622400 217262 622452 217268
rect 622412 210202 622440 217262
rect 622688 210202 622716 223994
rect 623320 214736 623372 214742
rect 623320 214678 623372 214684
rect 623332 210202 623360 214678
rect 623792 210202 623820 224470
rect 623962 218104 624018 218113
rect 623962 218039 624018 218048
rect 623976 214606 624004 218039
rect 623964 214600 624016 214606
rect 623964 214542 624016 214548
rect 624424 214464 624476 214470
rect 624424 214406 624476 214412
rect 624436 210202 624464 214406
rect 625264 210202 625292 224606
rect 625436 224392 625488 224398
rect 625436 224334 625488 224340
rect 625448 214606 625476 224334
rect 628748 224188 628800 224194
rect 628748 224130 628800 224136
rect 627092 223032 627144 223038
rect 627092 222974 627144 222980
rect 625620 222760 625672 222766
rect 625620 222702 625672 222708
rect 625436 214600 625488 214606
rect 625436 214542 625488 214548
rect 625632 210202 625660 222702
rect 626632 217592 626684 217598
rect 626632 217534 626684 217540
rect 626080 214600 626132 214606
rect 626080 214542 626132 214548
rect 626092 210202 626120 214542
rect 626644 210202 626672 217534
rect 627104 210202 627132 222974
rect 627920 222488 627972 222494
rect 627920 222430 627972 222436
rect 627932 210202 627960 222430
rect 628288 217456 628340 217462
rect 628288 217398 628340 217404
rect 628300 210202 628328 217398
rect 628760 210202 628788 224130
rect 629852 222352 629904 222358
rect 629852 222294 629904 222300
rect 629392 214464 629444 214470
rect 629392 214406 629444 214412
rect 629404 210202 629432 214406
rect 629864 210202 629892 222294
rect 630048 214606 630076 229066
rect 633716 227044 633768 227050
rect 633716 226986 633768 226992
rect 630864 225004 630916 225010
rect 630864 224946 630916 224952
rect 630678 218376 630734 218385
rect 630678 218311 630734 218320
rect 630036 214600 630088 214606
rect 630036 214542 630088 214548
rect 630692 210202 630720 218311
rect 630876 210338 630904 224946
rect 632704 222896 632756 222902
rect 632704 222838 632756 222844
rect 631508 222216 631560 222222
rect 631508 222158 631560 222164
rect 630876 210310 630996 210338
rect 630968 210202 630996 210310
rect 631520 210202 631548 222158
rect 632716 213042 632744 222838
rect 633440 221876 633492 221882
rect 633440 221818 633492 221824
rect 632888 214600 632940 214606
rect 632888 214542 632940 214548
rect 632704 213036 632756 213042
rect 632704 212978 632756 212984
rect 632900 210202 632928 214542
rect 633452 210202 633480 221818
rect 633728 210202 633756 226986
rect 634360 213036 634412 213042
rect 634360 212978 634412 212984
rect 634372 210202 634400 212978
rect 635108 210202 635136 277986
rect 635568 272406 635596 278052
rect 636292 277772 636344 277778
rect 636292 277714 636344 277720
rect 635556 272400 635608 272406
rect 635556 272342 635608 272348
rect 636304 229094 636332 277714
rect 636764 275466 636792 278052
rect 637592 278038 637974 278066
rect 636752 275460 636804 275466
rect 636752 275402 636804 275408
rect 637592 269822 637620 278038
rect 637764 277908 637816 277914
rect 637764 277850 637816 277856
rect 637580 269816 637632 269822
rect 637580 269758 637632 269764
rect 637776 229094 637804 277850
rect 639156 273970 639184 278052
rect 639144 273964 639196 273970
rect 639144 273906 639196 273912
rect 640352 272678 640380 278052
rect 640536 278038 641470 278066
rect 641732 278038 642666 278066
rect 640340 272672 640392 272678
rect 640340 272614 640392 272620
rect 640536 269958 640564 278038
rect 640524 269952 640576 269958
rect 640524 269894 640576 269900
rect 641732 268394 641760 278038
rect 643848 275330 643876 278052
rect 643836 275324 643888 275330
rect 643836 275266 643888 275272
rect 645044 271318 645072 278052
rect 645872 278038 646254 278066
rect 647252 278038 647450 278066
rect 645032 271312 645084 271318
rect 645032 271254 645084 271260
rect 641720 268388 641772 268394
rect 641720 268330 641772 268336
rect 645872 261526 645900 278038
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 647252 246362 647280 278038
rect 647240 246356 647292 246362
rect 647240 246298 647292 246304
rect 648632 242214 648660 278052
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 636304 229066 636516 229094
rect 637776 229066 638172 229094
rect 636488 210202 636516 229066
rect 638144 210202 638172 229066
rect 650642 225040 650698 225049
rect 650642 224975 650698 224984
rect 648620 220244 648672 220250
rect 648620 220186 648672 220192
rect 645858 219872 645914 219881
rect 645858 219807 645914 219816
rect 644940 215960 644992 215966
rect 644940 215902 644992 215908
rect 643836 213376 643888 213382
rect 643836 213318 643888 213324
rect 641720 212696 641772 212702
rect 641720 212638 641772 212644
rect 639880 212560 639932 212566
rect 639880 212502 639932 212508
rect 639892 210202 639920 212502
rect 641732 210202 641760 212638
rect 643848 210202 643876 213318
rect 644952 210202 644980 215902
rect 645872 213926 645900 219807
rect 648434 218648 648490 218657
rect 648434 218583 648490 218592
rect 648252 216708 648304 216714
rect 648252 216650 648304 216656
rect 646320 214600 646372 214606
rect 646320 214542 646372 214548
rect 645860 213920 645912 213926
rect 645860 213862 645912 213868
rect 645492 213240 645544 213246
rect 645492 213182 645544 213188
rect 645504 210202 645532 213182
rect 646332 210202 646360 214542
rect 646504 213920 646556 213926
rect 646504 213862 646556 213868
rect 614500 210174 614836 210202
rect 614960 210174 615388 210202
rect 615696 210174 615940 210202
rect 616064 210174 616492 210202
rect 616892 210174 617044 210202
rect 617168 210174 617596 210202
rect 617812 210174 618148 210202
rect 618456 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620112 210174 620356 210202
rect 620572 210174 620908 210202
rect 621124 210174 621460 210202
rect 621584 210174 622012 210202
rect 622412 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623792 210174 624220 210202
rect 624436 210174 624772 210202
rect 625264 210174 625324 210202
rect 625632 210174 625876 210202
rect 626092 210174 626428 210202
rect 626644 210174 626980 210202
rect 627104 210174 627532 210202
rect 627932 210174 628084 210202
rect 628300 210174 628636 210202
rect 628760 210174 629188 210202
rect 629404 210174 629740 210202
rect 629864 210174 630292 210202
rect 630692 210174 630844 210202
rect 630968 210174 631396 210202
rect 631520 210174 631948 210202
rect 632900 210174 633052 210202
rect 633452 210174 633604 210202
rect 633728 210174 634156 210202
rect 634372 210174 634708 210202
rect 635108 210174 635260 210202
rect 636488 210174 636916 210202
rect 638144 210174 638572 210202
rect 639892 210174 640228 210202
rect 641732 210174 641884 210202
rect 643540 210174 643876 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646360 210202
rect 646516 210202 646544 213862
rect 648264 210202 648292 216650
rect 646516 210174 646852 210202
rect 647956 210174 648292 210202
rect 648448 210202 648476 218583
rect 648632 213926 648660 220186
rect 650656 216714 650684 224975
rect 651288 222896 651340 222902
rect 651288 222838 651340 222844
rect 651102 217288 651158 217297
rect 651102 217223 651158 217232
rect 650644 216708 650696 216714
rect 650644 216650 650696 216656
rect 648620 213920 648672 213926
rect 648620 213862 648672 213868
rect 649264 213920 649316 213926
rect 649264 213862 649316 213868
rect 649276 210202 649304 213862
rect 650460 212764 650512 212770
rect 650460 212706 650512 212712
rect 650472 210202 650500 212706
rect 648448 210174 648508 210202
rect 649276 210174 649612 210202
rect 650164 210174 650500 210202
rect 651116 210202 651144 217223
rect 651300 212770 651328 222838
rect 651470 221504 651526 221513
rect 651470 221439 651526 221448
rect 651288 212764 651340 212770
rect 651288 212706 651340 212712
rect 651484 210202 651512 221439
rect 651116 210174 651268 210202
rect 651484 210174 651820 210202
rect 600700 209902 601036 209930
rect 652036 209574 652064 282095
rect 652220 233918 652248 287026
rect 652390 280392 652446 280401
rect 652390 280327 652446 280336
rect 652208 233912 652260 233918
rect 652208 233854 652260 233860
rect 652404 226953 652432 280327
rect 652588 279449 652616 287026
rect 652574 279440 652630 279449
rect 652574 279375 652630 279384
rect 658936 268161 658964 296686
rect 660592 293865 660620 298114
rect 664444 294024 664496 294030
rect 664444 293966 664496 293972
rect 660578 293856 660634 293865
rect 660578 293791 660634 293800
rect 660304 292596 660356 292602
rect 660304 292538 660356 292544
rect 658922 268152 658978 268161
rect 658922 268087 658978 268096
rect 660316 232558 660344 292538
rect 663064 289876 663116 289882
rect 663064 289818 663116 289824
rect 663076 232694 663104 289818
rect 664456 247761 664484 293966
rect 667572 287088 667624 287094
rect 667572 287030 667624 287036
rect 667388 285728 667440 285734
rect 667388 285670 667440 285676
rect 666560 282940 666612 282946
rect 666560 282882 666612 282888
rect 664442 247752 664498 247761
rect 664442 247687 664498 247696
rect 666572 245721 666600 282882
rect 667204 280220 667256 280226
rect 667204 280162 667256 280168
rect 666558 245712 666614 245721
rect 666558 245647 666614 245656
rect 663064 232688 663116 232694
rect 663064 232630 663116 232636
rect 660304 232552 660356 232558
rect 660304 232494 660356 232500
rect 662512 231464 662564 231470
rect 662512 231406 662564 231412
rect 662328 229764 662380 229770
rect 662328 229706 662380 229712
rect 660948 229492 661000 229498
rect 660948 229434 661000 229440
rect 652390 226944 652446 226953
rect 652390 226879 652446 226888
rect 658922 226400 658978 226409
rect 658922 226335 658978 226344
rect 656162 225584 656218 225593
rect 656162 225519 656218 225528
rect 652758 225312 652814 225321
rect 652758 225247 652814 225256
rect 652772 220250 652800 225247
rect 654782 223952 654838 223961
rect 654782 223887 654838 223896
rect 653402 222864 653458 222873
rect 653402 222799 653458 222808
rect 652760 220244 652812 220250
rect 652760 220186 652812 220192
rect 653220 213852 653272 213858
rect 653220 213794 653272 213800
rect 653232 210202 653260 213794
rect 653416 213382 653444 222799
rect 654138 220416 654194 220425
rect 654138 220351 654194 220360
rect 653770 217560 653826 217569
rect 653770 217495 653826 217504
rect 653404 213376 653456 213382
rect 653404 213318 653456 213324
rect 653784 210202 653812 217495
rect 654152 212974 654180 220351
rect 654796 213858 654824 223887
rect 656176 214606 656204 225519
rect 657542 223680 657598 223689
rect 657542 223615 657598 223624
rect 656806 218920 656862 218929
rect 656806 218855 656862 218864
rect 656164 214600 656216 214606
rect 656164 214542 656216 214548
rect 654784 213852 654836 213858
rect 654784 213794 654836 213800
rect 656532 213444 656584 213450
rect 656532 213386 656584 213392
rect 654600 213172 654652 213178
rect 654600 213114 654652 213120
rect 654140 212968 654192 212974
rect 654140 212910 654192 212916
rect 654612 210202 654640 213114
rect 654784 212968 654836 212974
rect 654784 212910 654836 212916
rect 652924 210174 653260 210202
rect 653476 210174 653812 210202
rect 654580 210174 654640 210202
rect 654796 210202 654824 212910
rect 656544 210202 656572 213386
rect 656820 210202 656848 218855
rect 657556 213178 657584 223615
rect 658936 215966 658964 226335
rect 660762 221776 660818 221785
rect 660762 221711 660818 221720
rect 658924 215960 658976 215966
rect 658924 215902 658976 215908
rect 659566 215384 659622 215393
rect 659566 215319 659622 215328
rect 658188 214736 658240 214742
rect 658188 214678 658240 214684
rect 657544 213172 657596 213178
rect 657544 213114 657596 213120
rect 658200 210202 658228 214678
rect 658738 213208 658794 213217
rect 658738 213143 658794 213152
rect 658752 210202 658780 213143
rect 659580 210202 659608 215319
rect 660394 214568 660450 214577
rect 660394 214503 660450 214512
rect 660408 210202 660436 214503
rect 660776 213314 660804 221711
rect 660764 213308 660816 213314
rect 660764 213250 660816 213256
rect 660960 210202 660988 229434
rect 662142 228576 662198 228585
rect 662142 228511 662198 228520
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662156 210202 662184 228511
rect 662340 210202 662368 229706
rect 662524 229498 662552 231406
rect 665088 231192 665140 231198
rect 665088 231134 665140 231140
rect 664902 230344 664958 230353
rect 664902 230279 664958 230288
rect 662512 229492 662564 229498
rect 662512 229434 662564 229440
rect 663706 229120 663762 229129
rect 663706 229055 663762 229064
rect 663524 226364 663576 226370
rect 663524 226306 663576 226312
rect 663156 213920 663208 213926
rect 663156 213862 663208 213868
rect 663168 210202 663196 213862
rect 663536 210202 663564 226306
rect 663720 213926 663748 229055
rect 664626 215656 664682 215665
rect 664626 215591 664682 215600
rect 663708 213920 663760 213926
rect 663708 213862 663760 213868
rect 664640 213450 664668 215591
rect 664628 213444 664680 213450
rect 664628 213386 664680 213392
rect 664260 212764 664312 212770
rect 664260 212706 664312 212712
rect 664272 210202 664300 212706
rect 664916 210202 664944 230279
rect 665100 212770 665128 231134
rect 665272 230648 665324 230654
rect 665272 230590 665324 230596
rect 665284 226370 665312 230590
rect 665272 226364 665324 226370
rect 665272 226306 665324 226312
rect 666468 225072 666520 225078
rect 666468 225014 666520 225020
rect 665822 223136 665878 223145
rect 665822 223071 665878 223080
rect 665836 214742 665864 223071
rect 666480 222902 666508 225014
rect 666836 224664 666888 224670
rect 666836 224606 666888 224612
rect 666468 222896 666520 222902
rect 666468 222838 666520 222844
rect 666848 221513 666876 224606
rect 667020 223848 667072 223854
rect 667020 223790 667072 223796
rect 666834 221504 666890 221513
rect 666834 221439 666890 221448
rect 667032 220425 667060 223790
rect 667018 220416 667074 220425
rect 667018 220351 667074 220360
rect 666834 219464 666890 219473
rect 666834 219399 666890 219408
rect 666650 215928 666706 215937
rect 666650 215863 666706 215872
rect 665824 214736 665876 214742
rect 665824 214678 665876 214684
rect 665088 212764 665140 212770
rect 665088 212706 665140 212712
rect 654796 210174 655132 210202
rect 656236 210174 656572 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659548 210174 659608 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662184 210202
rect 662308 210174 662368 210202
rect 662860 210174 663196 210202
rect 663412 210174 663564 210202
rect 663964 210174 664300 210202
rect 664516 210174 664944 210202
rect 632152 209568 632204 209574
rect 652024 209568 652076 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652024 209510 652076 209516
rect 632164 209494 632500 209510
rect 666664 198529 666692 215863
rect 666650 198520 666706 198529
rect 666650 198455 666706 198464
rect 666848 175001 666876 219399
rect 667018 217968 667074 217977
rect 667018 217903 667074 217912
rect 667032 188873 667060 217903
rect 667018 188864 667074 188873
rect 667018 188799 667074 188808
rect 666834 174992 666890 175001
rect 666834 174927 666890 174936
rect 667216 132569 667244 280162
rect 667400 180305 667428 285670
rect 667584 181393 667612 287030
rect 668952 264512 669004 264518
rect 668952 264454 669004 264460
rect 668124 264376 668176 264382
rect 668124 264318 668176 264324
rect 667940 264240 667992 264246
rect 667940 264182 667992 264188
rect 667756 224460 667808 224466
rect 667756 224402 667808 224408
rect 667768 224233 667796 224402
rect 667754 224224 667810 224233
rect 667754 224159 667810 224168
rect 667756 223984 667808 223990
rect 667756 223926 667808 223932
rect 667768 223689 667796 223926
rect 667754 223680 667810 223689
rect 667754 223615 667810 223624
rect 667756 223168 667808 223174
rect 667754 223136 667756 223145
rect 667808 223136 667810 223145
rect 667754 223071 667810 223080
rect 667756 209092 667808 209098
rect 667756 209034 667808 209040
rect 667570 181384 667626 181393
rect 667570 181319 667626 181328
rect 667386 180296 667442 180305
rect 667386 180231 667442 180240
rect 667768 133113 667796 209034
rect 667952 184521 667980 264182
rect 668136 194313 668164 264318
rect 668766 232520 668822 232529
rect 668766 232455 668822 232464
rect 668400 231328 668452 231334
rect 668400 231270 668452 231276
rect 668412 199209 668440 231270
rect 668584 229900 668636 229906
rect 668584 229842 668636 229848
rect 668596 222194 668624 229842
rect 668596 222166 668716 222194
rect 668688 219434 668716 222166
rect 668596 219406 668716 219434
rect 668398 199200 668454 199209
rect 668398 199135 668454 199144
rect 668122 194304 668178 194313
rect 668122 194239 668178 194248
rect 668398 191720 668454 191729
rect 668398 191655 668454 191664
rect 667938 184512 667994 184521
rect 667938 184447 667994 184456
rect 668216 178016 668268 178022
rect 668214 177984 668216 177993
rect 668268 177984 668270 177993
rect 668214 177919 668270 177928
rect 668032 175092 668084 175098
rect 668032 175034 668084 175040
rect 668044 174729 668072 175034
rect 668030 174720 668086 174729
rect 668030 174655 668086 174664
rect 667940 169720 667992 169726
rect 667938 169688 667940 169697
rect 667992 169688 667994 169697
rect 667938 169623 667994 169632
rect 667940 165096 667992 165102
rect 667940 165038 667992 165044
rect 667952 164937 667980 165038
rect 667938 164928 667994 164937
rect 667938 164863 667994 164872
rect 668216 160064 668268 160070
rect 668214 160032 668216 160041
rect 668268 160032 668270 160041
rect 668214 159967 668270 159976
rect 668216 155576 668268 155582
rect 668216 155518 668268 155524
rect 668228 155145 668256 155518
rect 668214 155136 668270 155145
rect 668214 155071 668270 155080
rect 668412 135561 668440 191655
rect 668596 138825 668624 219406
rect 668780 163305 668808 232455
rect 668964 189417 668992 264454
rect 669226 250200 669282 250209
rect 669226 250135 669282 250144
rect 669240 247761 669268 250135
rect 669226 247752 669282 247761
rect 669226 247687 669282 247696
rect 669134 231160 669190 231169
rect 669134 231095 669190 231104
rect 669148 204105 669176 231095
rect 669274 223440 669326 223446
rect 669272 223408 669274 223417
rect 669326 223408 669328 223417
rect 669272 223343 669328 223352
rect 669424 216617 669452 347239
rect 669870 302016 669926 302025
rect 669870 301951 669926 301960
rect 669688 234660 669740 234666
rect 669688 234602 669740 234608
rect 669700 224954 669728 234602
rect 669700 224926 669820 224954
rect 669596 223644 669648 223650
rect 669596 223586 669648 223592
rect 669410 216608 669466 216617
rect 669410 216543 669466 216552
rect 669608 215665 669636 223586
rect 669594 215656 669650 215665
rect 669594 215591 669650 215600
rect 669792 215294 669820 224926
rect 669700 215266 669820 215294
rect 669410 215112 669466 215121
rect 669410 215047 669466 215056
rect 669134 204096 669190 204105
rect 669134 204031 669190 204040
rect 669424 202881 669452 215047
rect 669410 202872 669466 202881
rect 669410 202807 669466 202816
rect 669134 198792 669190 198801
rect 669134 198727 669190 198736
rect 668950 189408 669006 189417
rect 668950 189343 669006 189352
rect 668952 184884 669004 184890
rect 668952 184826 669004 184832
rect 668766 163296 668822 163305
rect 668766 163231 668822 163240
rect 668766 162480 668822 162489
rect 668766 162415 668822 162424
rect 668780 148617 668808 162415
rect 668766 148608 668822 148617
rect 668766 148543 668822 148552
rect 668768 145784 668820 145790
rect 668768 145726 668820 145732
rect 668780 145353 668808 145726
rect 668766 145344 668822 145353
rect 668766 145279 668822 145288
rect 668582 138816 668638 138825
rect 668582 138751 668638 138760
rect 668398 135552 668454 135561
rect 668398 135487 668454 135496
rect 668766 135144 668822 135153
rect 668766 135079 668822 135088
rect 667940 133816 667992 133822
rect 667938 133784 667940 133793
rect 667992 133784 667994 133793
rect 667938 133719 667994 133728
rect 667754 133104 667810 133113
rect 667754 133039 667810 133048
rect 667202 132560 667258 132569
rect 667202 132495 667258 132504
rect 668492 130824 668544 130830
rect 668492 130766 668544 130772
rect 668504 130665 668532 130766
rect 668490 130656 668546 130665
rect 668490 130591 668546 130600
rect 668032 129736 668084 129742
rect 668032 129678 668084 129684
rect 668044 129033 668072 129678
rect 668030 129024 668086 129033
rect 668030 128959 668086 128968
rect 668582 127800 668638 127809
rect 668582 127735 668638 127744
rect 667940 108860 667992 108866
rect 667940 108802 667992 108808
rect 667952 107817 667980 108802
rect 667938 107808 667994 107817
rect 667938 107743 667994 107752
rect 668400 106208 668452 106214
rect 668398 106176 668400 106185
rect 668452 106176 668454 106185
rect 668398 106111 668454 106120
rect 668596 102921 668624 127735
rect 668780 119241 668808 135079
rect 668964 125769 668992 184826
rect 669148 143721 669176 198727
rect 669502 172408 669558 172417
rect 669502 172343 669558 172352
rect 669516 166994 669544 172343
rect 669700 169726 669728 215266
rect 669688 169720 669740 169726
rect 669688 169662 669740 169668
rect 669516 166966 669636 166994
rect 669608 150385 669636 166966
rect 669594 150376 669650 150385
rect 669594 150311 669650 150320
rect 669134 143712 669190 143721
rect 669134 143647 669190 143656
rect 669884 133822 669912 301951
rect 670330 262168 670386 262177
rect 670330 262103 670386 262112
rect 670146 258496 670202 258505
rect 670146 258431 670202 258440
rect 670160 234614 670188 258431
rect 670344 236201 670372 262103
rect 670330 236192 670386 236201
rect 670330 236127 670386 236136
rect 670160 234586 670464 234614
rect 670240 234524 670292 234530
rect 670240 234466 670292 234472
rect 670252 233322 670280 234466
rect 670252 233294 670372 233322
rect 670056 233028 670108 233034
rect 670056 232970 670108 232976
rect 670068 165102 670096 232970
rect 670344 222194 670372 233294
rect 670160 222166 670372 222194
rect 670160 218498 670188 222166
rect 670160 218482 670280 218498
rect 670160 218476 670292 218482
rect 670160 218470 670240 218476
rect 670240 218418 670292 218424
rect 670436 218346 670464 234586
rect 670528 222194 670556 392527
rect 670974 295760 671030 295769
rect 670974 295695 671030 295704
rect 670988 293865 671016 295695
rect 670974 293856 671030 293865
rect 670974 293791 671030 293800
rect 671356 278730 671384 570386
rect 671988 570172 672040 570178
rect 671988 570114 672040 570120
rect 671802 559736 671858 559745
rect 671802 559671 671858 559680
rect 671620 533112 671672 533118
rect 671620 533054 671672 533060
rect 671632 489326 671660 533054
rect 671620 489320 671672 489326
rect 671620 489262 671672 489268
rect 671816 483206 671844 559671
rect 671804 483200 671856 483206
rect 671804 483142 671856 483148
rect 672000 454866 672028 570114
rect 672184 455870 672212 640306
rect 672448 629740 672500 629746
rect 672448 629682 672500 629688
rect 672460 619614 672488 629682
rect 672632 624504 672684 624510
rect 672630 624472 672632 624481
rect 672684 624472 672686 624481
rect 672630 624407 672686 624416
rect 672632 623824 672684 623830
rect 672630 623792 672632 623801
rect 672684 623792 672686 623801
rect 672630 623727 672686 623736
rect 672632 623280 672684 623286
rect 672630 623248 672632 623257
rect 672684 623248 672686 623257
rect 672630 623183 672686 623192
rect 672632 622464 672684 622470
rect 672630 622432 672632 622441
rect 672684 622432 672686 622441
rect 672630 622367 672686 622376
rect 672448 619608 672500 619614
rect 672448 619550 672500 619556
rect 672354 604480 672410 604489
rect 672354 604415 672410 604424
rect 672368 528766 672396 604415
rect 672538 597408 672594 597417
rect 672538 597343 672594 597352
rect 672356 528760 672408 528766
rect 672356 528702 672408 528708
rect 672552 528154 672580 597343
rect 672828 573753 672856 649159
rect 672998 648816 673054 648825
rect 672998 648751 673054 648760
rect 672814 573744 672870 573753
rect 672814 573679 672870 573688
rect 673012 573345 673040 648751
rect 673196 630674 673224 683086
rect 673104 630646 673224 630674
rect 673104 625002 673132 630646
rect 673288 629746 673316 696895
rect 673472 682938 673500 727246
rect 673656 717614 673684 736906
rect 673564 717586 673684 717614
rect 673564 683114 673592 717586
rect 673748 707577 673776 782614
rect 673920 780020 673972 780026
rect 673920 779962 673972 779968
rect 673932 760394 673960 779962
rect 674852 779714 674880 785182
rect 675128 784638 675418 784666
rect 675128 784310 675156 784638
rect 675116 784304 675168 784310
rect 675116 784246 675168 784252
rect 675392 784168 675444 784174
rect 675392 784110 675444 784116
rect 675404 783972 675432 784110
rect 675128 783346 675418 783374
rect 675128 782678 675156 783346
rect 675116 782672 675168 782678
rect 675116 782614 675168 782620
rect 675300 782536 675352 782542
rect 675300 782478 675352 782484
rect 675312 781402 675340 782478
rect 675312 781374 675432 781402
rect 675024 781108 675076 781114
rect 675024 781050 675076 781056
rect 675036 780994 675064 781050
rect 674944 780966 675064 780994
rect 674944 779906 674972 780966
rect 675404 780844 675432 781374
rect 675312 780422 675432 780450
rect 675312 780314 675340 780422
rect 675128 780286 675340 780314
rect 675404 780300 675432 780422
rect 675128 780026 675156 780286
rect 675116 780020 675168 780026
rect 675116 779962 675168 779968
rect 674944 779878 675248 779906
rect 675220 779714 675248 779878
rect 674852 779686 675156 779714
rect 675220 779686 675340 779714
rect 674378 779376 674434 779385
rect 674378 779311 674434 779320
rect 673840 760366 673960 760394
rect 673840 720508 673868 760366
rect 674012 735140 674064 735146
rect 674012 735082 674064 735088
rect 674024 727274 674052 735082
rect 673932 727246 674052 727274
rect 673932 724514 673960 727246
rect 674392 726646 674420 779311
rect 674562 778832 674618 778841
rect 674562 778767 674618 778776
rect 674576 726782 674604 778767
rect 674932 778388 674984 778394
rect 674932 778330 674984 778336
rect 674944 777073 674972 778330
rect 674930 777064 674986 777073
rect 674930 776999 674986 777008
rect 674930 775704 674986 775713
rect 674930 775639 674932 775648
rect 674984 775639 674986 775648
rect 674932 775610 674984 775616
rect 675128 750734 675156 779686
rect 675312 778478 675340 779686
rect 675496 779385 675524 779688
rect 675482 779376 675538 779385
rect 675482 779311 675538 779320
rect 675496 778841 675524 779008
rect 675482 778832 675538 778841
rect 675482 778767 675538 778776
rect 675312 778450 675418 778478
rect 675404 777481 675432 777852
rect 675390 777472 675446 777481
rect 675390 777407 675446 777416
rect 675482 777064 675538 777073
rect 675300 777028 675352 777034
rect 675482 776999 675538 777008
rect 675300 776970 675352 776976
rect 675312 776914 675340 776970
rect 675220 776886 675340 776914
rect 675220 775350 675248 776886
rect 675496 776628 675524 776999
rect 675404 775713 675432 776016
rect 675390 775704 675446 775713
rect 675390 775639 675446 775648
rect 675220 775322 675418 775350
rect 675404 773650 675432 774180
rect 675312 773622 675432 773650
rect 675312 773430 675340 773622
rect 675300 773424 675352 773430
rect 675300 773366 675352 773372
rect 675036 750706 675156 750734
rect 674840 738608 674892 738614
rect 674840 738550 674892 738556
rect 674852 729994 674880 738550
rect 675036 736934 675064 750706
rect 675392 746632 675444 746638
rect 675392 746574 675444 746580
rect 675404 743852 675432 746574
rect 675206 743336 675262 743345
rect 675262 743294 675418 743322
rect 675206 743271 675262 743280
rect 675404 742490 675432 742696
rect 675392 742484 675444 742490
rect 675392 742426 675444 742432
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 675220 742002 675340 742030
rect 675404 742016 675432 742070
rect 675220 741198 675248 742002
rect 675208 741192 675260 741198
rect 675208 741134 675260 741140
rect 675220 740166 675418 740194
rect 675220 738614 675248 740166
rect 675404 739158 675432 739636
rect 675392 739152 675444 739158
rect 675392 739094 675444 739100
rect 675404 738750 675432 739024
rect 675392 738744 675444 738750
rect 675392 738686 675444 738692
rect 675208 738608 675260 738614
rect 675208 738550 675260 738556
rect 675220 738330 675418 738358
rect 675220 738177 675248 738330
rect 675206 738168 675262 738177
rect 675206 738103 675262 738112
rect 674760 729966 674880 729994
rect 674944 736906 675064 736934
rect 674760 729881 674788 729966
rect 674746 729872 674802 729881
rect 674746 729807 674802 729816
rect 674944 727410 674972 736906
rect 675116 736024 675168 736030
rect 675036 735972 675116 735978
rect 675036 735966 675168 735972
rect 675036 735950 675156 735966
rect 675036 735026 675064 735950
rect 675496 735729 675524 735896
rect 675482 735720 675538 735729
rect 675482 735655 675538 735664
rect 675404 735162 675432 735319
rect 675312 735146 675432 735162
rect 675300 735140 675432 735146
rect 675352 735134 675432 735140
rect 675300 735082 675352 735088
rect 675036 734998 675340 735026
rect 675116 734596 675168 734602
rect 675116 734538 675168 734544
rect 675128 731898 675156 734538
rect 675312 733493 675340 734998
rect 675496 734369 675524 734672
rect 675482 734360 675538 734369
rect 675482 734295 675538 734304
rect 675496 733825 675524 734031
rect 675482 733816 675538 733825
rect 675482 733751 675538 733760
rect 675312 733465 675418 733493
rect 675312 732822 675418 732850
rect 675312 732766 675340 732822
rect 675300 732760 675352 732766
rect 675300 732702 675352 732708
rect 675128 731870 675432 731898
rect 675404 731612 675432 731870
rect 674852 727382 674972 727410
rect 675036 731054 675248 731082
rect 674852 727258 674880 727382
rect 675036 727274 675064 731054
rect 675220 731014 675248 731054
rect 675220 730986 675418 731014
rect 675298 730824 675354 730833
rect 675298 730759 675354 730768
rect 675312 729298 675340 730759
rect 675496 730153 675524 730351
rect 675482 730144 675538 730153
rect 675482 730079 675538 730088
rect 675300 729292 675352 729298
rect 675300 729234 675352 729240
rect 675300 729088 675352 729094
rect 675300 729030 675352 729036
rect 674840 727252 674892 727258
rect 675036 727246 675156 727274
rect 674840 727194 674892 727200
rect 674564 726776 674616 726782
rect 674564 726718 674616 726724
rect 674380 726640 674432 726646
rect 674380 726582 674432 726588
rect 673932 724486 674052 724514
rect 674024 721857 674052 724486
rect 674010 721848 674066 721857
rect 674010 721783 674066 721792
rect 675128 721721 675156 727246
rect 675312 721750 675340 729030
rect 675496 728793 675524 729164
rect 675482 728784 675538 728793
rect 675482 728719 675538 728728
rect 681004 727252 681056 727258
rect 681004 727194 681056 727200
rect 675300 721744 675352 721750
rect 675114 721712 675170 721721
rect 675300 721686 675352 721692
rect 675114 721647 675170 721656
rect 675300 721268 675352 721274
rect 675300 721210 675352 721216
rect 675312 720866 675340 721210
rect 675300 720860 675352 720866
rect 675300 720802 675352 720808
rect 675300 720520 675352 720526
rect 673840 720480 674696 720508
rect 674010 719672 674066 719681
rect 674010 719607 674066 719616
rect 674024 714854 674052 719607
rect 673932 714826 674052 714854
rect 673734 707568 673790 707577
rect 673734 707503 673790 707512
rect 673734 706344 673790 706353
rect 673734 706279 673790 706288
rect 673748 705294 673776 706279
rect 673736 705288 673788 705294
rect 673736 705230 673788 705236
rect 673734 705120 673790 705129
rect 673734 705055 673790 705064
rect 673748 703866 673776 705055
rect 673736 703860 673788 703866
rect 673736 703802 673788 703808
rect 673736 701208 673788 701214
rect 673734 701176 673736 701185
rect 673788 701176 673790 701185
rect 673734 701111 673790 701120
rect 673734 692880 673790 692889
rect 673734 692815 673736 692824
rect 673788 692815 673790 692824
rect 673736 692786 673788 692792
rect 673734 690160 673790 690169
rect 673734 690095 673736 690104
rect 673788 690095 673790 690104
rect 673736 690066 673788 690072
rect 673736 688832 673788 688838
rect 673734 688800 673736 688809
rect 673788 688800 673790 688809
rect 673734 688735 673790 688744
rect 673734 688120 673790 688129
rect 673734 688055 673790 688064
rect 673564 683086 673684 683114
rect 673426 682910 673500 682938
rect 673426 682666 673454 682910
rect 673426 682638 673500 682666
rect 673472 682417 673500 682638
rect 673458 682408 673514 682417
rect 673458 682343 673514 682352
rect 673656 682258 673684 683086
rect 673564 682230 673684 682258
rect 673564 682009 673592 682230
rect 673550 682000 673606 682009
rect 673550 681935 673606 681944
rect 673550 671392 673606 671401
rect 673550 671327 673552 671336
rect 673604 671327 673606 671336
rect 673552 671298 673604 671304
rect 673552 671152 673604 671158
rect 673552 671094 673604 671100
rect 673564 670993 673592 671094
rect 673550 670984 673606 670993
rect 673550 670919 673606 670928
rect 673550 670576 673606 670585
rect 673550 670511 673606 670520
rect 673564 670410 673592 670511
rect 673552 670404 673604 670410
rect 673552 670346 673604 670352
rect 673552 670268 673604 670274
rect 673552 670210 673604 670216
rect 673564 669769 673592 670210
rect 673550 669760 673606 669769
rect 673550 669695 673606 669704
rect 673550 668944 673606 668953
rect 673550 668879 673606 668888
rect 673564 668710 673592 668879
rect 673552 668704 673604 668710
rect 673552 668646 673604 668652
rect 673552 668568 673604 668574
rect 673550 668536 673552 668545
rect 673604 668536 673606 668545
rect 673550 668471 673606 668480
rect 673550 668128 673606 668137
rect 673550 668063 673606 668072
rect 673564 667962 673592 668063
rect 673552 667956 673604 667962
rect 673552 667898 673604 667904
rect 673550 667720 673606 667729
rect 673550 667655 673606 667664
rect 673564 667350 673592 667655
rect 673552 667344 673604 667350
rect 673552 667286 673604 667292
rect 673552 667208 673604 667214
rect 673552 667150 673604 667156
rect 673564 666913 673592 667150
rect 673550 666904 673606 666913
rect 673550 666839 673606 666848
rect 673550 666632 673606 666641
rect 673550 666567 673552 666576
rect 673604 666567 673606 666576
rect 673552 666538 673604 666544
rect 673552 665304 673604 665310
rect 673550 665272 673552 665281
rect 673604 665272 673606 665281
rect 673550 665207 673606 665216
rect 673550 664456 673606 664465
rect 673550 664391 673552 664400
rect 673604 664391 673606 664400
rect 673552 664362 673604 664368
rect 673552 663944 673604 663950
rect 673552 663886 673604 663892
rect 673564 663785 673592 663886
rect 673550 663776 673606 663785
rect 673550 663711 673606 663720
rect 673550 643512 673606 643521
rect 673550 643447 673606 643456
rect 673564 642649 673592 643447
rect 673564 642621 673684 642649
rect 673458 641744 673514 641753
rect 673458 641679 673514 641688
rect 673276 629740 673328 629746
rect 673276 629682 673328 629688
rect 673276 626136 673328 626142
rect 673274 626104 673276 626113
rect 673328 626104 673330 626113
rect 673274 626039 673330 626048
rect 673276 625456 673328 625462
rect 673274 625424 673276 625433
rect 673328 625424 673330 625433
rect 673274 625359 673330 625368
rect 673276 625184 673328 625190
rect 673274 625152 673276 625161
rect 673328 625152 673330 625161
rect 673274 625087 673330 625096
rect 673104 624974 673224 625002
rect 673196 621382 673224 624974
rect 673184 621376 673236 621382
rect 673184 621318 673236 621324
rect 673274 621208 673330 621217
rect 673274 621143 673276 621152
rect 673328 621143 673330 621152
rect 673276 621114 673328 621120
rect 673274 618216 673330 618225
rect 673274 618151 673330 618160
rect 673288 617506 673316 618151
rect 673276 617500 673328 617506
rect 673276 617442 673328 617448
rect 673274 607336 673330 607345
rect 673274 607271 673330 607280
rect 672998 573336 673054 573345
rect 672998 573271 673054 573280
rect 673090 560144 673146 560153
rect 673090 560079 673146 560088
rect 672906 555248 672962 555257
rect 672906 555183 672962 555192
rect 672724 532772 672776 532778
rect 672724 532714 672776 532720
rect 672540 528148 672592 528154
rect 672540 528090 672592 528096
rect 672736 490113 672764 532714
rect 672722 490104 672778 490113
rect 672722 490039 672778 490048
rect 672632 489932 672684 489938
rect 672632 489874 672684 489880
rect 672448 489660 672500 489666
rect 672448 489602 672500 489608
rect 672172 455864 672224 455870
rect 672172 455806 672224 455812
rect 672000 454850 672120 454866
rect 672000 454844 672132 454850
rect 672000 454838 672080 454844
rect 672080 454786 672132 454792
rect 672264 453960 672316 453966
rect 672262 453928 672264 453937
rect 672316 453928 672318 453937
rect 672262 453863 672318 453872
rect 672460 401985 672488 489602
rect 672644 402529 672672 489874
rect 672920 486033 672948 555183
rect 672906 486024 672962 486033
rect 672906 485959 672962 485968
rect 673104 484809 673132 560079
rect 673288 530097 673316 607271
rect 673472 594561 673500 641679
rect 673656 625154 673684 642621
rect 673564 625126 673684 625154
rect 673564 598934 673592 625126
rect 673748 617409 673776 688055
rect 673932 662017 673960 714826
rect 674668 707198 674696 720480
rect 675300 720462 675352 720468
rect 675312 712065 675340 720462
rect 675298 712056 675354 712065
rect 675298 711991 675354 712000
rect 681016 710841 681044 727194
rect 683396 726776 683448 726782
rect 683396 726718 683448 726724
rect 682382 726608 682438 726617
rect 682382 726543 682438 726552
rect 682396 711249 682424 726543
rect 682382 711240 682438 711249
rect 682382 711175 682438 711184
rect 681002 710832 681058 710841
rect 681002 710767 681058 710776
rect 674656 707192 674708 707198
rect 676036 707192 676088 707198
rect 674656 707134 674708 707140
rect 676034 707160 676036 707169
rect 676088 707160 676090 707169
rect 676034 707095 676090 707104
rect 683408 706761 683436 726718
rect 684040 726640 684092 726646
rect 684040 726582 684092 726588
rect 684052 707985 684080 726582
rect 684222 726336 684278 726345
rect 684222 726271 684278 726280
rect 684236 709617 684264 726271
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 684222 709608 684278 709617
rect 684222 709543 684278 709552
rect 684038 707976 684094 707985
rect 684038 707911 684094 707920
rect 683394 706752 683450 706761
rect 683394 706687 683450 706696
rect 683118 705528 683174 705537
rect 683118 705463 683174 705472
rect 674286 705392 674342 705401
rect 683132 705362 683160 705463
rect 674286 705327 674288 705336
rect 674340 705327 674342 705336
rect 683120 705356 683172 705362
rect 674288 705298 674340 705304
rect 683120 705298 683172 705304
rect 675114 701176 675170 701185
rect 675114 701111 675170 701120
rect 675128 698889 675156 701111
rect 675128 698861 675418 698889
rect 675128 698329 675418 698337
rect 675114 698320 675418 698329
rect 675170 698309 675418 698320
rect 675114 698255 675170 698264
rect 675128 697666 675418 697694
rect 675128 696969 675156 697666
rect 675114 696960 675170 696969
rect 675114 696895 675170 696904
rect 675496 696833 675524 697035
rect 675482 696824 675538 696833
rect 675482 696759 675538 696768
rect 675114 695872 675170 695881
rect 675114 695807 675170 695816
rect 675128 695209 675156 695807
rect 675128 695181 675418 695209
rect 675312 694742 675432 694770
rect 675114 694648 675170 694657
rect 675312 694634 675340 694742
rect 675170 694606 675340 694634
rect 675404 694620 675432 694742
rect 675114 694583 675170 694592
rect 674576 693994 675418 694022
rect 674288 693048 674340 693054
rect 674288 692990 674340 692996
rect 674102 689888 674158 689897
rect 674102 689823 674158 689832
rect 674116 683114 674144 689823
rect 674300 688129 674328 692990
rect 674576 692774 674604 693994
rect 675496 693138 675524 693328
rect 675404 693110 675524 693138
rect 675404 693054 675432 693110
rect 675392 693048 675444 693054
rect 675392 692990 675444 692996
rect 675114 692880 675170 692889
rect 675114 692815 675170 692824
rect 674484 692746 674604 692774
rect 674484 688378 674512 692746
rect 675128 690894 675156 692815
rect 675128 690866 675418 690894
rect 675128 690322 675340 690350
rect 674930 690160 674986 690169
rect 674930 690095 674986 690104
rect 674944 689330 674972 690095
rect 675128 689897 675156 690322
rect 675312 690282 675340 690322
rect 675404 690282 675432 690336
rect 675312 690254 675432 690282
rect 675114 689888 675170 689897
rect 675114 689823 675170 689832
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 675128 689642 675340 689670
rect 675404 689656 675432 689710
rect 675128 689489 675156 689642
rect 675114 689480 675170 689489
rect 675114 689415 675170 689424
rect 674944 689302 675064 689330
rect 674840 689036 674892 689042
rect 674840 688978 674892 688984
rect 674852 688922 674880 688978
rect 674760 688894 674880 688922
rect 675036 688922 675064 689302
rect 675220 689042 675418 689058
rect 675208 689036 675418 689042
rect 675260 689030 675418 689036
rect 675208 688978 675260 688984
rect 675036 688894 675156 688922
rect 674484 688350 674604 688378
rect 674286 688120 674342 688129
rect 674286 688055 674342 688064
rect 674576 687970 674604 688350
rect 674484 687942 674604 687970
rect 674116 683086 674236 683114
rect 673918 662008 673974 662017
rect 673918 661943 673974 661952
rect 674012 661632 674064 661638
rect 674010 661600 674012 661609
rect 674064 661600 674066 661609
rect 674010 661535 674066 661544
rect 674010 661192 674066 661201
rect 674010 661127 674012 661136
rect 674064 661127 674066 661136
rect 674012 661098 674064 661104
rect 674010 660240 674066 660249
rect 674010 660175 674012 660184
rect 674064 660175 674066 660184
rect 674012 660146 674064 660152
rect 674010 659968 674066 659977
rect 674010 659903 674066 659912
rect 674024 659734 674052 659903
rect 674012 659728 674064 659734
rect 674012 659670 674064 659676
rect 674010 655616 674066 655625
rect 674010 655551 674012 655560
rect 674064 655551 674066 655560
rect 674012 655522 674064 655528
rect 674208 654134 674236 683086
rect 674208 654106 674420 654134
rect 674194 644600 674250 644609
rect 674194 644535 674250 644544
rect 674208 640334 674236 644535
rect 674392 640334 674420 654106
rect 674024 640306 674236 640334
rect 674300 640306 674420 640334
rect 674024 625154 674052 640306
rect 674300 636886 674328 640306
rect 674484 637022 674512 687942
rect 674760 683114 674788 688894
rect 674930 688800 674986 688809
rect 674930 688735 674986 688744
rect 674944 687698 674972 688735
rect 675128 688514 675156 688894
rect 675128 688486 675340 688514
rect 675312 688378 675340 688486
rect 675404 688378 675432 688500
rect 675312 688350 675432 688378
rect 675114 687848 675170 687857
rect 675170 687806 675418 687834
rect 675114 687783 675170 687792
rect 674944 687670 675156 687698
rect 675128 686678 675156 687670
rect 675128 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675114 686216 675170 686225
rect 675114 686151 675170 686160
rect 675128 685998 675156 686151
rect 675128 685970 675418 685998
rect 674930 685808 674986 685817
rect 674930 685743 674986 685752
rect 674944 684706 674972 685743
rect 675114 685536 675170 685545
rect 675114 685471 675170 685480
rect 675128 685386 675156 685471
rect 675128 685358 675340 685386
rect 675312 685250 675340 685358
rect 675404 685250 675432 685372
rect 675312 685222 675432 685250
rect 674944 684678 675432 684706
rect 675404 684148 675432 684678
rect 675114 684040 675170 684049
rect 675114 683975 675170 683984
rect 674668 683086 674788 683114
rect 674472 637016 674524 637022
rect 674472 636958 674524 636964
rect 674288 636880 674340 636886
rect 674288 636822 674340 636828
rect 674288 625184 674340 625190
rect 673840 625126 674052 625154
rect 674286 625152 674288 625161
rect 674340 625152 674342 625161
rect 673840 619290 673868 625126
rect 674286 625087 674342 625096
rect 674012 623960 674064 623966
rect 674010 623928 674012 623937
rect 674064 623928 674066 623937
rect 674010 623863 674066 623872
rect 674288 623892 674340 623898
rect 674288 623834 674340 623840
rect 674300 623665 674328 623834
rect 674286 623656 674342 623665
rect 674286 623591 674342 623600
rect 674668 623082 674696 683086
rect 674840 682440 674892 682446
rect 674838 682408 674840 682417
rect 674892 682408 674894 682417
rect 674838 682343 674894 682352
rect 675128 676433 675156 683975
rect 675298 683768 675354 683777
rect 675298 683703 675354 683712
rect 675114 676424 675170 676433
rect 675114 676359 675170 676368
rect 674840 666664 674892 666670
rect 674838 666632 674840 666641
rect 674892 666632 674894 666641
rect 674838 666567 674894 666576
rect 675312 666505 675340 683703
rect 684130 682680 684186 682689
rect 684130 682615 684186 682624
rect 675484 682576 675536 682582
rect 675484 682518 675536 682524
rect 683212 682576 683264 682582
rect 683212 682518 683264 682524
rect 675496 682009 675524 682518
rect 675482 682000 675538 682009
rect 675482 681935 675538 681944
rect 676034 667312 676090 667321
rect 676034 667247 676090 667256
rect 676048 666670 676076 667247
rect 676036 666664 676088 666670
rect 676036 666606 676088 666612
rect 675298 666496 675354 666505
rect 675298 666431 675354 666440
rect 676034 664864 676090 664873
rect 676034 664799 676090 664808
rect 676048 663814 676076 664799
rect 674840 663808 674892 663814
rect 674838 663776 674840 663785
rect 676036 663808 676088 663814
rect 674892 663776 674894 663785
rect 683224 663785 683252 682518
rect 683488 682440 683540 682446
rect 683488 682382 683540 682388
rect 676036 663750 676088 663756
rect 683210 663776 683266 663785
rect 674838 663711 674894 663720
rect 683210 663711 683266 663720
rect 683500 662969 683528 682382
rect 684144 666233 684172 682615
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 684130 666224 684186 666233
rect 684130 666159 684186 666168
rect 683486 662960 683542 662969
rect 683486 662895 683542 662904
rect 674838 660240 674894 660249
rect 674838 660175 674894 660184
rect 674852 659870 674880 660175
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 683132 659870 683160 660039
rect 674840 659864 674892 659870
rect 674840 659806 674892 659812
rect 683120 659864 683172 659870
rect 683120 659806 683172 659812
rect 675114 655616 675170 655625
rect 675114 655551 675170 655560
rect 675128 653698 675156 655551
rect 675128 653670 675418 653698
rect 675404 652905 675432 653140
rect 675390 652896 675446 652905
rect 675390 652831 675446 652840
rect 675312 652582 675432 652610
rect 675114 652488 675170 652497
rect 675312 652474 675340 652582
rect 675170 652446 675340 652474
rect 675404 652460 675432 652582
rect 675114 652423 675170 652432
rect 674852 651834 675418 651862
rect 674852 643838 674880 651834
rect 674944 649998 675340 650026
rect 674944 644042 674972 649998
rect 675312 649994 675340 649998
rect 675404 649994 675432 650012
rect 675312 649966 675432 649994
rect 675404 649233 675432 649468
rect 675390 649224 675446 649233
rect 675390 649159 675446 649168
rect 675114 648816 675170 648825
rect 675170 648774 675418 648802
rect 675114 648751 675170 648760
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 675114 645824 675170 645833
rect 675114 645759 675170 645768
rect 675128 645674 675156 645759
rect 675128 645646 675418 645674
rect 675312 645102 675418 645130
rect 675312 644609 675340 645102
rect 675298 644600 675354 644609
rect 675298 644535 675354 644544
rect 675404 644337 675432 644475
rect 675390 644328 675446 644337
rect 675390 644263 675446 644272
rect 674944 644014 675248 644042
rect 674806 643822 674880 643838
rect 674794 643816 674880 643822
rect 674846 643810 674880 643816
rect 675220 643770 675248 644014
rect 674794 643758 674846 643764
rect 674944 643742 675248 643770
rect 675312 643810 675418 643838
rect 674944 643634 674972 643742
rect 674760 643606 674972 643634
rect 674760 639962 674788 643606
rect 675312 643521 675340 643810
rect 675574 643648 675630 643657
rect 675574 643583 675630 643592
rect 675298 643512 675354 643521
rect 675298 643447 675354 643456
rect 674932 643408 674984 643414
rect 674932 643350 674984 643356
rect 674944 640370 674972 643350
rect 675588 643280 675616 643583
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675206 641472 675262 641481
rect 675262 641430 675418 641458
rect 675206 641407 675262 641416
rect 675220 640781 675418 640809
rect 675220 640490 675248 640781
rect 675208 640484 675260 640490
rect 675208 640426 675260 640432
rect 674944 640342 675248 640370
rect 675024 640144 675076 640150
rect 675024 640086 675076 640092
rect 674760 639934 674972 639962
rect 674944 635526 674972 639934
rect 675036 637650 675064 640086
rect 675036 637622 675156 637650
rect 674932 635520 674984 635526
rect 674932 635462 674984 635468
rect 674656 623076 674708 623082
rect 674656 623018 674708 623024
rect 674288 622668 674340 622674
rect 674288 622610 674340 622616
rect 674012 622600 674064 622606
rect 674300 622554 674328 622610
rect 674064 622548 674328 622554
rect 674012 622542 674328 622548
rect 674024 622526 674328 622542
rect 674288 622464 674340 622470
rect 674286 622432 674288 622441
rect 674340 622432 674342 622441
rect 674286 622367 674342 622376
rect 674288 621444 674340 621450
rect 674288 621386 674340 621392
rect 674012 621376 674064 621382
rect 674300 621330 674328 621386
rect 674064 621324 674328 621330
rect 674012 621318 674328 621324
rect 674024 621302 674328 621318
rect 674010 621072 674066 621081
rect 674010 621007 674012 621016
rect 674064 621007 674066 621016
rect 674012 620978 674064 620984
rect 674012 620832 674064 620838
rect 674288 620832 674340 620838
rect 674064 620780 674288 620786
rect 674012 620774 674340 620780
rect 674024 620758 674328 620774
rect 674012 620288 674064 620294
rect 674064 620236 674328 620242
rect 674012 620230 674328 620236
rect 674024 620214 674328 620230
rect 674300 620158 674328 620214
rect 674288 620152 674340 620158
rect 674288 620094 674340 620100
rect 674288 619948 674340 619954
rect 674288 619890 674340 619896
rect 674300 619834 674328 619890
rect 674024 619806 674328 619834
rect 674024 619750 674052 619806
rect 674012 619744 674064 619750
rect 674012 619686 674064 619692
rect 674012 619608 674064 619614
rect 674064 619556 674328 619562
rect 674012 619550 674328 619556
rect 674024 619546 674328 619550
rect 674024 619540 674340 619546
rect 674024 619534 674288 619540
rect 674288 619482 674340 619488
rect 673840 619262 673960 619290
rect 673734 617400 673790 617409
rect 673734 617335 673790 617344
rect 673932 616978 673960 619262
rect 674288 617160 674340 617166
rect 673840 616950 673960 616978
rect 674024 617108 674288 617114
rect 674024 617102 674340 617108
rect 674024 617086 674328 617102
rect 673840 601694 673868 616950
rect 674024 616894 674052 617086
rect 674012 616888 674064 616894
rect 674012 616830 674064 616836
rect 674012 615664 674064 615670
rect 674064 615612 674328 615618
rect 674012 615606 674328 615612
rect 674024 615590 674328 615606
rect 674300 615534 674328 615590
rect 674288 615528 674340 615534
rect 674288 615470 674340 615476
rect 674010 614952 674066 614961
rect 674010 614887 674012 614896
rect 674064 614887 674066 614896
rect 674012 614858 674064 614864
rect 674012 611380 674064 611386
rect 674288 611380 674340 611386
rect 674064 611328 674288 611354
rect 675128 611354 675156 637622
rect 675220 625154 675248 640342
rect 675404 639826 675432 640152
rect 675312 639798 675432 639826
rect 675312 631394 675340 639798
rect 675496 638625 675524 638928
rect 675482 638616 675538 638625
rect 675482 638551 675538 638560
rect 681002 637528 681058 637537
rect 681002 637463 681058 637472
rect 675668 635520 675720 635526
rect 675668 635462 675720 635468
rect 675680 631417 675708 635462
rect 675482 631408 675538 631417
rect 675312 631366 675482 631394
rect 675482 631343 675538 631352
rect 675666 631408 675722 631417
rect 675666 631343 675722 631352
rect 676218 625696 676274 625705
rect 676218 625631 676274 625640
rect 676232 625190 676260 625631
rect 676220 625184 676272 625190
rect 675220 625126 675340 625154
rect 676220 625126 676272 625132
rect 675312 617137 675340 625126
rect 676218 624472 676274 624481
rect 676218 624407 676274 624416
rect 676232 623898 676260 624407
rect 676220 623892 676272 623898
rect 676220 623834 676272 623840
rect 676402 622840 676458 622849
rect 676402 622775 676458 622784
rect 676034 622704 676090 622713
rect 676034 622639 676036 622648
rect 676088 622639 676090 622648
rect 676036 622610 676088 622616
rect 676416 622470 676444 622775
rect 676404 622464 676456 622470
rect 676404 622406 676456 622412
rect 681016 622033 681044 637463
rect 683212 637016 683264 637022
rect 683212 636958 683264 636964
rect 681002 622024 681058 622033
rect 681002 621959 681058 621968
rect 676034 621480 676090 621489
rect 676034 621415 676036 621424
rect 676088 621415 676090 621424
rect 676036 621386 676088 621392
rect 676220 620832 676272 620838
rect 676218 620800 676220 620809
rect 676272 620800 676274 620809
rect 676218 620735 676274 620744
rect 676496 620152 676548 620158
rect 676496 620094 676548 620100
rect 676508 619993 676536 620094
rect 676218 619984 676274 619993
rect 676218 619919 676220 619928
rect 676272 619919 676274 619928
rect 676494 619984 676550 619993
rect 676494 619919 676550 619928
rect 676220 619890 676272 619896
rect 676218 619576 676274 619585
rect 676218 619511 676220 619520
rect 676272 619511 676274 619520
rect 676220 619482 676272 619488
rect 683224 618769 683252 636958
rect 683396 636880 683448 636886
rect 683396 636822 683448 636828
rect 683408 634814 683436 636822
rect 683408 634786 683620 634814
rect 683396 623076 683448 623082
rect 683396 623018 683448 623024
rect 683210 618760 683266 618769
rect 683210 618695 683266 618704
rect 676034 617808 676090 617817
rect 676034 617743 676090 617752
rect 676048 617166 676076 617743
rect 676036 617160 676088 617166
rect 675298 617128 675354 617137
rect 676036 617102 676088 617108
rect 675298 617063 675354 617072
rect 683408 616729 683436 623018
rect 683592 617137 683620 634786
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683578 617128 683634 617137
rect 683578 617063 683634 617072
rect 683394 616720 683450 616729
rect 683394 616655 683450 616664
rect 683120 615528 683172 615534
rect 683118 615496 683120 615505
rect 683172 615496 683174 615505
rect 683118 615431 683174 615440
rect 674012 611326 674340 611328
rect 674012 611322 674064 611326
rect 674288 611322 674340 611326
rect 674852 611326 675156 611354
rect 675392 611380 675444 611386
rect 674024 608666 674328 608682
rect 674012 608660 674340 608666
rect 674064 608654 674288 608660
rect 674012 608602 674064 608608
rect 674288 608602 674340 608608
rect 674472 603288 674524 603294
rect 674472 603230 674524 603236
rect 673748 601666 673868 601694
rect 673748 599162 673776 601666
rect 674012 600500 674064 600506
rect 674012 600442 674064 600448
rect 674024 600386 674052 600442
rect 674024 600370 674328 600386
rect 674024 600364 674340 600370
rect 674024 600358 674288 600364
rect 674288 600306 674340 600312
rect 674012 599548 674064 599554
rect 674012 599490 674064 599496
rect 674024 599434 674052 599490
rect 674024 599418 674328 599434
rect 674024 599412 674340 599418
rect 674024 599406 674288 599412
rect 674288 599354 674340 599360
rect 673748 599134 674420 599162
rect 674194 599040 674250 599049
rect 674194 598975 674250 598984
rect 673564 598906 673776 598934
rect 673458 594552 673514 594561
rect 673458 594487 673514 594496
rect 673748 594130 673776 598906
rect 673918 598632 673974 598641
rect 673918 598567 673974 598576
rect 673472 594102 673776 594130
rect 673472 586514 673500 594102
rect 673932 592034 673960 598567
rect 673748 592006 673960 592034
rect 673472 586486 673592 586514
rect 673564 581369 673592 586486
rect 673550 581360 673606 581369
rect 673550 581295 673606 581304
rect 673550 580680 673606 580689
rect 673550 580615 673606 580624
rect 673564 579698 673592 580615
rect 673552 579692 673604 579698
rect 673552 579634 673604 579640
rect 673552 574592 673604 574598
rect 673550 574560 673552 574569
rect 673604 574560 673606 574569
rect 673550 574495 673606 574504
rect 673552 574320 673604 574326
rect 673552 574262 673604 574268
rect 673564 574161 673592 574262
rect 673550 574152 673606 574161
rect 673550 574087 673606 574096
rect 673550 570480 673606 570489
rect 673550 570415 673552 570424
rect 673604 570415 673606 570424
rect 673552 570386 673604 570392
rect 673552 565888 673604 565894
rect 673550 565856 673552 565865
rect 673604 565856 673606 565865
rect 673550 565791 673606 565800
rect 673550 564496 673606 564505
rect 673550 564431 673552 564440
rect 673604 564431 673606 564440
rect 673552 564402 673604 564408
rect 673550 554840 673606 554849
rect 673550 554775 673552 554784
rect 673604 554775 673606 554784
rect 673552 554746 673604 554752
rect 673550 553208 673606 553217
rect 673550 553143 673606 553152
rect 673274 530088 673330 530097
rect 673274 530023 673330 530032
rect 673368 528148 673420 528154
rect 673368 528090 673420 528096
rect 673380 527785 673408 528090
rect 673366 527776 673422 527785
rect 673366 527711 673422 527720
rect 673366 490512 673422 490521
rect 673366 490447 673422 490456
rect 673380 489938 673408 490447
rect 673368 489932 673420 489938
rect 673368 489874 673420 489880
rect 673090 484800 673146 484809
rect 673090 484735 673146 484744
rect 673564 482361 673592 553143
rect 673748 540818 673776 592006
rect 674208 591410 674236 598975
rect 674392 592034 674420 599134
rect 673840 591382 674236 591410
rect 674300 592006 674420 592034
rect 673840 567194 673868 591382
rect 674300 588606 674328 592006
rect 674288 588600 674340 588606
rect 674288 588542 674340 588548
rect 674484 586514 674512 603230
rect 674656 599616 674708 599622
rect 674656 599558 674708 599564
rect 674300 586486 674512 586514
rect 674010 581088 674066 581097
rect 674010 581023 674012 581032
rect 674064 581023 674066 581032
rect 674012 580994 674064 581000
rect 674010 580272 674066 580281
rect 674010 580207 674066 580216
rect 674024 580038 674052 580207
rect 674012 580032 674064 580038
rect 674012 579974 674064 579980
rect 674012 579896 674064 579902
rect 674010 579864 674012 579873
rect 674064 579864 674066 579873
rect 674010 579799 674066 579808
rect 674010 579456 674066 579465
rect 674010 579391 674012 579400
rect 674064 579391 674066 579400
rect 674012 579362 674064 579368
rect 674012 579080 674064 579086
rect 674010 579048 674012 579057
rect 674064 579048 674066 579057
rect 674010 578983 674066 578992
rect 674010 578640 674066 578649
rect 674010 578575 674012 578584
rect 674064 578575 674066 578584
rect 674012 578546 674064 578552
rect 674010 578232 674066 578241
rect 674010 578167 674012 578176
rect 674064 578167 674066 578176
rect 674012 578138 674064 578144
rect 674010 577824 674066 577833
rect 674010 577759 674012 577768
rect 674064 577759 674066 577768
rect 674012 577730 674064 577736
rect 674012 577448 674064 577454
rect 674010 577416 674012 577425
rect 674064 577416 674066 577425
rect 674010 577351 674066 577360
rect 674010 577008 674066 577017
rect 674010 576943 674012 576952
rect 674064 576943 674066 576952
rect 674012 576914 674064 576920
rect 674010 574968 674066 574977
rect 674010 574903 674066 574912
rect 674024 574122 674052 574903
rect 674012 574116 674064 574122
rect 674012 574058 674064 574064
rect 674010 572520 674066 572529
rect 674010 572455 674066 572464
rect 674024 572286 674052 572455
rect 674012 572280 674064 572286
rect 674012 572222 674064 572228
rect 674010 572112 674066 572121
rect 674010 572047 674066 572056
rect 674024 571606 674052 572047
rect 674012 571600 674064 571606
rect 674012 571542 674064 571548
rect 674010 570888 674066 570897
rect 674010 570823 674066 570832
rect 674024 570178 674052 570823
rect 674012 570172 674064 570178
rect 674012 570114 674064 570120
rect 674010 569664 674066 569673
rect 674010 569599 674066 569608
rect 674024 568614 674052 569599
rect 674012 568608 674064 568614
rect 674012 568550 674064 568556
rect 673840 567166 673960 567194
rect 673932 547369 673960 567166
rect 674102 558376 674158 558385
rect 674102 558311 674158 558320
rect 673918 547360 673974 547369
rect 673918 547295 673974 547304
rect 674116 543734 674144 558311
rect 674300 543734 674328 586486
rect 674470 581360 674526 581369
rect 674470 581295 674526 581304
rect 674484 571606 674512 581295
rect 674472 571600 674524 571606
rect 674472 571542 674524 571548
rect 674470 552120 674526 552129
rect 674470 552055 674526 552064
rect 673840 543706 674144 543734
rect 674208 543706 674328 543734
rect 673840 540954 673868 543706
rect 673840 540938 673960 540954
rect 673840 540932 673972 540938
rect 673840 540926 673920 540932
rect 673920 540874 673972 540880
rect 673748 540790 673960 540818
rect 673736 540660 673788 540666
rect 673736 540602 673788 540608
rect 673748 540546 673776 540602
rect 673656 540518 673776 540546
rect 673656 518894 673684 540518
rect 673932 539050 673960 540790
rect 673748 539022 673960 539050
rect 673748 528554 673776 539022
rect 674208 538914 674236 543706
rect 673840 538886 674236 538914
rect 673840 534018 673868 538886
rect 674012 535832 674064 535838
rect 674064 535780 674328 535786
rect 674012 535774 674328 535780
rect 674024 535770 674328 535774
rect 674024 535764 674340 535770
rect 674024 535758 674288 535764
rect 674288 535706 674340 535712
rect 674288 535560 674340 535566
rect 674024 535508 674288 535514
rect 674024 535502 674340 535508
rect 674024 535498 674328 535502
rect 674012 535492 674328 535498
rect 674064 535486 674328 535492
rect 674012 535434 674064 535440
rect 674012 535016 674064 535022
rect 674064 534964 674328 534970
rect 674012 534958 674328 534964
rect 674024 534954 674328 534958
rect 674024 534948 674340 534954
rect 674024 534942 674288 534948
rect 674288 534890 674340 534896
rect 674288 534472 674340 534478
rect 674024 534420 674288 534426
rect 674024 534414 674340 534420
rect 674024 534410 674328 534414
rect 674012 534404 674328 534410
rect 674064 534398 674328 534404
rect 674012 534346 674064 534352
rect 674288 534336 674340 534342
rect 674024 534284 674288 534290
rect 674024 534278 674340 534284
rect 674024 534274 674328 534278
rect 674012 534268 674328 534274
rect 674064 534262 674328 534268
rect 674012 534210 674064 534216
rect 674024 534138 674328 534154
rect 674012 534132 674340 534138
rect 674064 534126 674288 534132
rect 674012 534074 674064 534080
rect 674288 534074 674340 534080
rect 673840 533990 674328 534018
rect 674300 533390 674328 533990
rect 674288 533384 674340 533390
rect 674288 533326 674340 533332
rect 674012 533112 674064 533118
rect 674288 533112 674340 533118
rect 674064 533060 674288 533066
rect 674012 533054 674340 533060
rect 674024 533038 674328 533054
rect 674288 532976 674340 532982
rect 674024 532924 674288 532930
rect 674024 532918 674340 532924
rect 674024 532914 674328 532918
rect 674012 532908 674328 532914
rect 674064 532902 674328 532908
rect 674012 532850 674064 532856
rect 674288 532840 674340 532846
rect 674024 532788 674288 532794
rect 674024 532782 674340 532788
rect 674024 532778 674328 532782
rect 674012 532772 674328 532778
rect 674064 532766 674328 532772
rect 674012 532714 674064 532720
rect 674024 532234 674328 532250
rect 674024 532228 674340 532234
rect 674024 532222 674288 532228
rect 674024 532166 674052 532222
rect 674288 532170 674340 532176
rect 674012 532160 674064 532166
rect 674012 532102 674064 532108
rect 674288 532092 674340 532098
rect 674024 532040 674288 532046
rect 674024 532034 674340 532040
rect 674024 532030 674328 532034
rect 674012 532024 674328 532030
rect 674064 532018 674328 532024
rect 674012 531966 674064 531972
rect 674288 531752 674340 531758
rect 674024 531700 674288 531706
rect 674024 531694 674340 531700
rect 674024 531678 674328 531694
rect 674024 531486 674052 531678
rect 674012 531480 674064 531486
rect 674012 531422 674064 531428
rect 674024 529990 674328 530006
rect 674012 529984 674340 529990
rect 674064 529978 674288 529984
rect 674012 529926 674064 529932
rect 674288 529926 674340 529932
rect 674288 529372 674340 529378
rect 674288 529314 674340 529320
rect 674300 529258 674328 529314
rect 674024 529230 674328 529258
rect 674024 529174 674052 529230
rect 674012 529168 674064 529174
rect 674012 529110 674064 529116
rect 674288 529032 674340 529038
rect 674024 528980 674288 528986
rect 674024 528974 674340 528980
rect 674024 528970 674328 528974
rect 674012 528964 674328 528970
rect 674064 528958 674328 528964
rect 674012 528906 674064 528912
rect 674024 528766 674328 528782
rect 674012 528760 674340 528766
rect 674064 528754 674288 528760
rect 674012 528702 674064 528708
rect 674288 528702 674340 528708
rect 673748 528526 674328 528554
rect 674300 526386 674328 528526
rect 674288 526380 674340 526386
rect 674288 526322 674340 526328
rect 674012 525088 674064 525094
rect 674012 525030 674064 525036
rect 674024 524600 674052 525030
rect 674288 524612 674340 524618
rect 674024 524572 674288 524600
rect 674288 524554 674340 524560
rect 673656 518866 674144 518894
rect 674116 499574 674144 518866
rect 674116 499546 674328 499574
rect 674300 495038 674328 499546
rect 674288 495032 674340 495038
rect 674288 494974 674340 494980
rect 673826 492144 673882 492153
rect 673826 492079 673882 492088
rect 673840 491502 673868 492079
rect 674288 491700 674340 491706
rect 674288 491642 674340 491648
rect 674012 491632 674064 491638
rect 674300 491586 674328 491642
rect 674064 491580 674328 491586
rect 674012 491574 674328 491580
rect 674024 491558 674328 491574
rect 673828 491496 673880 491502
rect 673828 491438 673880 491444
rect 674012 491360 674064 491366
rect 674010 491328 674012 491337
rect 674064 491328 674066 491337
rect 674010 491263 674066 491272
rect 674012 490952 674064 490958
rect 674010 490920 674012 490929
rect 674064 490920 674066 490929
rect 674010 490855 674066 490864
rect 674010 489696 674066 489705
rect 674010 489631 674012 489640
rect 674064 489631 674066 489640
rect 674012 489602 674064 489608
rect 674012 489320 674064 489326
rect 674010 489288 674012 489297
rect 674064 489288 674066 489297
rect 674010 489223 674066 489232
rect 674012 488504 674064 488510
rect 674010 488472 674012 488481
rect 674064 488472 674066 488481
rect 674010 488407 674066 488416
rect 674288 486804 674340 486810
rect 674288 486746 674340 486752
rect 674300 486690 674328 486746
rect 674024 486662 674328 486690
rect 674024 485858 674052 486662
rect 674012 485852 674064 485858
rect 674012 485794 674064 485800
rect 674288 485172 674340 485178
rect 674288 485114 674340 485120
rect 674300 485058 674328 485114
rect 674024 485030 674328 485058
rect 674024 484430 674052 485030
rect 674012 484424 674064 484430
rect 674012 484366 674064 484372
rect 674484 484022 674512 552055
rect 674668 526794 674696 599558
rect 674852 590646 674880 611326
rect 675392 611322 675444 611328
rect 675404 608668 675432 611322
rect 675116 608660 675168 608666
rect 675116 608602 675168 608608
rect 675128 606846 675156 608602
rect 675312 608110 675418 608138
rect 675312 607345 675340 608110
rect 675482 607744 675538 607753
rect 675482 607679 675538 607688
rect 675496 607479 675524 607679
rect 675298 607336 675354 607345
rect 675298 607271 675354 607280
rect 675128 606818 675418 606846
rect 674944 604982 675418 605010
rect 674944 592770 674972 604982
rect 675114 604480 675170 604489
rect 675170 604438 675418 604466
rect 675114 604415 675170 604424
rect 675312 603894 675432 603922
rect 675312 603786 675340 603894
rect 675128 603758 675340 603786
rect 675404 603772 675432 603894
rect 675128 603294 675156 603758
rect 675116 603288 675168 603294
rect 675116 603230 675168 603236
rect 675128 603146 675418 603174
rect 675128 602993 675156 603146
rect 675114 602984 675170 602993
rect 675114 602919 675170 602928
rect 675390 600944 675446 600953
rect 675390 600879 675446 600888
rect 675404 600644 675432 600879
rect 675116 600364 675168 600370
rect 675116 600306 675168 600312
rect 675128 598278 675156 600306
rect 675312 600222 675432 600250
rect 675312 599622 675340 600222
rect 675404 600100 675432 600222
rect 675300 599616 675352 599622
rect 675300 599558 675352 599564
rect 675300 599412 675352 599418
rect 675300 599354 675352 599360
rect 675312 598466 675340 599354
rect 675496 599049 675524 599488
rect 675482 599040 675538 599049
rect 675482 598975 675538 598984
rect 675496 598641 675524 598808
rect 675482 598632 675538 598641
rect 675482 598567 675538 598576
rect 675300 598460 675352 598466
rect 675300 598402 675352 598408
rect 675128 598250 675418 598278
rect 675300 598188 675352 598194
rect 675300 598130 675352 598136
rect 675312 596442 675340 598130
rect 675496 597417 675524 597652
rect 675482 597408 675538 597417
rect 675482 597343 675538 597352
rect 675312 596414 675418 596442
rect 675404 595377 675432 595816
rect 675390 595368 675446 595377
rect 675390 595303 675446 595312
rect 675220 595122 675418 595150
rect 675220 594833 675248 595122
rect 675206 594824 675262 594833
rect 675206 594759 675262 594768
rect 675206 594552 675262 594561
rect 675206 594487 675262 594496
rect 675220 593314 675248 594487
rect 675404 593473 675432 593980
rect 675390 593464 675446 593473
rect 675390 593399 675446 593408
rect 675220 593286 675340 593314
rect 674944 592742 675156 592770
rect 674840 590640 674892 590646
rect 674840 590582 674892 590588
rect 674930 590472 674986 590481
rect 674930 590407 674986 590416
rect 674944 589274 674972 590407
rect 674944 589246 675064 589274
rect 674840 570512 674892 570518
rect 674838 570480 674840 570489
rect 674892 570480 674894 570489
rect 674838 570415 674894 570424
rect 675036 567194 675064 589246
rect 675128 586514 675156 592742
rect 675312 592686 675340 593286
rect 675482 593192 675538 593201
rect 675482 593127 675538 593136
rect 675300 592680 675352 592686
rect 675300 592622 675352 592628
rect 675128 586486 675248 586514
rect 675220 586265 675248 586486
rect 675206 586256 675262 586265
rect 675206 586191 675262 586200
rect 675496 570518 675524 593127
rect 683396 592680 683448 592686
rect 683396 592622 683448 592628
rect 681002 591696 681058 591705
rect 681002 591631 681058 591640
rect 681016 575657 681044 591631
rect 682384 590640 682436 590646
rect 682384 590582 682436 590588
rect 682396 576473 682424 590582
rect 682382 576464 682438 576473
rect 682382 576399 682438 576408
rect 681002 575648 681058 575657
rect 681002 575583 681058 575592
rect 683408 573209 683436 592622
rect 684222 591288 684278 591297
rect 684222 591223 684278 591232
rect 684040 588600 684092 588606
rect 684040 588542 684092 588548
rect 683394 573200 683450 573209
rect 683394 573135 683450 573144
rect 684052 571985 684080 588542
rect 684236 576065 684264 591223
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 684222 576056 684278 576065
rect 684222 575991 684278 576000
rect 684038 571976 684094 571985
rect 684038 571911 684094 571920
rect 676220 571600 676272 571606
rect 676218 571568 676220 571577
rect 676272 571568 676274 571577
rect 676218 571503 676274 571512
rect 675484 570512 675536 570518
rect 675484 570454 675536 570460
rect 683120 570512 683172 570518
rect 683120 570454 683172 570460
rect 683132 570353 683160 570454
rect 683118 570344 683174 570353
rect 683118 570279 683174 570288
rect 674944 567166 675064 567194
rect 674944 554933 674972 567166
rect 675390 565856 675446 565865
rect 675390 565791 675446 565800
rect 675114 564496 675170 564505
rect 675114 564431 675170 564440
rect 675128 562918 675156 564431
rect 675404 563448 675432 565791
rect 675312 562958 675432 562986
rect 675312 562918 675340 562958
rect 675128 562890 675340 562918
rect 675404 562904 675432 562958
rect 675114 562320 675170 562329
rect 675170 562278 675418 562306
rect 675114 562255 675170 562264
rect 675390 561912 675446 561921
rect 675390 561847 675446 561856
rect 675404 561612 675432 561847
rect 674760 554905 674972 554933
rect 675128 559830 675432 559858
rect 674760 554690 674788 554905
rect 674760 554662 674880 554690
rect 674852 545902 674880 554662
rect 675128 553432 675156 559830
rect 675404 559776 675432 559830
rect 675298 559736 675354 559745
rect 675298 559671 675354 559680
rect 675312 557954 675340 559671
rect 675482 559464 675538 559473
rect 675482 559399 675538 559408
rect 675496 559232 675524 559399
rect 675496 558385 675524 558620
rect 675482 558376 675538 558385
rect 675482 558311 675538 558320
rect 675312 557926 675418 557954
rect 675298 557560 675354 557569
rect 675298 557495 675354 557504
rect 675312 556186 675340 557495
rect 675220 556158 675340 556186
rect 675220 554933 675248 556158
rect 675404 555257 675432 555492
rect 675390 555248 675446 555257
rect 675390 555183 675446 555192
rect 675220 554905 675418 554933
rect 675298 554840 675354 554849
rect 675298 554775 675354 554784
rect 675128 553404 675248 553432
rect 675220 551818 675248 553404
rect 675312 553093 675340 554775
rect 675772 553897 675800 554268
rect 675758 553888 675814 553897
rect 675758 553823 675814 553832
rect 675588 553489 675616 553656
rect 675574 553480 675630 553489
rect 675574 553415 675630 553424
rect 675312 553065 675418 553093
rect 675404 552129 675432 552432
rect 675390 552120 675446 552129
rect 675390 552055 675446 552064
rect 675208 551812 675260 551818
rect 675208 551754 675260 551760
rect 675208 551608 675260 551614
rect 675208 551550 675260 551556
rect 675390 551576 675446 551585
rect 675220 550202 675248 551550
rect 675390 551511 675446 551520
rect 675404 551239 675432 551511
rect 675036 550174 675248 550202
rect 675312 550582 675418 550610
rect 675036 549114 675064 550174
rect 675312 549506 675340 550582
rect 675496 549681 675524 549951
rect 675482 549672 675538 549681
rect 675482 549607 675538 549616
rect 675300 549500 675352 549506
rect 675300 549442 675352 549448
rect 675036 549086 675248 549114
rect 675024 548820 675076 548826
rect 675024 548762 675076 548768
rect 675036 545986 675064 548762
rect 675036 545958 675156 545986
rect 674840 545896 674892 545902
rect 674840 545838 674892 545844
rect 674930 545728 674986 545737
rect 674930 545663 674986 545672
rect 674656 526788 674708 526794
rect 674656 526730 674708 526736
rect 674944 500954 674972 545663
rect 675128 503674 675156 545958
rect 675220 540974 675248 549086
rect 675772 548321 675800 548760
rect 675758 548312 675814 548321
rect 675758 548247 675814 548256
rect 677414 547632 677470 547641
rect 677414 547567 677470 547576
rect 675574 547360 675630 547369
rect 675574 547295 675630 547304
rect 675588 547194 675616 547295
rect 675576 547188 675628 547194
rect 675576 547130 675628 547136
rect 675220 540946 675340 540974
rect 675116 503668 675168 503674
rect 675116 503610 675168 503616
rect 675312 503538 675340 540946
rect 676218 535936 676274 535945
rect 676218 535871 676274 535880
rect 676036 535764 676088 535770
rect 676034 535732 676036 535741
rect 676088 535732 676090 535741
rect 676034 535667 676090 535676
rect 676232 535566 676260 535871
rect 676220 535560 676272 535566
rect 676220 535502 676272 535508
rect 676218 535120 676274 535129
rect 676218 535055 676274 535064
rect 676036 534948 676088 534954
rect 676034 534916 676036 534925
rect 676088 534916 676090 534925
rect 676034 534851 676090 534860
rect 676034 534508 676090 534517
rect 676034 534443 676036 534452
rect 676088 534443 676090 534452
rect 676036 534414 676088 534420
rect 676232 534342 676260 535055
rect 676220 534336 676272 534342
rect 676220 534278 676272 534284
rect 676036 534132 676088 534138
rect 676034 534100 676036 534109
rect 676088 534100 676090 534109
rect 676034 534035 676090 534044
rect 676402 533488 676458 533497
rect 676402 533423 676458 533432
rect 676034 533284 676090 533293
rect 676034 533219 676090 533228
rect 676048 532982 676076 533219
rect 676220 533112 676272 533118
rect 676218 533080 676220 533089
rect 676272 533080 676274 533089
rect 676218 533015 676274 533024
rect 676036 532976 676088 532982
rect 676036 532918 676088 532924
rect 676416 532846 676444 533423
rect 676404 532840 676456 532846
rect 676404 532782 676456 532788
rect 676218 532264 676274 532273
rect 676218 532199 676274 532208
rect 676404 532228 676456 532234
rect 676232 532098 676260 532199
rect 676404 532170 676456 532176
rect 676220 532092 676272 532098
rect 676034 532060 676090 532069
rect 676220 532034 676272 532040
rect 676034 531995 676090 532004
rect 676048 531758 676076 531995
rect 676416 531865 676444 532170
rect 676402 531856 676458 531865
rect 676402 531791 676458 531800
rect 676036 531752 676088 531758
rect 676036 531694 676088 531700
rect 676034 530020 676090 530029
rect 676034 529955 676036 529964
rect 676088 529955 676090 529964
rect 676036 529926 676088 529932
rect 676218 529408 676274 529417
rect 676218 529343 676220 529352
rect 676272 529343 676274 529352
rect 676220 529314 676272 529320
rect 676220 529032 676272 529038
rect 676218 529000 676220 529009
rect 676272 529000 676274 529009
rect 676218 528935 676274 528944
rect 676034 528796 676090 528805
rect 676034 528731 676036 528740
rect 676088 528731 676090 528740
rect 676036 528702 676088 528708
rect 676036 526788 676088 526794
rect 676034 526756 676036 526765
rect 676088 526756 676090 526765
rect 676034 526691 676090 526700
rect 676036 526380 676088 526386
rect 676034 526348 676036 526357
rect 676088 526348 676090 526357
rect 676034 526283 676090 526292
rect 675484 520260 675536 520266
rect 675484 520202 675536 520208
rect 675300 503532 675352 503538
rect 675300 503474 675352 503480
rect 674932 500948 674984 500954
rect 674932 500890 674984 500896
rect 674656 495032 674708 495038
rect 674656 494974 674708 494980
rect 674668 484401 674696 494974
rect 674654 484392 674710 484401
rect 674654 484327 674710 484336
rect 674472 484016 674524 484022
rect 674472 483958 674524 483964
rect 674012 483200 674064 483206
rect 674010 483168 674012 483177
rect 674064 483168 674066 483177
rect 674010 483103 674066 483112
rect 673550 482352 673606 482361
rect 673550 482287 673606 482296
rect 674024 480418 674328 480434
rect 674012 480412 674340 480418
rect 674064 480406 674288 480412
rect 674012 480354 674064 480360
rect 674288 480354 674340 480360
rect 673274 455424 673330 455433
rect 673274 455359 673276 455368
rect 673328 455359 673330 455368
rect 673276 455330 673328 455336
rect 673386 455288 673442 455297
rect 673386 455223 673388 455232
rect 673440 455223 673442 455232
rect 673506 455252 673558 455258
rect 673388 455194 673440 455200
rect 673506 455194 673558 455200
rect 673274 455152 673330 455161
rect 673518 455138 673546 455194
rect 673330 455110 673546 455138
rect 673274 455087 673330 455096
rect 674288 454912 674340 454918
rect 672814 454880 672870 454889
rect 672814 454815 672870 454824
rect 674286 454880 674288 454889
rect 674340 454880 674342 454889
rect 674286 454815 674342 454824
rect 672828 454510 672856 454815
rect 675496 454646 675524 520202
rect 675668 518832 675720 518838
rect 675668 518774 675720 518780
rect 673046 454640 673098 454646
rect 673044 454608 673046 454617
rect 674288 454640 674340 454646
rect 673098 454608 673100 454617
rect 673044 454543 673100 454552
rect 674286 454608 674288 454617
rect 675484 454640 675536 454646
rect 674340 454608 674342 454617
rect 675484 454582 675536 454588
rect 674286 454543 674342 454552
rect 672816 454504 672868 454510
rect 672816 454446 672868 454452
rect 675680 454374 675708 518774
rect 676034 491736 676090 491745
rect 676034 491671 676036 491680
rect 676088 491671 676090 491680
rect 676036 491642 676088 491648
rect 676034 486840 676090 486849
rect 676034 486775 676036 486784
rect 676088 486775 676090 486784
rect 676036 486746 676088 486752
rect 676034 485208 676090 485217
rect 676034 485143 676036 485152
rect 676088 485143 676090 485152
rect 676036 485114 676088 485120
rect 676036 484016 676088 484022
rect 676034 483984 676036 483993
rect 676088 483984 676090 483993
rect 676034 483919 676090 483928
rect 677428 483002 677456 547567
rect 683212 547188 683264 547194
rect 683212 547130 683264 547136
rect 681002 546816 681058 546825
rect 681002 546751 681058 546760
rect 681016 530641 681044 546751
rect 682384 545896 682436 545902
rect 682384 545838 682436 545844
rect 682396 531457 682424 545838
rect 682382 531448 682438 531457
rect 682382 531383 682438 531392
rect 681002 530632 681058 530641
rect 681002 530567 681058 530576
rect 683224 527785 683252 547130
rect 683394 547088 683450 547097
rect 683394 547023 683450 547032
rect 683210 527776 683266 527785
rect 683210 527711 683266 527720
rect 683408 527377 683436 547023
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683580 533384 683632 533390
rect 683580 533326 683632 533332
rect 683592 528601 683620 533326
rect 683578 528592 683634 528601
rect 683578 528527 683634 528536
rect 683394 527368 683450 527377
rect 683394 527303 683450 527312
rect 677874 525736 677930 525745
rect 677874 525671 677930 525680
rect 677888 518838 677916 525671
rect 683118 524920 683174 524929
rect 683118 524855 683174 524864
rect 683132 524618 683160 524855
rect 683120 524612 683172 524618
rect 683120 524554 683172 524560
rect 678978 524512 679034 524521
rect 678978 524447 679034 524456
rect 678992 520266 679020 524447
rect 678980 520260 679032 520266
rect 678980 520202 679032 520208
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683394 503704 683450 503713
rect 679624 503668 679676 503674
rect 683394 503639 683450 503648
rect 679624 503610 679676 503616
rect 679636 487257 679664 503610
rect 681004 503532 681056 503538
rect 681004 503474 681056 503480
rect 679622 487248 679678 487257
rect 679622 487183 679678 487192
rect 681016 486441 681044 503474
rect 683210 500984 683266 500993
rect 681188 500948 681240 500954
rect 683210 500919 683266 500928
rect 681188 500890 681240 500896
rect 681200 487665 681228 500890
rect 681186 487656 681242 487665
rect 681186 487591 681242 487600
rect 681002 486432 681058 486441
rect 681002 486367 681058 486376
rect 683224 483585 683252 500919
rect 683408 485625 683436 503639
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683394 485616 683450 485625
rect 683394 485551 683450 485560
rect 683210 483576 683266 483585
rect 683210 483511 683266 483520
rect 676220 482996 676272 483002
rect 676220 482938 676272 482944
rect 677416 482996 677468 483002
rect 677416 482938 677468 482944
rect 676034 482760 676090 482769
rect 676232 482746 676260 482938
rect 676090 482718 676260 482746
rect 676034 482695 676090 482704
rect 680358 481944 680414 481953
rect 680358 481879 680414 481888
rect 675850 480720 675906 480729
rect 675850 480655 675906 480664
rect 675864 454918 675892 480655
rect 680372 476134 680400 481879
rect 683118 481128 683174 481137
rect 683118 481063 683174 481072
rect 683132 480418 683160 481063
rect 683120 480412 683172 480418
rect 683120 480354 683172 480360
rect 676036 476128 676088 476134
rect 676036 476070 676088 476076
rect 680360 476128 680412 476134
rect 680360 476070 680412 476076
rect 675852 454912 675904 454918
rect 675852 454854 675904 454860
rect 672954 454368 673006 454374
rect 672952 454336 672954 454345
rect 674288 454368 674340 454374
rect 673006 454336 673008 454345
rect 672952 454271 673008 454280
rect 674286 454336 674288 454345
rect 675668 454368 675720 454374
rect 674340 454336 674342 454345
rect 675668 454310 675720 454316
rect 674286 454271 674342 454280
rect 676048 453966 676076 476070
rect 674288 453960 674340 453966
rect 674286 453928 674288 453937
rect 676036 453960 676088 453966
rect 674340 453928 674342 453937
rect 676036 453902 676088 453908
rect 674286 453863 674342 453872
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 676218 403336 676274 403345
rect 674564 403300 674616 403306
rect 676218 403271 676220 403280
rect 674564 403242 674616 403248
rect 676272 403271 676274 403280
rect 676220 403242 676272 403248
rect 672630 402520 672686 402529
rect 672630 402455 672686 402464
rect 672446 401976 672502 401985
rect 672446 401911 672502 401920
rect 673182 401704 673238 401713
rect 673182 401639 673238 401648
rect 672814 399664 672870 399673
rect 672814 399599 672870 399608
rect 672630 393952 672686 393961
rect 672630 393887 672686 393896
rect 671894 393680 671950 393689
rect 671894 393615 671950 393624
rect 671710 348936 671766 348945
rect 671710 348871 671766 348880
rect 671724 331265 671752 348871
rect 671710 331256 671766 331265
rect 671710 331191 671766 331200
rect 671526 302288 671582 302297
rect 671526 302223 671582 302232
rect 671344 278724 671396 278730
rect 671344 278666 671396 278672
rect 671540 263594 671568 302223
rect 671710 278624 671766 278633
rect 671710 278559 671712 278568
rect 671764 278559 671766 278568
rect 671712 278530 671764 278536
rect 671710 263800 671766 263809
rect 671710 263735 671766 263744
rect 671724 263594 671752 263735
rect 671908 263594 671936 393615
rect 672644 376281 672672 393887
rect 672630 376272 672686 376281
rect 672630 376207 672686 376216
rect 672354 357096 672410 357105
rect 672354 357031 672410 357040
rect 672170 350160 672226 350169
rect 672170 350095 672226 350104
rect 672184 335889 672212 350095
rect 672170 335880 672226 335889
rect 672170 335815 672226 335824
rect 672368 312497 672396 357031
rect 672538 356280 672594 356289
rect 672538 356215 672594 356224
rect 672354 312488 672410 312497
rect 672354 312423 672410 312432
rect 672552 311681 672580 356215
rect 672828 355065 672856 399599
rect 672998 395040 673054 395049
rect 672998 394975 673054 394984
rect 673012 381041 673040 394975
rect 672998 381032 673054 381041
rect 672998 380967 673054 380976
rect 673196 357513 673224 401639
rect 673918 401432 673974 401441
rect 673918 401367 673974 401376
rect 673366 400480 673422 400489
rect 673366 400415 673422 400424
rect 673182 357504 673238 357513
rect 673182 357439 673238 357448
rect 673380 355881 673408 400415
rect 673734 395720 673790 395729
rect 673734 395655 673790 395664
rect 673748 375465 673776 395655
rect 673734 375456 673790 375465
rect 673734 375391 673790 375400
rect 673932 356561 673960 401367
rect 674576 396681 674604 403242
rect 676586 402928 676642 402937
rect 676586 402863 676642 402872
rect 674838 402248 674894 402257
rect 674838 402183 674894 402192
rect 674852 401713 674880 402183
rect 674838 401704 674894 401713
rect 674838 401639 674894 401648
rect 676600 400897 676628 402863
rect 676586 400888 676642 400897
rect 676586 400823 676642 400832
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 676048 398886 676076 399327
rect 674932 398880 674984 398886
rect 674932 398822 674984 398828
rect 676036 398880 676088 398886
rect 676036 398822 676088 398828
rect 674746 397352 674802 397361
rect 674746 397287 674802 397296
rect 674562 396672 674618 396681
rect 674562 396607 674618 396616
rect 674564 396092 674616 396098
rect 674564 396034 674616 396040
rect 674380 394324 674432 394330
rect 674380 394266 674432 394272
rect 674392 393938 674420 394266
rect 674208 393910 674420 393938
rect 674208 380746 674236 393910
rect 674576 393314 674604 396034
rect 674760 393314 674788 397287
rect 674944 393314 674972 398822
rect 679622 398440 679678 398449
rect 679622 398375 679678 398384
rect 676218 398032 676274 398041
rect 676218 397967 676274 397976
rect 676034 396128 676090 396137
rect 676034 396063 676036 396072
rect 676088 396063 676090 396072
rect 676036 396034 676088 396040
rect 676232 395758 676260 397967
rect 678242 397624 678298 397633
rect 678242 397559 678298 397568
rect 675208 395752 675260 395758
rect 675208 395694 675260 395700
rect 676220 395752 676272 395758
rect 676220 395694 676272 395700
rect 674392 393286 674604 393314
rect 674668 393286 674788 393314
rect 674852 393286 674972 393314
rect 674392 382226 674420 393286
rect 674380 382220 674432 382226
rect 674380 382162 674432 382168
rect 674208 380718 674420 380746
rect 674392 378146 674420 380718
rect 674380 378140 674432 378146
rect 674380 378082 674432 378088
rect 674668 371566 674696 393286
rect 674852 384810 674880 393286
rect 675220 386458 675248 395694
rect 676218 394360 676274 394369
rect 676218 394295 676220 394304
rect 676272 394295 676274 394304
rect 676220 394266 676272 394272
rect 678256 387705 678284 397559
rect 678242 387696 678298 387705
rect 678242 387631 678298 387640
rect 679636 386782 679664 398375
rect 679624 386776 679676 386782
rect 679624 386718 679676 386724
rect 675036 386430 675248 386458
rect 674840 384804 674892 384810
rect 674840 384746 674892 384752
rect 675036 384690 675064 386430
rect 674944 384662 675064 384690
rect 675128 386261 675418 386289
rect 674944 382582 674972 384662
rect 675128 382945 675156 386261
rect 675484 386028 675536 386034
rect 675484 385970 675536 385976
rect 675496 385696 675524 385970
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675392 384804 675444 384810
rect 675392 384746 675444 384752
rect 675404 384435 675432 384746
rect 675114 382936 675170 382945
rect 675114 382871 675170 382880
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 674944 382554 675340 382582
rect 675404 382568 675432 382622
rect 675758 382256 675814 382265
rect 675116 382220 675168 382226
rect 675758 382191 675814 382200
rect 675116 382162 675168 382168
rect 675128 381426 675156 382162
rect 675772 382024 675800 382191
rect 675128 381398 675418 381426
rect 675390 381032 675446 381041
rect 675390 380967 675446 380976
rect 675404 380732 675432 380967
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675116 378140 675168 378146
rect 675116 378082 675168 378088
rect 675128 377754 675156 378082
rect 675128 377726 675340 377754
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675114 375456 675170 375465
rect 675114 375391 675170 375400
rect 675128 375238 675156 375391
rect 675128 375210 675418 375238
rect 675758 373688 675814 373697
rect 675758 373623 675814 373632
rect 675772 373388 675800 373623
rect 675404 372473 675432 372776
rect 675390 372464 675446 372473
rect 675390 372399 675446 372408
rect 674668 371538 675418 371566
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 674470 358320 674526 358329
rect 674470 358255 674526 358264
rect 673918 356552 673974 356561
rect 673918 356487 673974 356496
rect 673366 355872 673422 355881
rect 673366 355807 673422 355816
rect 673274 355464 673330 355473
rect 673274 355399 673330 355408
rect 672814 355056 672870 355065
rect 672814 354991 672870 355000
rect 673090 353424 673146 353433
rect 673090 353359 673146 353368
rect 672906 349752 672962 349761
rect 672906 349687 672962 349696
rect 672722 348528 672778 348537
rect 672722 348463 672778 348472
rect 672538 311672 672594 311681
rect 672538 311607 672594 311616
rect 672538 305552 672594 305561
rect 672538 305487 672594 305496
rect 672172 288448 672224 288454
rect 672172 288390 672224 288396
rect 671540 263566 671660 263594
rect 671724 263566 671844 263594
rect 671908 263566 672028 263594
rect 671632 260834 671660 263566
rect 671448 260806 671660 260834
rect 671250 259584 671306 259593
rect 671250 259519 671306 259528
rect 670698 257272 670754 257281
rect 670698 257207 670754 257216
rect 670712 224954 670740 257207
rect 671264 251174 671292 259519
rect 671448 251174 671476 260806
rect 671618 256320 671674 256329
rect 671618 256255 671674 256264
rect 671172 251146 671292 251174
rect 671356 251146 671476 251174
rect 671172 245585 671200 251146
rect 671158 245576 671214 245585
rect 671158 245511 671214 245520
rect 671356 245426 671384 251146
rect 671632 246022 671660 256255
rect 671816 251174 671844 263566
rect 671816 251146 671936 251174
rect 671908 249794 671936 251146
rect 671816 249766 671936 249794
rect 671620 246016 671672 246022
rect 671620 245958 671672 245964
rect 671356 245398 671568 245426
rect 671252 236904 671304 236910
rect 671252 236846 671304 236852
rect 671068 235952 671120 235958
rect 671068 235894 671120 235900
rect 670884 233912 670936 233918
rect 670882 233880 670884 233889
rect 670936 233880 670938 233889
rect 670882 233815 670938 233824
rect 670884 232892 670936 232898
rect 670884 232834 670936 232840
rect 670712 224926 670832 224954
rect 670528 222166 670648 222194
rect 670424 218340 670476 218346
rect 670424 218282 670476 218288
rect 670620 218249 670648 222166
rect 670606 218240 670662 218249
rect 670606 218175 670662 218184
rect 670608 218068 670660 218074
rect 670608 218010 670660 218016
rect 670424 217796 670476 217802
rect 670424 217738 670476 217744
rect 670240 217388 670292 217394
rect 670240 217330 670292 217336
rect 670252 212534 670280 217330
rect 670436 216594 670464 217738
rect 670620 217394 670648 218010
rect 670608 217388 670660 217394
rect 670608 217330 670660 217336
rect 670160 212506 670280 212534
rect 670344 216566 670464 216594
rect 670160 186314 670188 212506
rect 670344 186314 670372 216566
rect 670514 216472 670570 216481
rect 670514 216407 670570 216416
rect 670528 198257 670556 216407
rect 670804 215294 670832 224926
rect 670712 215266 670832 215294
rect 670514 198248 670570 198257
rect 670514 198183 670570 198192
rect 670160 186286 670280 186314
rect 670344 186286 670464 186314
rect 670056 165096 670108 165102
rect 670056 165038 670108 165044
rect 670252 157334 670280 186286
rect 670436 175098 670464 186286
rect 670712 184890 670740 215266
rect 670896 186314 670924 232834
rect 670896 186286 671016 186314
rect 670700 184884 670752 184890
rect 670700 184826 670752 184832
rect 670792 178016 670844 178022
rect 670790 177984 670792 177993
rect 670844 177984 670846 177993
rect 670790 177919 670846 177928
rect 670988 176654 671016 186286
rect 670896 176626 671016 176654
rect 670424 175092 670476 175098
rect 670424 175034 670476 175040
rect 670422 171184 670478 171193
rect 670422 171119 670478 171128
rect 670160 157306 670280 157334
rect 669872 133816 669924 133822
rect 669872 133758 669924 133764
rect 669962 130928 670018 130937
rect 669962 130863 670018 130872
rect 668950 125760 669006 125769
rect 668950 125695 669006 125704
rect 668766 119232 668822 119241
rect 668766 119167 668822 119176
rect 668950 118824 669006 118833
rect 668950 118759 669006 118768
rect 668768 116884 668820 116890
rect 668768 116826 668820 116832
rect 668780 112713 668808 116826
rect 668964 114345 668992 118759
rect 668950 114336 669006 114345
rect 668950 114271 669006 114280
rect 668766 112704 668822 112713
rect 668766 112639 668822 112648
rect 669976 108866 670004 130863
rect 670160 129742 670188 157306
rect 670436 155961 670464 171119
rect 670606 170368 670662 170377
rect 670606 170303 670662 170312
rect 670422 155952 670478 155961
rect 670422 155887 670478 155896
rect 670620 147665 670648 170303
rect 670896 166994 670924 176626
rect 670804 166966 670924 166994
rect 670804 160070 670832 166966
rect 670792 160064 670844 160070
rect 670792 160006 670844 160012
rect 671080 157334 671108 235894
rect 671264 186314 671292 236846
rect 671540 234614 671568 245398
rect 671816 245392 671844 249766
rect 671632 245364 671844 245392
rect 671632 240122 671660 245364
rect 671632 240094 671752 240122
rect 671724 238649 671752 240094
rect 671710 238640 671766 238649
rect 671710 238575 671766 238584
rect 671712 236564 671764 236570
rect 671712 236506 671764 236512
rect 671540 234586 671660 234614
rect 671436 234252 671488 234258
rect 671436 234194 671488 234200
rect 671448 224954 671476 234194
rect 671356 224926 671476 224954
rect 671356 215294 671384 224926
rect 671632 224210 671660 234586
rect 671608 224182 671660 224210
rect 671724 224210 671752 236506
rect 672000 234614 672028 263566
rect 672184 246265 672212 288390
rect 672552 285569 672580 305487
rect 672538 285560 672594 285569
rect 672538 285495 672594 285504
rect 672356 284368 672408 284374
rect 672356 284310 672408 284316
rect 672170 246256 672226 246265
rect 672170 246191 672226 246200
rect 672172 246016 672224 246022
rect 672172 245958 672224 245964
rect 672184 240281 672212 245958
rect 672170 240272 672226 240281
rect 672170 240207 672226 240216
rect 672172 237040 672224 237046
rect 672172 236982 672224 236988
rect 672184 236230 672212 236982
rect 672172 236224 672224 236230
rect 672172 236166 672224 236172
rect 671908 234586 672028 234614
rect 671908 231985 671936 234586
rect 672080 233300 672132 233306
rect 672080 233242 672132 233248
rect 671894 231976 671950 231985
rect 671894 231911 671950 231920
rect 672092 226930 672120 233242
rect 672368 227089 672396 284310
rect 672736 282914 672764 348463
rect 672920 335617 672948 349687
rect 673104 340785 673132 353359
rect 673090 340776 673146 340785
rect 673090 340711 673146 340720
rect 672906 335608 672962 335617
rect 672906 335543 672962 335552
rect 672906 325000 672962 325009
rect 672906 324935 672962 324944
rect 672644 282886 672764 282914
rect 672644 273254 672672 282886
rect 672920 278633 672948 324935
rect 673288 310865 673316 355399
rect 673734 352608 673790 352617
rect 673734 352543 673790 352552
rect 673550 349344 673606 349353
rect 673550 349279 673606 349288
rect 673564 332761 673592 349279
rect 673748 333985 673776 352543
rect 673918 352200 673974 352209
rect 673918 352135 673974 352144
rect 673734 333976 673790 333985
rect 673734 333911 673790 333920
rect 673550 332752 673606 332761
rect 673550 332687 673606 332696
rect 673932 326913 673960 352135
rect 674286 351384 674342 351393
rect 674286 351319 674342 351328
rect 674300 338065 674328 351319
rect 674484 351121 674512 358255
rect 675942 357912 675998 357921
rect 675942 357847 675998 357856
rect 675956 356833 675984 357847
rect 675942 356824 675998 356833
rect 675942 356759 675998 356768
rect 674654 354648 674710 354657
rect 674654 354583 674710 354592
rect 674470 351112 674526 351121
rect 674470 351047 674526 351056
rect 674470 350568 674526 350577
rect 674470 350503 674526 350512
rect 674286 338056 674342 338065
rect 674286 337991 674342 338000
rect 674484 331090 674512 350503
rect 674472 331084 674524 331090
rect 674472 331026 674524 331032
rect 673918 326904 673974 326913
rect 673918 326839 673974 326848
rect 674380 312044 674432 312050
rect 674380 311986 674432 311992
rect 673918 311264 673974 311273
rect 673918 311199 673974 311208
rect 673274 310856 673330 310865
rect 673274 310791 673330 310800
rect 673366 309496 673422 309505
rect 673366 309431 673422 309440
rect 673182 304328 673238 304337
rect 673182 304263 673238 304272
rect 673196 287881 673224 304263
rect 673182 287872 673238 287881
rect 673182 287807 673238 287816
rect 672906 278624 672962 278633
rect 672906 278559 672962 278568
rect 672644 273226 672764 273254
rect 672538 265296 672594 265305
rect 672538 265231 672594 265240
rect 672354 227080 672410 227089
rect 672354 227015 672410 227024
rect 672552 226930 672580 265231
rect 672736 234614 672764 273226
rect 673182 266112 673238 266121
rect 673182 266047 673238 266056
rect 673196 263594 673224 266047
rect 673380 265033 673408 309431
rect 673550 305960 673606 305969
rect 673550 305895 673606 305904
rect 673564 291553 673592 305895
rect 673932 302234 673960 311199
rect 673932 302206 674144 302234
rect 673826 291816 673882 291825
rect 673826 291751 673882 291760
rect 673550 291544 673606 291553
rect 673550 291479 673606 291488
rect 673642 287600 673698 287609
rect 673642 287535 673698 287544
rect 673366 265024 673422 265033
rect 673366 264959 673422 264968
rect 673458 264480 673514 264489
rect 673458 264415 673514 264424
rect 673472 263594 673500 264415
rect 673656 263594 673684 287535
rect 673840 268161 673868 291751
rect 673826 268152 673882 268161
rect 673826 268087 673882 268096
rect 674116 266665 674144 302206
rect 674392 267481 674420 311986
rect 674668 310049 674696 354583
rect 676034 350976 676090 350985
rect 676034 350911 676090 350920
rect 676048 346633 676076 350911
rect 676034 346624 676090 346633
rect 676034 346559 676090 346568
rect 674944 341074 675418 341102
rect 674944 338745 674972 341074
rect 675114 340776 675170 340785
rect 675114 340711 675170 340720
rect 675128 340558 675156 340711
rect 675128 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340232 675814 340241
rect 675758 340167 675814 340176
rect 675772 339864 675800 340167
rect 675482 339416 675538 339425
rect 675482 339351 675538 339360
rect 675496 339252 675524 339351
rect 674930 338736 674986 338745
rect 674930 338671 674986 338680
rect 675114 338056 675170 338065
rect 675114 337991 675170 338000
rect 675128 336857 675156 337991
rect 675758 337920 675814 337929
rect 675758 337855 675814 337864
rect 675772 337416 675800 337855
rect 675128 336829 675418 336857
rect 675758 336560 675814 336569
rect 675758 336495 675814 336504
rect 675772 336192 675800 336495
rect 674930 335880 674986 335889
rect 674930 335815 674986 335824
rect 674944 331889 674972 335815
rect 675114 335608 675170 335617
rect 675170 335566 675340 335594
rect 675114 335543 675170 335552
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 675312 335430 675432 335458
rect 675114 333976 675170 333985
rect 675114 333911 675170 333920
rect 675128 333078 675156 333911
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 674944 331861 675418 331889
rect 675114 331256 675170 331265
rect 675170 331214 675418 331242
rect 675114 331191 675170 331200
rect 675116 331084 675168 331090
rect 675116 331026 675168 331032
rect 675128 330049 675156 331026
rect 675128 330021 675418 330049
rect 675312 328222 675432 328250
rect 675312 328182 675340 328222
rect 675220 328154 675340 328182
rect 675404 328168 675432 328222
rect 675022 327992 675078 328001
rect 675022 327927 675078 327936
rect 675036 325009 675064 327927
rect 675220 325689 675248 328154
rect 675390 327992 675446 328001
rect 675390 327927 675446 327936
rect 675404 327556 675432 327927
rect 675390 326904 675446 326913
rect 675390 326839 675446 326848
rect 675404 326332 675432 326839
rect 675206 325680 675262 325689
rect 675206 325615 675262 325624
rect 675022 325000 675078 325009
rect 675022 324935 675078 324944
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676218 313984 676274 313993
rect 676218 313919 676274 313928
rect 674838 312896 674894 312905
rect 674838 312831 674894 312840
rect 674852 311953 674880 312831
rect 675482 312080 675538 312089
rect 675482 312015 675484 312024
rect 675536 312015 675538 312024
rect 675484 311986 675536 311992
rect 674838 311944 674894 311953
rect 674838 311879 674894 311888
rect 675482 310448 675538 310457
rect 675482 310383 675538 310392
rect 674654 310040 674710 310049
rect 674654 309975 674710 309984
rect 675496 309874 675524 310383
rect 674748 309868 674800 309874
rect 674748 309810 674800 309816
rect 675484 309868 675536 309874
rect 675484 309810 675536 309816
rect 674760 309134 674788 309810
rect 675942 309768 675998 309777
rect 676232 309754 676260 313919
rect 675998 309726 676260 309754
rect 675942 309703 675998 309712
rect 674484 309106 674788 309134
rect 674484 292618 674512 309106
rect 675114 308408 675170 308417
rect 675114 308343 675170 308352
rect 674930 308000 674986 308009
rect 674930 307935 674986 307944
rect 674654 303920 674710 303929
rect 674654 303855 674710 303864
rect 674668 299554 674696 303855
rect 674576 299526 674696 299554
rect 674576 297514 674604 299526
rect 674748 297832 674800 297838
rect 674800 297780 674880 297786
rect 674748 297774 674880 297780
rect 674760 297758 674880 297774
rect 674576 297486 674788 297514
rect 674484 292590 674696 292618
rect 674378 267472 674434 267481
rect 674378 267407 674434 267416
rect 674286 267064 674342 267073
rect 674286 266999 674342 267008
rect 674102 266656 674158 266665
rect 674102 266591 674158 266600
rect 674300 263594 674328 266999
rect 674668 265849 674696 292590
rect 674760 286226 674788 297486
rect 674852 288062 674880 297758
rect 674944 292414 674972 307935
rect 675128 299474 675156 308343
rect 676034 307592 676090 307601
rect 676090 307550 676444 307578
rect 676034 307527 676090 307536
rect 676034 307184 676090 307193
rect 676090 307142 676260 307170
rect 676034 307119 676090 307128
rect 676232 306406 676260 307142
rect 676220 306400 676272 306406
rect 676220 306342 676272 306348
rect 676416 304910 676444 307550
rect 678242 306776 678298 306785
rect 678242 306711 678298 306720
rect 676864 306400 676916 306406
rect 676864 306342 676916 306348
rect 675852 304904 675904 304910
rect 675852 304846 675904 304852
rect 676404 304904 676456 304910
rect 676404 304846 676456 304852
rect 675864 302234 675892 304846
rect 676586 304736 676642 304745
rect 676586 304671 676642 304680
rect 676034 303512 676090 303521
rect 676034 303447 676090 303456
rect 675496 302206 675892 302234
rect 675128 299446 675248 299474
rect 675220 297378 675248 299446
rect 675496 297838 675524 302206
rect 676048 302025 676076 303447
rect 676034 302016 676090 302025
rect 676034 301951 676090 301960
rect 676600 301617 676628 304671
rect 676586 301608 676642 301617
rect 676586 301543 676642 301552
rect 675484 297832 675536 297838
rect 675484 297774 675536 297780
rect 676036 297628 676088 297634
rect 676036 297570 676088 297576
rect 675852 297492 675904 297498
rect 675852 297434 675904 297440
rect 675864 297378 675892 297434
rect 675128 297350 675248 297378
rect 675312 297350 675892 297378
rect 675128 295542 675156 297350
rect 675312 296206 675340 297350
rect 676048 296585 676076 297570
rect 676876 297401 676904 306342
rect 678256 297498 678284 306711
rect 678978 306368 679034 306377
rect 678978 306303 679034 306312
rect 678992 297634 679020 306303
rect 678980 297628 679032 297634
rect 678980 297570 679032 297576
rect 678244 297492 678296 297498
rect 678244 297434 678296 297440
rect 676862 297392 676918 297401
rect 676862 297327 676918 297336
rect 676034 296576 676090 296585
rect 676034 296511 676090 296520
rect 675300 296200 675352 296206
rect 675300 296142 675352 296148
rect 675588 295769 675616 296072
rect 675574 295760 675630 295769
rect 675574 295695 675630 295704
rect 675128 295514 675418 295542
rect 675300 295452 675352 295458
rect 675300 295394 675352 295400
rect 675312 295066 675340 295394
rect 675312 295038 675432 295066
rect 675404 294879 675432 295038
rect 675758 294672 675814 294681
rect 675758 294607 675814 294616
rect 675772 294236 675800 294607
rect 674944 292386 675418 292414
rect 675574 292224 675630 292233
rect 675574 292159 675630 292168
rect 675588 291856 675616 292159
rect 675390 291544 675446 291553
rect 675390 291479 675446 291488
rect 675404 291176 675432 291479
rect 675758 291000 675814 291009
rect 675758 290935 675814 290944
rect 675772 290564 675800 290935
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674852 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675312 286334 675432 286362
rect 675312 286226 675340 286334
rect 674760 286198 675340 286226
rect 675404 286212 675432 286334
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675758 282704 675814 282713
rect 675758 282639 675814 282648
rect 675772 282554 675800 282639
rect 675312 282540 675800 282554
rect 675312 282526 675786 282540
rect 674838 278352 674894 278361
rect 674838 278287 674894 278296
rect 674852 273873 674880 278287
rect 675312 277409 675340 282526
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 676862 279440 676918 279449
rect 676862 279375 676918 279384
rect 675482 278080 675538 278089
rect 675482 278015 675538 278024
rect 675298 277400 675354 277409
rect 675298 277335 675354 277344
rect 674838 273864 674894 273873
rect 674838 273799 674894 273808
rect 674654 265840 674710 265849
rect 674654 265775 674710 265784
rect 675114 264752 675170 264761
rect 675114 264687 675170 264696
rect 673196 263566 673316 263594
rect 673472 263566 673592 263594
rect 673656 263566 673776 263594
rect 674300 263566 674420 263594
rect 673090 263392 673146 263401
rect 673090 263327 673146 263336
rect 672906 259312 672962 259321
rect 672906 259247 672962 259256
rect 672920 242729 672948 259247
rect 673104 250753 673132 263327
rect 673090 250744 673146 250753
rect 673090 250679 673146 250688
rect 673090 249656 673146 249665
rect 673090 249591 673146 249600
rect 673104 245313 673132 249591
rect 673090 245304 673146 245313
rect 673090 245239 673146 245248
rect 672906 242720 672962 242729
rect 672906 242655 672962 242664
rect 673288 241641 673316 263566
rect 673564 241913 673592 263566
rect 673748 246265 673776 263566
rect 674194 260944 674250 260953
rect 673840 260902 674194 260930
rect 673840 250050 673868 260902
rect 674194 260879 674250 260888
rect 674392 260250 674420 263566
rect 674654 262576 674710 262585
rect 674654 262511 674710 262520
rect 674024 260222 674420 260250
rect 673840 250022 673960 250050
rect 673734 246256 673790 246265
rect 673734 246191 673790 246200
rect 673932 246106 673960 250022
rect 673840 246078 673960 246106
rect 673840 245857 673868 246078
rect 673826 245848 673882 245857
rect 673826 245783 673882 245792
rect 674024 244274 674052 260222
rect 674194 260128 674250 260137
rect 674194 260063 674250 260072
rect 674208 253934 674236 260063
rect 674378 258904 674434 258913
rect 674378 258839 674434 258848
rect 674208 253906 674328 253934
rect 674300 244274 674328 253906
rect 673932 244246 674052 244274
rect 674208 244246 674328 244274
rect 674392 244274 674420 258839
rect 674392 244246 674512 244274
rect 673550 241904 673606 241913
rect 673550 241839 673606 241848
rect 673274 241632 673330 241641
rect 673274 241567 673330 241576
rect 672954 236768 673006 236774
rect 672952 236736 672954 236745
rect 673006 236736 673008 236745
rect 672952 236671 673008 236680
rect 673184 236496 673236 236502
rect 673236 236444 673868 236450
rect 673184 236438 673868 236444
rect 673196 236422 673868 236438
rect 673092 236224 673144 236230
rect 673144 236172 673776 236178
rect 673092 236166 673776 236172
rect 673104 236150 673776 236166
rect 673414 235884 673466 235890
rect 673414 235826 673466 235832
rect 673426 235770 673454 235826
rect 672908 235748 672960 235754
rect 673426 235742 673684 235770
rect 672908 235690 672960 235696
rect 672920 234614 672948 235690
rect 673368 235000 673420 235006
rect 672644 234586 672764 234614
rect 672828 234586 672948 234614
rect 673012 234948 673368 234954
rect 673012 234942 673420 234948
rect 673012 234926 673408 234942
rect 672644 231854 672672 234586
rect 672828 232914 672856 234586
rect 673012 233034 673040 234926
rect 673184 234864 673236 234870
rect 673184 234806 673236 234812
rect 673460 234864 673512 234870
rect 673460 234806 673512 234812
rect 673196 233306 673224 234806
rect 673184 233300 673236 233306
rect 673184 233242 673236 233248
rect 673472 233238 673500 234806
rect 673460 233232 673512 233238
rect 673460 233174 673512 233180
rect 673656 233050 673684 235742
rect 673000 233028 673052 233034
rect 673000 232970 673052 232976
rect 673564 233022 673684 233050
rect 672828 232898 672948 232914
rect 672828 232892 672960 232898
rect 672828 232886 672908 232892
rect 672908 232834 672960 232840
rect 673564 232529 673592 233022
rect 673550 232520 673606 232529
rect 673550 232455 673606 232464
rect 672644 231826 672764 231854
rect 672736 229906 672764 231826
rect 673184 230988 673236 230994
rect 673184 230930 673236 230936
rect 672724 229900 672776 229906
rect 672724 229842 672776 229848
rect 673196 229770 673224 230930
rect 673460 230240 673512 230246
rect 673460 230182 673512 230188
rect 673184 229764 673236 229770
rect 673184 229706 673236 229712
rect 672816 229628 672868 229634
rect 672816 229570 672868 229576
rect 672828 227202 672856 229570
rect 673276 229424 673328 229430
rect 673276 229366 673328 229372
rect 672828 227174 672948 227202
rect 672092 226902 672304 226930
rect 672460 226914 672580 226930
rect 671896 225684 671948 225690
rect 671896 225626 671948 225632
rect 671908 225049 671936 225626
rect 672156 225344 672208 225350
rect 672032 225312 672088 225321
rect 672156 225286 672208 225292
rect 672032 225247 672034 225256
rect 672086 225247 672088 225256
rect 672034 225218 672086 225224
rect 672168 225185 672196 225286
rect 672154 225176 672210 225185
rect 672154 225111 672210 225120
rect 671894 225040 671950 225049
rect 671894 224975 671950 224984
rect 671820 224800 671872 224806
rect 671818 224768 671820 224777
rect 671872 224768 671874 224777
rect 671818 224703 671874 224712
rect 671724 224182 671844 224210
rect 671482 224120 671534 224126
rect 671480 224088 671482 224097
rect 671534 224088 671536 224097
rect 671480 224023 671536 224032
rect 671608 223938 671636 224182
rect 671540 223910 671636 223938
rect 671356 215266 671476 215294
rect 671448 190454 671476 215266
rect 671172 186286 671292 186314
rect 671356 190426 671476 190454
rect 671172 176654 671200 186286
rect 671356 177993 671384 190426
rect 671342 177984 671398 177993
rect 671342 177919 671398 177928
rect 671172 176626 671292 176654
rect 670988 157306 671108 157334
rect 670988 155666 671016 157306
rect 670804 155638 671016 155666
rect 670804 155582 670832 155638
rect 670792 155576 670844 155582
rect 670792 155518 670844 155524
rect 671264 151814 671292 176626
rect 670804 151786 671292 151814
rect 670606 147656 670662 147665
rect 670606 147591 670662 147600
rect 670804 145790 670832 151786
rect 670792 145784 670844 145790
rect 670792 145726 670844 145732
rect 671540 138014 671568 223910
rect 671816 215294 671844 224182
rect 672078 224088 672134 224097
rect 672078 224023 672134 224032
rect 672092 217569 672120 224023
rect 672078 217560 672134 217569
rect 672078 217495 672134 217504
rect 672078 216200 672134 216209
rect 672078 216135 672134 216144
rect 672092 215665 672120 216135
rect 672078 215656 672134 215665
rect 672078 215591 672134 215600
rect 671724 215266 671844 215294
rect 671724 150113 671752 215266
rect 672078 214160 672134 214169
rect 672078 214095 672134 214104
rect 672092 199753 672120 214095
rect 672078 199744 672134 199753
rect 672078 199679 672134 199688
rect 672276 176654 672304 226902
rect 672448 226908 672580 226914
rect 672500 226902 672580 226908
rect 672448 226850 672500 226856
rect 672724 226432 672776 226438
rect 672722 226400 672724 226409
rect 672776 226400 672778 226409
rect 672722 226335 672778 226344
rect 672604 226160 672656 226166
rect 672602 226128 672604 226137
rect 672656 226128 672658 226137
rect 672602 226063 672658 226072
rect 672492 225992 672548 226001
rect 672492 225927 672494 225936
rect 672546 225927 672548 225936
rect 672494 225898 672546 225904
rect 672380 225752 672432 225758
rect 672378 225720 672380 225729
rect 672432 225720 672434 225729
rect 672378 225655 672434 225664
rect 672446 220280 672502 220289
rect 672446 220215 672502 220224
rect 672460 215294 672488 220215
rect 672630 217968 672686 217977
rect 672630 217903 672686 217912
rect 672644 215294 672672 217903
rect 672920 215294 672948 227174
rect 673288 227089 673316 229366
rect 673472 228585 673500 230182
rect 673458 228576 673514 228585
rect 673458 228511 673514 228520
rect 673552 228404 673604 228410
rect 673552 228346 673604 228352
rect 673274 227080 673330 227089
rect 673274 227015 673330 227024
rect 673092 226908 673144 226914
rect 673092 226850 673144 226856
rect 673104 220697 673132 226850
rect 673564 226817 673592 228346
rect 673550 226808 673606 226817
rect 673550 226743 673606 226752
rect 673276 226568 673328 226574
rect 673276 226510 673328 226516
rect 673288 222873 673316 226510
rect 673748 224954 673776 236150
rect 673656 224926 673776 224954
rect 673458 224768 673514 224777
rect 673458 224703 673514 224712
rect 673274 222864 673330 222873
rect 673274 222799 673330 222808
rect 673274 221096 673330 221105
rect 673274 221031 673330 221040
rect 673090 220688 673146 220697
rect 673090 220623 673146 220632
rect 673090 217424 673146 217433
rect 673090 217359 673146 217368
rect 673104 216481 673132 217359
rect 673090 216472 673146 216481
rect 673090 216407 673146 216416
rect 673090 216200 673146 216209
rect 673090 216135 673146 216144
rect 673104 215294 673132 216135
rect 672368 215266 672488 215294
rect 672552 215266 672672 215294
rect 672736 215266 672948 215294
rect 673012 215266 673132 215294
rect 672368 190454 672396 215266
rect 672552 213217 672580 215266
rect 672736 213625 672764 215266
rect 672722 213616 672778 213625
rect 672722 213551 672778 213560
rect 672814 213344 672870 213353
rect 672814 213279 672870 213288
rect 672538 213208 672594 213217
rect 672538 213143 672594 213152
rect 672630 212120 672686 212129
rect 672630 212055 672686 212064
rect 672368 190426 672488 190454
rect 672184 176626 672304 176654
rect 671986 172000 672042 172009
rect 671986 171935 672042 171944
rect 671710 150104 671766 150113
rect 671710 150039 671766 150048
rect 672000 144945 672028 171935
rect 672184 168065 672212 176626
rect 672460 175681 672488 190426
rect 672446 175672 672502 175681
rect 672446 175607 672502 175616
rect 672354 168328 672410 168337
rect 672354 168263 672410 168272
rect 672170 168056 672226 168065
rect 672170 167991 672226 168000
rect 672368 167634 672396 168263
rect 672184 167606 672396 167634
rect 671986 144936 672042 144945
rect 671986 144871 672042 144880
rect 670804 137986 671568 138014
rect 670804 130830 670832 137986
rect 672184 135153 672212 167606
rect 672354 166968 672410 166977
rect 672354 166903 672410 166912
rect 672170 135144 672226 135153
rect 672170 135079 672226 135088
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670792 130824 670844 130830
rect 670792 130766 670844 130772
rect 670148 129736 670200 129742
rect 670148 129678 670200 129684
rect 670606 122496 670662 122505
rect 670606 122431 670662 122440
rect 670620 116890 670648 122431
rect 670608 116884 670660 116890
rect 670608 116826 670660 116832
rect 671356 109034 671384 131679
rect 671526 129296 671582 129305
rect 671526 129231 671582 129240
rect 671540 109034 671568 129231
rect 672078 123312 672134 123321
rect 672078 123247 672134 123256
rect 672092 118833 672120 123247
rect 672078 118824 672134 118833
rect 672078 118759 672134 118768
rect 672368 115841 672396 166903
rect 672644 120873 672672 212055
rect 672828 124137 672856 213279
rect 673012 201385 673040 215266
rect 672998 201376 673054 201385
rect 672998 201311 673054 201320
rect 672998 200832 673054 200841
rect 672998 200767 673054 200776
rect 673012 190454 673040 200767
rect 673288 197985 673316 221031
rect 673472 216889 673500 224703
rect 673458 216880 673514 216889
rect 673458 216815 673514 216824
rect 673458 216608 673514 216617
rect 673458 216543 673514 216552
rect 673472 215393 673500 216543
rect 673458 215384 673514 215393
rect 673458 215319 673514 215328
rect 673274 197976 673330 197985
rect 673274 197911 673330 197920
rect 673012 190426 673132 190454
rect 673104 181529 673132 190426
rect 673090 181520 673146 181529
rect 673090 181455 673146 181464
rect 673366 176896 673422 176905
rect 673366 176831 673422 176840
rect 672998 169144 673054 169153
rect 672998 169079 673054 169088
rect 673012 168858 673040 169079
rect 672920 168830 673040 168858
rect 672920 157334 672948 168830
rect 673090 168736 673146 168745
rect 673090 168671 673146 168680
rect 673104 166994 673132 168671
rect 673012 166966 673132 166994
rect 673012 164234 673040 166966
rect 673380 164234 673408 176831
rect 673656 176654 673684 224926
rect 673840 215294 673868 236422
rect 673932 233322 673960 244246
rect 674208 242185 674236 244246
rect 674194 242176 674250 242185
rect 674194 242111 674250 242120
rect 674484 241097 674512 244246
rect 674668 243545 674696 262511
rect 674838 260536 674894 260545
rect 674838 260471 674894 260480
rect 674852 256329 674880 260471
rect 674838 256320 674894 256329
rect 674838 256255 674894 256264
rect 674838 254960 674894 254969
rect 674838 254895 674894 254904
rect 674852 249762 674880 254895
rect 675128 253934 675156 264687
rect 675496 258097 675524 278015
rect 676876 268569 676904 279375
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 676862 268560 676918 268569
rect 676862 268495 676918 268504
rect 676218 268152 676274 268161
rect 676218 268087 676274 268096
rect 676232 267753 676260 268087
rect 676218 267744 676274 267753
rect 676218 267679 676274 267688
rect 676402 264072 676458 264081
rect 676402 264007 676458 264016
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 259570 676260 262783
rect 675680 259542 676260 259570
rect 675482 258088 675538 258097
rect 675482 258023 675538 258032
rect 675036 253906 675156 253934
rect 674840 249756 674892 249762
rect 674840 249698 674892 249704
rect 675036 248962 675064 253906
rect 675680 251410 675708 259542
rect 676416 258738 676444 264007
rect 675852 258732 675904 258738
rect 675852 258674 675904 258680
rect 676404 258732 676456 258738
rect 676404 258674 676456 258680
rect 675864 254969 675892 258674
rect 675850 254960 675906 254969
rect 675850 254895 675906 254904
rect 674760 248934 675064 248962
rect 675128 251382 675708 251410
rect 674760 246213 674788 248934
rect 675128 248418 675156 251382
rect 675312 251110 675432 251138
rect 675312 250209 675340 251110
rect 675404 251056 675432 251110
rect 675482 250744 675538 250753
rect 675482 250679 675538 250688
rect 675496 250512 675524 250679
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675298 250200 675354 250209
rect 675298 250135 675354 250144
rect 675482 250064 675538 250073
rect 675036 248390 675156 248418
rect 675220 250022 675482 250050
rect 675036 247994 675064 248390
rect 675024 247988 675076 247994
rect 675024 247930 675076 247936
rect 675220 247874 675248 250022
rect 675482 249999 675538 250008
rect 675772 249900 675800 250271
rect 675484 249756 675536 249762
rect 675484 249698 675536 249704
rect 675496 249220 675524 249698
rect 675036 247846 675248 247874
rect 675392 247852 675444 247858
rect 675036 246378 675064 247846
rect 675392 247794 675444 247800
rect 675404 247384 675432 247794
rect 675772 246673 675800 246840
rect 675758 246664 675814 246673
rect 675758 246599 675814 246608
rect 675036 246350 675156 246378
rect 674760 246185 674880 246213
rect 674852 245410 674880 246185
rect 675128 245970 675156 246350
rect 675036 245942 675156 245970
rect 675220 246185 675418 246213
rect 674840 245404 674892 245410
rect 674840 245346 674892 245352
rect 675036 245290 675064 245942
rect 675220 245857 675248 246185
rect 675206 245848 675262 245857
rect 675206 245783 675262 245792
rect 675206 245576 675262 245585
rect 675262 245534 675418 245562
rect 675206 245511 675262 245520
rect 675208 245404 675260 245410
rect 675208 245346 675260 245352
rect 674852 245262 675064 245290
rect 674654 243536 674710 243545
rect 674654 243471 674710 243480
rect 674470 241088 674526 241097
rect 674470 241023 674526 241032
rect 674852 237289 674880 245262
rect 675022 241632 675078 241641
rect 675022 241567 675078 241576
rect 674838 237280 674894 237289
rect 674838 237215 674894 237224
rect 674194 236736 674250 236745
rect 674194 236671 674250 236680
rect 674088 234728 674140 234734
rect 674088 234670 674140 234676
rect 674100 234614 674128 234670
rect 674100 234586 674144 234614
rect 674116 234274 674144 234586
rect 674100 234258 674144 234274
rect 674088 234252 674144 234258
rect 674140 234246 674144 234252
rect 674088 234194 674140 234200
rect 673932 233294 674144 233322
rect 673966 233232 674018 233238
rect 674018 233180 674052 233186
rect 673966 233174 674052 233180
rect 673978 233158 674052 233174
rect 674024 222194 674052 233158
rect 674116 226930 674144 233294
rect 674208 231854 674236 236671
rect 674380 232688 674432 232694
rect 674378 232656 674380 232665
rect 674432 232656 674434 232665
rect 674378 232591 674434 232600
rect 674564 232552 674616 232558
rect 674564 232494 674616 232500
rect 674576 232393 674604 232494
rect 674562 232384 674618 232393
rect 674562 232319 674618 232328
rect 674208 231826 674604 231854
rect 674332 230072 674388 230081
rect 674332 230007 674388 230016
rect 674346 229838 674374 230007
rect 674452 229968 674504 229974
rect 674452 229910 674504 229916
rect 674334 229832 674386 229838
rect 674334 229774 674386 229780
rect 674464 229650 674492 229910
rect 674464 229622 674512 229650
rect 674484 229265 674512 229622
rect 674576 229378 674604 231826
rect 674840 231464 674892 231470
rect 674840 231406 674892 231412
rect 674852 230858 674880 231406
rect 674840 230852 674892 230858
rect 674840 230794 674892 230800
rect 674674 230344 674730 230353
rect 674674 230279 674676 230288
rect 674728 230279 674730 230288
rect 674676 230250 674728 230256
rect 674576 229350 674696 229378
rect 674470 229256 674526 229265
rect 674470 229191 674526 229200
rect 674116 226902 674328 226930
rect 674300 222465 674328 226902
rect 674286 222456 674342 222465
rect 674286 222391 674342 222400
rect 674668 222194 674696 229350
rect 674838 226128 674894 226137
rect 674838 226063 674894 226072
rect 674024 222166 674144 222194
rect 673012 164206 673224 164234
rect 672920 157306 673132 157334
rect 673104 152697 673132 157306
rect 673196 154574 673224 164206
rect 673288 164206 673408 164234
rect 673472 176626 673684 176654
rect 673748 215266 673868 215294
rect 673288 159338 673316 164206
rect 673472 162489 673500 176626
rect 673748 171850 673776 215266
rect 673918 214432 673974 214441
rect 673918 214367 673974 214376
rect 673932 177313 673960 214367
rect 673918 177304 673974 177313
rect 673918 177239 673974 177248
rect 673918 174448 673974 174457
rect 673918 174383 673974 174392
rect 673932 171986 673960 174383
rect 674116 172961 674144 222166
rect 674208 222166 674696 222194
rect 674208 220130 674236 222166
rect 674852 221785 674880 226063
rect 674838 221776 674894 221785
rect 674838 221711 674894 221720
rect 675036 221513 675064 241567
rect 675220 234614 675248 245346
rect 675390 243536 675446 243545
rect 675390 243471 675446 243480
rect 675404 243071 675432 243471
rect 675482 242720 675538 242729
rect 675482 242655 675538 242664
rect 675496 242519 675524 242655
rect 675390 242176 675446 242185
rect 675390 242111 675446 242120
rect 675404 241876 675432 242111
rect 675404 241097 675432 241231
rect 675390 241088 675446 241097
rect 675390 241023 675446 241032
rect 675390 240272 675446 240281
rect 675390 240207 675446 240216
rect 675404 240040 675432 240207
rect 675390 238640 675446 238649
rect 675390 238575 675446 238584
rect 675404 238204 675432 238575
rect 675496 237289 675524 237524
rect 675482 237280 675538 237289
rect 675482 237215 675538 237224
rect 675496 236201 675524 236368
rect 675482 236192 675538 236201
rect 675482 236127 675538 236136
rect 675482 235512 675538 235521
rect 675482 235447 675538 235456
rect 675220 234586 675340 234614
rect 675022 221504 675078 221513
rect 675022 221439 675078 221448
rect 674208 220102 674604 220130
rect 674576 215294 674604 220102
rect 675114 219056 675170 219065
rect 675114 218991 675170 219000
rect 674930 218240 674986 218249
rect 674930 218175 674986 218184
rect 674300 215266 674604 215294
rect 674102 172952 674158 172961
rect 674102 172887 674158 172896
rect 673932 171958 674236 171986
rect 673748 171822 674144 171850
rect 673734 170776 673790 170785
rect 673734 170711 673790 170720
rect 673748 164234 673776 170711
rect 674116 170626 674144 171822
rect 673656 164206 673776 164234
rect 673932 170598 674144 170626
rect 673458 162480 673514 162489
rect 673458 162415 673514 162424
rect 673656 162330 673684 164206
rect 673564 162302 673684 162330
rect 673288 159310 673408 159338
rect 673196 154546 673316 154574
rect 673090 152688 673146 152697
rect 673090 152623 673146 152632
rect 673288 151814 673316 154546
rect 673196 151786 673316 151814
rect 673196 151337 673224 151786
rect 673182 151328 673238 151337
rect 673182 151263 673238 151272
rect 673380 132161 673408 159310
rect 673564 156505 673592 162302
rect 673932 162194 673960 170598
rect 673656 162166 673960 162194
rect 673656 158930 673684 162166
rect 674208 161922 674236 171958
rect 673932 161894 674236 161922
rect 673656 158902 673776 158930
rect 673748 158817 673776 158902
rect 673734 158808 673790 158817
rect 673734 158743 673790 158752
rect 673550 156496 673606 156505
rect 673550 156431 673606 156440
rect 673366 132152 673422 132161
rect 673366 132087 673422 132096
rect 673932 129713 673960 161894
rect 674102 161800 674158 161809
rect 674102 161735 674158 161744
rect 673918 129704 673974 129713
rect 673918 129639 673974 129648
rect 673366 126576 673422 126585
rect 673366 126511 673422 126520
rect 673182 124944 673238 124953
rect 673182 124879 673238 124888
rect 672814 124128 672870 124137
rect 672814 124063 672870 124072
rect 673196 123162 673224 124879
rect 673196 123134 673316 123162
rect 673090 123040 673146 123049
rect 673090 122975 673146 122984
rect 672630 120864 672686 120873
rect 672630 120799 672686 120808
rect 672906 120728 672962 120737
rect 672906 120663 672962 120672
rect 672354 115832 672410 115841
rect 672354 115767 672410 115776
rect 672920 111081 672948 120663
rect 672906 111072 672962 111081
rect 672906 111007 672962 111016
rect 673104 109034 673132 122975
rect 673288 109034 673316 123134
rect 670804 109006 671384 109034
rect 671448 109006 671568 109034
rect 673012 109006 673132 109034
rect 673196 109006 673316 109034
rect 669964 108860 670016 108866
rect 669964 108802 670016 108808
rect 670804 106214 670832 109006
rect 670792 106208 670844 106214
rect 670792 106150 670844 106156
rect 671448 104802 671476 109006
rect 673012 106185 673040 109006
rect 672998 106176 673054 106185
rect 672998 106111 673054 106120
rect 670804 104774 671476 104802
rect 670804 104718 670832 104774
rect 668768 104712 668820 104718
rect 668768 104654 668820 104660
rect 670792 104712 670844 104718
rect 673196 104689 673224 109006
rect 670792 104654 670844 104660
rect 673182 104680 673238 104689
rect 668780 104553 668808 104654
rect 673182 104615 673238 104624
rect 668766 104544 668822 104553
rect 668766 104479 668822 104488
rect 668582 102912 668638 102921
rect 668582 102847 668638 102856
rect 673380 101017 673408 126511
rect 673918 124536 673974 124545
rect 673918 124471 673974 124480
rect 673932 107001 673960 124471
rect 674116 117473 674144 161735
rect 674300 153241 674328 215266
rect 674470 214976 674526 214985
rect 674470 214911 674526 214920
rect 674484 197169 674512 214911
rect 674654 213752 674710 213761
rect 674654 213687 674710 213696
rect 674668 205634 674696 213687
rect 674944 210746 674972 218175
rect 675128 215294 675156 218991
rect 674576 205606 674696 205634
rect 674760 210718 674972 210746
rect 675036 215266 675156 215294
rect 674576 202874 674604 205606
rect 674760 205057 674788 210718
rect 675036 208298 675064 215266
rect 675312 212537 675340 234586
rect 675496 228585 675524 235447
rect 675852 233912 675904 233918
rect 675850 233880 675852 233889
rect 678244 233912 678296 233918
rect 675904 233880 675906 233889
rect 678244 233854 678296 233860
rect 675850 233815 675906 233824
rect 675852 232688 675904 232694
rect 675850 232656 675852 232665
rect 675904 232656 675906 232665
rect 675850 232591 675906 232600
rect 676036 232552 676088 232558
rect 676036 232494 676088 232500
rect 676048 232393 676076 232494
rect 676034 232384 676090 232393
rect 676034 232319 676090 232328
rect 676494 230208 676550 230217
rect 676494 230143 676550 230152
rect 675482 228576 675538 228585
rect 675482 228511 675538 228520
rect 675482 225720 675538 225729
rect 675482 225655 675538 225664
rect 675496 219881 675524 225655
rect 675850 225176 675906 225185
rect 675850 225111 675906 225120
rect 675864 224954 675892 225111
rect 675680 224926 675892 224954
rect 675482 219872 675538 219881
rect 675482 219807 675538 219816
rect 675482 218648 675538 218657
rect 675680 218634 675708 224926
rect 676034 221912 676090 221921
rect 676034 221847 676090 221856
rect 675538 218606 675708 218634
rect 675482 218583 675538 218592
rect 675852 218000 675904 218006
rect 675666 217968 675722 217977
rect 675722 217948 675852 217954
rect 675722 217942 675904 217948
rect 675722 217926 675892 217942
rect 675666 217903 675722 217912
rect 675852 215688 675904 215694
rect 675666 215656 675722 215665
rect 675722 215636 675852 215642
rect 675722 215630 675904 215636
rect 675722 215614 675892 215630
rect 675666 215591 675722 215600
rect 675852 215008 675904 215014
rect 675680 214956 675852 214962
rect 675680 214950 675904 214956
rect 675680 214934 675892 214950
rect 675680 214713 675708 214934
rect 676048 214826 676076 221847
rect 676508 215014 676536 230143
rect 676770 227080 676826 227089
rect 676770 227015 676826 227024
rect 676784 218006 676812 227015
rect 676954 226808 677010 226817
rect 676954 226743 677010 226752
rect 676772 218000 676824 218006
rect 676772 217942 676824 217948
rect 676968 215694 676996 226743
rect 678256 223825 678284 233854
rect 683212 232688 683264 232694
rect 683212 232630 683264 232636
rect 678242 223816 678298 223825
rect 678242 223751 678298 223760
rect 683224 222737 683252 232630
rect 683396 232552 683448 232558
rect 683396 232494 683448 232500
rect 683408 223145 683436 232494
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683394 223136 683450 223145
rect 683394 223071 683450 223080
rect 683210 222728 683266 222737
rect 683210 222663 683266 222672
rect 676956 215688 677008 215694
rect 676956 215630 677008 215636
rect 676496 215008 676548 215014
rect 676496 214950 676548 214956
rect 675864 214798 676076 214826
rect 675666 214704 675722 214713
rect 675666 214639 675722 214648
rect 675864 214441 675892 214798
rect 676034 214568 676090 214577
rect 676034 214503 676090 214512
rect 675850 214432 675906 214441
rect 675850 214367 675906 214376
rect 675298 212528 675354 212537
rect 675298 212463 675354 212472
rect 676048 211449 676076 214503
rect 676034 211440 676090 211449
rect 676034 211375 676090 211384
rect 674944 208270 675064 208298
rect 674944 205714 674972 208270
rect 675114 206952 675170 206961
rect 675114 206887 675170 206896
rect 675128 205889 675156 206887
rect 675128 205861 675418 205889
rect 674944 205686 675156 205714
rect 674746 205048 674802 205057
rect 674746 204983 674802 204992
rect 674930 204232 674986 204241
rect 674930 204167 674986 204176
rect 674944 202881 674972 204167
rect 675128 204049 675156 205686
rect 675404 205057 675432 205323
rect 675390 205048 675446 205057
rect 675390 204983 675446 204992
rect 675404 204241 675432 204680
rect 675390 204232 675446 204241
rect 675390 204167 675446 204176
rect 675128 204021 675418 204049
rect 674576 202846 674788 202874
rect 674470 197160 674526 197169
rect 674470 197095 674526 197104
rect 674760 196058 674788 202846
rect 674930 202872 674986 202881
rect 674930 202807 674986 202816
rect 675758 202736 675814 202745
rect 675758 202671 675814 202680
rect 675772 202195 675800 202671
rect 675496 201385 675524 201620
rect 675482 201376 675538 201385
rect 675482 201311 675538 201320
rect 675128 200994 675418 201022
rect 674930 199744 674986 199753
rect 674930 199679 674986 199688
rect 674944 197350 674972 199679
rect 675128 198529 675156 200994
rect 675772 200025 675800 200328
rect 675758 200016 675814 200025
rect 675758 199951 675814 199960
rect 675114 198520 675170 198529
rect 675114 198455 675170 198464
rect 675482 198248 675538 198257
rect 675482 198183 675538 198192
rect 675496 197880 675524 198183
rect 674944 197322 675248 197350
rect 675220 197282 675248 197322
rect 675404 197282 675432 197336
rect 675220 197254 675432 197282
rect 675390 197160 675446 197169
rect 675390 197095 675446 197104
rect 675404 196656 675432 197095
rect 674760 196030 675418 196058
rect 675772 194585 675800 194820
rect 675758 194576 675814 194585
rect 675758 194511 675814 194520
rect 675758 193216 675814 193225
rect 675758 193151 675814 193160
rect 675772 192984 675800 193151
rect 675666 192808 675722 192817
rect 675666 192743 675722 192752
rect 675680 192372 675708 192743
rect 675128 191134 675418 191162
rect 675128 188873 675156 191134
rect 676034 189136 676090 189145
rect 676034 189071 676090 189080
rect 675114 188864 675170 188873
rect 675114 188799 675170 188808
rect 675850 180296 675906 180305
rect 675850 180231 675906 180240
rect 675864 177721 675892 180231
rect 675850 177712 675906 177721
rect 675850 177647 675906 177656
rect 676048 176654 676076 189071
rect 676218 181248 676274 181257
rect 676218 181183 676274 181192
rect 676232 178945 676260 181183
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 676218 178936 676274 178945
rect 676218 178871 676274 178880
rect 675680 176626 676076 176654
rect 674746 176080 674802 176089
rect 674746 176015 674802 176024
rect 674562 175264 674618 175273
rect 674562 175199 674618 175208
rect 674576 173894 674604 175199
rect 674760 174162 674788 176015
rect 674392 173866 674604 173894
rect 674668 174134 674788 174162
rect 674392 166994 674420 173866
rect 674392 166966 674512 166994
rect 674286 153232 674342 153241
rect 674286 153167 674342 153176
rect 674484 130529 674512 166966
rect 674668 131345 674696 174134
rect 674838 174040 674894 174049
rect 674838 173975 674894 173984
rect 674852 159066 674880 173975
rect 675680 167521 675708 176626
rect 681002 173632 681058 173641
rect 681002 173567 681058 173576
rect 676034 173224 676090 173233
rect 676090 173182 676260 173210
rect 676034 173159 676090 173168
rect 676232 169674 676260 173182
rect 676586 169960 676642 169969
rect 676586 169895 676642 169904
rect 675864 169646 676260 169674
rect 675666 167512 675722 167521
rect 675666 167447 675722 167456
rect 675864 166994 675892 169646
rect 675680 166966 675892 166994
rect 675206 162072 675262 162081
rect 675206 162007 675262 162016
rect 675220 159678 675248 162007
rect 675680 161786 675708 166966
rect 676600 166433 676628 169895
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 675852 164212 675904 164218
rect 675852 164154 675904 164160
rect 675864 162081 675892 164154
rect 681016 162761 681044 173567
rect 682382 171592 682438 171601
rect 682382 171527 682438 171536
rect 682396 164218 682424 171527
rect 683118 167920 683174 167929
rect 683118 167855 683174 167864
rect 682384 164212 682436 164218
rect 682384 164154 682436 164160
rect 681002 162752 681058 162761
rect 681002 162687 681058 162696
rect 683132 162081 683160 167855
rect 675850 162072 675906 162081
rect 675850 162007 675906 162016
rect 683118 162072 683174 162081
rect 683118 162007 683174 162016
rect 675312 161758 675708 161786
rect 675312 160290 675340 161758
rect 675482 161528 675538 161537
rect 675482 161463 675538 161472
rect 675496 160888 675524 161463
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675220 159650 675418 159678
rect 674852 159038 675340 159066
rect 675312 158930 675340 159038
rect 675404 158930 675432 159052
rect 675312 158902 675432 158930
rect 675772 157049 675800 157216
rect 675758 157040 675814 157049
rect 675758 156975 675814 156984
rect 675128 156629 675418 156657
rect 675128 155961 675156 156629
rect 675298 156496 675354 156505
rect 675298 156431 675354 156440
rect 675312 156006 675340 156431
rect 675312 155978 675418 156006
rect 675114 155952 675170 155961
rect 675114 155887 675170 155896
rect 675758 155816 675814 155825
rect 675758 155751 675814 155760
rect 675772 155380 675800 155751
rect 674944 152850 675418 152878
rect 674944 150385 674972 152850
rect 675114 152688 675170 152697
rect 675114 152623 675170 152632
rect 675128 152334 675156 152623
rect 675128 152306 675418 152334
rect 675772 151473 675800 151675
rect 675758 151464 675814 151473
rect 675758 151399 675814 151408
rect 675114 151328 675170 151337
rect 675114 151263 675170 151272
rect 675128 151042 675156 151263
rect 675128 151014 675418 151042
rect 674930 150376 674986 150385
rect 674930 150311 674986 150320
rect 675128 149821 675418 149849
rect 675128 147665 675156 149821
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675114 147656 675170 147665
rect 675114 147591 675170 147600
rect 675390 147656 675446 147665
rect 675390 147591 675446 147600
rect 675404 147356 675432 147591
rect 675312 146254 675432 146282
rect 675312 146146 675340 146254
rect 675128 146118 675340 146146
rect 675404 146132 675432 146254
rect 675128 144945 675156 146118
rect 675114 144936 675170 144945
rect 675114 144871 675170 144880
rect 675850 134600 675906 134609
rect 675850 134535 675906 134544
rect 675864 133958 675892 134535
rect 675852 133952 675904 133958
rect 675852 133894 675904 133900
rect 676496 133952 676548 133958
rect 676496 133894 676548 133900
rect 676508 133113 676536 133894
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676494 133104 676550 133113
rect 676494 133039 676550 133048
rect 674654 131336 674710 131345
rect 674654 131271 674710 131280
rect 674470 130520 674526 130529
rect 674470 130455 674526 130464
rect 676218 130248 676274 130257
rect 676218 130183 676274 130192
rect 675022 128888 675078 128897
rect 675022 128823 675078 128832
rect 674378 128480 674434 128489
rect 674378 128415 674434 128424
rect 674102 117464 674158 117473
rect 674102 117399 674158 117408
rect 673918 106992 673974 107001
rect 673918 106927 673974 106936
rect 674392 102830 674420 128415
rect 674654 124128 674710 124137
rect 674654 124063 674710 124072
rect 674668 105822 674696 124063
rect 674838 123720 674894 123729
rect 674838 123655 674894 123664
rect 674852 123049 674880 123655
rect 674838 123040 674894 123049
rect 674838 122975 674894 122984
rect 675036 122834 675064 128823
rect 676232 127809 676260 130183
rect 676218 127800 676274 127809
rect 676218 127735 676274 127744
rect 676402 127800 676458 127809
rect 676402 127735 676458 127744
rect 676416 125458 676444 127735
rect 679622 126168 679678 126177
rect 679622 126103 679678 126112
rect 675852 125452 675904 125458
rect 674852 122806 675064 122834
rect 675496 125412 675852 125440
rect 674852 113846 674880 122806
rect 675206 117056 675262 117065
rect 675206 116991 675262 117000
rect 675220 114493 675248 116991
rect 675496 115934 675524 125412
rect 675852 125394 675904 125400
rect 676404 125452 676456 125458
rect 676404 125394 676456 125400
rect 679636 118522 679664 126103
rect 682382 125352 682438 125361
rect 682382 125287 682438 125296
rect 675852 118516 675904 118522
rect 675852 118458 675904 118464
rect 679624 118516 679676 118522
rect 679624 118458 679676 118464
rect 675864 117065 675892 118458
rect 682396 117337 682424 125287
rect 682382 117328 682438 117337
rect 682382 117263 682438 117272
rect 675850 117056 675906 117065
rect 675850 116991 675906 117000
rect 675312 115906 675524 115934
rect 675312 115138 675340 115906
rect 675482 115832 675538 115841
rect 675482 115767 675538 115776
rect 675496 115668 675524 115767
rect 675312 115110 675418 115138
rect 675220 114465 675418 114493
rect 674852 113818 675418 113846
rect 675758 112432 675814 112441
rect 675758 112367 675814 112376
rect 675772 111996 675800 112367
rect 675758 111752 675814 111761
rect 675758 111687 675814 111696
rect 675772 111452 675800 111687
rect 675758 111344 675814 111353
rect 675758 111279 675814 111288
rect 675772 110772 675800 111279
rect 675758 110392 675814 110401
rect 675758 110327 675814 110336
rect 675772 110160 675800 110327
rect 675758 108216 675814 108225
rect 675758 108151 675814 108160
rect 675772 107644 675800 108151
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106185 675156 107086
rect 675390 106992 675446 107001
rect 675390 106927 675446 106936
rect 675404 106488 675432 106927
rect 675114 106176 675170 106185
rect 675114 106111 675170 106120
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 674668 105794 675340 105822
rect 675404 105808 675432 105862
rect 675114 104680 675170 104689
rect 675170 104638 675340 104666
rect 675114 104615 675170 104624
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 674392 102802 675340 102830
rect 675312 102762 675340 102802
rect 675404 102762 675432 102816
rect 675312 102734 675432 102762
rect 675404 101969 675432 102136
rect 675390 101960 675446 101969
rect 675390 101895 675446 101904
rect 673366 101008 673422 101017
rect 673366 100943 673422 100952
rect 675114 101008 675170 101017
rect 675170 100966 675340 100994
rect 675114 100943 675170 100952
rect 675312 100858 675340 100966
rect 675404 100858 675432 100980
rect 675312 100830 675432 100858
rect 595272 100014 595608 100042
rect 596344 100014 596496 100042
rect 595272 99142 595300 100014
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 595272 93854 595300 99078
rect 596180 96960 596232 96966
rect 596180 96902 596232 96908
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 596192 54398 596220 96902
rect 596468 55214 596496 100014
rect 596744 100014 597080 100042
rect 596744 96966 596772 100014
rect 597802 99770 597830 100028
rect 598216 100014 598552 100042
rect 599136 100014 599288 100042
rect 599688 100014 600024 100042
rect 600516 100014 600760 100042
rect 601160 100014 601496 100042
rect 601712 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 597802 99742 597876 99770
rect 596732 96960 596784 96966
rect 596732 96902 596784 96908
rect 597652 96960 597704 96966
rect 597652 96902 597704 96908
rect 596456 55208 596508 55214
rect 596456 55150 596508 55156
rect 597664 54942 597692 96902
rect 597848 55078 597876 99742
rect 598216 96966 598244 100014
rect 598204 96960 598256 96966
rect 598204 96902 598256 96908
rect 598940 96960 598992 96966
rect 598940 96902 598992 96908
rect 598952 56030 598980 96902
rect 598940 56024 598992 56030
rect 598940 55966 598992 55972
rect 597836 55072 597888 55078
rect 597836 55014 597888 55020
rect 597652 54936 597704 54942
rect 597652 54878 597704 54884
rect 599136 54806 599164 100014
rect 599688 96966 599716 100014
rect 599676 96960 599728 96966
rect 599676 96902 599728 96908
rect 600320 96960 600372 96966
rect 600320 96902 600372 96908
rect 600332 57254 600360 96902
rect 600320 57248 600372 57254
rect 600320 57190 600372 57196
rect 600516 55894 600544 100014
rect 601160 96966 601188 100014
rect 601148 96960 601200 96966
rect 601148 96902 601200 96908
rect 601712 72486 601740 100014
rect 602356 84194 602384 100014
rect 601896 84166 602384 84194
rect 601700 72480 601752 72486
rect 601700 72422 601752 72428
rect 601896 58682 601924 84166
rect 603092 60042 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 604426 99742 604500 99770
rect 604472 68338 604500 99742
rect 605484 97306 605512 100014
rect 605472 97300 605524 97306
rect 605472 97242 605524 97248
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606956 92886 606984 100014
rect 607128 96960 607180 96966
rect 607128 96902 607180 96908
rect 606944 92880 606996 92886
rect 606944 92822 606996 92828
rect 607140 75206 607168 96902
rect 607692 95946 607720 100014
rect 607680 95940 607732 95946
rect 607680 95882 607732 95888
rect 608520 84182 608548 100014
rect 609164 94518 609192 100014
rect 609152 94512 609204 94518
rect 609152 94454 609204 94460
rect 609900 85406 609928 100014
rect 610636 96762 610664 100014
rect 611050 99770 611078 100028
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613884 100042
rect 611050 99742 611124 99770
rect 610624 96756 610676 96762
rect 610624 96698 610676 96704
rect 611096 96082 611124 99742
rect 611912 97300 611964 97306
rect 611912 97242 611964 97248
rect 611268 96756 611320 96762
rect 611268 96698 611320 96704
rect 611084 96076 611136 96082
rect 611084 96018 611136 96024
rect 611280 93158 611308 96698
rect 611924 93854 611952 97242
rect 612108 96898 612136 100014
rect 612660 97442 612688 100014
rect 612648 97436 612700 97442
rect 612648 97378 612700 97384
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 611924 93826 612044 93854
rect 611268 93152 611320 93158
rect 611268 93094 611320 93100
rect 610072 92880 610124 92886
rect 610072 92822 610124 92828
rect 610084 88330 610112 92822
rect 610072 88324 610124 88330
rect 610072 88266 610124 88272
rect 609888 85400 609940 85406
rect 609888 85342 609940 85348
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 612016 76566 612044 93826
rect 612660 80850 612688 96834
rect 612648 80844 612700 80850
rect 612648 80786 612700 80792
rect 613856 79490 613884 100014
rect 613994 99770 614022 100028
rect 614744 100014 615264 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613994 99742 614068 99770
rect 613844 79484 613896 79490
rect 613844 79426 613896 79432
rect 614040 79354 614068 99742
rect 615236 93854 615264 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 616524 95062 616552 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616512 95056 616564 95062
rect 616512 94998 616564 95004
rect 615236 93826 615448 93854
rect 614028 79348 614080 79354
rect 614028 79290 614080 79296
rect 612004 76560 612056 76566
rect 612004 76502 612056 76508
rect 615420 75342 615448 93826
rect 616800 76702 616828 96902
rect 617260 96898 617288 100014
rect 617248 96892 617300 96898
rect 617248 96834 617300 96840
rect 617996 92478 618024 100014
rect 618732 97986 618760 100014
rect 618720 97980 618772 97986
rect 618720 97922 618772 97928
rect 618904 97436 618956 97442
rect 618904 97378 618956 97384
rect 618168 96892 618220 96898
rect 618168 96834 618220 96840
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91050 618208 96834
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 616788 76696 616840 76702
rect 616788 76638 616840 76644
rect 618916 75478 618944 97378
rect 619560 93838 619588 100014
rect 620204 97850 620232 100014
rect 620192 97844 620244 97850
rect 620192 97786 620244 97792
rect 620940 95198 620968 100014
rect 621676 97578 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 621664 97572 621716 97578
rect 621664 97514 621716 97520
rect 623148 97442 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 623136 97436 623188 97442
rect 623136 97378 623188 97384
rect 624620 97034 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633296 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 625080 99074 625108 99742
rect 625068 99068 625120 99074
rect 625068 99010 625120 99016
rect 625804 97980 625856 97986
rect 625804 97922 625856 97928
rect 625620 97844 625672 97850
rect 625620 97786 625672 97792
rect 624608 97028 624660 97034
rect 624608 96970 624660 96976
rect 622308 96076 622360 96082
rect 622308 96018 622360 96024
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620284 94512 620336 94518
rect 620284 94454 620336 94460
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 619272 93152 619324 93158
rect 619272 93094 619324 93100
rect 619284 86358 619312 93094
rect 619272 86352 619324 86358
rect 619272 86294 619324 86300
rect 620296 85542 620324 94454
rect 622320 88194 622348 96018
rect 624976 95940 625028 95946
rect 624976 95882 625028 95888
rect 622952 95056 623004 95062
rect 622952 94998 623004 95004
rect 622964 89622 622992 94998
rect 622952 89616 623004 89622
rect 622952 89558 623004 89564
rect 624988 88777 625016 95882
rect 625632 93673 625660 97786
rect 625618 93664 625674 93673
rect 625618 93599 625674 93608
rect 625816 92041 625844 97922
rect 626092 97306 626120 100014
rect 626080 97300 626132 97306
rect 626080 97242 626132 97248
rect 626828 97170 626856 100014
rect 627564 97850 627592 100014
rect 628300 98938 628328 100014
rect 628288 98932 628340 98938
rect 628288 98874 628340 98880
rect 629036 98802 629064 100014
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 629772 97986 629800 100014
rect 630508 98666 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98660 630548 98666
rect 630496 98602 630548 98608
rect 629760 97980 629812 97986
rect 629760 97922 629812 97928
rect 627552 97844 627604 97850
rect 627552 97786 627604 97792
rect 629300 97572 629352 97578
rect 629300 97514 629352 97520
rect 626816 97164 626868 97170
rect 626816 97106 626868 97112
rect 629312 95826 629340 97514
rect 630784 95826 630812 99282
rect 631048 98252 631100 98258
rect 631048 98194 631100 98200
rect 631060 97850 631088 98194
rect 631048 97844 631100 97850
rect 631048 97786 631100 97792
rect 631244 96354 631272 100014
rect 631980 97850 632008 100014
rect 631968 97844 632020 97850
rect 631968 97786 632020 97792
rect 632716 97714 632744 100014
rect 632704 97708 632756 97714
rect 632704 97650 632756 97656
rect 633268 97442 633296 100014
rect 633440 99204 633492 99210
rect 633440 99146 633492 99152
rect 632060 97436 632112 97442
rect 632060 97378 632112 97384
rect 633256 97436 633308 97442
rect 633256 97378 633308 97384
rect 631232 96348 631284 96354
rect 631232 96290 631284 96296
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 632072 95826 632100 97378
rect 633452 95826 633480 99146
rect 634188 97578 634216 100014
rect 634176 97572 634228 97578
rect 634176 97514 634228 97520
rect 634740 96898 634768 100014
rect 635568 97034 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635004 97028 635056 97034
rect 635004 96970 635056 96976
rect 635556 97028 635608 97034
rect 635556 96970 635608 96976
rect 634728 96892 634780 96898
rect 634728 96834 634780 96840
rect 635016 95826 635044 96970
rect 632072 95798 632224 95826
rect 633452 95798 633696 95826
rect 635016 95798 635168 95826
rect 635752 95441 635780 100014
rect 636292 99068 636344 99074
rect 636292 99010 636344 99016
rect 636304 95826 636332 99010
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96218 637620 99742
rect 637764 97300 637816 97306
rect 637764 97242 637816 97248
rect 637580 96212 637632 96218
rect 637580 96154 637632 96160
rect 637776 95826 637804 97242
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 638604 95742 638632 100014
rect 639018 99770 639046 100028
rect 639768 100014 640104 100042
rect 639018 99742 639092 99770
rect 639064 96490 639092 99742
rect 639236 97164 639288 97170
rect 639236 97106 639288 97112
rect 639052 96484 639104 96490
rect 639052 96426 639104 96432
rect 639248 95826 639276 97106
rect 639248 95798 639584 95826
rect 638592 95736 638644 95742
rect 638592 95678 638644 95684
rect 640076 95606 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640536 96626 640564 99742
rect 640708 98184 640760 98190
rect 640708 98126 640760 98132
rect 640524 96620 640576 96626
rect 640524 96562 640576 96568
rect 640720 95826 640748 98126
rect 640720 95798 641056 95826
rect 640064 95600 640116 95606
rect 640064 95542 640116 95548
rect 641548 95470 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 642008 96529 642036 99742
rect 642180 98932 642232 98938
rect 642180 98874 642232 98880
rect 641994 96520 642050 96529
rect 641994 96455 642050 96464
rect 642192 95826 642220 98874
rect 643020 97306 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 643434 99742 643508 99770
rect 643008 97300 643060 97306
rect 643008 97242 643060 97248
rect 643480 95878 643508 99742
rect 643652 98796 643704 98802
rect 643652 98738 643704 98744
rect 643468 95872 643520 95878
rect 642192 95798 642528 95826
rect 643468 95814 643520 95820
rect 643664 95826 643692 98738
rect 644308 97170 644336 100014
rect 644906 99770 644934 100028
rect 645656 100014 645808 100042
rect 644906 99742 644980 99770
rect 644296 97164 644348 97170
rect 644296 97106 644348 97112
rect 644952 96014 644980 99742
rect 645308 98048 645360 98054
rect 645308 97990 645360 97996
rect 645124 96484 645176 96490
rect 645124 96426 645176 96432
rect 644940 96008 644992 96014
rect 644940 95950 644992 95956
rect 643664 95798 644000 95826
rect 645136 95470 645164 96426
rect 645320 95826 645348 97990
rect 645780 96626 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648476 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651328 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 645768 96620 645820 96626
rect 645768 96562 645820 96568
rect 646424 96490 646452 99742
rect 647160 98802 647188 99742
rect 647148 98796 647200 98802
rect 647148 98738 647200 98744
rect 646596 98660 646648 98666
rect 646596 98602 646648 98608
rect 646412 96484 646464 96490
rect 646412 96426 646464 96432
rect 646608 95826 646636 98602
rect 647516 97844 647568 97850
rect 647516 97786 647568 97792
rect 647148 96348 647200 96354
rect 647148 96290 647200 96296
rect 645320 95798 645472 95826
rect 646608 95798 646944 95826
rect 641536 95464 641588 95470
rect 635738 95432 635794 95441
rect 641536 95406 641588 95412
rect 645124 95464 645176 95470
rect 645124 95406 645176 95412
rect 635738 95367 635794 95376
rect 626448 95192 626500 95198
rect 626448 95134 626500 95140
rect 626460 94489 626488 95134
rect 647160 95033 647188 96290
rect 647332 95736 647384 95742
rect 647332 95678 647384 95684
rect 647146 95024 647202 95033
rect 647146 94959 647202 94968
rect 626446 94480 626502 94489
rect 626446 94415 626502 94424
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 626460 92857 626488 93774
rect 626446 92848 626502 92857
rect 626446 92783 626502 92792
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626460 91225 626488 92414
rect 647344 92410 647372 95678
rect 647528 92449 647556 97786
rect 648252 97708 648304 97714
rect 648252 97650 648304 97656
rect 647700 97028 647752 97034
rect 647700 96970 647752 96976
rect 647712 95130 647740 96970
rect 647884 96756 647936 96762
rect 647884 96698 647936 96704
rect 647896 95742 647924 96698
rect 647884 95736 647936 95742
rect 647884 95678 647936 95684
rect 647884 95600 647936 95606
rect 647884 95542 647936 95548
rect 647700 95124 647752 95130
rect 647700 95066 647752 95072
rect 647514 92440 647570 92449
rect 647332 92404 647384 92410
rect 647514 92375 647570 92384
rect 647332 92346 647384 92352
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 625252 89616 625304 89622
rect 625250 89584 625252 89593
rect 625304 89584 625306 89593
rect 625250 89519 625306 89528
rect 624974 88768 625030 88777
rect 624974 88703 625030 88712
rect 625160 88324 625212 88330
rect 625160 88266 625212 88272
rect 622308 88188 622360 88194
rect 622308 88130 622360 88136
rect 625172 87961 625200 88266
rect 625344 88188 625396 88194
rect 625344 88130 625396 88136
rect 625158 87952 625214 87961
rect 625158 87887 625214 87896
rect 625356 87145 625384 88130
rect 625342 87136 625398 87145
rect 625342 87071 625398 87080
rect 647896 86630 647924 95542
rect 648264 89593 648292 97650
rect 648250 89584 648306 89593
rect 648250 89519 648306 89528
rect 648448 87038 648476 100014
rect 648620 97436 648672 97442
rect 648620 97378 648672 97384
rect 648632 92546 648660 97378
rect 648908 96354 648936 100014
rect 648896 96348 648948 96354
rect 648896 96290 648948 96296
rect 649540 96008 649592 96014
rect 649540 95950 649592 95956
rect 649264 95872 649316 95878
rect 649264 95814 649316 95820
rect 648804 95124 648856 95130
rect 648804 95066 648856 95072
rect 648620 92540 648672 92546
rect 648620 92482 648672 92488
rect 648436 87032 648488 87038
rect 648436 86974 648488 86980
rect 647884 86624 647936 86630
rect 647884 86566 647936 86572
rect 625160 86352 625212 86358
rect 625158 86320 625160 86329
rect 625212 86320 625214 86329
rect 625158 86255 625214 86264
rect 620284 85536 620336 85542
rect 625344 85536 625396 85542
rect 620284 85478 620336 85484
rect 625158 85504 625214 85513
rect 625344 85478 625396 85484
rect 625158 85439 625214 85448
rect 625172 85338 625200 85439
rect 625160 85332 625212 85338
rect 625160 85274 625212 85280
rect 625356 84697 625384 85478
rect 625342 84688 625398 84697
rect 625342 84623 625398 84632
rect 625160 84176 625212 84182
rect 625160 84118 625212 84124
rect 625172 83881 625200 84118
rect 625158 83872 625214 83881
rect 625158 83807 625214 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 80986 628788 83263
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 80980 628800 80986
rect 628748 80922 628800 80928
rect 629220 80034 629248 81631
rect 632808 80974 633144 81002
rect 642456 80980 642508 80986
rect 629208 80028 629260 80034
rect 629208 79970 629260 79976
rect 631048 77988 631100 77994
rect 631048 77930 631100 77936
rect 628472 77784 628524 77790
rect 628472 77726 628524 77732
rect 624422 77344 624478 77353
rect 624422 77279 624478 77288
rect 625804 77308 625856 77314
rect 618904 75472 618956 75478
rect 618904 75414 618956 75420
rect 615408 75336 615460 75342
rect 615408 75278 615460 75284
rect 607128 75200 607180 75206
rect 607128 75142 607180 75148
rect 604460 68332 604512 68338
rect 604460 68274 604512 68280
rect 603080 60036 603132 60042
rect 603080 59978 603132 59984
rect 601884 58676 601936 58682
rect 601884 58618 601936 58624
rect 600504 55888 600556 55894
rect 600504 55830 600556 55836
rect 599124 54800 599176 54806
rect 599124 54742 599176 54748
rect 624436 54670 624464 77279
rect 625804 77250 625856 77256
rect 624424 54664 624476 54670
rect 624424 54606 624476 54612
rect 625816 54534 625844 77250
rect 628484 75290 628512 77726
rect 631060 77314 631088 77930
rect 632808 77790 632836 80974
rect 643080 80974 643140 81002
rect 642456 80922 642508 80928
rect 636752 80708 636804 80714
rect 636752 80650 636804 80656
rect 633440 80028 633492 80034
rect 633440 79970 633492 79976
rect 633452 78130 633480 79970
rect 633898 78568 633954 78577
rect 633898 78503 633954 78512
rect 633440 78124 633492 78130
rect 633440 78066 633492 78072
rect 632796 77784 632848 77790
rect 632796 77726 632848 77732
rect 633912 77353 633940 78503
rect 633898 77344 633954 77353
rect 631048 77308 631100 77314
rect 633898 77279 633954 77288
rect 631048 77250 631100 77256
rect 631060 75290 631088 77250
rect 633912 75290 633940 77279
rect 636764 75290 636792 80650
rect 639602 78160 639658 78169
rect 639602 78095 639658 78104
rect 639616 75290 639644 78095
rect 642468 75290 642496 80922
rect 643112 77994 643140 80974
rect 647424 80844 647476 80850
rect 647424 80786 647476 80792
rect 645952 79484 646004 79490
rect 645952 79426 646004 79432
rect 645308 78124 645360 78130
rect 645308 78066 645360 78072
rect 643100 77988 643152 77994
rect 643100 77930 643152 77936
rect 645320 75290 645348 78066
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 645964 64874 645992 79426
rect 646504 79348 646556 79354
rect 646504 79290 646556 79296
rect 646320 76696 646372 76702
rect 646320 76638 646372 76644
rect 646136 75200 646188 75206
rect 646136 75142 646188 75148
rect 646148 74225 646176 75142
rect 646134 74216 646190 74225
rect 646134 74151 646190 74160
rect 646332 71777 646360 76638
rect 646318 71768 646374 71777
rect 646318 71703 646374 71712
rect 646516 67153 646544 79290
rect 646872 75336 646924 75342
rect 646872 75278 646924 75284
rect 646884 74534 646912 75278
rect 646884 74506 647280 74534
rect 647252 68921 647280 74506
rect 647238 68912 647294 68921
rect 647238 68847 647294 68856
rect 646502 67144 646558 67153
rect 646502 67079 646558 67088
rect 647436 64874 647464 80786
rect 648620 75472 648672 75478
rect 648620 75414 648672 75420
rect 645964 64846 646176 64874
rect 646148 64433 646176 64846
rect 647252 64846 647464 64874
rect 646134 64424 646190 64433
rect 646134 64359 646190 64368
rect 647252 59265 647280 64846
rect 648632 62121 648660 75414
rect 648618 62112 648674 62121
rect 648618 62047 648674 62056
rect 647238 59256 647294 59265
rect 647238 59191 647294 59200
rect 648816 57361 648844 95066
rect 649276 86766 649304 95814
rect 649552 93974 649580 95950
rect 649540 93968 649592 93974
rect 649540 93910 649592 93916
rect 649736 88806 649764 100014
rect 650380 97578 650408 100014
rect 650368 97572 650420 97578
rect 650368 97514 650420 97520
rect 650552 97436 650604 97442
rect 650552 97378 650604 97384
rect 650368 96892 650420 96898
rect 650368 96834 650420 96840
rect 649908 96076 649960 96082
rect 649908 96018 649960 96024
rect 649920 95334 649948 96018
rect 649908 95328 649960 95334
rect 649908 95270 649960 95276
rect 650000 92540 650052 92546
rect 650000 92482 650052 92488
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 650012 87145 650040 92482
rect 649998 87136 650054 87145
rect 649998 87071 650054 87080
rect 649264 86760 649316 86766
rect 649264 86702 649316 86708
rect 650380 82249 650408 96834
rect 650564 84697 650592 97378
rect 651300 93566 651328 100014
rect 651852 97714 651880 100014
rect 651840 97708 651892 97714
rect 651840 97650 651892 97656
rect 652588 96490 652616 100014
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 652576 96484 652628 96490
rect 652576 96426 652628 96432
rect 651840 95464 651892 95470
rect 651840 95406 651892 95412
rect 651288 93560 651340 93566
rect 651288 93502 651340 93508
rect 651852 90710 651880 95406
rect 651840 90704 651892 90710
rect 651840 90646 651892 90652
rect 652036 86358 652064 96426
rect 653324 95674 653352 100014
rect 653968 96898 653996 100014
rect 653956 96892 654008 96898
rect 653956 96834 654008 96840
rect 654796 96762 654824 100014
rect 655440 97850 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97844 655480 97850
rect 655428 97786 655480 97792
rect 655244 96892 655296 96898
rect 655244 96834 655296 96840
rect 654784 96756 654836 96762
rect 654784 96698 654836 96704
rect 653312 95668 653364 95674
rect 653312 95610 653364 95616
rect 655256 94217 655284 96834
rect 655428 96756 655480 96762
rect 655428 96698 655480 96704
rect 655242 94208 655298 94217
rect 655242 94143 655298 94152
rect 655440 93854 655468 96698
rect 655256 93826 655468 93854
rect 654324 92404 654376 92410
rect 654324 92346 654376 92352
rect 654336 91497 654364 92346
rect 654322 91488 654378 91497
rect 654322 91423 654378 91432
rect 655256 88330 655284 93826
rect 655428 93560 655480 93566
rect 655428 93502 655480 93508
rect 655440 93401 655468 93502
rect 655426 93392 655482 93401
rect 655426 93327 655482 93336
rect 655428 90704 655480 90710
rect 655426 90672 655428 90681
rect 655480 90672 655482 90681
rect 655426 90607 655482 90616
rect 655808 89865 655836 100014
rect 656820 97306 656848 100014
rect 656532 97300 656584 97306
rect 656532 97242 656584 97248
rect 656808 97300 656860 97306
rect 656808 97242 656860 97248
rect 656544 96762 656572 97242
rect 656716 96892 656768 96898
rect 656716 96834 656768 96840
rect 656532 96756 656584 96762
rect 656532 96698 656584 96704
rect 656348 96620 656400 96626
rect 656348 96562 656400 96568
rect 656164 93968 656216 93974
rect 656164 93910 656216 93916
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 656176 86494 656204 93910
rect 656360 88670 656388 96562
rect 656348 88664 656400 88670
rect 656348 88606 656400 88612
rect 656728 86902 656756 96834
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 658108 99742 658182 99770
rect 658108 97442 658136 99742
rect 658280 97572 658332 97578
rect 658280 97514 658332 97520
rect 658096 97436 658148 97442
rect 658096 97378 658148 97384
rect 658292 95132 658320 97514
rect 658832 97164 658884 97170
rect 658832 97106 658884 97112
rect 658844 95132 658872 97106
rect 659212 97034 659240 100014
rect 659948 97986 659976 100014
rect 660132 100014 660376 100042
rect 659936 97980 659988 97986
rect 659936 97922 659988 97928
rect 659568 97708 659620 97714
rect 659568 97650 659620 97656
rect 659200 97028 659252 97034
rect 659200 96970 659252 96976
rect 659580 95132 659608 97650
rect 660132 96898 660160 100014
rect 661960 98796 662012 98802
rect 661960 98738 662012 98744
rect 661408 97300 661460 97306
rect 661408 97242 661460 97248
rect 660120 96892 660172 96898
rect 660120 96834 660172 96840
rect 660120 96756 660172 96762
rect 660120 96698 660172 96704
rect 660132 95132 660160 96698
rect 660672 96212 660724 96218
rect 660672 96154 660724 96160
rect 660684 95132 660712 96154
rect 661420 95132 661448 97242
rect 661972 95132 662000 98738
rect 665180 97980 665232 97986
rect 665180 97922 665232 97928
rect 662512 97844 662564 97850
rect 662512 97786 662564 97792
rect 662524 95132 662552 97786
rect 663064 97436 663116 97442
rect 663064 97378 663116 97384
rect 663076 95132 663104 97378
rect 663892 97028 663944 97034
rect 663892 96970 663944 96976
rect 663708 96076 663760 96082
rect 663708 96018 663760 96024
rect 663720 95962 663748 96018
rect 663720 95934 663840 95962
rect 663812 92970 663840 95934
rect 663720 92942 663840 92970
rect 663720 92857 663748 92942
rect 663706 92848 663762 92857
rect 663706 92783 663762 92792
rect 663904 88806 663932 96970
rect 664168 96348 664220 96354
rect 664168 96290 664220 96296
rect 664180 89865 664208 96290
rect 664352 95668 664404 95674
rect 664352 95610 664404 95616
rect 664166 89856 664222 89865
rect 664166 89791 664222 89800
rect 664364 89049 664392 95610
rect 665192 93401 665220 97922
rect 665548 96484 665600 96490
rect 665548 96426 665600 96432
rect 665364 95940 665416 95946
rect 665364 95882 665416 95888
rect 665178 93392 665234 93401
rect 665178 93327 665234 93336
rect 665376 91769 665404 95882
rect 665362 91760 665418 91769
rect 665362 91695 665418 91704
rect 665560 90681 665588 96426
rect 665546 90672 665602 90681
rect 665546 90607 665602 90616
rect 664350 89040 664406 89049
rect 664350 88975 664406 88984
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 663892 88800 663944 88806
rect 663892 88742 663944 88748
rect 661986 88726 662368 88742
rect 657452 88664 657504 88670
rect 657504 88612 657754 88618
rect 657452 88606 657754 88612
rect 657464 88590 657754 88606
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656716 86896 656768 86902
rect 656716 86838 656768 86844
rect 656164 86488 656216 86494
rect 656164 86430 656216 86436
rect 657188 86358 657216 88196
rect 659580 86902 659608 88196
rect 659568 86896 659620 86902
rect 659568 86838 659620 86844
rect 660132 86630 660160 88196
rect 660120 86624 660172 86630
rect 660120 86566 660172 86572
rect 660684 86494 660712 88196
rect 661420 86766 661448 88196
rect 662524 87038 662552 88196
rect 662512 87032 662564 87038
rect 662512 86974 662564 86980
rect 661408 86760 661460 86766
rect 661408 86702 661460 86708
rect 660672 86488 660724 86494
rect 660672 86430 660724 86436
rect 652024 86352 652076 86358
rect 652024 86294 652076 86300
rect 657176 86352 657228 86358
rect 657176 86294 657228 86300
rect 650550 84688 650606 84697
rect 650550 84623 650606 84632
rect 650366 82240 650422 82249
rect 650366 82175 650422 82184
rect 662420 76560 662472 76566
rect 662420 76502 662472 76508
rect 648802 57352 648858 57361
rect 648802 57287 648858 57296
rect 625804 54528 625856 54534
rect 625804 54470 625856 54476
rect 596180 54392 596232 54398
rect 596180 54334 596232 54340
rect 592684 51740 592736 51746
rect 592684 51682 592736 51688
rect 661590 48510 661646 48519
rect 661590 48445 661646 48454
rect 553674 48104 553730 48113
rect 553674 48039 553730 48048
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 46744 465318 46753
rect 465262 46679 465318 46688
rect 661604 45554 661632 48445
rect 662432 47433 662460 76502
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661420 45526 661632 45554
rect 464342 44160 464398 44169
rect 464342 44095 464398 44104
rect 471058 43480 471114 43489
rect 471058 43415 471114 43424
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 464160 42764 464212 42770
rect 464160 42706 464212 42712
rect 463056 42492 463108 42498
rect 463988 42486 464050 42514
rect 463056 42434 463108 42440
rect 461950 42256 462006 42265
rect 464022 42228 464050 42486
rect 465828 42364 465856 43143
rect 461950 42191 462006 42200
rect 471072 42106 471100 43415
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42228 518848 42735
rect 661420 42187 661448 45526
rect 661408 42181 661460 42187
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 661408 42123 661460 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 426900 41472 426952 41478
rect 426900 41414 426952 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 40352 141754 40361
rect 141698 40287 141754 40296
rect 141712 39984 141740 40287
<< via2 >>
rect 185030 1002088 185086 1002144
rect 82174 1001952 82230 1002008
rect 133694 1001972 133750 1002008
rect 133694 1001952 133696 1001972
rect 133696 1001952 133748 1001972
rect 133748 1001952 133750 1001972
rect 81346 983456 81402 983512
rect 483018 1001952 483074 1002008
rect 534998 1001952 535054 1002008
rect 232962 997328 233018 997384
rect 240138 997192 240194 997248
rect 235906 990936 235962 990992
rect 238666 984000 238722 984056
rect 285402 997328 285458 997384
rect 292578 997328 292634 997384
rect 286966 987944 287022 988000
rect 235906 983728 235962 983784
rect 240138 983728 240194 983784
rect 286966 983728 287022 983784
rect 184938 983456 184994 983512
rect 132498 982504 132554 982560
rect 387522 997328 387578 997384
rect 389178 990936 389234 990992
rect 404358 997328 404414 997384
rect 292578 983728 292634 983784
rect 391938 983456 391994 983512
rect 394422 983492 394424 983512
rect 394424 983492 394476 983512
rect 394476 983492 394478 983512
rect 394422 983456 394478 983492
rect 399758 983456 399814 983512
rect 636198 1001952 636254 1002008
rect 535458 983728 535514 983784
rect 636198 983728 636254 983784
rect 483846 982524 483902 982560
rect 483846 982504 483848 982524
rect 483848 982504 483900 982524
rect 483900 982504 483902 982524
rect 289726 980872 289782 980928
rect 30102 960200 30158 960256
rect 651378 959132 651434 959168
rect 651378 959112 651380 959132
rect 651380 959112 651432 959132
rect 651432 959112 651434 959132
rect 677414 959132 677470 959168
rect 677414 959112 677416 959132
rect 677416 959112 677468 959132
rect 677468 959112 677470 959132
rect 63406 958976 63462 959032
rect 676034 897116 676090 897152
rect 676034 897096 676036 897116
rect 676036 897096 676088 897116
rect 676088 897096 676090 897116
rect 651470 868536 651526 868592
rect 675850 896688 675906 896744
rect 676034 896280 676090 896336
rect 652022 867584 652078 867640
rect 651470 866224 651526 866280
rect 651378 865172 651380 865192
rect 651380 865172 651432 865192
rect 651432 865172 651434 865192
rect 651378 865136 651434 865172
rect 651470 863812 651472 863832
rect 651472 863812 651524 863832
rect 651524 863812 651526 863832
rect 651470 863776 651526 863812
rect 651470 862280 651526 862336
rect 35622 817944 35678 818000
rect 35806 817264 35862 817320
rect 35438 816856 35494 816912
rect 35806 816040 35862 816096
rect 35622 815224 35678 815280
rect 35806 814408 35862 814464
rect 41326 813592 41382 813648
rect 40958 812776 41014 812832
rect 37922 811552 37978 811608
rect 34518 811144 34574 811200
rect 32586 810736 32642 810792
rect 31022 809920 31078 809976
rect 32586 802440 32642 802496
rect 36542 809512 36598 809568
rect 41326 812368 41382 812424
rect 41142 811960 41198 812016
rect 41970 810328 42026 810384
rect 41786 809920 41842 809976
rect 41326 809104 41382 809160
rect 41786 808696 41842 808752
rect 41142 808288 41198 808344
rect 41326 807492 41382 807528
rect 41326 807472 41328 807492
rect 41328 807472 41380 807492
rect 41380 807472 41382 807492
rect 41142 806656 41198 806712
rect 41326 806248 41382 806304
rect 41970 805568 42026 805624
rect 41786 805160 41842 805216
rect 40498 800708 40500 800728
rect 40500 800708 40552 800728
rect 40552 800708 40554 800728
rect 40498 800672 40554 800708
rect 39762 800536 39818 800592
rect 42154 800944 42210 801000
rect 42154 797272 42210 797328
rect 41786 796184 41842 796240
rect 41786 794824 41842 794880
rect 42154 794416 42210 794472
rect 41786 793056 41842 793112
rect 41786 790608 41842 790664
rect 41786 789384 41842 789440
rect 42246 789112 42302 789168
rect 42430 788704 42486 788760
rect 42246 788160 42302 788216
rect 35806 774696 35862 774752
rect 35254 773880 35310 773936
rect 35622 773472 35678 773528
rect 35438 773064 35494 773120
rect 35806 773100 35808 773120
rect 35808 773100 35860 773120
rect 35860 773100 35862 773120
rect 35806 773064 35862 773100
rect 41510 773064 41566 773120
rect 35622 772248 35678 772304
rect 40314 772248 40370 772304
rect 35806 771860 35862 771896
rect 35806 771840 35808 771860
rect 35808 771840 35860 771860
rect 35860 771840 35862 771860
rect 35806 771452 35862 771488
rect 35806 771432 35808 771452
rect 35808 771432 35860 771452
rect 35860 771432 35862 771452
rect 39946 771432 40002 771488
rect 35438 771024 35494 771080
rect 35622 770616 35678 770672
rect 35806 770208 35862 770264
rect 40314 770208 40370 770264
rect 35622 769392 35678 769448
rect 35806 768576 35862 768632
rect 35162 768168 35218 768224
rect 32402 767760 32458 767816
rect 33782 766944 33838 767000
rect 35806 767352 35862 767408
rect 35806 766536 35862 766592
rect 35622 765720 35678 765776
rect 35806 764496 35862 764552
rect 35622 764088 35678 764144
rect 35806 763680 35862 763736
rect 35806 762864 35862 762920
rect 39394 764496 39450 764552
rect 39946 764088 40002 764144
rect 39946 763272 40002 763328
rect 39946 758276 39948 758296
rect 39948 758276 40000 758296
rect 40000 758276 40002 758296
rect 39946 758240 40002 758276
rect 39670 757968 39726 758024
rect 36542 757696 36598 757752
rect 41786 757016 41842 757072
rect 41878 756608 41934 756664
rect 42614 758240 42670 758296
rect 42430 757968 42486 758024
rect 41878 754160 41934 754216
rect 42062 754024 42118 754080
rect 42154 753480 42210 753536
rect 42062 752936 42118 752992
rect 42062 751576 42118 751632
rect 42062 751168 42118 751224
rect 42062 750352 42118 750408
rect 41786 746680 41842 746736
rect 42982 753480 43038 753536
rect 42890 752936 42946 752992
rect 42614 745728 42670 745784
rect 42246 745456 42302 745512
rect 42614 745048 42670 745104
rect 40406 732264 40462 732320
rect 40038 731584 40094 731640
rect 35438 731312 35494 731368
rect 35806 730904 35862 730960
rect 35622 730496 35678 730552
rect 35438 729680 35494 729736
rect 35806 730088 35862 730144
rect 35622 729272 35678 729328
rect 35806 728864 35862 728920
rect 35806 728456 35862 728512
rect 35438 728048 35494 728104
rect 42982 731584 43038 731640
rect 41694 731076 41696 731096
rect 41696 731076 41748 731096
rect 41748 731076 41750 731096
rect 41694 731040 41750 731076
rect 41694 728184 41750 728240
rect 41694 727776 41750 727832
rect 43074 727776 43130 727832
rect 35622 727640 35678 727696
rect 35806 727232 35862 727288
rect 41142 726824 41198 726880
rect 41326 726416 41382 726472
rect 40958 725600 41014 725656
rect 41786 725600 41842 725656
rect 32402 725192 32458 725248
rect 31666 723968 31722 724024
rect 35162 724784 35218 724840
rect 37278 724376 37334 724432
rect 39302 723152 39358 723208
rect 37278 716896 37334 716952
rect 40590 715808 40646 715864
rect 41786 722336 41842 722392
rect 41786 718528 41842 718584
rect 42890 721112 42946 721168
rect 40958 714856 41014 714912
rect 39302 714176 39358 714232
rect 42430 715808 42486 715864
rect 42338 714856 42394 714912
rect 42246 714312 42302 714368
rect 42154 710776 42210 710832
rect 41786 709824 41842 709880
rect 42062 708464 42118 708520
rect 41786 707104 41842 707160
rect 42430 706288 42486 706344
rect 41786 704248 41842 704304
rect 42062 703024 42118 703080
rect 42614 703024 42670 703080
rect 41878 700440 41934 700496
rect 42522 701800 42578 701856
rect 42522 701528 42578 701584
rect 35438 688336 35494 688392
rect 35806 687656 35862 687712
rect 41694 687540 41750 687576
rect 41694 687520 41696 687540
rect 41696 687520 41748 687540
rect 41748 687520 41750 687540
rect 35622 687248 35678 687304
rect 35438 686840 35494 686896
rect 41694 687148 41696 687168
rect 41696 687148 41748 687168
rect 41748 687148 41750 687168
rect 41694 687112 41750 687148
rect 35806 686432 35862 686488
rect 35806 686024 35862 686080
rect 35806 685616 35862 685672
rect 35622 685208 35678 685264
rect 35806 684800 35862 684856
rect 41694 684684 41750 684720
rect 41694 684664 41696 684684
rect 41696 684664 41748 684684
rect 41748 684664 41750 684684
rect 35622 684392 35678 684448
rect 35438 683984 35494 684040
rect 41694 683848 41750 683904
rect 35806 683168 35862 683224
rect 41694 683068 41696 683088
rect 41696 683068 41748 683088
rect 41748 683068 41750 683088
rect 41694 683032 41750 683068
rect 35622 682760 35678 682816
rect 35162 681944 35218 682000
rect 33046 681536 33102 681592
rect 31022 680720 31078 680776
rect 33782 681128 33838 681184
rect 35806 682352 35862 682408
rect 41694 681400 41750 681456
rect 41694 680992 41750 681048
rect 35806 680312 35862 680368
rect 41694 680176 41750 680232
rect 35806 679904 35862 679960
rect 35622 679496 35678 679552
rect 41694 679396 41696 679416
rect 41696 679396 41748 679416
rect 41748 679396 41750 679416
rect 41694 679360 41750 679396
rect 35806 679124 35808 679144
rect 35808 679124 35860 679144
rect 35860 679124 35862 679144
rect 35806 679088 35862 679124
rect 41694 678988 41696 679008
rect 41696 678988 41748 679008
rect 41748 678988 41750 679008
rect 41694 678952 41750 678988
rect 42706 680992 42762 681048
rect 41694 678544 41750 678600
rect 33782 672696 33838 672752
rect 42246 672560 42302 672616
rect 41970 668480 42026 668536
rect 42062 667664 42118 667720
rect 42062 667120 42118 667176
rect 42062 666576 42118 666632
rect 41786 665080 41842 665136
rect 41786 663992 41842 664048
rect 41786 658280 41842 658336
rect 41786 657192 41842 657248
rect 42522 658552 42578 658608
rect 35806 644680 35862 644736
rect 38566 644272 38622 644328
rect 35346 643864 35402 643920
rect 35530 643456 35586 643512
rect 35806 643492 35808 643512
rect 35808 643492 35860 643512
rect 35860 643492 35862 643512
rect 35806 643456 35862 643492
rect 35438 642640 35494 642696
rect 35806 642640 35862 642696
rect 35622 642232 35678 642288
rect 35806 641416 35862 641472
rect 35622 641008 35678 641064
rect 35806 640600 35862 640656
rect 41142 641008 41198 641064
rect 40866 640192 40922 640248
rect 34426 639784 34482 639840
rect 39394 639784 39450 639840
rect 35530 639376 35586 639432
rect 35806 639376 35862 639432
rect 35622 638560 35678 638616
rect 32402 637744 32458 637800
rect 35162 637336 35218 637392
rect 32402 629856 32458 629912
rect 35806 638152 35862 638208
rect 35806 636928 35862 636984
rect 35530 636520 35586 636576
rect 35806 636520 35862 636576
rect 35806 635704 35862 635760
rect 35806 634480 35862 634536
rect 35806 633664 35862 633720
rect 39118 636148 39120 636168
rect 39120 636148 39172 636168
rect 39172 636148 39174 636168
rect 39118 636112 39174 636148
rect 40038 636556 40040 636576
rect 40040 636556 40092 636576
rect 40092 636556 40094 636576
rect 40038 636520 40094 636556
rect 39578 635704 39634 635760
rect 40130 634072 40186 634128
rect 41602 633256 41658 633312
rect 40590 632848 40646 632904
rect 40038 630808 40094 630864
rect 42062 633256 42118 633312
rect 39302 629176 39358 629232
rect 39394 628668 39396 628688
rect 39396 628668 39448 628688
rect 39448 628668 39450 628688
rect 39394 628632 39450 628668
rect 41786 627408 41842 627464
rect 41786 627136 41842 627192
rect 42614 632848 42670 632904
rect 42614 628632 42670 628688
rect 42154 624552 42210 624608
rect 41786 621968 41842 622024
rect 42154 621968 42210 622024
rect 41786 620744 41842 620800
rect 42338 615712 42394 615768
rect 42614 615440 42670 615496
rect 41878 613400 41934 613456
rect 43074 684664 43130 684720
rect 43074 634072 43130 634128
rect 42890 614216 42946 614272
rect 42246 612348 42248 612368
rect 42248 612348 42300 612368
rect 42300 612348 42302 612368
rect 42246 612312 42302 612348
rect 43626 797272 43682 797328
rect 43442 772248 43498 772304
rect 44270 771432 44326 771488
rect 43626 770208 43682 770264
rect 43442 753752 43498 753808
rect 43902 754024 43958 754080
rect 45098 773064 45154 773120
rect 44454 764496 44510 764552
rect 44638 764088 44694 764144
rect 44454 753480 44510 753536
rect 44914 763272 44970 763328
rect 44638 751168 44694 751224
rect 44270 728184 44326 728240
rect 43810 723560 43866 723616
rect 43626 720296 43682 720352
rect 43626 710776 43682 710832
rect 43442 683848 43498 683904
rect 43442 677864 43498 677920
rect 44730 721520 44786 721576
rect 44730 708464 44786 708520
rect 44454 680176 44510 680232
rect 44270 679360 44326 679416
rect 43810 678544 43866 678600
rect 43994 677048 44050 677104
rect 44086 667664 44142 667720
rect 44270 666576 44326 666632
rect 44730 678952 44786 679008
rect 44730 667120 44786 667176
rect 44546 641008 44602 641064
rect 44362 639784 44418 639840
rect 43810 636520 43866 636576
rect 43626 630808 43682 630864
rect 43442 611088 43498 611144
rect 44178 636112 44234 636168
rect 43994 635704 44050 635760
rect 44178 624552 44234 624608
rect 44178 621968 44234 622024
rect 44086 614216 44142 614272
rect 43764 611768 43820 611824
rect 43994 611360 44050 611416
rect 43626 610680 43682 610736
rect 40314 601976 40370 602032
rect 35806 601724 35862 601760
rect 35806 601704 35808 601724
rect 35808 601704 35860 601724
rect 35860 601704 35862 601724
rect 35162 595754 35218 595810
rect 33046 595176 33102 595232
rect 31022 594360 31078 594416
rect 33782 593544 33838 593600
rect 35622 591912 35678 591968
rect 35806 591504 35862 591560
rect 39946 601296 40002 601352
rect 40130 600888 40186 600944
rect 37922 594530 37978 594586
rect 36542 589600 36598 589656
rect 45282 751576 45338 751632
rect 45098 732264 45154 732320
rect 46202 731040 46258 731096
rect 45098 722744 45154 722800
rect 45466 687520 45522 687576
rect 45098 683032 45154 683088
rect 46202 687112 46258 687168
rect 45098 640192 45154 640248
rect 44730 611108 44786 611144
rect 44730 611088 44732 611108
rect 44732 611088 44784 611108
rect 44784 611088 44786 611108
rect 44730 610716 44732 610736
rect 44732 610716 44784 610736
rect 44784 610716 44786 610736
rect 44730 610680 44786 610716
rect 44546 600480 44602 600536
rect 44638 600072 44694 600128
rect 44454 599664 44510 599720
rect 42890 597624 42946 597680
rect 40958 596808 41014 596864
rect 41142 596400 41198 596456
rect 41326 595754 41382 595810
rect 41694 595756 41696 595776
rect 41696 595756 41748 595776
rect 41748 595756 41750 595776
rect 41694 595720 41750 595756
rect 41694 594532 41696 594552
rect 41696 594532 41748 594552
rect 41748 594532 41750 594552
rect 41694 594496 41750 594532
rect 41694 592048 41750 592104
rect 39762 589328 39818 589384
rect 37922 585112 37978 585168
rect 41694 590416 41750 590472
rect 43074 596944 43130 597000
rect 40590 585928 40646 585984
rect 40406 585656 40462 585712
rect 42430 585928 42486 585984
rect 39854 584568 39910 584624
rect 41786 580216 41842 580272
rect 42246 580216 42302 580272
rect 41970 578856 42026 578912
rect 42246 578448 42302 578504
rect 41786 577768 41842 577824
rect 42246 575864 42302 575920
rect 41970 573824 42026 573880
rect 42614 573280 42670 573336
rect 42062 571512 42118 571568
rect 42430 571376 42486 571432
rect 41786 570152 41842 570208
rect 39854 559000 39910 559056
rect 42798 559000 42854 559056
rect 35806 558048 35862 558104
rect 35806 555600 35862 555656
rect 35806 554804 35862 554840
rect 44362 593136 44418 593192
rect 43258 590416 43314 590472
rect 43442 589328 43498 589384
rect 40498 558728 40554 558784
rect 43074 558728 43130 558784
rect 35806 554784 35808 554804
rect 35808 554784 35860 554804
rect 35860 554784 35862 554804
rect 35622 554376 35678 554432
rect 35806 553560 35862 553616
rect 37922 553352 37978 553408
rect 29642 551928 29698 551984
rect 41694 553016 41750 553072
rect 43166 553016 43222 553072
rect 41326 552336 41382 552392
rect 41694 551792 41750 551848
rect 41142 551112 41198 551168
rect 42062 550160 42118 550216
rect 40498 549480 40554 549536
rect 39210 547440 39266 547496
rect 41326 548256 41382 548312
rect 41786 549888 41842 549944
rect 41694 547712 41750 547768
rect 41510 545536 41566 545592
rect 40498 545264 40554 545320
rect 42798 549072 42854 549128
rect 39210 543632 39266 543688
rect 37922 542272 37978 542328
rect 42614 539552 42670 539608
rect 42430 538192 42486 538248
rect 42062 537376 42118 537432
rect 42062 536968 42118 537024
rect 42614 536968 42670 537024
rect 42062 535608 42118 535664
rect 41786 535200 41842 535256
rect 42706 536696 42762 536752
rect 42706 535608 42762 535664
rect 42430 533840 42486 533896
rect 42706 533568 42762 533624
rect 42246 533296 42302 533352
rect 42522 532616 42578 532672
rect 42614 530032 42670 530088
rect 42706 528944 42762 529000
rect 42706 528672 42762 528728
rect 42890 527176 42946 527232
rect 35806 430072 35862 430128
rect 35806 428440 35862 428496
rect 43166 427352 43222 427408
rect 42154 427080 42210 427136
rect 41970 426536 42026 426592
rect 42890 426536 42946 426592
rect 40958 426400 41014 426456
rect 39302 425584 39358 425640
rect 32770 424768 32826 424824
rect 34518 424360 34574 424416
rect 33782 423952 33838 424008
rect 41142 425992 41198 426048
rect 41786 422320 41842 422376
rect 41326 419872 41382 419928
rect 41326 418784 41382 418840
rect 41786 418512 41842 418568
rect 42154 421504 42210 421560
rect 43074 425176 43130 425232
rect 42154 418240 42210 418296
rect 40958 417696 41014 417752
rect 39302 415248 39358 415304
rect 33782 414568 33838 414624
rect 41786 413480 41842 413536
rect 41786 413072 41842 413128
rect 42246 409808 42302 409864
rect 42062 408040 42118 408096
rect 42430 407224 42486 407280
rect 41786 406952 41842 407008
rect 41786 406680 41842 406736
rect 42430 404912 42486 404968
rect 42246 404504 42302 404560
rect 42338 402872 42394 402928
rect 41786 400016 41842 400072
rect 41786 399336 41842 399392
rect 41970 398792 42026 398848
rect 42154 395664 42210 395720
rect 41326 387096 41382 387152
rect 41142 386688 41198 386744
rect 40958 385872 41014 385928
rect 41142 385872 41198 385928
rect 41142 383016 41198 383072
rect 40038 382200 40094 382256
rect 40958 382200 41014 382256
rect 35438 381792 35494 381848
rect 33966 380976 34022 381032
rect 39302 381384 39358 381440
rect 35806 379344 35862 379400
rect 35806 378156 35808 378176
rect 35808 378156 35860 378176
rect 35860 378156 35862 378176
rect 35806 378120 35862 378156
rect 35806 376488 35862 376544
rect 35806 376080 35862 376136
rect 35438 374584 35494 374640
rect 41326 382608 41382 382664
rect 41142 381792 41198 381848
rect 41326 379772 41382 379808
rect 41326 379752 41328 379772
rect 41328 379752 41380 379772
rect 41380 379752 41382 379772
rect 41510 379772 41566 379808
rect 41510 379752 41512 379772
rect 41512 379752 41564 379772
rect 41564 379752 41566 379772
rect 40038 379344 40094 379400
rect 42982 417696 43038 417752
rect 42798 385600 42854 385656
rect 43258 385192 43314 385248
rect 41878 381520 41934 381576
rect 42890 380704 42946 380760
rect 41694 378156 41696 378176
rect 41696 378156 41748 378176
rect 41748 378156 41750 378176
rect 41694 378120 41750 378156
rect 40406 376896 40462 376952
rect 41786 364792 41842 364848
rect 41786 364112 41842 364168
rect 42062 363568 42118 363624
rect 42706 363024 42762 363080
rect 42430 362208 42486 362264
rect 41786 360032 41842 360088
rect 42154 359896 42210 359952
rect 42430 358944 42486 359000
rect 41878 358672 41934 358728
rect 41786 356904 41842 356960
rect 43074 376896 43130 376952
rect 42430 355952 42486 356008
rect 41878 355680 41934 355736
rect 44362 579672 44418 579728
rect 44914 599256 44970 599312
rect 44638 559272 44694 559328
rect 44546 556824 44602 556880
rect 44362 555192 44418 555248
rect 43994 551792 44050 551848
rect 43810 550704 43866 550760
rect 43626 547712 43682 547768
rect 44178 548664 44234 548720
rect 44178 536832 44234 536888
rect 43994 533840 44050 533896
rect 43810 533568 43866 533624
rect 45098 598848 45154 598904
rect 45282 598032 45338 598088
rect 45098 580216 45154 580272
rect 44914 556416 44970 556472
rect 45006 556008 45062 556064
rect 44730 537376 44786 537432
rect 44822 527176 44878 527232
rect 44822 430888 44878 430944
rect 44546 429664 44602 429720
rect 44638 429256 44694 429312
rect 44362 428032 44418 428088
rect 44454 427624 44510 427680
rect 44270 426808 44326 426864
rect 43810 422728 43866 422784
rect 43994 421096 44050 421152
rect 43810 409808 43866 409864
rect 43994 408040 44050 408096
rect 45190 551520 45246 551576
rect 45374 550432 45430 550488
rect 45374 539552 45430 539608
rect 45190 528944 45246 529000
rect 45006 428848 45062 428904
rect 45098 423136 45154 423192
rect 45466 420688 45522 420744
rect 45282 407224 45338 407280
rect 45098 402872 45154 402928
rect 44638 386416 44694 386472
rect 44454 384784 44510 384840
rect 45098 384376 45154 384432
rect 44270 383968 44326 384024
rect 44914 382200 44970 382256
rect 44638 380296 44694 380352
rect 43810 379752 43866 379808
rect 43994 378120 44050 378176
rect 44270 377440 44326 377496
rect 43994 363568 44050 363624
rect 43810 359896 43866 359952
rect 43626 354728 43682 354784
rect 43442 354184 43498 354240
rect 44638 358944 44694 359000
rect 44638 355952 44694 356008
rect 44454 354456 44510 354512
rect 44730 354184 44786 354240
rect 44270 353096 44326 353152
rect 40222 345480 40278 345536
rect 43258 345480 43314 345536
rect 35806 344256 35862 344312
rect 35622 343848 35678 343904
rect 33046 343440 33102 343496
rect 35806 342252 35808 342272
rect 35808 342252 35860 342272
rect 35860 342252 35862 342272
rect 35806 342216 35862 342252
rect 39854 342216 39910 342272
rect 44914 343304 44970 343360
rect 39854 341808 39910 341864
rect 40038 341808 40094 341864
rect 35806 341400 35862 341456
rect 35806 341028 35808 341048
rect 35808 341028 35860 341048
rect 35860 341028 35862 341048
rect 35806 340992 35862 341028
rect 39486 340992 39542 341048
rect 35530 339768 35586 339824
rect 35806 339768 35862 339824
rect 35806 336096 35862 336152
rect 35806 334464 35862 334520
rect 40222 341420 40278 341456
rect 40222 341400 40224 341420
rect 40224 341400 40276 341420
rect 40276 341400 40278 341420
rect 45282 383560 45338 383616
rect 40222 340992 40278 341048
rect 45098 340992 45154 341048
rect 45650 363024 45706 363080
rect 45834 354728 45890 354784
rect 45650 354340 45706 354376
rect 45650 354320 45652 354340
rect 45652 354320 45704 354340
rect 45704 354320 45706 354340
rect 45466 353640 45522 353696
rect 45466 353404 45468 353424
rect 45468 353404 45520 353424
rect 45520 353404 45522 353424
rect 45466 353368 45522 353404
rect 45420 353132 45422 353152
rect 45422 353132 45474 353152
rect 45474 353132 45476 353152
rect 45420 353096 45476 353132
rect 45466 341420 45522 341456
rect 45466 341400 45468 341420
rect 45468 341400 45520 341420
rect 45520 341400 45522 341420
rect 40038 340584 40094 340640
rect 45282 340584 45338 340640
rect 39670 340176 39726 340232
rect 39854 340176 39910 340232
rect 39670 339768 39726 339824
rect 45650 339224 45706 339280
rect 45466 337592 45522 337648
rect 39486 337320 39542 337376
rect 38658 336504 38714 336560
rect 43994 334600 44050 334656
rect 44270 334600 44326 334656
rect 40222 334464 40278 334520
rect 43074 334464 43130 334520
rect 39762 332832 39818 332888
rect 42890 332832 42946 332888
rect 37922 331200 37978 331256
rect 41786 324808 41842 324864
rect 42246 324264 42302 324320
rect 41786 321136 41842 321192
rect 41786 319912 41842 319968
rect 42246 319912 42302 319968
rect 42614 320592 42670 320648
rect 42430 319368 42486 319424
rect 41786 317328 41842 317384
rect 42430 316376 42486 316432
rect 41786 315968 41842 316024
rect 41786 313656 41842 313712
rect 42430 313112 42486 313168
rect 42430 312840 42486 312896
rect 42154 312568 42210 312624
rect 42154 311752 42210 311808
rect 41326 301552 41382 301608
rect 41142 300872 41198 300928
rect 42154 298696 42210 298752
rect 42338 297336 42394 297392
rect 43166 297064 43222 297120
rect 41142 296384 41198 296440
rect 42798 295976 42854 296032
rect 41326 295160 41382 295216
rect 33782 294752 33838 294808
rect 32402 293936 32458 293992
rect 41326 293528 41382 293584
rect 39946 290264 40002 290320
rect 32402 284824 32458 284880
rect 42430 281424 42486 281480
rect 42062 278432 42118 278488
rect 42154 277888 42210 277944
rect 41786 277072 41842 277128
rect 42982 293120 43038 293176
rect 43350 292712 43406 292768
rect 42614 275848 42670 275904
rect 41786 274216 41842 274272
rect 42338 273128 42394 273184
rect 41786 272992 41842 273048
rect 41786 272312 41842 272368
rect 41786 270408 41842 270464
rect 41786 269728 41842 269784
rect 42154 267688 42210 267744
rect 43442 277888 43498 277944
rect 43626 273128 43682 273184
rect 43442 269728 43498 269784
rect 35806 257080 35862 257136
rect 40498 257080 40554 257136
rect 43350 257080 43406 257136
rect 35622 256264 35678 256320
rect 40222 256264 40278 256320
rect 42982 256264 43038 256320
rect 35806 255856 35862 255912
rect 39578 255484 39580 255504
rect 39580 255484 39632 255504
rect 39632 255484 39634 255504
rect 39578 255448 39634 255484
rect 35806 254224 35862 254280
rect 39854 254224 39910 254280
rect 43074 255448 43130 255504
rect 42890 254224 42946 254280
rect 35622 253408 35678 253464
rect 35806 253000 35862 253056
rect 35806 252184 35862 252240
rect 35806 250552 35862 250608
rect 35806 247696 35862 247752
rect 39762 245656 39818 245712
rect 41694 246472 41750 246528
rect 42062 240080 42118 240136
rect 41970 238448 42026 238504
rect 42338 238040 42394 238096
rect 41786 236544 41842 236600
rect 41786 234640 41842 234696
rect 42338 233824 42394 233880
rect 42430 232192 42486 232248
rect 42430 231784 42486 231840
rect 42430 231512 42486 231568
rect 42154 230424 42210 230480
rect 41970 227296 42026 227352
rect 42430 225664 42486 225720
rect 41694 224440 41750 224496
rect 35530 217912 35586 217968
rect 39946 216416 40002 216472
rect 39578 216144 39634 216200
rect 35530 214240 35586 214296
rect 35806 214240 35862 214296
rect 35622 213424 35678 213480
rect 35806 213016 35862 213072
rect 42614 224848 42670 224904
rect 42154 223488 42210 223544
rect 43442 246472 43498 246528
rect 43258 245656 43314 245712
rect 43074 216416 43130 216472
rect 42890 216144 42946 216200
rect 44270 319912 44326 319968
rect 45282 320592 45338 320648
rect 45282 312840 45338 312896
rect 45650 312568 45706 312624
rect 45466 311752 45522 311808
rect 45190 300464 45246 300520
rect 44362 299648 44418 299704
rect 44178 298968 44234 299024
rect 44638 298016 44694 298072
rect 44362 256808 44418 256864
rect 44178 255992 44234 256048
rect 45006 292576 45062 292632
rect 45466 292576 45522 292632
rect 45190 291488 45246 291544
rect 45006 281424 45062 281480
rect 45190 278432 45246 278488
rect 44822 258032 44878 258088
rect 44638 255176 44694 255232
rect 44270 254768 44326 254824
rect 43994 231104 44050 231160
rect 35806 210160 35862 210216
rect 35622 209344 35678 209400
rect 35806 208936 35862 208992
rect 40406 208936 40462 208992
rect 42890 208936 42946 208992
rect 35806 208548 35862 208584
rect 35806 208528 35808 208548
rect 35808 208528 35860 208548
rect 35860 208528 35862 208548
rect 40038 208120 40094 208176
rect 35806 207304 35862 207360
rect 35806 205264 35862 205320
rect 35806 204448 35862 204504
rect 40590 206896 40646 206952
rect 42706 206896 42762 206952
rect 41510 204484 41512 204504
rect 41512 204484 41564 204504
rect 41564 204484 41566 204504
rect 41510 204448 41566 204484
rect 41694 204040 41750 204096
rect 35806 203632 35862 203688
rect 39946 203632 40002 203688
rect 37922 198736 37978 198792
rect 44914 253952 44970 254008
rect 44546 251504 44602 251560
rect 44730 250280 44786 250336
rect 44546 240080 44602 240136
rect 45558 252728 45614 252784
rect 45098 249056 45154 249112
rect 44638 230424 44694 230480
rect 44270 212064 44326 212120
rect 45006 231512 45062 231568
rect 45834 248648 45890 248704
rect 46018 248240 46074 248296
rect 46018 233144 46074 233200
rect 45834 231784 45890 231840
rect 46938 578176 46994 578232
rect 47582 558456 47638 558512
rect 47582 489912 47638 489968
rect 46386 376080 46442 376136
rect 46938 338816 46994 338872
rect 47122 337864 47178 337920
rect 47122 324264 47178 324320
rect 46938 313112 46994 313168
rect 47766 430480 47822 430536
rect 47766 387640 47822 387696
rect 47766 354320 47822 354376
rect 47582 290672 47638 290728
rect 46386 257624 46442 257680
rect 47214 251912 47270 251968
rect 46938 251096 46994 251152
rect 45558 225664 45614 225720
rect 47398 247016 47454 247072
rect 47398 238448 47454 238504
rect 47214 232192 47270 232248
rect 46938 224848 46994 224904
rect 44822 211248 44878 211304
rect 44454 208392 44510 208448
rect 44178 207712 44234 207768
rect 43718 204448 43774 204504
rect 43442 204040 43498 204096
rect 43258 203632 43314 203688
rect 42430 197240 42486 197296
rect 41970 195608 42026 195664
rect 41786 195200 41842 195256
rect 42246 194928 42302 194984
rect 41786 193432 41842 193488
rect 42062 191528 42118 191584
rect 42430 190440 42486 190496
rect 42246 187584 42302 187640
rect 41786 186360 41842 186416
rect 41786 185952 41842 186008
rect 43718 190440 43774 190496
rect 42430 183504 42486 183560
rect 42246 183232 42302 183288
rect 42062 180784 42118 180840
rect 43902 183504 43958 183560
rect 44638 205944 44694 206000
rect 44454 197240 44510 197296
rect 44822 205128 44878 205184
rect 46202 204856 46258 204912
rect 44822 191528 44878 191584
rect 44638 187584 44694 187640
rect 44178 183232 44234 183288
rect 47766 247424 47822 247480
rect 49330 418784 49386 418840
rect 49146 334056 49202 334112
rect 62210 790472 62266 790528
rect 62118 789148 62120 789168
rect 62120 789148 62172 789168
rect 62172 789148 62174 789168
rect 62118 789112 62174 789148
rect 62118 787344 62174 787400
rect 62302 786120 62358 786176
rect 62118 784896 62174 784952
rect 51722 538192 51778 538248
rect 51446 404912 51502 404968
rect 51078 395664 51134 395720
rect 51078 362208 51134 362264
rect 51906 353640 51962 353696
rect 50526 291080 50582 291136
rect 55862 611632 55918 611688
rect 53102 264696 53158 264752
rect 57242 278024 57298 278080
rect 57426 275848 57482 275904
rect 62118 746136 62174 746192
rect 62118 744096 62174 744152
rect 62118 743724 62120 743744
rect 62120 743724 62172 743744
rect 62172 743724 62174 743744
rect 62118 743688 62174 743724
rect 62118 742364 62120 742384
rect 62120 742364 62172 742384
rect 62172 742364 62174 742384
rect 62118 742328 62174 742364
rect 62118 704384 62174 704440
rect 62118 703296 62174 703352
rect 61382 699624 61438 699680
rect 62210 697992 62266 698048
rect 62118 660900 62120 660920
rect 62120 660900 62172 660920
rect 62172 660900 62174 660920
rect 62118 660864 62174 660900
rect 61382 659504 61438 659560
rect 62118 658280 62174 658336
rect 62118 656512 62174 656568
rect 62118 655288 62174 655344
rect 60002 278296 60058 278352
rect 62118 616528 62174 616584
rect 62118 614624 62174 614680
rect 61382 613808 61438 613864
rect 62118 612620 62120 612640
rect 62120 612620 62172 612640
rect 62172 612620 62174 612640
rect 62118 612584 62174 612620
rect 60186 277344 60242 277400
rect 60370 267688 60426 267744
rect 62486 590008 62542 590064
rect 62118 574776 62174 574832
rect 62118 573552 62174 573608
rect 62486 569880 62542 569936
rect 62486 556688 62542 556744
rect 62118 531120 62174 531176
rect 62302 530576 62358 530632
rect 62118 528572 62120 528592
rect 62120 528572 62172 528592
rect 62172 528572 62174 528592
rect 62118 528536 62174 528572
rect 62486 527992 62542 528048
rect 62118 527076 62120 527096
rect 62120 527076 62172 527096
rect 62172 527076 62174 527096
rect 62118 527040 62174 527076
rect 62486 427080 62542 427136
rect 62118 404096 62174 404152
rect 62118 402600 62174 402656
rect 62118 400560 62174 400616
rect 62486 400152 62542 400208
rect 62118 399336 62174 399392
rect 62118 398248 62174 398304
rect 62486 385872 62542 385928
rect 62118 360848 62174 360904
rect 62118 359760 62174 359816
rect 62118 357720 62174 357776
rect 62486 357312 62542 357368
rect 62118 355988 62120 356008
rect 62120 355988 62172 356008
rect 62172 355988 62174 356008
rect 62118 355952 62174 355988
rect 62486 341672 62542 341728
rect 61566 319368 61622 319424
rect 62118 317364 62120 317384
rect 62120 317364 62172 317384
rect 62172 317364 62174 317384
rect 62118 317328 62174 317364
rect 61566 315968 61622 316024
rect 62118 314764 62174 314800
rect 62118 314744 62120 314764
rect 62120 314744 62172 314764
rect 62172 314744 62174 314764
rect 62302 314064 62358 314120
rect 62486 312976 62542 313032
rect 62486 297336 62542 297392
rect 62118 295704 62174 295760
rect 62118 294092 62174 294128
rect 62118 294072 62120 294092
rect 62120 294072 62172 294092
rect 62172 294072 62174 294092
rect 62302 292712 62358 292768
rect 62118 292460 62174 292496
rect 62118 292440 62120 292460
rect 62120 292440 62172 292460
rect 62172 292440 62174 292460
rect 62486 290944 62542 291000
rect 62210 288496 62266 288552
rect 62394 287136 62450 287192
rect 62118 285912 62174 285968
rect 62118 283192 62174 283248
rect 62118 280880 62174 280936
rect 62394 269728 62450 269784
rect 58622 223488 58678 223544
rect 56046 217912 56102 217968
rect 62946 787072 63002 787128
rect 651470 778368 651526 778424
rect 652022 777008 652078 777064
rect 651470 776056 651526 776112
rect 651378 775276 651380 775296
rect 651380 775276 651432 775296
rect 651432 775276 651434 775296
rect 651378 775240 651434 775276
rect 651470 774172 651526 774208
rect 651470 774152 651472 774172
rect 651472 774152 651524 774172
rect 651524 774152 651526 774172
rect 651470 773336 651526 773392
rect 62946 747632 63002 747688
rect 63038 741784 63094 741840
rect 651470 734168 651526 734224
rect 652666 732808 652722 732864
rect 651470 731720 651526 731776
rect 651378 731076 651380 731096
rect 651380 731076 651432 731096
rect 651432 731076 651434 731096
rect 651378 731040 651434 731076
rect 651470 729816 651526 729872
rect 651470 728492 651472 728512
rect 651472 728492 651524 728512
rect 651524 728492 651526 728512
rect 651470 728456 651526 728492
rect 62946 701256 63002 701312
rect 63130 700848 63186 700904
rect 651470 689424 651526 689480
rect 651654 688744 651710 688800
rect 651470 687384 651526 687440
rect 651470 686704 651526 686760
rect 651470 685208 651526 685264
rect 652574 684392 652630 684448
rect 62946 657600 63002 657656
rect 651470 643184 651526 643240
rect 652022 641824 652078 641880
rect 651470 640736 651526 640792
rect 651378 640092 651380 640112
rect 651380 640092 651432 640112
rect 651432 640092 651434 640112
rect 651378 640056 651434 640092
rect 651470 638560 651526 638616
rect 651654 638152 651710 638208
rect 63130 618024 63186 618080
rect 62946 612040 63002 612096
rect 64142 611360 64198 611416
rect 63314 595720 63370 595776
rect 63130 594088 63186 594144
rect 62946 590688 63002 590744
rect 63314 571104 63370 571160
rect 63130 568520 63186 568576
rect 63314 550160 63370 550216
rect 63314 525680 63370 525736
rect 63314 381520 63370 381576
rect 63314 354456 63370 354512
rect 63130 341400 63186 341456
rect 63406 332560 63462 332616
rect 63130 311752 63186 311808
rect 63130 298696 63186 298752
rect 63130 289720 63186 289776
rect 63222 284552 63278 284608
rect 62854 282104 62910 282160
rect 63130 280336 63186 280392
rect 62946 278840 63002 278896
rect 62670 224168 62726 224224
rect 651470 597896 651526 597952
rect 651470 596672 651526 596728
rect 651470 595312 651526 595368
rect 651654 595040 651710 595096
rect 651470 594088 651526 594144
rect 651470 592864 651526 592920
rect 651470 553424 651526 553480
rect 651654 552064 651710 552120
rect 651470 551112 651526 551168
rect 651378 550332 651380 550352
rect 651380 550332 651432 550352
rect 651432 550332 651434 550352
rect 651378 550296 651434 550332
rect 651470 549228 651526 549264
rect 651470 549208 651472 549228
rect 651472 549208 651524 549228
rect 651524 549208 651526 549228
rect 651470 548392 651526 548448
rect 64326 353368 64382 353424
rect 667662 698264 667718 698320
rect 667478 645768 667534 645824
rect 667294 600888 667350 600944
rect 668214 687792 668270 687848
rect 668858 730088 668914 730144
rect 669594 735664 669650 735720
rect 669410 728728 669466 728784
rect 669042 689424 669098 689480
rect 671250 733760 671306 733816
rect 670882 695816 670938 695872
rect 669778 685752 669834 685808
rect 668766 594768 668822 594824
rect 668582 562264 668638 562320
rect 668950 593408 669006 593464
rect 669594 644272 669650 644328
rect 670606 685480 670662 685536
rect 671986 713224 672042 713280
rect 671986 712408 672042 712464
rect 675850 895464 675906 895520
rect 676034 894648 676090 894704
rect 675850 893832 675906 893888
rect 676034 893016 676090 893072
rect 676034 892608 676090 892664
rect 676034 891384 676090 891440
rect 675298 890976 675354 891032
rect 676034 890160 676090 890216
rect 676034 889344 676090 889400
rect 676034 888956 676090 888992
rect 676034 888936 676036 888956
rect 676036 888936 676088 888956
rect 676088 888936 676090 888956
rect 676034 888548 676090 888584
rect 676034 888528 676036 888548
rect 676036 888528 676088 888548
rect 676088 888528 676090 888548
rect 676034 887324 676090 887360
rect 676034 887304 676036 887324
rect 676036 887304 676088 887324
rect 676088 887304 676090 887324
rect 676034 886916 676090 886952
rect 676034 886896 676036 886916
rect 676036 886896 676088 886916
rect 676088 886896 676090 886916
rect 679622 891792 679678 891848
rect 675666 878464 675722 878520
rect 676034 885692 676090 885728
rect 676034 885672 676036 885692
rect 676036 885672 676088 885692
rect 676088 885672 676090 885692
rect 678242 889752 678298 889808
rect 681002 890568 681058 890624
rect 683118 888120 683174 888176
rect 681002 880640 681058 880696
rect 683118 880368 683174 880424
rect 675206 877104 675262 877160
rect 674838 874656 674894 874712
rect 675482 874656 675538 874712
rect 675574 874112 675630 874168
rect 675758 873024 675814 873080
rect 675022 872752 675078 872808
rect 675390 870440 675446 870496
rect 675298 865680 675354 865736
rect 675758 865408 675814 865464
rect 675666 865000 675722 865056
rect 675758 788024 675814 788080
rect 675114 786664 675170 786720
rect 675390 786664 675446 786720
rect 673274 777416 673330 777472
rect 672538 713632 672594 713688
rect 672446 669976 672502 670032
rect 673458 734304 673514 734360
rect 673274 716488 673330 716544
rect 673274 716080 673330 716136
rect 673090 715708 673092 715728
rect 673092 715708 673144 715728
rect 673144 715708 673146 715728
rect 673090 715672 673146 715708
rect 673090 715300 673092 715320
rect 673092 715300 673144 715320
rect 673144 715300 673146 715320
rect 673090 715264 673146 715300
rect 673090 714992 673146 715048
rect 673274 714484 673276 714504
rect 673276 714484 673328 714504
rect 673328 714484 673330 714504
rect 673274 714448 673330 714484
rect 673274 714040 673330 714096
rect 673274 712816 673330 712872
rect 673274 711592 673330 711648
rect 673274 710368 673330 710424
rect 673090 709996 673092 710016
rect 673092 709996 673144 710016
rect 673144 709996 673146 710016
rect 673090 709960 673146 709996
rect 673274 709180 673276 709200
rect 673276 709180 673328 709200
rect 673328 709180 673330 709200
rect 673274 709144 673330 709180
rect 673274 708736 673330 708792
rect 672814 708328 672870 708384
rect 673274 705372 673276 705392
rect 673276 705372 673328 705392
rect 673328 705372 673330 705392
rect 673274 705336 673330 705372
rect 672630 669432 672686 669488
rect 672262 663992 672318 664048
rect 673274 696904 673330 696960
rect 673090 686160 673146 686216
rect 672906 662904 672962 662960
rect 671250 645496 671306 645552
rect 671250 641416 671306 641472
rect 671986 652432 672042 652488
rect 671710 647808 671766 647864
rect 671342 638560 671398 638616
rect 671434 624144 671490 624200
rect 670422 551520 670478 551576
rect 670422 549616 670478 549672
rect 669778 455368 669834 455424
rect 670974 607688 671030 607744
rect 672814 649168 672870 649224
rect 670606 455096 670662 455152
rect 657542 403280 657598 403336
rect 652022 400832 652078 400888
rect 651470 373224 651526 373280
rect 652206 396616 652262 396672
rect 654782 382880 654838 382936
rect 652206 373904 652262 373960
rect 652022 372136 652078 372192
rect 670514 392536 670570 392592
rect 651470 370640 651526 370696
rect 655518 366288 655574 366344
rect 654782 358536 654838 358592
rect 652022 356632 652078 356688
rect 651378 328072 651434 328128
rect 652390 351056 652446 351112
rect 653402 338680 653458 338736
rect 652390 329704 652446 329760
rect 652022 326848 652078 326904
rect 651378 325644 651434 325680
rect 669410 347248 669466 347304
rect 651378 325624 651380 325644
rect 651380 325624 651432 325644
rect 651432 325624 651434 325644
rect 653402 313248 653458 313304
rect 652298 309848 652354 309904
rect 651378 303320 651434 303376
rect 658922 311888 658978 311944
rect 652298 302096 652354 302152
rect 651470 300600 651526 300656
rect 651470 298696 651526 298752
rect 652390 297472 652446 297528
rect 652206 296812 652262 296848
rect 652206 296792 652208 296812
rect 652208 296792 652260 296812
rect 652260 296792 652262 296812
rect 651654 295296 651710 295352
rect 651470 294208 651526 294264
rect 651470 292984 651526 293040
rect 651654 291760 651710 291816
rect 652114 291488 652170 291544
rect 651470 290400 651526 290456
rect 651654 289176 651710 289232
rect 651470 288632 651526 288688
rect 651654 287680 651710 287736
rect 651470 287408 651526 287464
rect 651470 285912 651526 285968
rect 651470 284688 651526 284744
rect 651470 283328 651526 283384
rect 652022 282104 652078 282160
rect 651470 280880 651526 280936
rect 136638 270444 136640 270464
rect 136640 270444 136692 270464
rect 136692 270444 136694 270464
rect 136638 270408 136694 270444
rect 137834 270444 137836 270464
rect 137836 270444 137888 270464
rect 137888 270444 137890 270464
rect 137834 270408 137890 270444
rect 459374 272620 459376 272640
rect 459376 272620 459428 272640
rect 459428 272620 459430 272640
rect 459374 272584 459430 272620
rect 464710 272312 464766 272368
rect 466090 272584 466146 272640
rect 470690 272484 470692 272504
rect 470692 272484 470744 272504
rect 470744 272484 470746 272504
rect 470690 272448 470746 272484
rect 470598 271904 470654 271960
rect 478050 271904 478106 271960
rect 479522 271904 479578 271960
rect 483018 271904 483074 271960
rect 500866 272176 500922 272232
rect 501602 271904 501658 271960
rect 504546 272212 504548 272232
rect 504548 272212 504600 272232
rect 504600 272212 504602 272232
rect 504546 272176 504602 272212
rect 504546 271940 504548 271960
rect 504548 271940 504600 271960
rect 504600 271940 504602 271960
rect 504546 271904 504602 271940
rect 509238 269864 509294 269920
rect 509146 269456 509202 269512
rect 509882 269492 509884 269512
rect 509884 269492 509936 269512
rect 509936 269492 509938 269512
rect 509882 269456 509938 269492
rect 516506 269864 516562 269920
rect 530398 270136 530454 270192
rect 534078 270136 534134 270192
rect 536378 272856 536434 272912
rect 538126 272892 538128 272912
rect 538128 272892 538180 272912
rect 538180 272892 538182 272912
rect 538126 272856 538182 272892
rect 537942 272584 537998 272640
rect 538218 272312 538274 272368
rect 539322 273944 539378 274000
rect 538678 272620 538680 272640
rect 538680 272620 538732 272640
rect 538732 272620 538734 272640
rect 538678 272584 538734 272620
rect 537850 269900 537852 269920
rect 537852 269900 537904 269920
rect 537904 269900 537906 269920
rect 537850 269864 537906 269900
rect 538310 269864 538366 269920
rect 545946 273964 546002 274000
rect 545946 273944 545948 273964
rect 545948 273944 546000 273964
rect 546000 273944 546002 273964
rect 547694 272312 547750 272368
rect 547510 272076 547512 272096
rect 547512 272076 547564 272096
rect 547564 272076 547566 272096
rect 547510 272040 547566 272076
rect 547878 272040 547934 272096
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 554502 255604 554558 255640
rect 554502 255584 554504 255604
rect 554504 255584 554556 255604
rect 554556 255584 554558 255604
rect 554410 253408 554466 253464
rect 554134 251252 554190 251288
rect 554134 251232 554136 251252
rect 554136 251232 554188 251252
rect 554188 251232 554190 251252
rect 554042 249056 554098 249112
rect 553858 246880 553914 246936
rect 553490 244704 553546 244760
rect 553674 242528 553730 242584
rect 553766 236000 553822 236056
rect 63130 224440 63186 224496
rect 62946 223488 63002 223544
rect 118422 222264 118478 222320
rect 132498 218340 132554 218376
rect 132498 218320 132500 218340
rect 132500 218320 132552 218340
rect 132552 218320 132554 218340
rect 140042 229064 140098 229120
rect 136638 227860 136694 227896
rect 136638 227840 136640 227860
rect 136640 227840 136692 227860
rect 136692 227840 136694 227860
rect 136730 223896 136786 223952
rect 136730 218320 136786 218376
rect 141514 227860 141570 227896
rect 141514 227840 141516 227860
rect 141516 227840 141568 227860
rect 141568 227840 141570 227860
rect 143538 229064 143594 229120
rect 141606 226500 141662 226536
rect 141606 226480 141608 226500
rect 141608 226480 141660 226500
rect 141660 226480 141662 226500
rect 142250 226500 142306 226536
rect 142250 226480 142252 226500
rect 142252 226480 142304 226500
rect 142304 226480 142306 226500
rect 142618 225972 142620 225992
rect 142620 225972 142672 225992
rect 142672 225972 142674 225992
rect 142618 225936 142674 225972
rect 142250 223896 142306 223952
rect 142434 223896 142490 223952
rect 142158 223252 142166 223272
rect 142166 223252 142214 223272
rect 142158 223216 142214 223252
rect 141974 222844 141976 222864
rect 141976 222844 142028 222864
rect 142028 222844 142030 222864
rect 141974 222808 142030 222844
rect 142434 222808 142490 222864
rect 141974 222264 142030 222320
rect 142112 220924 142168 220960
rect 142112 220904 142114 220924
rect 142114 220904 142166 220924
rect 142166 220904 142168 220924
rect 142434 218476 142490 218512
rect 142434 218456 142436 218476
rect 142436 218456 142488 218476
rect 142488 218456 142490 218476
rect 144642 230424 144698 230480
rect 144458 229764 144514 229800
rect 144458 229744 144460 229764
rect 144460 229744 144512 229764
rect 144512 229744 144514 229764
rect 145838 229356 145894 229392
rect 145838 229336 145840 229356
rect 145840 229336 145892 229356
rect 145892 229336 145894 229356
rect 146114 227976 146170 228032
rect 145930 222944 145986 223000
rect 147126 227976 147182 228032
rect 148138 229744 148194 229800
rect 147954 229336 148010 229392
rect 148138 229220 148194 229256
rect 148138 229200 148140 229220
rect 148140 229200 148192 229220
rect 148192 229200 148194 229220
rect 147126 222980 147128 223000
rect 147128 222980 147180 223000
rect 147180 222980 147182 223000
rect 147126 222944 147182 222980
rect 148874 225392 148930 225448
rect 148506 220924 148562 220960
rect 148506 220904 148508 220924
rect 148508 220904 148560 220924
rect 148560 220904 148562 220924
rect 146574 218456 146630 218512
rect 151082 230424 151138 230480
rect 150346 229472 150402 229528
rect 149794 225936 149850 225992
rect 149518 223216 149574 223272
rect 150990 229200 151046 229256
rect 151450 226208 151506 226264
rect 150714 220516 150770 220552
rect 150714 220496 150716 220516
rect 150716 220496 150768 220516
rect 150768 220496 150770 220516
rect 151634 224440 151690 224496
rect 151634 223896 151690 223952
rect 152370 224440 152426 224496
rect 151910 220516 151966 220552
rect 151910 220496 151912 220516
rect 151912 220496 151964 220516
rect 151964 220496 151966 220516
rect 152186 220108 152242 220144
rect 152186 220088 152188 220108
rect 152188 220088 152240 220108
rect 152240 220088 152242 220108
rect 151818 219816 151874 219872
rect 155590 227024 155646 227080
rect 154394 220124 154396 220144
rect 154396 220124 154448 220144
rect 154448 220124 154450 220144
rect 154394 220088 154450 220124
rect 156786 230036 156842 230072
rect 156786 230016 156788 230036
rect 156788 230016 156840 230036
rect 156840 230016 156842 230036
rect 157614 230172 157670 230208
rect 157614 230152 157616 230172
rect 157616 230152 157668 230172
rect 157668 230152 157670 230172
rect 157430 230036 157486 230072
rect 157430 230016 157432 230036
rect 157432 230016 157484 230036
rect 157484 230016 157486 230036
rect 156786 229764 156842 229800
rect 156786 229744 156788 229764
rect 156788 229744 156840 229764
rect 156840 229744 156842 229764
rect 157982 229628 158038 229664
rect 157982 229608 157984 229628
rect 157984 229608 158036 229628
rect 158036 229608 158038 229628
rect 157338 227432 157394 227488
rect 157522 227024 157578 227080
rect 157154 226208 157210 226264
rect 156602 225800 156658 225856
rect 157154 225392 157210 225448
rect 156326 219816 156382 219872
rect 157614 222012 157670 222048
rect 157614 221992 157616 222012
rect 157616 221992 157668 222012
rect 157668 221992 157670 222012
rect 157430 221584 157486 221640
rect 158166 225800 158222 225856
rect 158350 222012 158406 222048
rect 158350 221992 158352 222012
rect 158352 221992 158404 222012
rect 158404 221992 158406 222012
rect 158166 221584 158222 221640
rect 159362 228812 159418 228848
rect 159362 228792 159364 228812
rect 159364 228792 159416 228812
rect 159416 228792 159418 228812
rect 160006 228384 160062 228440
rect 160650 220924 160706 220960
rect 161018 221176 161074 221232
rect 160650 220904 160652 220924
rect 160652 220904 160704 220924
rect 160704 220904 160706 220924
rect 162306 230152 162362 230208
rect 162490 229336 162546 229392
rect 162490 228792 162546 228848
rect 162306 221196 162362 221232
rect 162306 221176 162308 221196
rect 162308 221176 162360 221196
rect 162360 221176 162362 221196
rect 166814 228384 166870 228440
rect 166538 227432 166594 227488
rect 164514 220924 164570 220960
rect 164514 220904 164516 220924
rect 164516 220904 164568 220924
rect 164568 220904 164570 220924
rect 166814 222012 166870 222048
rect 166814 221992 166816 222012
rect 166816 221992 166868 222012
rect 166868 221992 166870 222012
rect 166998 222012 167054 222048
rect 166998 221992 167000 222012
rect 167000 221992 167052 222012
rect 167052 221992 167054 222012
rect 169574 227160 169630 227216
rect 170770 227452 170826 227488
rect 170770 227432 170772 227452
rect 170772 227432 170824 227452
rect 170824 227432 170826 227452
rect 171690 227432 171746 227488
rect 171092 227160 171148 227216
rect 172242 222400 172298 222456
rect 171414 221312 171470 221368
rect 171966 221332 172022 221368
rect 171966 221312 171968 221332
rect 171968 221312 172020 221332
rect 172020 221312 172022 221332
rect 173162 228792 173218 228848
rect 175186 227588 175242 227624
rect 175186 227568 175188 227588
rect 175188 227568 175240 227588
rect 175240 227568 175242 227588
rect 176106 228812 176162 228848
rect 176106 228792 176108 228812
rect 176108 228792 176160 228812
rect 176160 228792 176162 228812
rect 175922 227296 175978 227352
rect 175830 222420 175886 222456
rect 175830 222400 175832 222420
rect 175832 222400 175884 222420
rect 175884 222400 175886 222420
rect 177210 227568 177266 227624
rect 176750 227316 176806 227352
rect 176750 227296 176752 227316
rect 176752 227296 176804 227316
rect 176804 227296 176806 227316
rect 176566 221876 176622 221912
rect 176566 221856 176568 221876
rect 176568 221856 176620 221876
rect 176620 221856 176622 221876
rect 177394 221856 177450 221912
rect 176566 220632 176622 220688
rect 180798 220904 180854 220960
rect 181074 220652 181130 220688
rect 181074 220632 181076 220652
rect 181076 220632 181128 220652
rect 181128 220632 181130 220652
rect 185398 229880 185454 229936
rect 186042 229880 186098 229936
rect 185030 220904 185086 220960
rect 185858 220768 185914 220824
rect 190412 220788 190468 220824
rect 190412 220768 190414 220788
rect 190414 220768 190466 220788
rect 190466 220768 190468 220788
rect 190274 219972 190330 220008
rect 193034 228928 193090 228984
rect 190274 219952 190276 219972
rect 190276 219952 190328 219972
rect 190328 219952 190330 219972
rect 190642 219952 190698 220008
rect 195426 228948 195482 228984
rect 195426 228928 195428 228948
rect 195428 228928 195480 228948
rect 195480 228928 195482 228948
rect 221830 226752 221886 226808
rect 223118 226772 223174 226808
rect 223118 226752 223120 226772
rect 223120 226752 223172 226772
rect 223172 226752 223174 226772
rect 486974 220224 487030 220280
rect 487802 218048 487858 218104
rect 488814 217096 488870 217152
rect 492954 219680 493010 219736
rect 493690 219680 493746 219736
rect 494702 218320 494758 218376
rect 495162 217096 495218 217152
rect 500958 217232 501014 217288
rect 510986 217504 511042 217560
rect 513562 220904 513618 220960
rect 515770 221176 515826 221232
rect 515126 219952 515182 220008
rect 520186 219408 520242 219464
rect 520002 217504 520058 217560
rect 522578 221448 522634 221504
rect 531502 217504 531558 217560
rect 532514 217504 532570 217560
rect 542450 224476 542452 224496
rect 542452 224476 542504 224496
rect 542504 224476 542506 224496
rect 542450 224440 542506 224476
rect 543186 224440 543242 224496
rect 548062 224748 548064 224768
rect 548064 224748 548116 224768
rect 548116 224748 548118 224768
rect 548062 224712 548118 224748
rect 545762 221720 545818 221776
rect 549994 224712 550050 224768
rect 550454 224712 550510 224768
rect 549258 221720 549314 221776
rect 547418 218728 547474 218784
rect 548614 218748 548670 218784
rect 548614 218728 548616 218748
rect 548616 218728 548668 218748
rect 548668 218728 548670 218748
rect 554502 240352 554558 240408
rect 554318 238176 554374 238232
rect 554410 233824 554466 233880
rect 554870 224440 554926 224496
rect 556066 224440 556122 224496
rect 553306 222264 553362 222320
rect 556986 221892 556988 221912
rect 556988 221892 557040 221912
rect 557040 221892 557042 221912
rect 556986 221856 557042 221892
rect 557998 224576 558054 224632
rect 557354 222264 557410 222320
rect 557538 221856 557594 221912
rect 559378 222028 559380 222048
rect 559380 222028 559432 222048
rect 559432 222028 559434 222048
rect 559378 221992 559434 222028
rect 560298 218592 560354 218648
rect 562138 224748 562140 224768
rect 562140 224748 562192 224768
rect 562192 224748 562194 224768
rect 562138 224712 562194 224748
rect 563702 224712 563758 224768
rect 561494 221992 561550 222048
rect 560758 217504 560814 217560
rect 560942 217504 560998 217560
rect 563702 221720 563758 221776
rect 561770 220516 561826 220552
rect 561770 220496 561772 220516
rect 561772 220496 561824 220516
rect 561824 220496 561826 220516
rect 563150 220516 563206 220552
rect 563150 220496 563152 220516
rect 563152 220496 563204 220516
rect 563204 220496 563206 220516
rect 561678 218592 561734 218648
rect 563012 219020 563068 219056
rect 563012 219000 563014 219020
rect 563014 219000 563066 219020
rect 563066 219000 563068 219020
rect 563150 217504 563206 217560
rect 565634 220496 565690 220552
rect 564806 217776 564862 217832
rect 567658 218728 567714 218784
rect 568302 218748 568358 218784
rect 568302 218728 568304 218748
rect 568304 218728 568356 218748
rect 568356 218728 568358 218748
rect 569958 220496 570014 220552
rect 572626 221720 572682 221776
rect 572534 219136 572590 219192
rect 574742 219136 574798 219192
rect 572534 218864 572590 218920
rect 571890 217776 571946 217832
rect 572074 217776 572130 217832
rect 574374 217776 574430 217832
rect 572534 217504 572590 217560
rect 574190 217504 574246 217560
rect 53286 215056 53342 215112
rect 575478 216688 575534 216744
rect 51722 180784 51778 180840
rect 591486 224168 591542 224224
rect 578882 213968 578938 214024
rect 578514 211656 578570 211712
rect 579526 209788 579528 209808
rect 579528 209788 579580 209808
rect 579580 209788 579582 209808
rect 579526 209752 579582 209788
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 578238 166912 578294 166968
rect 579526 164464 579582 164520
rect 579342 162696 579398 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153992 578386 154048
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147464 579582 147520
rect 578606 140528 578662 140584
rect 578606 138760 578662 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 579526 142976 579582 143032
rect 578882 136584 578938 136640
rect 579526 134408 579582 134464
rect 579066 132232 579122 132288
rect 578882 129648 578938 129704
rect 579526 127880 579582 127936
rect 578330 125296 578386 125352
rect 578422 123564 578424 123584
rect 578424 123564 578476 123584
rect 578476 123564 578478 123584
rect 578422 123528 578478 123564
rect 578882 121352 578938 121408
rect 578514 118396 578516 118416
rect 578516 118396 578568 118416
rect 578568 118396 578570 118416
rect 578514 118360 578570 118396
rect 578330 108296 578386 108352
rect 578606 99220 578608 99240
rect 578608 99220 578660 99240
rect 578660 99220 578662 99240
rect 578606 99184 578662 99220
rect 578330 97416 578386 97472
rect 578514 93064 578570 93120
rect 579526 116900 579528 116920
rect 579528 116900 579580 116920
rect 579580 116900 579582 116920
rect 579526 116864 579582 116900
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579526 112512 579582 112568
rect 579342 110100 579344 110120
rect 579344 110100 579396 110120
rect 579396 110100 579398 110120
rect 579342 110064 579398 110100
rect 579066 105848 579122 105904
rect 579526 103264 579582 103320
rect 579526 101632 579582 101688
rect 579526 95004 579528 95024
rect 579528 95004 579580 95024
rect 579580 95004 579582 95024
rect 579526 94968 579582 95004
rect 579066 90888 579122 90944
rect 579526 88068 579528 88088
rect 579528 88068 579580 88088
rect 579580 88068 579582 88088
rect 579526 88032 579582 88068
rect 579342 86400 579398 86456
rect 579158 83952 579214 84008
rect 579066 82184 579122 82240
rect 578882 80008 578938 80064
rect 578238 75520 578294 75576
rect 579526 77832 579582 77888
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589462 204720 589518 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589646 170448 589702 170504
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589278 157412 589334 157448
rect 589278 157392 589280 157412
rect 589280 157392 589332 157412
rect 589332 157392 589334 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 590014 150864 590070 150920
rect 589462 149232 589518 149288
rect 588542 147600 588598 147656
rect 589462 145968 589518 146024
rect 589462 144336 589518 144392
rect 589830 142704 589886 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590382 134544 590438 134600
rect 589462 132912 589518 132968
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 588542 129648 588598 129704
rect 581642 77832 581698 77888
rect 579066 73072 579122 73128
rect 576122 54984 576178 55040
rect 579066 71168 579122 71224
rect 580262 54712 580318 54768
rect 578882 54440 578938 54496
rect 589462 128016 589518 128072
rect 589922 126384 589978 126440
rect 589462 124752 589518 124808
rect 589462 123120 589518 123176
rect 590014 121488 590070 121544
rect 589646 119856 589702 119912
rect 589462 116592 589518 116648
rect 590106 118224 590162 118280
rect 589462 113328 589518 113384
rect 590290 114960 590346 115016
rect 589462 111696 589518 111752
rect 589278 110064 589334 110120
rect 589462 108432 589518 108488
rect 589830 106800 589886 106856
rect 589462 105168 589518 105224
rect 588726 103536 588782 103592
rect 589462 101904 589518 101960
rect 577502 54168 577558 54224
rect 459834 53624 459890 53680
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 464158 53352 464214 53408
rect 464710 53352 464766 53408
rect 471794 53508 471850 53544
rect 471794 53488 471796 53508
rect 471796 53488 471848 53508
rect 471848 53488 471850 53508
rect 473542 53508 473598 53544
rect 473542 53488 473544 53508
rect 473544 53488 473596 53508
rect 473596 53488 473598 53508
rect 130382 44240 130438 44296
rect 458178 46960 458234 47016
rect 522946 47776 523002 47832
rect 132406 44276 132408 44296
rect 132408 44276 132460 44296
rect 132460 44276 132462 44296
rect 132406 44240 132462 44276
rect 458362 46688 458418 46744
rect 142618 44240 142674 44296
rect 255870 44104 255926 44160
rect 361762 43832 361818 43888
rect 440238 43852 440294 43888
rect 440238 43832 440240 43852
rect 440240 43832 440292 43852
rect 440292 43832 440294 43852
rect 441066 43852 441122 43888
rect 441066 43832 441068 43852
rect 441068 43832 441120 43852
rect 441120 43832 441122 43852
rect 415582 42336 415638 42392
rect 365074 41792 365130 41848
rect 416686 41792 416742 41848
rect 419906 41792 419962 41848
rect 446218 42200 446274 42256
rect 446218 41520 446274 41576
rect 460110 44104 460166 44160
rect 461030 44376 461086 44432
rect 460846 43424 460902 43480
rect 461766 42880 461822 42936
rect 462870 44376 462926 44432
rect 462686 43152 462742 43208
rect 463790 44376 463846 44432
rect 463974 42880 464030 42936
rect 465078 46960 465134 47016
rect 549994 48864 550050 48920
rect 591486 101632 591542 101688
rect 600870 221176 600926 221232
rect 599490 220904 599546 220960
rect 595166 217232 595222 217288
rect 595718 216960 595774 217016
rect 599030 215600 599086 215656
rect 611634 220224 611690 220280
rect 612738 219680 612794 219736
rect 618258 221448 618314 221504
rect 617154 219952 617210 220008
rect 617798 215872 617854 215928
rect 618442 219408 618498 219464
rect 621110 215328 621166 215384
rect 623962 218048 624018 218104
rect 630678 218320 630734 218376
rect 650642 224984 650698 225040
rect 645858 219816 645914 219872
rect 648434 218592 648490 218648
rect 651102 217232 651158 217288
rect 651470 221448 651526 221504
rect 652390 280336 652446 280392
rect 652574 279384 652630 279440
rect 660578 293800 660634 293856
rect 658922 268096 658978 268152
rect 664442 247696 664498 247752
rect 666558 245656 666614 245712
rect 652390 226888 652446 226944
rect 658922 226344 658978 226400
rect 656162 225528 656218 225584
rect 652758 225256 652814 225312
rect 654782 223896 654838 223952
rect 653402 222808 653458 222864
rect 654138 220360 654194 220416
rect 653770 217504 653826 217560
rect 657542 223624 657598 223680
rect 656806 218864 656862 218920
rect 660762 221720 660818 221776
rect 659566 215328 659622 215384
rect 658738 213152 658794 213208
rect 660394 214512 660450 214568
rect 662142 228520 662198 228576
rect 661498 213424 661554 213480
rect 664902 230288 664958 230344
rect 663706 229064 663762 229120
rect 664626 215600 664682 215656
rect 665822 223080 665878 223136
rect 666834 221448 666890 221504
rect 667018 220360 667074 220416
rect 666834 219408 666890 219464
rect 666650 215872 666706 215928
rect 666650 198464 666706 198520
rect 667018 217912 667074 217968
rect 667018 188808 667074 188864
rect 666834 174936 666890 174992
rect 667754 224168 667810 224224
rect 667754 223624 667810 223680
rect 667754 223116 667756 223136
rect 667756 223116 667808 223136
rect 667808 223116 667810 223136
rect 667754 223080 667810 223116
rect 667570 181328 667626 181384
rect 667386 180240 667442 180296
rect 668766 232464 668822 232520
rect 668398 199144 668454 199200
rect 668122 194248 668178 194304
rect 668398 191664 668454 191720
rect 667938 184456 667994 184512
rect 668214 177964 668216 177984
rect 668216 177964 668268 177984
rect 668268 177964 668270 177984
rect 668214 177928 668270 177964
rect 668030 174664 668086 174720
rect 667938 169668 667940 169688
rect 667940 169668 667992 169688
rect 667992 169668 667994 169688
rect 667938 169632 667994 169668
rect 667938 164872 667994 164928
rect 668214 160012 668216 160032
rect 668216 160012 668268 160032
rect 668268 160012 668270 160032
rect 668214 159976 668270 160012
rect 668214 155080 668270 155136
rect 669226 250144 669282 250200
rect 669226 247696 669282 247752
rect 669134 231104 669190 231160
rect 669272 223388 669274 223408
rect 669274 223388 669326 223408
rect 669326 223388 669328 223408
rect 669272 223352 669328 223388
rect 669870 301960 669926 302016
rect 669410 216552 669466 216608
rect 669594 215600 669650 215656
rect 669410 215056 669466 215112
rect 669134 204040 669190 204096
rect 669410 202816 669466 202872
rect 669134 198736 669190 198792
rect 668950 189352 669006 189408
rect 668766 163240 668822 163296
rect 668766 162424 668822 162480
rect 668766 148552 668822 148608
rect 668766 145288 668822 145344
rect 668582 138760 668638 138816
rect 668398 135496 668454 135552
rect 668766 135088 668822 135144
rect 667938 133764 667940 133784
rect 667940 133764 667992 133784
rect 667992 133764 667994 133784
rect 667938 133728 667994 133764
rect 667754 133048 667810 133104
rect 667202 132504 667258 132560
rect 668490 130600 668546 130656
rect 668030 128968 668086 129024
rect 668582 127744 668638 127800
rect 667938 107752 667994 107808
rect 668398 106156 668400 106176
rect 668400 106156 668452 106176
rect 668452 106156 668454 106176
rect 668398 106120 668454 106156
rect 669502 172352 669558 172408
rect 669594 150320 669650 150376
rect 669134 143656 669190 143712
rect 670330 262112 670386 262168
rect 670146 258440 670202 258496
rect 670330 236136 670386 236192
rect 670974 295704 671030 295760
rect 670974 293800 671030 293856
rect 671802 559680 671858 559736
rect 672630 624452 672632 624472
rect 672632 624452 672684 624472
rect 672684 624452 672686 624472
rect 672630 624416 672686 624452
rect 672630 623772 672632 623792
rect 672632 623772 672684 623792
rect 672684 623772 672686 623792
rect 672630 623736 672686 623772
rect 672630 623228 672632 623248
rect 672632 623228 672684 623248
rect 672684 623228 672686 623248
rect 672630 623192 672686 623228
rect 672630 622412 672632 622432
rect 672632 622412 672684 622432
rect 672684 622412 672686 622432
rect 672630 622376 672686 622412
rect 672354 604424 672410 604480
rect 672538 597352 672594 597408
rect 672998 648760 673054 648816
rect 672814 573688 672870 573744
rect 674378 779320 674434 779376
rect 674562 778776 674618 778832
rect 674930 777008 674986 777064
rect 674930 775668 674986 775704
rect 674930 775648 674932 775668
rect 674932 775648 674984 775668
rect 674984 775648 674986 775668
rect 675482 779320 675538 779376
rect 675482 778776 675538 778832
rect 675390 777416 675446 777472
rect 675482 777008 675538 777064
rect 675390 775648 675446 775704
rect 675206 743280 675262 743336
rect 675206 738112 675262 738168
rect 674746 729816 674802 729872
rect 675482 735664 675538 735720
rect 675482 734304 675538 734360
rect 675482 733760 675538 733816
rect 675298 730768 675354 730824
rect 675482 730088 675538 730144
rect 674010 721792 674066 721848
rect 675482 728728 675538 728784
rect 675114 721656 675170 721712
rect 674010 719616 674066 719672
rect 673734 707512 673790 707568
rect 673734 706288 673790 706344
rect 673734 705064 673790 705120
rect 673734 701156 673736 701176
rect 673736 701156 673788 701176
rect 673788 701156 673790 701176
rect 673734 701120 673790 701156
rect 673734 692844 673790 692880
rect 673734 692824 673736 692844
rect 673736 692824 673788 692844
rect 673788 692824 673790 692844
rect 673734 690124 673790 690160
rect 673734 690104 673736 690124
rect 673736 690104 673788 690124
rect 673788 690104 673790 690124
rect 673734 688780 673736 688800
rect 673736 688780 673788 688800
rect 673788 688780 673790 688800
rect 673734 688744 673790 688780
rect 673734 688064 673790 688120
rect 673458 682352 673514 682408
rect 673550 681944 673606 682000
rect 673550 671356 673606 671392
rect 673550 671336 673552 671356
rect 673552 671336 673604 671356
rect 673604 671336 673606 671356
rect 673550 670928 673606 670984
rect 673550 670520 673606 670576
rect 673550 669704 673606 669760
rect 673550 668888 673606 668944
rect 673550 668516 673552 668536
rect 673552 668516 673604 668536
rect 673604 668516 673606 668536
rect 673550 668480 673606 668516
rect 673550 668072 673606 668128
rect 673550 667664 673606 667720
rect 673550 666848 673606 666904
rect 673550 666596 673606 666632
rect 673550 666576 673552 666596
rect 673552 666576 673604 666596
rect 673604 666576 673606 666596
rect 673550 665252 673552 665272
rect 673552 665252 673604 665272
rect 673604 665252 673606 665272
rect 673550 665216 673606 665252
rect 673550 664420 673606 664456
rect 673550 664400 673552 664420
rect 673552 664400 673604 664420
rect 673604 664400 673606 664420
rect 673550 663720 673606 663776
rect 673550 643456 673606 643512
rect 673458 641688 673514 641744
rect 673274 626084 673276 626104
rect 673276 626084 673328 626104
rect 673328 626084 673330 626104
rect 673274 626048 673330 626084
rect 673274 625404 673276 625424
rect 673276 625404 673328 625424
rect 673328 625404 673330 625424
rect 673274 625368 673330 625404
rect 673274 625132 673276 625152
rect 673276 625132 673328 625152
rect 673328 625132 673330 625152
rect 673274 625096 673330 625132
rect 673274 621172 673330 621208
rect 673274 621152 673276 621172
rect 673276 621152 673328 621172
rect 673328 621152 673330 621172
rect 673274 618160 673330 618216
rect 673274 607280 673330 607336
rect 672998 573280 673054 573336
rect 673090 560088 673146 560144
rect 672906 555192 672962 555248
rect 672722 490048 672778 490104
rect 672262 453908 672264 453928
rect 672264 453908 672316 453928
rect 672316 453908 672318 453928
rect 672262 453872 672318 453908
rect 672906 485968 672962 486024
rect 675298 712000 675354 712056
rect 682382 726552 682438 726608
rect 682382 711184 682438 711240
rect 681002 710776 681058 710832
rect 676034 707140 676036 707160
rect 676036 707140 676088 707160
rect 676088 707140 676090 707160
rect 676034 707104 676090 707140
rect 684222 726280 684278 726336
rect 684222 709552 684278 709608
rect 684038 707920 684094 707976
rect 683394 706696 683450 706752
rect 683118 705472 683174 705528
rect 674286 705356 674342 705392
rect 674286 705336 674288 705356
rect 674288 705336 674340 705356
rect 674340 705336 674342 705356
rect 675114 701120 675170 701176
rect 675114 698264 675170 698320
rect 675114 696904 675170 696960
rect 675482 696768 675538 696824
rect 675114 695816 675170 695872
rect 675114 694592 675170 694648
rect 674102 689832 674158 689888
rect 675114 692824 675170 692880
rect 674930 690104 674986 690160
rect 675114 689832 675170 689888
rect 675114 689424 675170 689480
rect 674286 688064 674342 688120
rect 673918 661952 673974 662008
rect 674010 661580 674012 661600
rect 674012 661580 674064 661600
rect 674064 661580 674066 661600
rect 674010 661544 674066 661580
rect 674010 661156 674066 661192
rect 674010 661136 674012 661156
rect 674012 661136 674064 661156
rect 674064 661136 674066 661156
rect 674010 660204 674066 660240
rect 674010 660184 674012 660204
rect 674012 660184 674064 660204
rect 674064 660184 674066 660204
rect 674010 659912 674066 659968
rect 674010 655580 674066 655616
rect 674010 655560 674012 655580
rect 674012 655560 674064 655580
rect 674064 655560 674066 655580
rect 674194 644544 674250 644600
rect 674930 688744 674986 688800
rect 675114 687792 675170 687848
rect 675114 686160 675170 686216
rect 674930 685752 674986 685808
rect 675114 685480 675170 685536
rect 675114 683984 675170 684040
rect 674286 625132 674288 625152
rect 674288 625132 674340 625152
rect 674340 625132 674342 625152
rect 674286 625096 674342 625132
rect 674010 623908 674012 623928
rect 674012 623908 674064 623928
rect 674064 623908 674066 623928
rect 674010 623872 674066 623908
rect 674286 623600 674342 623656
rect 674838 682388 674840 682408
rect 674840 682388 674892 682408
rect 674892 682388 674894 682408
rect 674838 682352 674894 682388
rect 675298 683712 675354 683768
rect 675114 676368 675170 676424
rect 674838 666612 674840 666632
rect 674840 666612 674892 666632
rect 674892 666612 674894 666632
rect 674838 666576 674894 666612
rect 684130 682624 684186 682680
rect 675482 681944 675538 682000
rect 676034 667256 676090 667312
rect 675298 666440 675354 666496
rect 676034 664808 676090 664864
rect 674838 663756 674840 663776
rect 674840 663756 674892 663776
rect 674892 663756 674894 663776
rect 674838 663720 674894 663756
rect 683210 663720 683266 663776
rect 684130 666168 684186 666224
rect 683486 662904 683542 662960
rect 674838 660184 674894 660240
rect 683118 660048 683174 660104
rect 675114 655560 675170 655616
rect 675390 652840 675446 652896
rect 675114 652432 675170 652488
rect 675390 649168 675446 649224
rect 675114 648760 675170 648816
rect 675390 647808 675446 647864
rect 675114 645768 675170 645824
rect 675298 644544 675354 644600
rect 675390 644272 675446 644328
rect 675574 643592 675630 643648
rect 675298 643456 675354 643512
rect 675298 641688 675354 641744
rect 675206 641416 675262 641472
rect 674286 622412 674288 622432
rect 674288 622412 674340 622432
rect 674340 622412 674342 622432
rect 674286 622376 674342 622412
rect 674010 621036 674066 621072
rect 674010 621016 674012 621036
rect 674012 621016 674064 621036
rect 674064 621016 674066 621036
rect 673734 617344 673790 617400
rect 674010 614916 674066 614952
rect 674010 614896 674012 614916
rect 674012 614896 674064 614916
rect 674064 614896 674066 614916
rect 675482 638560 675538 638616
rect 681002 637472 681058 637528
rect 675482 631352 675538 631408
rect 675666 631352 675722 631408
rect 676218 625640 676274 625696
rect 676218 624416 676274 624472
rect 676402 622784 676458 622840
rect 676034 622668 676090 622704
rect 676034 622648 676036 622668
rect 676036 622648 676088 622668
rect 676088 622648 676090 622668
rect 681002 621968 681058 622024
rect 676034 621444 676090 621480
rect 676034 621424 676036 621444
rect 676036 621424 676088 621444
rect 676088 621424 676090 621444
rect 676218 620780 676220 620800
rect 676220 620780 676272 620800
rect 676272 620780 676274 620800
rect 676218 620744 676274 620780
rect 676218 619948 676274 619984
rect 676218 619928 676220 619948
rect 676220 619928 676272 619948
rect 676272 619928 676274 619948
rect 676494 619928 676550 619984
rect 676218 619540 676274 619576
rect 676218 619520 676220 619540
rect 676220 619520 676272 619540
rect 676272 619520 676274 619540
rect 683210 618704 683266 618760
rect 676034 617752 676090 617808
rect 675298 617072 675354 617128
rect 683578 617072 683634 617128
rect 683394 616664 683450 616720
rect 683118 615476 683120 615496
rect 683120 615476 683172 615496
rect 683172 615476 683174 615496
rect 683118 615440 683174 615476
rect 674194 598984 674250 599040
rect 673458 594496 673514 594552
rect 673918 598576 673974 598632
rect 673550 581304 673606 581360
rect 673550 580624 673606 580680
rect 673550 574540 673552 574560
rect 673552 574540 673604 574560
rect 673604 574540 673606 574560
rect 673550 574504 673606 574540
rect 673550 574096 673606 574152
rect 673550 570444 673606 570480
rect 673550 570424 673552 570444
rect 673552 570424 673604 570444
rect 673604 570424 673606 570444
rect 673550 565836 673552 565856
rect 673552 565836 673604 565856
rect 673604 565836 673606 565856
rect 673550 565800 673606 565836
rect 673550 564460 673606 564496
rect 673550 564440 673552 564460
rect 673552 564440 673604 564460
rect 673604 564440 673606 564460
rect 673550 554804 673606 554840
rect 673550 554784 673552 554804
rect 673552 554784 673604 554804
rect 673604 554784 673606 554804
rect 673550 553152 673606 553208
rect 673274 530032 673330 530088
rect 673366 527720 673422 527776
rect 673366 490456 673422 490512
rect 673090 484744 673146 484800
rect 674010 581052 674066 581088
rect 674010 581032 674012 581052
rect 674012 581032 674064 581052
rect 674064 581032 674066 581052
rect 674010 580216 674066 580272
rect 674010 579844 674012 579864
rect 674012 579844 674064 579864
rect 674064 579844 674066 579864
rect 674010 579808 674066 579844
rect 674010 579420 674066 579456
rect 674010 579400 674012 579420
rect 674012 579400 674064 579420
rect 674064 579400 674066 579420
rect 674010 579028 674012 579048
rect 674012 579028 674064 579048
rect 674064 579028 674066 579048
rect 674010 578992 674066 579028
rect 674010 578604 674066 578640
rect 674010 578584 674012 578604
rect 674012 578584 674064 578604
rect 674064 578584 674066 578604
rect 674010 578196 674066 578232
rect 674010 578176 674012 578196
rect 674012 578176 674064 578196
rect 674064 578176 674066 578196
rect 674010 577788 674066 577824
rect 674010 577768 674012 577788
rect 674012 577768 674064 577788
rect 674064 577768 674066 577788
rect 674010 577396 674012 577416
rect 674012 577396 674064 577416
rect 674064 577396 674066 577416
rect 674010 577360 674066 577396
rect 674010 576972 674066 577008
rect 674010 576952 674012 576972
rect 674012 576952 674064 576972
rect 674064 576952 674066 576972
rect 674010 574912 674066 574968
rect 674010 572464 674066 572520
rect 674010 572056 674066 572112
rect 674010 570832 674066 570888
rect 674010 569608 674066 569664
rect 674102 558320 674158 558376
rect 673918 547304 673974 547360
rect 674470 581304 674526 581360
rect 674470 552064 674526 552120
rect 673826 492088 673882 492144
rect 674010 491308 674012 491328
rect 674012 491308 674064 491328
rect 674064 491308 674066 491328
rect 674010 491272 674066 491308
rect 674010 490900 674012 490920
rect 674012 490900 674064 490920
rect 674064 490900 674066 490920
rect 674010 490864 674066 490900
rect 674010 489660 674066 489696
rect 674010 489640 674012 489660
rect 674012 489640 674064 489660
rect 674064 489640 674066 489660
rect 674010 489268 674012 489288
rect 674012 489268 674064 489288
rect 674064 489268 674066 489288
rect 674010 489232 674066 489268
rect 674010 488452 674012 488472
rect 674012 488452 674064 488472
rect 674064 488452 674066 488472
rect 674010 488416 674066 488452
rect 675482 607688 675538 607744
rect 675298 607280 675354 607336
rect 675114 604424 675170 604480
rect 675114 602928 675170 602984
rect 675390 600888 675446 600944
rect 675482 598984 675538 599040
rect 675482 598576 675538 598632
rect 675482 597352 675538 597408
rect 675390 595312 675446 595368
rect 675206 594768 675262 594824
rect 675206 594496 675262 594552
rect 675390 593408 675446 593464
rect 674930 590416 674986 590472
rect 674838 570460 674840 570480
rect 674840 570460 674892 570480
rect 674892 570460 674894 570480
rect 674838 570424 674894 570460
rect 675482 593136 675538 593192
rect 675206 586200 675262 586256
rect 681002 591640 681058 591696
rect 682382 576408 682438 576464
rect 681002 575592 681058 575648
rect 684222 591232 684278 591288
rect 683394 573144 683450 573200
rect 684222 576000 684278 576056
rect 684038 571920 684094 571976
rect 676218 571548 676220 571568
rect 676220 571548 676272 571568
rect 676272 571548 676274 571568
rect 676218 571512 676274 571548
rect 683118 570288 683174 570344
rect 675390 565800 675446 565856
rect 675114 564440 675170 564496
rect 675114 562264 675170 562320
rect 675390 561856 675446 561912
rect 675298 559680 675354 559736
rect 675482 559408 675538 559464
rect 675482 558320 675538 558376
rect 675298 557504 675354 557560
rect 675390 555192 675446 555248
rect 675298 554784 675354 554840
rect 675758 553832 675814 553888
rect 675574 553424 675630 553480
rect 675390 552064 675446 552120
rect 675390 551520 675446 551576
rect 675482 549616 675538 549672
rect 674930 545672 674986 545728
rect 675758 548256 675814 548312
rect 677414 547576 677470 547632
rect 675574 547304 675630 547360
rect 676218 535880 676274 535936
rect 676034 535712 676036 535732
rect 676036 535712 676088 535732
rect 676088 535712 676090 535732
rect 676034 535676 676090 535712
rect 676218 535064 676274 535120
rect 676034 534896 676036 534916
rect 676036 534896 676088 534916
rect 676088 534896 676090 534916
rect 676034 534860 676090 534896
rect 676034 534472 676090 534508
rect 676034 534452 676036 534472
rect 676036 534452 676088 534472
rect 676088 534452 676090 534472
rect 676034 534080 676036 534100
rect 676036 534080 676088 534100
rect 676088 534080 676090 534100
rect 676034 534044 676090 534080
rect 676402 533432 676458 533488
rect 676034 533228 676090 533284
rect 676218 533060 676220 533080
rect 676220 533060 676272 533080
rect 676272 533060 676274 533080
rect 676218 533024 676274 533060
rect 676218 532208 676274 532264
rect 676034 532004 676090 532060
rect 676402 531800 676458 531856
rect 676034 529984 676090 530020
rect 676034 529964 676036 529984
rect 676036 529964 676088 529984
rect 676088 529964 676090 529984
rect 676218 529372 676274 529408
rect 676218 529352 676220 529372
rect 676220 529352 676272 529372
rect 676272 529352 676274 529372
rect 676218 528980 676220 529000
rect 676220 528980 676272 529000
rect 676272 528980 676274 529000
rect 676218 528944 676274 528980
rect 676034 528760 676090 528796
rect 676034 528740 676036 528760
rect 676036 528740 676088 528760
rect 676088 528740 676090 528760
rect 676034 526736 676036 526756
rect 676036 526736 676088 526756
rect 676088 526736 676090 526756
rect 676034 526700 676090 526736
rect 676034 526328 676036 526348
rect 676036 526328 676088 526348
rect 676088 526328 676090 526348
rect 676034 526292 676090 526328
rect 674654 484336 674710 484392
rect 674010 483148 674012 483168
rect 674012 483148 674064 483168
rect 674064 483148 674066 483168
rect 674010 483112 674066 483148
rect 673550 482296 673606 482352
rect 673274 455388 673330 455424
rect 673274 455368 673276 455388
rect 673276 455368 673328 455388
rect 673328 455368 673330 455388
rect 673386 455252 673442 455288
rect 673386 455232 673388 455252
rect 673388 455232 673440 455252
rect 673440 455232 673442 455252
rect 673274 455096 673330 455152
rect 672814 454824 672870 454880
rect 674286 454860 674288 454880
rect 674288 454860 674340 454880
rect 674340 454860 674342 454880
rect 674286 454824 674342 454860
rect 673044 454588 673046 454608
rect 673046 454588 673098 454608
rect 673098 454588 673100 454608
rect 673044 454552 673100 454588
rect 674286 454588 674288 454608
rect 674288 454588 674340 454608
rect 674340 454588 674342 454608
rect 674286 454552 674342 454588
rect 676034 491700 676090 491736
rect 676034 491680 676036 491700
rect 676036 491680 676088 491700
rect 676088 491680 676090 491700
rect 676034 486804 676090 486840
rect 676034 486784 676036 486804
rect 676036 486784 676088 486804
rect 676088 486784 676090 486804
rect 676034 485172 676090 485208
rect 676034 485152 676036 485172
rect 676036 485152 676088 485172
rect 676088 485152 676090 485172
rect 676034 483964 676036 483984
rect 676036 483964 676088 483984
rect 676088 483964 676090 483984
rect 676034 483928 676090 483964
rect 681002 546760 681058 546816
rect 682382 531392 682438 531448
rect 681002 530576 681058 530632
rect 683394 547032 683450 547088
rect 683210 527720 683266 527776
rect 683578 528536 683634 528592
rect 683394 527312 683450 527368
rect 677874 525680 677930 525736
rect 683118 524864 683174 524920
rect 678978 524456 679034 524512
rect 683394 503648 683450 503704
rect 679622 487192 679678 487248
rect 683210 500928 683266 500984
rect 681186 487600 681242 487656
rect 681002 486376 681058 486432
rect 683394 485560 683450 485616
rect 683210 483520 683266 483576
rect 676034 482704 676090 482760
rect 680358 481888 680414 481944
rect 675850 480664 675906 480720
rect 683118 481072 683174 481128
rect 672952 454316 672954 454336
rect 672954 454316 673006 454336
rect 673006 454316 673008 454336
rect 672952 454280 673008 454316
rect 674286 454316 674288 454336
rect 674288 454316 674340 454336
rect 674340 454316 674342 454336
rect 674286 454280 674342 454316
rect 674286 453908 674288 453928
rect 674288 453908 674340 453928
rect 674340 453908 674342 453928
rect 674286 453872 674342 453908
rect 676218 403300 676274 403336
rect 676218 403280 676220 403300
rect 676220 403280 676272 403300
rect 676272 403280 676274 403300
rect 672630 402464 672686 402520
rect 672446 401920 672502 401976
rect 673182 401648 673238 401704
rect 672814 399608 672870 399664
rect 672630 393896 672686 393952
rect 671894 393624 671950 393680
rect 671710 348880 671766 348936
rect 671710 331200 671766 331256
rect 671526 302232 671582 302288
rect 671710 278588 671766 278624
rect 671710 278568 671712 278588
rect 671712 278568 671764 278588
rect 671764 278568 671766 278588
rect 671710 263744 671766 263800
rect 672630 376216 672686 376272
rect 672354 357040 672410 357096
rect 672170 350104 672226 350160
rect 672170 335824 672226 335880
rect 672538 356224 672594 356280
rect 672354 312432 672410 312488
rect 672998 394984 673054 395040
rect 672998 380976 673054 381032
rect 673918 401376 673974 401432
rect 673366 400424 673422 400480
rect 673182 357448 673238 357504
rect 673734 395664 673790 395720
rect 673734 375400 673790 375456
rect 676586 402872 676642 402928
rect 674838 402192 674894 402248
rect 674838 401648 674894 401704
rect 676586 400832 676642 400888
rect 676034 399336 676090 399392
rect 674746 397296 674802 397352
rect 674562 396616 674618 396672
rect 679622 398384 679678 398440
rect 676218 397976 676274 398032
rect 676034 396092 676090 396128
rect 676034 396072 676036 396092
rect 676036 396072 676088 396092
rect 676088 396072 676090 396092
rect 678242 397568 678298 397624
rect 676218 394324 676274 394360
rect 676218 394304 676220 394324
rect 676220 394304 676272 394324
rect 676272 394304 676274 394324
rect 678242 387640 678298 387696
rect 675758 384920 675814 384976
rect 675114 382880 675170 382936
rect 675758 382200 675814 382256
rect 675390 380976 675446 381032
rect 675758 378664 675814 378720
rect 675758 377304 675814 377360
rect 675390 376216 675446 376272
rect 675114 375400 675170 375456
rect 675758 373632 675814 373688
rect 675390 372408 675446 372464
rect 674470 358264 674526 358320
rect 673918 356496 673974 356552
rect 673366 355816 673422 355872
rect 673274 355408 673330 355464
rect 672814 355000 672870 355056
rect 673090 353368 673146 353424
rect 672906 349696 672962 349752
rect 672722 348472 672778 348528
rect 672538 311616 672594 311672
rect 672538 305496 672594 305552
rect 671250 259528 671306 259584
rect 670698 257216 670754 257272
rect 671618 256264 671674 256320
rect 671158 245520 671214 245576
rect 670882 233860 670884 233880
rect 670884 233860 670936 233880
rect 670936 233860 670938 233880
rect 670882 233824 670938 233860
rect 670606 218184 670662 218240
rect 670514 216416 670570 216472
rect 670514 198192 670570 198248
rect 670790 177964 670792 177984
rect 670792 177964 670844 177984
rect 670844 177964 670846 177984
rect 670790 177928 670846 177964
rect 670422 171128 670478 171184
rect 669962 130872 670018 130928
rect 668950 125704 669006 125760
rect 668766 119176 668822 119232
rect 668950 118768 669006 118824
rect 668950 114280 669006 114336
rect 668766 112648 668822 112704
rect 670606 170312 670662 170368
rect 670422 155896 670478 155952
rect 671710 238584 671766 238640
rect 672538 285504 672594 285560
rect 672170 246200 672226 246256
rect 672170 240216 672226 240272
rect 671894 231920 671950 231976
rect 673090 340720 673146 340776
rect 672906 335552 672962 335608
rect 672906 324944 672962 325000
rect 673734 352552 673790 352608
rect 673550 349288 673606 349344
rect 673918 352144 673974 352200
rect 673734 333920 673790 333976
rect 673550 332696 673606 332752
rect 674286 351328 674342 351384
rect 675942 357856 675998 357912
rect 675942 356768 675998 356824
rect 674654 354592 674710 354648
rect 674470 351056 674526 351112
rect 674470 350512 674526 350568
rect 674286 338000 674342 338056
rect 673918 326848 673974 326904
rect 673918 311208 673974 311264
rect 673274 310800 673330 310856
rect 673366 309440 673422 309496
rect 673182 304272 673238 304328
rect 673182 287816 673238 287872
rect 672906 278568 672962 278624
rect 672538 265240 672594 265296
rect 672354 227024 672410 227080
rect 673182 266056 673238 266112
rect 673550 305904 673606 305960
rect 673826 291760 673882 291816
rect 673550 291488 673606 291544
rect 673642 287544 673698 287600
rect 673366 264968 673422 265024
rect 673458 264424 673514 264480
rect 673826 268096 673882 268152
rect 676034 350920 676090 350976
rect 676034 346568 676090 346624
rect 675114 340720 675170 340776
rect 675758 340176 675814 340232
rect 675482 339360 675538 339416
rect 674930 338680 674986 338736
rect 675114 338000 675170 338056
rect 675758 337864 675814 337920
rect 675758 336504 675814 336560
rect 674930 335824 674986 335880
rect 675114 335552 675170 335608
rect 675114 333920 675170 333976
rect 675114 332696 675170 332752
rect 675114 331200 675170 331256
rect 675022 327936 675078 327992
rect 675390 327936 675446 327992
rect 675390 326848 675446 326904
rect 675206 325624 675262 325680
rect 675022 324944 675078 325000
rect 676218 313928 676274 313984
rect 674838 312840 674894 312896
rect 675482 312044 675538 312080
rect 675482 312024 675484 312044
rect 675484 312024 675536 312044
rect 675536 312024 675538 312044
rect 674838 311888 674894 311944
rect 675482 310392 675538 310448
rect 674654 309984 674710 310040
rect 675942 309712 675998 309768
rect 675114 308352 675170 308408
rect 674930 307944 674986 308000
rect 674654 303864 674710 303920
rect 674378 267416 674434 267472
rect 674286 267008 674342 267064
rect 674102 266600 674158 266656
rect 676034 307536 676090 307592
rect 676034 307128 676090 307184
rect 678242 306720 678298 306776
rect 676586 304680 676642 304736
rect 676034 303456 676090 303512
rect 676034 301960 676090 302016
rect 676586 301552 676642 301608
rect 678978 306312 679034 306368
rect 676862 297336 676918 297392
rect 676034 296520 676090 296576
rect 675574 295704 675630 295760
rect 675758 294616 675814 294672
rect 675574 292168 675630 292224
rect 675390 291488 675446 291544
rect 675758 290944 675814 291000
rect 675114 287816 675170 287872
rect 675758 287000 675814 287056
rect 675114 285504 675170 285560
rect 675758 283600 675814 283656
rect 675758 282648 675814 282704
rect 674838 278296 674894 278352
rect 675666 281560 675722 281616
rect 676862 279384 676918 279440
rect 675482 278024 675538 278080
rect 675298 277344 675354 277400
rect 674838 273808 674894 273864
rect 674654 265784 674710 265840
rect 675114 264696 675170 264752
rect 673090 263336 673146 263392
rect 672906 259256 672962 259312
rect 673090 250688 673146 250744
rect 673090 249600 673146 249656
rect 673090 245248 673146 245304
rect 672906 242664 672962 242720
rect 674194 260888 674250 260944
rect 674654 262520 674710 262576
rect 673734 246200 673790 246256
rect 673826 245792 673882 245848
rect 674194 260072 674250 260128
rect 674378 258848 674434 258904
rect 673550 241848 673606 241904
rect 673274 241576 673330 241632
rect 672952 236716 672954 236736
rect 672954 236716 673006 236736
rect 673006 236716 673008 236736
rect 672952 236680 673008 236716
rect 673550 232464 673606 232520
rect 672032 225276 672088 225312
rect 672032 225256 672034 225276
rect 672034 225256 672086 225276
rect 672086 225256 672088 225276
rect 672154 225120 672210 225176
rect 671894 224984 671950 225040
rect 671818 224748 671820 224768
rect 671820 224748 671872 224768
rect 671872 224748 671874 224768
rect 671818 224712 671874 224748
rect 671480 224068 671482 224088
rect 671482 224068 671534 224088
rect 671534 224068 671536 224088
rect 671480 224032 671536 224068
rect 671342 177928 671398 177984
rect 670606 147600 670662 147656
rect 672078 224032 672134 224088
rect 672078 217504 672134 217560
rect 672078 216144 672134 216200
rect 672078 215600 672134 215656
rect 672078 214104 672134 214160
rect 672078 199688 672134 199744
rect 672722 226380 672724 226400
rect 672724 226380 672776 226400
rect 672776 226380 672778 226400
rect 672722 226344 672778 226380
rect 672602 226108 672604 226128
rect 672604 226108 672656 226128
rect 672656 226108 672658 226128
rect 672602 226072 672658 226108
rect 672492 225956 672548 225992
rect 672492 225936 672494 225956
rect 672494 225936 672546 225956
rect 672546 225936 672548 225956
rect 672378 225700 672380 225720
rect 672380 225700 672432 225720
rect 672432 225700 672434 225720
rect 672378 225664 672434 225700
rect 672446 220224 672502 220280
rect 672630 217912 672686 217968
rect 673458 228520 673514 228576
rect 673274 227024 673330 227080
rect 673550 226752 673606 226808
rect 673458 224712 673514 224768
rect 673274 222808 673330 222864
rect 673274 221040 673330 221096
rect 673090 220632 673146 220688
rect 673090 217368 673146 217424
rect 673090 216416 673146 216472
rect 673090 216144 673146 216200
rect 672722 213560 672778 213616
rect 672814 213288 672870 213344
rect 672538 213152 672594 213208
rect 672630 212064 672686 212120
rect 671986 171944 672042 172000
rect 671710 150048 671766 150104
rect 672446 175616 672502 175672
rect 672354 168272 672410 168328
rect 672170 168000 672226 168056
rect 671986 144880 672042 144936
rect 672354 166912 672410 166968
rect 672170 135088 672226 135144
rect 671342 131688 671398 131744
rect 670606 122440 670662 122496
rect 671526 129240 671582 129296
rect 672078 123256 672134 123312
rect 672078 118768 672134 118824
rect 672998 201320 673054 201376
rect 672998 200776 673054 200832
rect 673458 216824 673514 216880
rect 673458 216552 673514 216608
rect 673458 215328 673514 215384
rect 673274 197920 673330 197976
rect 673090 181464 673146 181520
rect 673366 176840 673422 176896
rect 672998 169088 673054 169144
rect 673090 168680 673146 168736
rect 674194 242120 674250 242176
rect 674838 260480 674894 260536
rect 674838 256264 674894 256320
rect 674838 254904 674894 254960
rect 676862 268504 676918 268560
rect 676218 268096 676274 268152
rect 676218 267688 676274 267744
rect 676402 264016 676458 264072
rect 676218 262792 676274 262848
rect 675482 258032 675538 258088
rect 675850 254904 675906 254960
rect 675482 250688 675538 250744
rect 675758 250280 675814 250336
rect 675298 250144 675354 250200
rect 675482 250008 675538 250064
rect 675758 246608 675814 246664
rect 675206 245792 675262 245848
rect 675206 245520 675262 245576
rect 674654 243480 674710 243536
rect 674470 241032 674526 241088
rect 675022 241576 675078 241632
rect 674838 237224 674894 237280
rect 674194 236680 674250 236736
rect 674378 232636 674380 232656
rect 674380 232636 674432 232656
rect 674432 232636 674434 232656
rect 674378 232600 674434 232636
rect 674562 232328 674618 232384
rect 674332 230016 674388 230072
rect 674674 230308 674730 230344
rect 674674 230288 674676 230308
rect 674676 230288 674728 230308
rect 674728 230288 674730 230308
rect 674470 229200 674526 229256
rect 674286 222400 674342 222456
rect 674838 226072 674894 226128
rect 673918 214376 673974 214432
rect 673918 177248 673974 177304
rect 673918 174392 673974 174448
rect 674838 221720 674894 221776
rect 675390 243480 675446 243536
rect 675482 242664 675538 242720
rect 675390 242120 675446 242176
rect 675390 241032 675446 241088
rect 675390 240216 675446 240272
rect 675390 238584 675446 238640
rect 675482 237224 675538 237280
rect 675482 236136 675538 236192
rect 675482 235456 675538 235512
rect 675022 221448 675078 221504
rect 675114 219000 675170 219056
rect 674930 218184 674986 218240
rect 674102 172896 674158 172952
rect 673734 170720 673790 170776
rect 673458 162424 673514 162480
rect 673090 152632 673146 152688
rect 673182 151272 673238 151328
rect 673734 158752 673790 158808
rect 673550 156440 673606 156496
rect 673366 132096 673422 132152
rect 674102 161744 674158 161800
rect 673918 129648 673974 129704
rect 673366 126520 673422 126576
rect 673182 124888 673238 124944
rect 672814 124072 672870 124128
rect 673090 122984 673146 123040
rect 672630 120808 672686 120864
rect 672906 120672 672962 120728
rect 672354 115776 672410 115832
rect 672906 111016 672962 111072
rect 672998 106120 673054 106176
rect 673182 104624 673238 104680
rect 668766 104488 668822 104544
rect 668582 102856 668638 102912
rect 673918 124480 673974 124536
rect 674470 214920 674526 214976
rect 674654 213696 674710 213752
rect 675850 233860 675852 233880
rect 675852 233860 675904 233880
rect 675904 233860 675906 233880
rect 675850 233824 675906 233860
rect 675850 232636 675852 232656
rect 675852 232636 675904 232656
rect 675904 232636 675906 232656
rect 675850 232600 675906 232636
rect 676034 232328 676090 232384
rect 676494 230152 676550 230208
rect 675482 228520 675538 228576
rect 675482 225664 675538 225720
rect 675850 225120 675906 225176
rect 675482 219816 675538 219872
rect 675482 218592 675538 218648
rect 676034 221856 676090 221912
rect 675666 217912 675722 217968
rect 675666 215600 675722 215656
rect 676770 227024 676826 227080
rect 676954 226752 677010 226808
rect 678242 223760 678298 223816
rect 683394 223080 683450 223136
rect 683210 222672 683266 222728
rect 675666 214648 675722 214704
rect 676034 214512 676090 214568
rect 675850 214376 675906 214432
rect 675298 212472 675354 212528
rect 676034 211384 676090 211440
rect 675114 206896 675170 206952
rect 674746 204992 674802 205048
rect 674930 204176 674986 204232
rect 675390 204992 675446 205048
rect 675390 204176 675446 204232
rect 674470 197104 674526 197160
rect 674930 202816 674986 202872
rect 675758 202680 675814 202736
rect 675482 201320 675538 201376
rect 674930 199688 674986 199744
rect 675758 199960 675814 200016
rect 675114 198464 675170 198520
rect 675482 198192 675538 198248
rect 675390 197104 675446 197160
rect 675758 194520 675814 194576
rect 675758 193160 675814 193216
rect 675666 192752 675722 192808
rect 676034 189080 676090 189136
rect 675114 188808 675170 188864
rect 675850 180240 675906 180296
rect 675850 177656 675906 177712
rect 676218 181192 676274 181248
rect 676218 178880 676274 178936
rect 674746 176024 674802 176080
rect 674562 175208 674618 175264
rect 674286 153176 674342 153232
rect 674838 173984 674894 174040
rect 681002 173576 681058 173632
rect 676034 173168 676090 173224
rect 676586 169904 676642 169960
rect 675666 167456 675722 167512
rect 675206 162016 675262 162072
rect 676586 166368 676642 166424
rect 682382 171536 682438 171592
rect 683118 167864 683174 167920
rect 681002 162696 681058 162752
rect 675850 162016 675906 162072
rect 683118 162016 683174 162072
rect 675482 161472 675538 161528
rect 675758 156984 675814 157040
rect 675298 156440 675354 156496
rect 675114 155896 675170 155952
rect 675758 155760 675814 155816
rect 675114 152632 675170 152688
rect 675758 151408 675814 151464
rect 675114 151272 675170 151328
rect 674930 150320 674986 150376
rect 675758 148416 675814 148472
rect 675114 147600 675170 147656
rect 675390 147600 675446 147656
rect 675114 144880 675170 144936
rect 675850 134544 675906 134600
rect 676494 133048 676550 133104
rect 674654 131280 674710 131336
rect 674470 130464 674526 130520
rect 676218 130192 676274 130248
rect 675022 128832 675078 128888
rect 674378 128424 674434 128480
rect 674102 117408 674158 117464
rect 673918 106936 673974 106992
rect 674654 124072 674710 124128
rect 674838 123664 674894 123720
rect 674838 122984 674894 123040
rect 676218 127744 676274 127800
rect 676402 127744 676458 127800
rect 679622 126112 679678 126168
rect 675206 117000 675262 117056
rect 682382 125296 682438 125352
rect 682382 117272 682438 117328
rect 675850 117000 675906 117056
rect 675482 115776 675538 115832
rect 675758 112376 675814 112432
rect 675758 111696 675814 111752
rect 675758 111288 675814 111344
rect 675758 110336 675814 110392
rect 675758 108160 675814 108216
rect 675390 106936 675446 106992
rect 675114 106120 675170 106176
rect 675114 104624 675170 104680
rect 675390 101904 675446 101960
rect 673366 100952 673422 101008
rect 675114 100952 675170 101008
rect 625618 93608 625674 93664
rect 637026 96872 637082 96928
rect 641994 96464 642050 96520
rect 635738 95376 635794 95432
rect 647146 94968 647202 95024
rect 626446 94424 626502 94480
rect 626446 92792 626502 92848
rect 625802 91976 625858 92032
rect 647514 92384 647570 92440
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 625250 89564 625252 89584
rect 625252 89564 625304 89584
rect 625304 89564 625306 89584
rect 625250 89528 625306 89564
rect 624974 88712 625030 88768
rect 625158 87896 625214 87952
rect 625342 87080 625398 87136
rect 648250 89528 648306 89584
rect 625158 86300 625160 86320
rect 625160 86300 625212 86320
rect 625212 86300 625214 86320
rect 625158 86264 625214 86300
rect 625158 85448 625214 85504
rect 625342 84632 625398 84688
rect 625158 83816 625214 83872
rect 628746 83272 628802 83328
rect 629206 81640 629262 81696
rect 624422 77288 624478 77344
rect 633898 78512 633954 78568
rect 633898 77288 633954 77344
rect 639602 78104 639658 78160
rect 646134 74160 646190 74216
rect 646318 71712 646374 71768
rect 647238 68856 647294 68912
rect 646502 67088 646558 67144
rect 646134 64368 646190 64424
rect 648618 62056 648674 62112
rect 647238 59200 647294 59256
rect 649998 87080 650054 87136
rect 655242 94152 655298 94208
rect 654322 91432 654378 91488
rect 655426 93336 655482 93392
rect 655426 90652 655428 90672
rect 655428 90652 655480 90672
rect 655480 90652 655482 90672
rect 655426 90616 655482 90652
rect 655794 89800 655850 89856
rect 663706 92792 663762 92848
rect 664166 89800 664222 89856
rect 665178 93336 665234 93392
rect 665362 91704 665418 91760
rect 665546 90616 665602 90672
rect 664350 88984 664406 89040
rect 650550 84632 650606 84688
rect 650366 82184 650422 82240
rect 648802 57296 648858 57352
rect 661590 48454 661646 48510
rect 553674 48048 553730 48104
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 545670 47232 545726 47288
rect 465262 46688 465318 46744
rect 662418 47368 662474 47424
rect 464342 44104 464398 44160
rect 471058 43424 471114 43480
rect 465814 43152 465870 43208
rect 461950 42200 462006 42256
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 40296 141754 40352
<< metal3 >>
rect 185025 1002146 185091 1002149
rect 185012 1002144 185091 1002146
rect 185012 1002088 185030 1002144
rect 185086 1002088 185091 1002144
rect 185012 1002086 185091 1002088
rect 185025 1002083 185091 1002086
rect 82169 1002010 82235 1002013
rect 133689 1002010 133755 1002013
rect 82156 1002008 82235 1002010
rect 82156 1001952 82174 1002008
rect 82230 1001952 82235 1002008
rect 82156 1001950 82235 1001952
rect 133676 1002008 133755 1002010
rect 133676 1001952 133694 1002008
rect 133750 1001952 133755 1002008
rect 133676 1001950 133755 1001952
rect 82169 1001947 82235 1001950
rect 133689 1001947 133755 1001950
rect 483013 1002010 483079 1002013
rect 534993 1002010 535059 1002013
rect 636193 1002010 636259 1002013
rect 483013 1002008 483092 1002010
rect 483013 1001952 483018 1002008
rect 483074 1001952 483092 1002008
rect 483013 1001950 483092 1001952
rect 534980 1002008 535059 1002010
rect 534980 1001952 534998 1002008
rect 535054 1001952 535059 1002008
rect 534980 1001950 535059 1001952
rect 636180 1002008 636259 1002010
rect 636180 1001952 636198 1002008
rect 636254 1001952 636259 1002008
rect 636180 1001950 636259 1001952
rect 483013 1001947 483079 1001950
rect 534993 1001947 535059 1001950
rect 636193 1001947 636259 1001950
rect 232957 997388 233023 997389
rect 232957 997384 233004 997388
rect 233068 997386 233074 997388
rect 232957 997328 232962 997384
rect 232957 997324 233004 997328
rect 233068 997326 233114 997386
rect 233068 997324 233074 997326
rect 232957 997323 233023 997324
rect 240133 997250 240199 997253
rect 240550 997250 240610 997628
rect 285397 997388 285463 997389
rect 285397 997384 285444 997388
rect 285508 997386 285514 997388
rect 292573 997386 292639 997389
rect 293174 997386 293234 997628
rect 404310 997389 404370 997628
rect 285397 997328 285402 997384
rect 285397 997324 285444 997328
rect 285508 997326 285554 997386
rect 292573 997384 293234 997386
rect 292573 997328 292578 997384
rect 292634 997328 293234 997384
rect 292573 997326 293234 997328
rect 387517 997388 387583 997389
rect 387517 997384 387564 997388
rect 387628 997386 387634 997388
rect 387517 997328 387522 997384
rect 285508 997324 285514 997326
rect 285397 997323 285463 997324
rect 292573 997323 292639 997326
rect 387517 997324 387564 997328
rect 387628 997326 387674 997386
rect 404310 997384 404419 997389
rect 404310 997328 404358 997384
rect 404414 997328 404419 997384
rect 404310 997326 404419 997328
rect 387628 997324 387634 997326
rect 387517 997323 387583 997324
rect 404353 997323 404419 997326
rect 240133 997248 240610 997250
rect 240133 997192 240138 997248
rect 240194 997192 240610 997248
rect 240133 997190 240610 997192
rect 240133 997187 240199 997190
rect 232998 990932 233004 990996
rect 233068 990994 233074 990996
rect 235901 990994 235967 990997
rect 233068 990992 235967 990994
rect 233068 990936 235906 990992
rect 235962 990936 235967 990992
rect 233068 990934 235967 990936
rect 233068 990932 233074 990934
rect 235901 990931 235967 990934
rect 387558 990932 387564 990996
rect 387628 990994 387634 990996
rect 389173 990994 389239 990997
rect 387628 990992 389239 990994
rect 387628 990936 389178 990992
rect 389234 990936 389239 990992
rect 387628 990934 389239 990936
rect 387628 990932 387634 990934
rect 389173 990931 389239 990934
rect 285438 987940 285444 988004
rect 285508 988002 285514 988004
rect 286961 988002 287027 988005
rect 285508 988000 287027 988002
rect 285508 987944 286966 988000
rect 287022 987944 287027 988000
rect 285508 987942 287027 987944
rect 285508 987940 285514 987942
rect 286961 987939 287027 987942
rect 238661 984058 238727 984061
rect 238661 984056 238770 984058
rect 238661 984000 238666 984056
rect 238722 984000 238770 984056
rect 238661 983995 238770 984000
rect 235901 983786 235967 983789
rect 235901 983784 236378 983786
rect 235901 983728 235906 983784
rect 235962 983728 236378 983784
rect 235901 983726 236378 983728
rect 235901 983723 235967 983726
rect 81341 983514 81407 983517
rect 184933 983514 184999 983517
rect 81341 983512 81604 983514
rect 81341 983456 81346 983512
rect 81402 983456 81604 983512
rect 81341 983454 81604 983456
rect 184933 983512 185564 983514
rect 184933 983456 184938 983512
rect 184994 983456 185564 983512
rect 236318 983484 236378 983726
rect 238710 983484 238770 983995
rect 240133 983786 240199 983789
rect 286961 983786 287027 983789
rect 292573 983786 292639 983789
rect 535453 983786 535519 983789
rect 636193 983786 636259 983789
rect 240133 983784 241346 983786
rect 240133 983728 240138 983784
rect 240194 983728 241346 983784
rect 240133 983726 241346 983728
rect 240133 983723 240199 983726
rect 241286 983484 241346 983726
rect 286961 983784 288082 983786
rect 286961 983728 286966 983784
rect 287022 983728 288082 983784
rect 286961 983726 288082 983728
rect 286961 983723 287027 983726
rect 288022 983484 288082 983726
rect 292573 983784 293234 983786
rect 292573 983728 292578 983784
rect 292634 983728 293234 983784
rect 292573 983726 293234 983728
rect 292573 983723 292639 983726
rect 293174 983484 293234 983726
rect 535453 983784 535562 983786
rect 535453 983728 535458 983784
rect 535514 983728 535562 983784
rect 535453 983723 535562 983728
rect 391933 983514 391999 983517
rect 394417 983514 394483 983517
rect 399753 983514 399819 983517
rect 391644 983512 391999 983514
rect 184933 983454 185564 983456
rect 391644 983456 391938 983512
rect 391994 983456 391999 983512
rect 391644 983454 391999 983456
rect 394220 983512 394483 983514
rect 394220 983456 394422 983512
rect 394478 983456 394483 983512
rect 394220 983454 394483 983456
rect 399556 983512 399819 983514
rect 399556 983456 399758 983512
rect 399814 983456 399819 983512
rect 535502 983484 535562 983723
rect 636150 983784 636259 983786
rect 636150 983728 636198 983784
rect 636254 983728 636259 983784
rect 636150 983723 636259 983728
rect 636150 983484 636210 983723
rect 399556 983454 399819 983456
rect 81341 983451 81407 983454
rect 184933 983451 184999 983454
rect 391933 983451 391999 983454
rect 394417 983451 394483 983454
rect 399753 983451 399819 983454
rect 132493 982562 132559 982565
rect 483841 982562 483907 982565
rect 132493 982560 133676 982562
rect 132493 982504 132498 982560
rect 132554 982504 133676 982560
rect 132493 982502 133676 982504
rect 483644 982560 483907 982562
rect 483644 982504 483846 982560
rect 483902 982504 483907 982560
rect 483644 982502 483907 982504
rect 132493 982499 132559 982502
rect 483841 982499 483907 982502
rect 289721 980930 289787 980933
rect 290414 980930 290474 981036
rect 289721 980928 290474 980930
rect 289721 980872 289726 980928
rect 289782 980872 290474 980928
rect 289721 980870 290474 980872
rect 289721 980867 289787 980870
rect 30097 960258 30163 960261
rect 30084 960256 30163 960258
rect 30084 960200 30102 960256
rect 30158 960200 30163 960256
rect 30084 960198 30163 960200
rect 30097 960195 30163 960198
rect 651373 959170 651439 959173
rect 649980 959168 651439 959170
rect 649980 959112 651378 959168
rect 651434 959112 651439 959168
rect 649980 959110 651439 959112
rect 651373 959107 651439 959110
rect 677409 959170 677475 959173
rect 677409 959168 677764 959170
rect 677409 959112 677414 959168
rect 677470 959112 677764 959168
rect 677409 959110 677764 959112
rect 677409 959107 677475 959110
rect 63401 959034 63467 959037
rect 63401 959032 64676 959034
rect 63401 958976 63406 959032
rect 63462 958976 64676 959032
rect 63401 958974 64676 958976
rect 63401 958971 63467 958974
rect 676029 897154 676095 897157
rect 676029 897152 676292 897154
rect 676029 897096 676034 897152
rect 676090 897096 676292 897152
rect 676029 897094 676292 897096
rect 676029 897091 676095 897094
rect 675845 896746 675911 896749
rect 675845 896744 676292 896746
rect 675845 896688 675850 896744
rect 675906 896688 676292 896744
rect 675845 896686 676292 896688
rect 675845 896683 675911 896686
rect 676029 896338 676095 896341
rect 676029 896336 676292 896338
rect 676029 896280 676034 896336
rect 676090 896280 676292 896336
rect 676029 896278 676292 896280
rect 676029 896275 676095 896278
rect 675845 895522 675911 895525
rect 675845 895520 676292 895522
rect 675845 895464 675850 895520
rect 675906 895464 676292 895520
rect 675845 895462 676292 895464
rect 675845 895459 675911 895462
rect 676029 894706 676095 894709
rect 676029 894704 676292 894706
rect 676029 894648 676034 894704
rect 676090 894648 676292 894704
rect 676029 894646 676292 894648
rect 676029 894643 676095 894646
rect 675845 893890 675911 893893
rect 675845 893888 676292 893890
rect 675845 893832 675850 893888
rect 675906 893832 676292 893888
rect 675845 893830 676292 893832
rect 675845 893827 675911 893830
rect 676029 893074 676095 893077
rect 676029 893072 676292 893074
rect 676029 893016 676034 893072
rect 676090 893016 676292 893072
rect 676029 893014 676292 893016
rect 676029 893011 676095 893014
rect 676029 892666 676095 892669
rect 676029 892664 676292 892666
rect 676029 892608 676034 892664
rect 676090 892608 676292 892664
rect 676029 892606 676292 892608
rect 676029 892603 676095 892606
rect 675886 892196 675892 892260
rect 675956 892258 675962 892260
rect 675956 892198 676292 892258
rect 675956 892196 675962 892198
rect 679617 891850 679683 891853
rect 679604 891848 679683 891850
rect 679604 891792 679622 891848
rect 679678 891792 679683 891848
rect 679604 891790 679683 891792
rect 679617 891787 679683 891790
rect 676029 891442 676095 891445
rect 676029 891440 676292 891442
rect 676029 891384 676034 891440
rect 676090 891384 676292 891440
rect 676029 891382 676292 891384
rect 676029 891379 676095 891382
rect 675293 891034 675359 891037
rect 675293 891032 676292 891034
rect 675293 890976 675298 891032
rect 675354 890976 676292 891032
rect 675293 890974 676292 890976
rect 675293 890971 675359 890974
rect 680997 890626 681063 890629
rect 680997 890624 681076 890626
rect 680997 890568 681002 890624
rect 681058 890568 681076 890624
rect 680997 890566 681076 890568
rect 680997 890563 681063 890566
rect 676029 890218 676095 890221
rect 676029 890216 676292 890218
rect 676029 890160 676034 890216
rect 676090 890160 676292 890216
rect 676029 890158 676292 890160
rect 676029 890155 676095 890158
rect 678237 889810 678303 889813
rect 678237 889808 678316 889810
rect 678237 889752 678242 889808
rect 678298 889752 678316 889808
rect 678237 889750 678316 889752
rect 678237 889747 678303 889750
rect 676029 889402 676095 889405
rect 676029 889400 676292 889402
rect 676029 889344 676034 889400
rect 676090 889344 676292 889400
rect 676029 889342 676292 889344
rect 676029 889339 676095 889342
rect 676029 888994 676095 888997
rect 676029 888992 676292 888994
rect 676029 888936 676034 888992
rect 676090 888936 676292 888992
rect 676029 888934 676292 888936
rect 676029 888931 676095 888934
rect 676029 888586 676095 888589
rect 676029 888584 676292 888586
rect 676029 888528 676034 888584
rect 676090 888528 676292 888584
rect 676029 888526 676292 888528
rect 676029 888523 676095 888526
rect 683113 888178 683179 888181
rect 683100 888176 683179 888178
rect 683100 888120 683118 888176
rect 683174 888120 683179 888176
rect 683100 888118 683179 888120
rect 683113 888115 683179 888118
rect 675886 887708 675892 887772
rect 675956 887770 675962 887772
rect 675956 887710 676292 887770
rect 675956 887708 675962 887710
rect 676029 887362 676095 887365
rect 676029 887360 676292 887362
rect 676029 887304 676034 887360
rect 676090 887304 676292 887360
rect 676029 887302 676292 887304
rect 676029 887299 676095 887302
rect 676029 886954 676095 886957
rect 676029 886952 676292 886954
rect 676029 886896 676034 886952
rect 676090 886896 676292 886952
rect 676029 886894 676292 886896
rect 676029 886891 676095 886894
rect 683070 886138 683130 886516
rect 675894 886108 683130 886138
rect 675894 886078 683100 886108
rect 675702 885804 675708 885868
rect 675772 885866 675778 885868
rect 675894 885866 675954 886078
rect 675772 885806 675954 885866
rect 675772 885804 675778 885806
rect 676029 885730 676095 885733
rect 676029 885728 676292 885730
rect 676029 885672 676034 885728
rect 676090 885672 676292 885728
rect 676029 885670 676292 885672
rect 676029 885667 676095 885670
rect 675518 880636 675524 880700
rect 675588 880698 675594 880700
rect 680997 880698 681063 880701
rect 675588 880696 681063 880698
rect 675588 880640 681002 880696
rect 681058 880640 681063 880696
rect 675588 880638 681063 880640
rect 675588 880636 675594 880638
rect 680997 880635 681063 880638
rect 676254 880364 676260 880428
rect 676324 880426 676330 880428
rect 683113 880426 683179 880429
rect 676324 880424 683179 880426
rect 676324 880368 683118 880424
rect 683174 880368 683179 880424
rect 676324 880366 683179 880368
rect 676324 880364 676330 880366
rect 683113 880363 683179 880366
rect 675334 878460 675340 878524
rect 675404 878522 675410 878524
rect 675661 878522 675727 878525
rect 675404 878520 675727 878522
rect 675404 878464 675666 878520
rect 675722 878464 675727 878520
rect 675404 878462 675727 878464
rect 675404 878460 675410 878462
rect 675661 878459 675727 878462
rect 675201 877164 675267 877165
rect 675150 877100 675156 877164
rect 675220 877162 675267 877164
rect 675220 877160 675312 877162
rect 675262 877104 675312 877160
rect 675220 877102 675312 877104
rect 675220 877100 675267 877102
rect 675201 877099 675267 877100
rect 674833 874714 674899 874717
rect 675477 874714 675543 874717
rect 674833 874712 675543 874714
rect 674833 874656 674838 874712
rect 674894 874656 675482 874712
rect 675538 874656 675543 874712
rect 674833 874654 675543 874656
rect 674833 874651 674899 874654
rect 675477 874651 675543 874654
rect 675334 874108 675340 874172
rect 675404 874170 675410 874172
rect 675569 874170 675635 874173
rect 675404 874168 675635 874170
rect 675404 874112 675574 874168
rect 675630 874112 675635 874168
rect 675404 874110 675635 874112
rect 675404 874108 675410 874110
rect 675569 874107 675635 874110
rect 675753 873082 675819 873085
rect 676254 873082 676260 873084
rect 675753 873080 676260 873082
rect 675753 873024 675758 873080
rect 675814 873024 676260 873080
rect 675753 873022 676260 873024
rect 675753 873019 675819 873022
rect 676254 873020 676260 873022
rect 676324 873020 676330 873084
rect 675017 872810 675083 872813
rect 676438 872810 676444 872812
rect 675017 872808 676444 872810
rect 675017 872752 675022 872808
rect 675078 872752 676444 872808
rect 675017 872750 676444 872752
rect 675017 872747 675083 872750
rect 676438 872748 676444 872750
rect 676508 872748 676514 872812
rect 675150 870436 675156 870500
rect 675220 870498 675226 870500
rect 675385 870498 675451 870501
rect 675220 870496 675451 870498
rect 675220 870440 675390 870496
rect 675446 870440 675451 870496
rect 675220 870438 675451 870440
rect 675220 870436 675226 870438
rect 675385 870435 675451 870438
rect 651465 868594 651531 868597
rect 649950 868592 651531 868594
rect 649950 868536 651470 868592
rect 651526 868536 651531 868592
rect 649950 868534 651531 868536
rect 649950 868246 650010 868534
rect 651465 868531 651531 868534
rect 652017 867642 652083 867645
rect 649950 867640 652083 867642
rect 649950 867584 652022 867640
rect 652078 867584 652083 867640
rect 649950 867582 652083 867584
rect 649950 867064 650010 867582
rect 652017 867579 652083 867582
rect 651465 866282 651531 866285
rect 649950 866280 651531 866282
rect 649950 866224 651470 866280
rect 651526 866224 651531 866280
rect 649950 866222 651531 866224
rect 649950 865882 650010 866222
rect 651465 866219 651531 866222
rect 675293 865738 675359 865741
rect 675702 865738 675708 865740
rect 675293 865736 675708 865738
rect 675293 865680 675298 865736
rect 675354 865680 675708 865736
rect 675293 865678 675708 865680
rect 675293 865675 675359 865678
rect 675702 865676 675708 865678
rect 675772 865676 675778 865740
rect 675753 865466 675819 865469
rect 676070 865466 676076 865468
rect 675753 865464 676076 865466
rect 675753 865408 675758 865464
rect 675814 865408 676076 865464
rect 675753 865406 676076 865408
rect 675753 865403 675819 865406
rect 676070 865404 676076 865406
rect 676140 865404 676146 865468
rect 651373 865194 651439 865197
rect 649950 865192 651439 865194
rect 649950 865136 651378 865192
rect 651434 865136 651439 865192
rect 649950 865134 651439 865136
rect 649950 864700 650010 865134
rect 651373 865131 651439 865134
rect 675661 865058 675727 865061
rect 675886 865058 675892 865060
rect 675661 865056 675892 865058
rect 675661 865000 675666 865056
rect 675722 865000 675892 865056
rect 675661 864998 675892 865000
rect 675661 864995 675727 864998
rect 675886 864996 675892 864998
rect 675956 864996 675962 865060
rect 651465 863834 651531 863837
rect 649766 863832 651531 863834
rect 649766 863776 651470 863832
rect 651526 863776 651531 863832
rect 649766 863774 651531 863776
rect 649766 863518 649826 863774
rect 651465 863771 651531 863774
rect 651465 862338 651531 862341
rect 649766 862336 651531 862338
rect 649766 862280 651470 862336
rect 651526 862280 651531 862336
rect 649766 862278 651531 862280
rect 651465 862275 651531 862278
rect 35617 818002 35683 818005
rect 35574 818000 35683 818002
rect 35574 817944 35622 818000
rect 35678 817944 35683 818000
rect 35574 817939 35683 817944
rect 35574 817700 35634 817939
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 35433 816914 35499 816917
rect 35420 816912 35499 816914
rect 35420 816856 35438 816912
rect 35494 816856 35499 816912
rect 35420 816854 35499 816856
rect 35433 816851 35499 816854
rect 35801 816098 35867 816101
rect 35788 816096 35867 816098
rect 35788 816040 35806 816096
rect 35862 816040 35867 816096
rect 35788 816038 35867 816040
rect 35801 816035 35867 816038
rect 35617 815282 35683 815285
rect 35604 815280 35683 815282
rect 35604 815224 35622 815280
rect 35678 815224 35683 815280
rect 35604 815222 35683 815224
rect 35617 815219 35683 815222
rect 35801 814466 35867 814469
rect 35788 814464 35867 814466
rect 35788 814408 35806 814464
rect 35862 814408 35867 814464
rect 35788 814406 35867 814408
rect 35801 814403 35867 814406
rect 41321 813650 41387 813653
rect 41308 813648 41387 813650
rect 41308 813592 41326 813648
rect 41382 813592 41387 813648
rect 41308 813590 41387 813592
rect 41321 813587 41387 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 40953 812834 41019 812837
rect 40940 812832 41019 812834
rect 40940 812776 40958 812832
rect 41014 812776 41019 812832
rect 40940 812774 41019 812776
rect 40953 812771 41019 812774
rect 41321 812426 41387 812429
rect 41308 812424 41387 812426
rect 41308 812368 41326 812424
rect 41382 812368 41387 812424
rect 41308 812366 41387 812368
rect 41321 812363 41387 812366
rect 41137 812018 41203 812021
rect 41124 812016 41203 812018
rect 41124 811960 41142 812016
rect 41198 811960 41203 812016
rect 41124 811958 41203 811960
rect 41137 811955 41203 811958
rect 37917 811610 37983 811613
rect 37917 811608 37996 811610
rect 37917 811552 37922 811608
rect 37978 811552 37996 811608
rect 37917 811550 37996 811552
rect 37917 811547 37983 811550
rect 34513 811202 34579 811205
rect 34500 811200 34579 811202
rect 34500 811144 34518 811200
rect 34574 811144 34579 811200
rect 34500 811142 34579 811144
rect 34513 811139 34579 811142
rect 32581 810794 32647 810797
rect 32581 810792 32660 810794
rect 32581 810736 32586 810792
rect 32642 810736 32660 810792
rect 32581 810734 32660 810736
rect 32581 810731 32647 810734
rect 41965 810386 42031 810389
rect 41492 810384 42031 810386
rect 41492 810328 41970 810384
rect 42026 810328 42031 810384
rect 41492 810326 42031 810328
rect 41965 810323 42031 810326
rect 31017 809978 31083 809981
rect 31004 809976 31083 809978
rect 31004 809920 31022 809976
rect 31078 809920 31083 809976
rect 31004 809918 31083 809920
rect 31017 809915 31083 809918
rect 41781 809980 41847 809981
rect 41781 809976 41828 809980
rect 41892 809978 41898 809980
rect 41781 809920 41786 809976
rect 41781 809916 41828 809920
rect 41892 809918 41938 809978
rect 41892 809916 41898 809918
rect 41781 809915 41847 809916
rect 36537 809570 36603 809573
rect 36524 809568 36603 809570
rect 36524 809512 36542 809568
rect 36598 809512 36603 809568
rect 36524 809510 36603 809512
rect 36537 809507 36603 809510
rect 41321 809162 41387 809165
rect 41308 809160 41387 809162
rect 41308 809104 41326 809160
rect 41382 809104 41387 809160
rect 41308 809102 41387 809104
rect 41321 809099 41387 809102
rect 41781 808754 41847 808757
rect 41492 808752 41847 808754
rect 41492 808696 41786 808752
rect 41842 808696 41847 808752
rect 41492 808694 41847 808696
rect 41781 808691 41847 808694
rect 41137 808346 41203 808349
rect 41124 808344 41203 808346
rect 41124 808288 41142 808344
rect 41198 808288 41203 808344
rect 41124 808286 41203 808288
rect 41137 808283 41203 808286
rect 41822 807938 41828 807940
rect 41492 807878 41828 807938
rect 41822 807876 41828 807878
rect 41892 807876 41898 807940
rect 41321 807530 41387 807533
rect 41308 807528 41387 807530
rect 41308 807472 41326 807528
rect 41382 807472 41387 807528
rect 41308 807470 41387 807472
rect 41321 807467 41387 807470
rect 41094 806717 41154 807092
rect 41094 806712 41203 806717
rect 41094 806684 41142 806712
rect 41124 806656 41142 806684
rect 41198 806656 41203 806712
rect 41124 806654 41203 806656
rect 41137 806651 41203 806654
rect 41321 806306 41387 806309
rect 41308 806304 41387 806306
rect 41308 806248 41326 806304
rect 41382 806248 41387 806304
rect 41308 806246 41387 806248
rect 41321 806243 41387 806246
rect 40534 805564 40540 805628
rect 40604 805626 40610 805628
rect 41965 805626 42031 805629
rect 40604 805624 42031 805626
rect 40604 805568 41970 805624
rect 42026 805568 42031 805624
rect 40604 805566 42031 805568
rect 40604 805564 40610 805566
rect 41965 805563 42031 805566
rect 40718 805156 40724 805220
rect 40788 805218 40794 805220
rect 41781 805218 41847 805221
rect 40788 805216 41847 805218
rect 40788 805160 41786 805216
rect 41842 805160 41847 805216
rect 40788 805158 41847 805160
rect 40788 805156 40794 805158
rect 41781 805155 41847 805158
rect 40902 804748 40908 804812
rect 40972 804810 40978 804812
rect 41822 804810 41828 804812
rect 40972 804750 41828 804810
rect 40972 804748 40978 804750
rect 41822 804748 41828 804750
rect 41892 804748 41898 804812
rect 32581 802498 32647 802501
rect 41822 802498 41828 802500
rect 32581 802496 41828 802498
rect 32581 802440 32586 802496
rect 32642 802440 41828 802496
rect 32581 802438 41828 802440
rect 32581 802435 32647 802438
rect 41822 802436 41828 802438
rect 41892 802436 41898 802500
rect 42149 801004 42215 801005
rect 42149 801000 42196 801004
rect 42260 801002 42266 801004
rect 42149 800944 42154 801000
rect 42149 800940 42196 800944
rect 42260 800942 42306 801002
rect 42260 800940 42266 800942
rect 42149 800939 42215 800940
rect 40493 800730 40559 800733
rect 41086 800730 41092 800732
rect 40493 800728 41092 800730
rect 40493 800672 40498 800728
rect 40554 800672 41092 800728
rect 40493 800670 41092 800672
rect 40493 800667 40559 800670
rect 41086 800668 41092 800670
rect 41156 800668 41162 800732
rect 39757 800594 39823 800597
rect 40350 800594 40356 800596
rect 39757 800592 40356 800594
rect 39757 800536 39762 800592
rect 39818 800536 40356 800592
rect 39757 800534 40356 800536
rect 39757 800531 39823 800534
rect 40350 800532 40356 800534
rect 40420 800532 40426 800596
rect 42149 797330 42215 797333
rect 43621 797330 43687 797333
rect 42149 797328 43687 797330
rect 42149 797272 42154 797328
rect 42210 797272 43626 797328
rect 43682 797272 43687 797328
rect 42149 797270 43687 797272
rect 42149 797267 42215 797270
rect 43621 797267 43687 797270
rect 41086 796180 41092 796244
rect 41156 796242 41162 796244
rect 41781 796242 41847 796245
rect 41156 796240 41847 796242
rect 41156 796184 41786 796240
rect 41842 796184 41847 796240
rect 41156 796182 41847 796184
rect 41156 796180 41162 796182
rect 41781 796179 41847 796182
rect 40902 794820 40908 794884
rect 40972 794882 40978 794884
rect 41781 794882 41847 794885
rect 40972 794880 41847 794882
rect 40972 794824 41786 794880
rect 41842 794824 41847 794880
rect 40972 794822 41847 794824
rect 40972 794820 40978 794822
rect 41781 794819 41847 794822
rect 42149 794476 42215 794477
rect 42149 794474 42196 794476
rect 42104 794472 42196 794474
rect 42104 794416 42154 794472
rect 42104 794414 42196 794416
rect 42149 794412 42196 794414
rect 42260 794412 42266 794476
rect 42149 794411 42215 794412
rect 40350 793052 40356 793116
rect 40420 793114 40426 793116
rect 41781 793114 41847 793117
rect 40420 793112 41847 793114
rect 40420 793056 41786 793112
rect 41842 793056 41847 793112
rect 40420 793054 41847 793056
rect 40420 793052 40426 793054
rect 41781 793051 41847 793054
rect 40718 790604 40724 790668
rect 40788 790666 40794 790668
rect 41781 790666 41847 790669
rect 40788 790664 41847 790666
rect 40788 790608 41786 790664
rect 41842 790608 41847 790664
rect 40788 790606 41847 790608
rect 40788 790604 40794 790606
rect 41781 790603 41847 790606
rect 62205 790530 62271 790533
rect 62205 790528 64706 790530
rect 62205 790472 62210 790528
rect 62266 790472 64706 790528
rect 62205 790470 64706 790472
rect 62205 790467 62271 790470
rect 64646 790304 64706 790470
rect 40534 789380 40540 789444
rect 40604 789442 40610 789444
rect 41781 789442 41847 789445
rect 40604 789440 41847 789442
rect 40604 789384 41786 789440
rect 41842 789384 41847 789440
rect 40604 789382 41847 789384
rect 40604 789380 40610 789382
rect 41781 789379 41847 789382
rect 41638 789108 41644 789172
rect 41708 789170 41714 789172
rect 42241 789170 42307 789173
rect 41708 789168 42307 789170
rect 41708 789112 42246 789168
rect 42302 789112 42307 789168
rect 41708 789110 42307 789112
rect 41708 789108 41714 789110
rect 42241 789107 42307 789110
rect 62113 789170 62179 789173
rect 62113 789168 64706 789170
rect 62113 789112 62118 789168
rect 62174 789112 64706 789168
rect 62113 789110 64706 789112
rect 62113 789107 62179 789110
rect 41822 788700 41828 788764
rect 41892 788762 41898 788764
rect 42425 788762 42491 788765
rect 41892 788760 42491 788762
rect 41892 788704 42430 788760
rect 42486 788704 42491 788760
rect 41892 788702 42491 788704
rect 41892 788700 41898 788702
rect 42425 788699 42491 788702
rect 41454 788156 41460 788220
rect 41524 788218 41530 788220
rect 42241 788218 42307 788221
rect 41524 788216 42307 788218
rect 41524 788160 42246 788216
rect 42302 788160 42307 788216
rect 41524 788158 42307 788160
rect 41524 788156 41530 788158
rect 42241 788155 42307 788158
rect 675753 788082 675819 788085
rect 676070 788082 676076 788084
rect 675753 788080 676076 788082
rect 675753 788024 675758 788080
rect 675814 788024 676076 788080
rect 675753 788022 676076 788024
rect 675753 788019 675819 788022
rect 676070 788020 676076 788022
rect 676140 788020 676146 788084
rect 62113 787402 62179 787405
rect 64646 787402 64706 787940
rect 62113 787400 64706 787402
rect 62113 787344 62118 787400
rect 62174 787344 64706 787400
rect 62113 787342 64706 787344
rect 62113 787339 62179 787342
rect 62941 787130 63007 787133
rect 62941 787128 64706 787130
rect 62941 787072 62946 787128
rect 63002 787072 64706 787128
rect 62941 787070 64706 787072
rect 62941 787067 63007 787070
rect 64646 786758 64706 787070
rect 674414 786660 674420 786724
rect 674484 786722 674490 786724
rect 675109 786722 675175 786725
rect 675385 786724 675451 786725
rect 675334 786722 675340 786724
rect 674484 786720 675175 786722
rect 674484 786664 675114 786720
rect 675170 786664 675175 786720
rect 674484 786662 675175 786664
rect 675294 786662 675340 786722
rect 675404 786720 675451 786724
rect 675446 786664 675451 786720
rect 674484 786660 674490 786662
rect 675109 786659 675175 786662
rect 675334 786660 675340 786662
rect 675404 786660 675451 786664
rect 675385 786659 675451 786660
rect 62297 786178 62363 786181
rect 62297 786176 64706 786178
rect 62297 786120 62302 786176
rect 62358 786120 64706 786176
rect 62297 786118 64706 786120
rect 62297 786115 62363 786118
rect 64646 785576 64706 786118
rect 62113 784954 62179 784957
rect 62113 784952 64706 784954
rect 62113 784896 62118 784952
rect 62174 784896 64706 784952
rect 62113 784894 64706 784896
rect 62113 784891 62179 784894
rect 64646 784394 64706 784894
rect 674373 779378 674439 779381
rect 675477 779378 675543 779381
rect 674373 779376 675543 779378
rect 674373 779320 674378 779376
rect 674434 779320 675482 779376
rect 675538 779320 675543 779376
rect 674373 779318 675543 779320
rect 674373 779315 674439 779318
rect 675477 779315 675543 779318
rect 674557 778834 674623 778837
rect 675477 778834 675543 778837
rect 674557 778832 675543 778834
rect 649950 778426 650010 778824
rect 674557 778776 674562 778832
rect 674618 778776 675482 778832
rect 675538 778776 675543 778832
rect 674557 778774 675543 778776
rect 674557 778771 674623 778774
rect 675477 778771 675543 778774
rect 651465 778426 651531 778429
rect 649950 778424 651531 778426
rect 649950 778368 651470 778424
rect 651526 778368 651531 778424
rect 649950 778366 651531 778368
rect 651465 778363 651531 778366
rect 649950 777066 650010 777642
rect 673269 777474 673335 777477
rect 675385 777474 675451 777477
rect 673269 777472 675451 777474
rect 673269 777416 673274 777472
rect 673330 777416 675390 777472
rect 675446 777416 675451 777472
rect 673269 777414 675451 777416
rect 673269 777411 673335 777414
rect 675385 777411 675451 777414
rect 652017 777066 652083 777069
rect 649950 777064 652083 777066
rect 649950 777008 652022 777064
rect 652078 777008 652083 777064
rect 649950 777006 652083 777008
rect 652017 777003 652083 777006
rect 674925 777066 674991 777069
rect 675477 777066 675543 777069
rect 674925 777064 675543 777066
rect 674925 777008 674930 777064
rect 674986 777008 675482 777064
rect 675538 777008 675543 777064
rect 674925 777006 675543 777008
rect 674925 777003 674991 777006
rect 675477 777003 675543 777006
rect 649950 776114 650010 776460
rect 651465 776114 651531 776117
rect 649950 776112 651531 776114
rect 649950 776056 651470 776112
rect 651526 776056 651531 776112
rect 649950 776054 651531 776056
rect 651465 776051 651531 776054
rect 674925 775706 674991 775709
rect 675385 775706 675451 775709
rect 674925 775704 675451 775706
rect 674925 775648 674930 775704
rect 674986 775648 675390 775704
rect 675446 775648 675451 775704
rect 674925 775646 675451 775648
rect 674925 775643 674991 775646
rect 675385 775643 675451 775646
rect 651373 775298 651439 775301
rect 649950 775296 651439 775298
rect 649950 775240 651378 775296
rect 651434 775240 651439 775296
rect 649950 775238 651439 775240
rect 651373 775235 651439 775238
rect 35801 774754 35867 774757
rect 35758 774752 35867 774754
rect 35758 774696 35806 774752
rect 35862 774696 35867 774752
rect 35758 774691 35867 774696
rect 35758 774452 35818 774691
rect 651465 774210 651531 774213
rect 649950 774208 651531 774210
rect 649950 774152 651470 774208
rect 651526 774152 651531 774208
rect 649950 774150 651531 774152
rect 649950 774096 650010 774150
rect 651465 774147 651531 774150
rect 35206 773941 35266 774044
rect 35206 773936 35315 773941
rect 35206 773880 35254 773936
rect 35310 773880 35315 773936
rect 35206 773878 35315 773880
rect 35249 773875 35315 773878
rect 35574 773533 35634 773636
rect 35574 773528 35683 773533
rect 35574 773472 35622 773528
rect 35678 773472 35683 773528
rect 35574 773470 35683 773472
rect 35617 773467 35683 773470
rect 651465 773394 651531 773397
rect 649950 773392 651531 773394
rect 649950 773336 651470 773392
rect 651526 773336 651531 773392
rect 649950 773334 651531 773336
rect 35758 773125 35818 773228
rect 35433 773122 35499 773125
rect 35390 773120 35499 773122
rect 35390 773064 35438 773120
rect 35494 773064 35499 773120
rect 35390 773059 35499 773064
rect 35758 773120 35867 773125
rect 35758 773064 35806 773120
rect 35862 773064 35867 773120
rect 35758 773062 35867 773064
rect 35801 773059 35867 773062
rect 41505 773122 41571 773125
rect 45093 773122 45159 773125
rect 41505 773120 45159 773122
rect 41505 773064 41510 773120
rect 41566 773064 45098 773120
rect 45154 773064 45159 773120
rect 41505 773062 45159 773064
rect 41505 773059 41571 773062
rect 45093 773059 45159 773062
rect 35390 772820 35450 773059
rect 649950 772914 650010 773334
rect 651465 773331 651531 773334
rect 35574 772309 35634 772412
rect 35574 772304 35683 772309
rect 35574 772248 35622 772304
rect 35678 772248 35683 772304
rect 35574 772246 35683 772248
rect 35617 772243 35683 772246
rect 40309 772306 40375 772309
rect 43437 772306 43503 772309
rect 40309 772304 43503 772306
rect 40309 772248 40314 772304
rect 40370 772248 43442 772304
rect 43498 772248 43503 772304
rect 40309 772246 43503 772248
rect 40309 772243 40375 772246
rect 43437 772243 43503 772246
rect 35758 771901 35818 772004
rect 35758 771896 35867 771901
rect 35758 771840 35806 771896
rect 35862 771840 35867 771896
rect 35758 771838 35867 771840
rect 35801 771835 35867 771838
rect 35758 771493 35818 771596
rect 35758 771488 35867 771493
rect 35758 771432 35806 771488
rect 35862 771432 35867 771488
rect 35758 771430 35867 771432
rect 35801 771427 35867 771430
rect 39941 771490 40007 771493
rect 44265 771490 44331 771493
rect 39941 771488 44331 771490
rect 39941 771432 39946 771488
rect 40002 771432 44270 771488
rect 44326 771432 44331 771488
rect 39941 771430 44331 771432
rect 39941 771427 40007 771430
rect 44265 771427 44331 771430
rect 35390 771085 35450 771188
rect 35390 771080 35499 771085
rect 35390 771024 35438 771080
rect 35494 771024 35499 771080
rect 35390 771022 35499 771024
rect 35433 771019 35499 771022
rect 35574 770677 35634 770780
rect 35574 770672 35683 770677
rect 35574 770616 35622 770672
rect 35678 770616 35683 770672
rect 35574 770614 35683 770616
rect 35617 770611 35683 770614
rect 35758 770269 35818 770372
rect 35758 770264 35867 770269
rect 35758 770208 35806 770264
rect 35862 770208 35867 770264
rect 35758 770206 35867 770208
rect 35801 770203 35867 770206
rect 40309 770266 40375 770269
rect 43621 770266 43687 770269
rect 40309 770264 43687 770266
rect 40309 770208 40314 770264
rect 40370 770208 43626 770264
rect 43682 770208 43687 770264
rect 40309 770206 43687 770208
rect 40309 770203 40375 770206
rect 43621 770203 43687 770206
rect 41462 769858 41522 769964
rect 41638 769858 41644 769860
rect 41462 769798 41644 769858
rect 41638 769796 41644 769798
rect 41708 769796 41714 769860
rect 35574 769453 35634 769556
rect 35574 769448 35683 769453
rect 35574 769392 35622 769448
rect 35678 769392 35683 769448
rect 35574 769390 35683 769392
rect 35617 769387 35683 769390
rect 41462 769044 41522 769148
rect 41454 768980 41460 769044
rect 41524 768980 41530 769044
rect 35758 768637 35818 768740
rect 35758 768632 35867 768637
rect 35758 768576 35806 768632
rect 35862 768576 35867 768632
rect 35758 768574 35867 768576
rect 35801 768571 35867 768574
rect 35206 768229 35266 768332
rect 35157 768224 35266 768229
rect 35157 768168 35162 768224
rect 35218 768168 35266 768224
rect 35157 768166 35266 768168
rect 35157 768163 35223 768166
rect 32446 767821 32506 767924
rect 32397 767816 32506 767821
rect 32397 767760 32402 767816
rect 32458 767760 32506 767816
rect 32397 767758 32506 767760
rect 32397 767755 32463 767758
rect 35758 767413 35818 767516
rect 35758 767408 35867 767413
rect 35758 767352 35806 767408
rect 35862 767352 35867 767408
rect 35758 767350 35867 767352
rect 35801 767347 35867 767350
rect 33734 767005 33794 767108
rect 33734 767000 33843 767005
rect 33734 766944 33782 767000
rect 33838 766944 33843 767000
rect 33734 766942 33843 766944
rect 33777 766939 33843 766942
rect 35801 766594 35867 766597
rect 40542 766596 40602 766700
rect 35758 766592 35867 766594
rect 35758 766536 35806 766592
rect 35862 766536 35867 766592
rect 35758 766531 35867 766536
rect 40534 766532 40540 766596
rect 40604 766532 40610 766596
rect 35758 766292 35818 766531
rect 35574 765781 35634 765884
rect 35574 765776 35683 765781
rect 35574 765720 35622 765776
rect 35678 765720 35683 765776
rect 35574 765718 35683 765720
rect 35617 765715 35683 765718
rect 40726 765372 40786 765476
rect 40718 765308 40724 765372
rect 40788 765308 40794 765372
rect 40910 764964 40970 765068
rect 40902 764900 40908 764964
rect 40972 764900 40978 764964
rect 35758 764557 35818 764660
rect 35758 764552 35867 764557
rect 35758 764496 35806 764552
rect 35862 764496 35867 764552
rect 35758 764494 35867 764496
rect 35801 764491 35867 764494
rect 39389 764554 39455 764557
rect 44449 764554 44515 764557
rect 39389 764552 44515 764554
rect 39389 764496 39394 764552
rect 39450 764496 44454 764552
rect 44510 764496 44515 764552
rect 39389 764494 44515 764496
rect 39389 764491 39455 764494
rect 44449 764491 44515 764494
rect 35574 764149 35634 764252
rect 35574 764144 35683 764149
rect 35574 764088 35622 764144
rect 35678 764088 35683 764144
rect 35574 764086 35683 764088
rect 35617 764083 35683 764086
rect 39941 764146 40007 764149
rect 44633 764146 44699 764149
rect 39941 764144 44699 764146
rect 39941 764088 39946 764144
rect 40002 764088 44638 764144
rect 44694 764088 44699 764144
rect 39941 764086 44699 764088
rect 39941 764083 40007 764086
rect 44633 764083 44699 764086
rect 35801 763738 35867 763741
rect 35758 763736 35867 763738
rect 35758 763680 35806 763736
rect 35862 763680 35867 763736
rect 35758 763675 35867 763680
rect 35758 763436 35818 763675
rect 39941 763330 40007 763333
rect 44909 763330 44975 763333
rect 39941 763328 44975 763330
rect 39941 763272 39946 763328
rect 40002 763272 44914 763328
rect 44970 763272 44975 763328
rect 39941 763270 44975 763272
rect 39941 763267 40007 763270
rect 44909 763267 44975 763270
rect 35758 762925 35818 763028
rect 35758 762920 35867 762925
rect 35758 762864 35806 762920
rect 35862 762864 35867 762920
rect 35758 762862 35867 762864
rect 35801 762859 35867 762862
rect 39941 758298 40007 758301
rect 42609 758298 42675 758301
rect 39941 758296 42675 758298
rect 39941 758240 39946 758296
rect 40002 758240 42614 758296
rect 42670 758240 42675 758296
rect 39941 758238 42675 758240
rect 39941 758235 40007 758238
rect 42609 758235 42675 758238
rect 39665 758026 39731 758029
rect 42425 758026 42491 758029
rect 39665 758024 42491 758026
rect 39665 757968 39670 758024
rect 39726 757968 42430 758024
rect 42486 757968 42491 758024
rect 39665 757966 42491 757968
rect 39665 757963 39731 757966
rect 42425 757963 42491 757966
rect 36537 757754 36603 757757
rect 41822 757754 41828 757756
rect 36537 757752 41828 757754
rect 36537 757696 36542 757752
rect 36598 757696 41828 757752
rect 36537 757694 41828 757696
rect 36537 757691 36603 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 41781 757074 41847 757077
rect 41781 757072 41890 757074
rect 41781 757016 41786 757072
rect 41842 757016 41890 757072
rect 41781 757011 41890 757016
rect 41830 756669 41890 757011
rect 41830 756664 41939 756669
rect 41830 756608 41878 756664
rect 41934 756608 41939 756664
rect 41830 756606 41939 756608
rect 41873 756603 41939 756606
rect 40902 754836 40908 754900
rect 40972 754898 40978 754900
rect 42006 754898 42012 754900
rect 40972 754838 42012 754898
rect 40972 754836 40978 754838
rect 42006 754836 42012 754838
rect 42076 754836 42082 754900
rect 40718 754156 40724 754220
rect 40788 754218 40794 754220
rect 41873 754218 41939 754221
rect 40788 754216 41939 754218
rect 40788 754160 41878 754216
rect 41934 754160 41939 754216
rect 40788 754158 41939 754160
rect 40788 754156 40794 754158
rect 41873 754155 41939 754158
rect 42057 754082 42123 754085
rect 43897 754082 43963 754085
rect 42057 754080 43963 754082
rect 42057 754024 42062 754080
rect 42118 754024 43902 754080
rect 43958 754024 43963 754080
rect 42057 754022 43963 754024
rect 42057 754019 42123 754022
rect 43897 754019 43963 754022
rect 43437 753810 43503 753813
rect 42198 753808 43503 753810
rect 42198 753752 43442 753808
rect 43498 753752 43503 753808
rect 42198 753750 43503 753752
rect 42198 753541 42258 753750
rect 43437 753747 43503 753750
rect 42149 753536 42258 753541
rect 42149 753480 42154 753536
rect 42210 753480 42258 753536
rect 42149 753478 42258 753480
rect 42977 753538 43043 753541
rect 44449 753538 44515 753541
rect 42977 753536 44515 753538
rect 42977 753480 42982 753536
rect 43038 753480 44454 753536
rect 44510 753480 44515 753536
rect 42977 753478 44515 753480
rect 42149 753475 42215 753478
rect 42977 753475 43043 753478
rect 44449 753475 44515 753478
rect 42057 752994 42123 752997
rect 42885 752994 42951 752997
rect 42057 752992 42951 752994
rect 42057 752936 42062 752992
rect 42118 752936 42890 752992
rect 42946 752936 42951 752992
rect 42057 752934 42951 752936
rect 42057 752931 42123 752934
rect 42885 752931 42951 752934
rect 42057 751634 42123 751637
rect 45277 751634 45343 751637
rect 42057 751632 45343 751634
rect 42057 751576 42062 751632
rect 42118 751576 45282 751632
rect 45338 751576 45343 751632
rect 42057 751574 45343 751576
rect 42057 751571 42123 751574
rect 45277 751571 45343 751574
rect 42057 751226 42123 751229
rect 44633 751226 44699 751229
rect 42057 751224 44699 751226
rect 42057 751168 42062 751224
rect 42118 751168 44638 751224
rect 44694 751168 44699 751224
rect 42057 751166 44699 751168
rect 42057 751163 42123 751166
rect 44633 751163 44699 751166
rect 42057 750412 42123 750413
rect 42006 750410 42012 750412
rect 41966 750350 42012 750410
rect 42076 750408 42123 750412
rect 42118 750352 42123 750408
rect 42006 750348 42012 750350
rect 42076 750348 42123 750352
rect 42057 750347 42123 750348
rect 62941 747690 63007 747693
rect 62941 747688 64706 747690
rect 62941 747632 62946 747688
rect 63002 747632 64706 747688
rect 62941 747630 64706 747632
rect 62941 747627 63007 747630
rect 64646 747082 64706 747630
rect 40534 746676 40540 746740
rect 40604 746738 40610 746740
rect 41781 746738 41847 746741
rect 40604 746736 41847 746738
rect 40604 746680 41786 746736
rect 41842 746680 41847 746736
rect 40604 746678 41847 746680
rect 40604 746676 40610 746678
rect 41781 746675 41847 746678
rect 62113 746194 62179 746197
rect 62113 746192 64706 746194
rect 62113 746136 62118 746192
rect 62174 746136 64706 746192
rect 62113 746134 64706 746136
rect 62113 746131 62179 746134
rect 64646 745900 64706 746134
rect 41822 745724 41828 745788
rect 41892 745786 41898 745788
rect 42609 745786 42675 745789
rect 41892 745784 42675 745786
rect 41892 745728 42614 745784
rect 42670 745728 42675 745784
rect 41892 745726 42675 745728
rect 41892 745724 41898 745726
rect 42609 745723 42675 745726
rect 41638 745452 41644 745516
rect 41708 745514 41714 745516
rect 42241 745514 42307 745517
rect 41708 745512 42307 745514
rect 41708 745456 42246 745512
rect 42302 745456 42307 745512
rect 41708 745454 42307 745456
rect 41708 745452 41714 745454
rect 42241 745451 42307 745454
rect 41454 745044 41460 745108
rect 41524 745106 41530 745108
rect 42609 745106 42675 745109
rect 41524 745104 42675 745106
rect 41524 745048 42614 745104
rect 42670 745048 42675 745104
rect 41524 745046 42675 745048
rect 41524 745044 41530 745046
rect 42609 745043 42675 745046
rect 62113 744154 62179 744157
rect 64646 744154 64706 744718
rect 62113 744152 64706 744154
rect 62113 744096 62118 744152
rect 62174 744096 64706 744152
rect 62113 744094 64706 744096
rect 62113 744091 62179 744094
rect 62113 743746 62179 743749
rect 62113 743744 64706 743746
rect 62113 743688 62118 743744
rect 62174 743688 64706 743744
rect 62113 743686 64706 743688
rect 62113 743683 62179 743686
rect 64646 743536 64706 743686
rect 674230 743276 674236 743340
rect 674300 743338 674306 743340
rect 675201 743338 675267 743341
rect 674300 743336 675267 743338
rect 674300 743280 675206 743336
rect 675262 743280 675267 743336
rect 674300 743278 675267 743280
rect 674300 743276 674306 743278
rect 675201 743275 675267 743278
rect 62113 742386 62179 742389
rect 62113 742384 64706 742386
rect 62113 742328 62118 742384
rect 62174 742328 64706 742384
rect 62113 742326 64706 742328
rect 62113 742323 62179 742326
rect 63033 741842 63099 741845
rect 63033 741840 64706 741842
rect 63033 741784 63038 741840
rect 63094 741784 64706 741840
rect 63033 741782 64706 741784
rect 63033 741779 63099 741782
rect 64646 741172 64706 741782
rect 674598 738108 674604 738172
rect 674668 738170 674674 738172
rect 675201 738170 675267 738173
rect 674668 738168 675267 738170
rect 674668 738112 675206 738168
rect 675262 738112 675267 738168
rect 674668 738110 675267 738112
rect 674668 738108 674674 738110
rect 675201 738107 675267 738110
rect 669589 735722 669655 735725
rect 675477 735722 675543 735725
rect 669589 735720 675543 735722
rect 669589 735664 669594 735720
rect 669650 735664 675482 735720
rect 675538 735664 675543 735720
rect 669589 735662 675543 735664
rect 669589 735659 669655 735662
rect 675477 735659 675543 735662
rect 649950 734226 650010 734402
rect 673453 734362 673519 734365
rect 675477 734362 675543 734365
rect 673453 734360 675543 734362
rect 673453 734304 673458 734360
rect 673514 734304 675482 734360
rect 675538 734304 675543 734360
rect 673453 734302 675543 734304
rect 673453 734299 673519 734302
rect 675477 734299 675543 734302
rect 651465 734226 651531 734229
rect 649950 734224 651531 734226
rect 649950 734168 651470 734224
rect 651526 734168 651531 734224
rect 649950 734166 651531 734168
rect 651465 734163 651531 734166
rect 671245 733818 671311 733821
rect 675477 733818 675543 733821
rect 671245 733816 675543 733818
rect 671245 733760 671250 733816
rect 671306 733760 675482 733816
rect 675538 733760 675543 733816
rect 671245 733758 675543 733760
rect 671245 733755 671311 733758
rect 675477 733755 675543 733758
rect 649950 732866 650010 733220
rect 652661 732866 652727 732869
rect 649950 732864 652727 732866
rect 649950 732808 652666 732864
rect 652722 732808 652727 732864
rect 649950 732806 652727 732808
rect 652661 732803 652727 732806
rect 40401 732322 40467 732325
rect 45093 732322 45159 732325
rect 40401 732320 45159 732322
rect 40401 732264 40406 732320
rect 40462 732264 45098 732320
rect 45154 732264 45159 732320
rect 40401 732262 45159 732264
rect 40401 732259 40467 732262
rect 45093 732259 45159 732262
rect 649950 731778 650010 732038
rect 651465 731778 651531 731781
rect 649950 731776 651531 731778
rect 649950 731720 651470 731776
rect 651526 731720 651531 731776
rect 649950 731718 651531 731720
rect 651465 731715 651531 731718
rect 40033 731642 40099 731645
rect 42977 731642 43043 731645
rect 40033 731640 43043 731642
rect 40033 731584 40038 731640
rect 40094 731584 42982 731640
rect 43038 731584 43043 731640
rect 40033 731582 43043 731584
rect 40033 731579 40099 731582
rect 42977 731579 43043 731582
rect 35433 731370 35499 731373
rect 35420 731368 35499 731370
rect 35420 731312 35438 731368
rect 35494 731312 35499 731368
rect 35420 731310 35499 731312
rect 35433 731307 35499 731310
rect 41689 731098 41755 731101
rect 46197 731098 46263 731101
rect 651373 731098 651439 731101
rect 41689 731096 46263 731098
rect 41689 731040 41694 731096
rect 41750 731040 46202 731096
rect 46258 731040 46263 731096
rect 41689 731038 46263 731040
rect 41689 731035 41755 731038
rect 46197 731035 46263 731038
rect 649950 731096 651439 731098
rect 649950 731040 651378 731096
rect 651434 731040 651439 731096
rect 649950 731038 651439 731040
rect 35801 730962 35867 730965
rect 35788 730960 35867 730962
rect 35788 730904 35806 730960
rect 35862 730904 35867 730960
rect 35788 730902 35867 730904
rect 35801 730899 35867 730902
rect 649950 730856 650010 731038
rect 651373 731035 651439 731038
rect 675293 730828 675359 730829
rect 675293 730826 675340 730828
rect 675248 730824 675340 730826
rect 675248 730768 675298 730824
rect 675248 730766 675340 730768
rect 675293 730764 675340 730766
rect 675404 730764 675410 730828
rect 675293 730763 675359 730764
rect 35617 730554 35683 730557
rect 35604 730552 35683 730554
rect 35604 730496 35622 730552
rect 35678 730496 35683 730552
rect 35604 730494 35683 730496
rect 35617 730491 35683 730494
rect 35801 730146 35867 730149
rect 35788 730144 35867 730146
rect 35788 730088 35806 730144
rect 35862 730088 35867 730144
rect 35788 730086 35867 730088
rect 35801 730083 35867 730086
rect 668853 730146 668919 730149
rect 675477 730146 675543 730149
rect 668853 730144 675543 730146
rect 668853 730088 668858 730144
rect 668914 730088 675482 730144
rect 675538 730088 675543 730144
rect 668853 730086 675543 730088
rect 668853 730083 668919 730086
rect 675477 730083 675543 730086
rect 651465 729874 651531 729877
rect 649950 729872 651531 729874
rect 649950 729816 651470 729872
rect 651526 729816 651531 729872
rect 649950 729814 651531 729816
rect 35433 729738 35499 729741
rect 35420 729736 35499 729738
rect 35420 729680 35438 729736
rect 35494 729680 35499 729736
rect 35420 729678 35499 729680
rect 35433 729675 35499 729678
rect 649950 729674 650010 729814
rect 651465 729811 651531 729814
rect 674741 729874 674807 729877
rect 676806 729874 676812 729876
rect 674741 729872 676812 729874
rect 674741 729816 674746 729872
rect 674802 729816 676812 729872
rect 674741 729814 676812 729816
rect 674741 729811 674807 729814
rect 676806 729812 676812 729814
rect 676876 729812 676882 729876
rect 35617 729330 35683 729333
rect 35604 729328 35683 729330
rect 35604 729272 35622 729328
rect 35678 729272 35683 729328
rect 35604 729270 35683 729272
rect 35617 729267 35683 729270
rect 35801 728922 35867 728925
rect 35788 728920 35867 728922
rect 35788 728864 35806 728920
rect 35862 728864 35867 728920
rect 35788 728862 35867 728864
rect 35801 728859 35867 728862
rect 669405 728786 669471 728789
rect 675477 728786 675543 728789
rect 669405 728784 675543 728786
rect 669405 728728 669410 728784
rect 669466 728728 675482 728784
rect 675538 728728 675543 728784
rect 669405 728726 675543 728728
rect 669405 728723 669471 728726
rect 675477 728723 675543 728726
rect 35801 728514 35867 728517
rect 651465 728514 651531 728517
rect 35788 728512 35867 728514
rect 35788 728456 35806 728512
rect 35862 728456 35867 728512
rect 35788 728454 35867 728456
rect 649950 728512 651531 728514
rect 649950 728456 651470 728512
rect 651526 728456 651531 728512
rect 649950 728454 651531 728456
rect 35801 728451 35867 728454
rect 651465 728451 651531 728454
rect 41689 728242 41755 728245
rect 44265 728242 44331 728245
rect 41689 728240 44331 728242
rect 41689 728184 41694 728240
rect 41750 728184 44270 728240
rect 44326 728184 44331 728240
rect 41689 728182 44331 728184
rect 41689 728179 41755 728182
rect 44265 728179 44331 728182
rect 35433 728106 35499 728109
rect 35420 728104 35499 728106
rect 35420 728048 35438 728104
rect 35494 728048 35499 728104
rect 35420 728046 35499 728048
rect 35433 728043 35499 728046
rect 41689 727834 41755 727837
rect 43069 727834 43135 727837
rect 41689 727832 43135 727834
rect 41689 727776 41694 727832
rect 41750 727776 43074 727832
rect 43130 727776 43135 727832
rect 41689 727774 43135 727776
rect 41689 727771 41755 727774
rect 43069 727771 43135 727774
rect 35617 727698 35683 727701
rect 35604 727696 35683 727698
rect 35604 727640 35622 727696
rect 35678 727640 35683 727696
rect 35604 727638 35683 727640
rect 35617 727635 35683 727638
rect 35801 727290 35867 727293
rect 35788 727288 35867 727290
rect 35788 727232 35806 727288
rect 35862 727232 35867 727288
rect 35788 727230 35867 727232
rect 35801 727227 35867 727230
rect 41137 726882 41203 726885
rect 41124 726880 41203 726882
rect 41124 726824 41142 726880
rect 41198 726824 41203 726880
rect 41124 726822 41203 726824
rect 41137 726819 41203 726822
rect 676070 726548 676076 726612
rect 676140 726610 676146 726612
rect 682377 726610 682443 726613
rect 676140 726608 682443 726610
rect 676140 726552 682382 726608
rect 682438 726552 682443 726608
rect 676140 726550 682443 726552
rect 676140 726548 676146 726550
rect 682377 726547 682443 726550
rect 41321 726474 41387 726477
rect 41308 726472 41387 726474
rect 41308 726416 41326 726472
rect 41382 726416 41387 726472
rect 41308 726414 41387 726416
rect 41321 726411 41387 726414
rect 674414 726276 674420 726340
rect 674484 726338 674490 726340
rect 684217 726338 684283 726341
rect 674484 726336 684283 726338
rect 674484 726280 684222 726336
rect 684278 726280 684283 726336
rect 674484 726278 684283 726280
rect 674484 726276 674490 726278
rect 684217 726275 684283 726278
rect 41324 726066 41844 726100
rect 41308 726040 41844 726066
rect 41308 726006 41384 726040
rect 41784 725932 41844 726040
rect 41784 725870 41828 725932
rect 41822 725868 41828 725870
rect 41892 725868 41898 725932
rect 40953 725658 41019 725661
rect 40940 725656 41019 725658
rect 40940 725600 40958 725656
rect 41014 725600 41019 725656
rect 40940 725598 41019 725600
rect 40953 725595 41019 725598
rect 41781 725660 41847 725661
rect 41781 725656 41828 725660
rect 41892 725658 41898 725660
rect 41781 725600 41786 725656
rect 41781 725596 41828 725600
rect 41892 725598 41938 725658
rect 41892 725596 41898 725598
rect 41781 725595 41847 725596
rect 32397 725250 32463 725253
rect 32397 725248 32476 725250
rect 32397 725192 32402 725248
rect 32458 725192 32476 725248
rect 32397 725190 32476 725192
rect 32397 725187 32463 725190
rect 35157 724842 35223 724845
rect 35157 724840 35236 724842
rect 35157 724784 35162 724840
rect 35218 724784 35236 724840
rect 35157 724782 35236 724784
rect 35157 724779 35223 724782
rect 37273 724434 37339 724437
rect 37260 724432 37339 724434
rect 37260 724376 37278 724432
rect 37334 724376 37339 724432
rect 37260 724374 37339 724376
rect 37273 724371 37339 724374
rect 31661 724026 31727 724029
rect 31661 724024 31740 724026
rect 31661 723968 31666 724024
rect 31722 723968 31740 724024
rect 31661 723966 31740 723968
rect 31661 723963 31727 723966
rect 43805 723618 43871 723621
rect 41492 723616 43871 723618
rect 41492 723560 43810 723616
rect 43866 723560 43871 723616
rect 41492 723558 43871 723560
rect 43805 723555 43871 723558
rect 39297 723210 39363 723213
rect 39284 723208 39363 723210
rect 39284 723152 39302 723208
rect 39358 723152 39363 723208
rect 39284 723150 39363 723152
rect 39297 723147 39363 723150
rect 45093 722802 45159 722805
rect 41492 722800 45159 722802
rect 41492 722744 45098 722800
rect 45154 722744 45159 722800
rect 41492 722742 45159 722744
rect 45093 722739 45159 722742
rect 41781 722394 41847 722397
rect 41492 722392 41847 722394
rect 41492 722336 41786 722392
rect 41842 722336 41847 722392
rect 41492 722334 41847 722336
rect 41781 722331 41847 722334
rect 40726 721772 40786 721956
rect 674005 721852 674071 721853
rect 674005 721848 674052 721852
rect 674116 721850 674122 721852
rect 674005 721792 674010 721848
rect 674005 721788 674052 721792
rect 674116 721790 674162 721850
rect 674116 721788 674122 721790
rect 674005 721787 674071 721788
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 675109 721716 675175 721717
rect 675109 721714 675156 721716
rect 675064 721712 675156 721714
rect 675064 721656 675114 721712
rect 675064 721654 675156 721656
rect 675109 721652 675156 721654
rect 675220 721652 675226 721716
rect 675109 721651 675175 721652
rect 44725 721578 44791 721581
rect 41492 721576 44791 721578
rect 41492 721520 44730 721576
rect 44786 721520 44791 721576
rect 41492 721518 44791 721520
rect 44725 721515 44791 721518
rect 42885 721170 42951 721173
rect 41492 721168 42951 721170
rect 41492 721112 42890 721168
rect 42946 721112 42951 721168
rect 41492 721110 42951 721112
rect 42885 721107 42951 721110
rect 43621 720354 43687 720357
rect 41492 720352 43687 720354
rect 41492 720296 43626 720352
rect 43682 720296 43687 720352
rect 41492 720294 43687 720296
rect 43621 720291 43687 720294
rect 674005 719676 674071 719677
rect 674005 719674 674052 719676
rect 673960 719672 674052 719674
rect 673960 719616 674010 719672
rect 673960 719614 674052 719616
rect 674005 719612 674052 719614
rect 674116 719612 674122 719676
rect 674005 719611 674071 719612
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41781 718586 41847 718589
rect 40604 718584 41847 718586
rect 40604 718528 41786 718584
rect 41842 718528 41847 718584
rect 40604 718526 41847 718528
rect 40604 718524 40610 718526
rect 41781 718523 41847 718526
rect 37273 716954 37339 716957
rect 41822 716954 41828 716956
rect 37273 716952 41828 716954
rect 37273 716896 37278 716952
rect 37334 716896 41828 716952
rect 37273 716894 41828 716896
rect 37273 716891 37339 716894
rect 41822 716892 41828 716894
rect 41892 716892 41898 716956
rect 673269 716546 673335 716549
rect 673269 716544 676292 716546
rect 673269 716488 673274 716544
rect 673330 716488 676292 716544
rect 673269 716486 676292 716488
rect 673269 716483 673335 716486
rect 673269 716138 673335 716141
rect 673269 716136 676292 716138
rect 673269 716080 673274 716136
rect 673330 716080 676292 716136
rect 673269 716078 676292 716080
rect 673269 716075 673335 716078
rect 40585 715866 40651 715869
rect 42425 715866 42491 715869
rect 40585 715864 42491 715866
rect 40585 715808 40590 715864
rect 40646 715808 42430 715864
rect 42486 715808 42491 715864
rect 40585 715806 42491 715808
rect 40585 715803 40651 715806
rect 42425 715803 42491 715806
rect 673085 715730 673151 715733
rect 673085 715728 676292 715730
rect 673085 715672 673090 715728
rect 673146 715672 676292 715728
rect 673085 715670 676292 715672
rect 673085 715667 673151 715670
rect 673085 715322 673151 715325
rect 673085 715320 676292 715322
rect 673085 715264 673090 715320
rect 673146 715264 676292 715320
rect 673085 715262 676292 715264
rect 673085 715259 673151 715262
rect 673085 715050 673151 715053
rect 673085 715048 676230 715050
rect 673085 714992 673090 715048
rect 673146 714992 676230 715048
rect 673085 714990 676230 714992
rect 673085 714987 673151 714990
rect 40953 714914 41019 714917
rect 42333 714914 42399 714917
rect 40953 714912 42399 714914
rect 40953 714856 40958 714912
rect 41014 714856 42338 714912
rect 42394 714856 42399 714912
rect 40953 714854 42399 714856
rect 676170 714914 676230 714990
rect 676170 714854 676292 714914
rect 40953 714851 41019 714854
rect 42333 714851 42399 714854
rect 673269 714506 673335 714509
rect 673269 714504 676292 714506
rect 673269 714448 673274 714504
rect 673330 714448 676292 714504
rect 673269 714446 676292 714448
rect 673269 714443 673335 714446
rect 42241 714372 42307 714373
rect 42190 714308 42196 714372
rect 42260 714370 42307 714372
rect 42260 714368 42352 714370
rect 42302 714312 42352 714368
rect 42260 714310 42352 714312
rect 42260 714308 42307 714310
rect 42241 714307 42307 714308
rect 39297 714234 39363 714237
rect 40350 714234 40356 714236
rect 39297 714232 40356 714234
rect 39297 714176 39302 714232
rect 39358 714176 40356 714232
rect 39297 714174 40356 714176
rect 39297 714171 39363 714174
rect 40350 714172 40356 714174
rect 40420 714172 40426 714236
rect 673269 714098 673335 714101
rect 673269 714096 676292 714098
rect 673269 714040 673274 714096
rect 673330 714040 676292 714096
rect 673269 714038 676292 714040
rect 673269 714035 673335 714038
rect 672533 713690 672599 713693
rect 672533 713688 676292 713690
rect 672533 713632 672538 713688
rect 672594 713632 676292 713688
rect 672533 713630 676292 713632
rect 672533 713627 672599 713630
rect 671981 713282 672047 713285
rect 671981 713280 676292 713282
rect 671981 713224 671986 713280
rect 672042 713224 676292 713280
rect 671981 713222 676292 713224
rect 671981 713219 672047 713222
rect 673269 712874 673335 712877
rect 673269 712872 676292 712874
rect 673269 712816 673274 712872
rect 673330 712816 676292 712872
rect 673269 712814 676292 712816
rect 673269 712811 673335 712814
rect 671981 712466 672047 712469
rect 671981 712464 676292 712466
rect 671981 712408 671986 712464
rect 672042 712408 676292 712464
rect 671981 712406 676292 712408
rect 671981 712403 672047 712406
rect 675293 712058 675359 712061
rect 675293 712056 676292 712058
rect 675293 712000 675298 712056
rect 675354 712000 676292 712056
rect 675293 711998 676292 712000
rect 675293 711995 675359 711998
rect 673269 711650 673335 711653
rect 673269 711648 676292 711650
rect 673269 711592 673274 711648
rect 673330 711592 676292 711648
rect 673269 711590 676292 711592
rect 673269 711587 673335 711590
rect 682377 711242 682443 711245
rect 682364 711240 682443 711242
rect 682364 711184 682382 711240
rect 682438 711184 682443 711240
rect 682364 711182 682443 711184
rect 682377 711179 682443 711182
rect 42149 710834 42215 710837
rect 43621 710834 43687 710837
rect 42149 710832 43687 710834
rect 42149 710776 42154 710832
rect 42210 710776 43626 710832
rect 43682 710776 43687 710832
rect 42149 710774 43687 710776
rect 42149 710771 42215 710774
rect 43621 710771 43687 710774
rect 680997 710834 681063 710837
rect 680997 710832 681076 710834
rect 680997 710776 681002 710832
rect 681058 710776 681076 710832
rect 680997 710774 681076 710776
rect 680997 710771 681063 710774
rect 673269 710426 673335 710429
rect 673269 710424 676292 710426
rect 673269 710368 673274 710424
rect 673330 710368 676292 710424
rect 673269 710366 676292 710368
rect 673269 710363 673335 710366
rect 673085 710018 673151 710021
rect 673085 710016 676292 710018
rect 673085 709960 673090 710016
rect 673146 709960 676292 710016
rect 673085 709958 676292 709960
rect 673085 709955 673151 709958
rect 40350 709820 40356 709884
rect 40420 709882 40426 709884
rect 41781 709882 41847 709885
rect 40420 709880 41847 709882
rect 40420 709824 41786 709880
rect 41842 709824 41847 709880
rect 40420 709822 41847 709824
rect 40420 709820 40426 709822
rect 41781 709819 41847 709822
rect 684217 709610 684283 709613
rect 684204 709608 684283 709610
rect 684204 709552 684222 709608
rect 684278 709552 684283 709608
rect 684204 709550 684283 709552
rect 684217 709547 684283 709550
rect 673269 709202 673335 709205
rect 673269 709200 676292 709202
rect 673269 709144 673274 709200
rect 673330 709144 676292 709200
rect 673269 709142 676292 709144
rect 673269 709139 673335 709142
rect 673269 708794 673335 708797
rect 673269 708792 676292 708794
rect 673269 708736 673274 708792
rect 673330 708736 676292 708792
rect 673269 708734 676292 708736
rect 673269 708731 673335 708734
rect 42057 708522 42123 708525
rect 44725 708522 44791 708525
rect 42057 708520 44791 708522
rect 42057 708464 42062 708520
rect 42118 708464 44730 708520
rect 44786 708464 44791 708520
rect 42057 708462 44791 708464
rect 42057 708459 42123 708462
rect 44725 708459 44791 708462
rect 672809 708386 672875 708389
rect 672809 708384 676292 708386
rect 672809 708328 672814 708384
rect 672870 708328 676292 708384
rect 672809 708326 676292 708328
rect 672809 708323 672875 708326
rect 684033 707978 684099 707981
rect 684020 707976 684099 707978
rect 684020 707920 684038 707976
rect 684094 707920 684099 707976
rect 684020 707918 684099 707920
rect 684033 707915 684099 707918
rect 673729 707570 673795 707573
rect 673729 707568 676292 707570
rect 673729 707512 673734 707568
rect 673790 707512 676292 707568
rect 673729 707510 676292 707512
rect 673729 707507 673795 707510
rect 40718 707100 40724 707164
rect 40788 707162 40794 707164
rect 41781 707162 41847 707165
rect 40788 707160 41847 707162
rect 40788 707104 41786 707160
rect 41842 707104 41847 707160
rect 40788 707102 41847 707104
rect 40788 707100 40794 707102
rect 41781 707099 41847 707102
rect 676029 707162 676095 707165
rect 676029 707160 676292 707162
rect 676029 707104 676034 707160
rect 676090 707104 676292 707160
rect 676029 707102 676292 707104
rect 676029 707099 676095 707102
rect 683389 706754 683455 706757
rect 683389 706752 683468 706754
rect 683389 706696 683394 706752
rect 683450 706696 683468 706752
rect 683389 706694 683468 706696
rect 683389 706691 683455 706694
rect 42190 706284 42196 706348
rect 42260 706346 42266 706348
rect 42425 706346 42491 706349
rect 42260 706344 42491 706346
rect 42260 706288 42430 706344
rect 42486 706288 42491 706344
rect 42260 706286 42491 706288
rect 42260 706284 42266 706286
rect 42425 706283 42491 706286
rect 673729 706346 673795 706349
rect 673729 706344 676292 706346
rect 673729 706288 673734 706344
rect 673790 706288 676292 706344
rect 673729 706286 676292 706288
rect 673729 706283 673795 706286
rect 677182 705530 677242 705908
rect 683113 705530 683179 705533
rect 677182 705528 683179 705530
rect 677182 705500 683118 705528
rect 677212 705472 683118 705500
rect 683174 705472 683179 705528
rect 677212 705470 683179 705472
rect 683113 705467 683179 705470
rect 673269 705394 673335 705397
rect 674281 705394 674347 705397
rect 673269 705392 674347 705394
rect 673269 705336 673274 705392
rect 673330 705336 674286 705392
rect 674342 705336 674347 705392
rect 673269 705334 674347 705336
rect 673269 705331 673335 705334
rect 674281 705331 674347 705334
rect 673729 705122 673795 705125
rect 673729 705120 676292 705122
rect 673729 705064 673734 705120
rect 673790 705064 676292 705120
rect 673729 705062 676292 705064
rect 673729 705059 673795 705062
rect 62113 704442 62179 704445
rect 62113 704440 64706 704442
rect 62113 704384 62118 704440
rect 62174 704384 64706 704440
rect 62113 704382 64706 704384
rect 62113 704379 62179 704382
rect 40534 704244 40540 704308
rect 40604 704306 40610 704308
rect 41781 704306 41847 704309
rect 40604 704304 41847 704306
rect 40604 704248 41786 704304
rect 41842 704248 41847 704304
rect 40604 704246 41847 704248
rect 40604 704244 40610 704246
rect 41781 704243 41847 704246
rect 64646 703860 64706 704382
rect 62113 703354 62179 703357
rect 62113 703352 64706 703354
rect 62113 703296 62118 703352
rect 62174 703296 64706 703352
rect 62113 703294 64706 703296
rect 62113 703291 62179 703294
rect 42057 703082 42123 703085
rect 42609 703082 42675 703085
rect 42057 703080 42675 703082
rect 42057 703024 42062 703080
rect 42118 703024 42614 703080
rect 42670 703024 42675 703080
rect 42057 703022 42675 703024
rect 42057 703019 42123 703022
rect 42609 703019 42675 703022
rect 64646 702678 64706 703294
rect 41822 701796 41828 701860
rect 41892 701858 41898 701860
rect 42517 701858 42583 701861
rect 41892 701856 42583 701858
rect 41892 701800 42522 701856
rect 42578 701800 42583 701856
rect 41892 701798 42583 701800
rect 41892 701796 41898 701798
rect 42517 701795 42583 701798
rect 41454 701524 41460 701588
rect 41524 701586 41530 701588
rect 42517 701586 42583 701589
rect 41524 701584 42583 701586
rect 41524 701528 42522 701584
rect 42578 701528 42583 701584
rect 41524 701526 42583 701528
rect 41524 701524 41530 701526
rect 42517 701523 42583 701526
rect 62941 701314 63007 701317
rect 64646 701314 64706 701496
rect 62941 701312 64706 701314
rect 62941 701256 62946 701312
rect 63002 701256 64706 701312
rect 62941 701254 64706 701256
rect 62941 701251 63007 701254
rect 673729 701178 673795 701181
rect 675109 701178 675175 701181
rect 673729 701176 675175 701178
rect 673729 701120 673734 701176
rect 673790 701120 675114 701176
rect 675170 701120 675175 701176
rect 673729 701118 675175 701120
rect 673729 701115 673795 701118
rect 675109 701115 675175 701118
rect 63125 700906 63191 700909
rect 63125 700904 64706 700906
rect 63125 700848 63130 700904
rect 63186 700848 64706 700904
rect 63125 700846 64706 700848
rect 63125 700843 63191 700846
rect 41873 700500 41939 700501
rect 41822 700498 41828 700500
rect 41782 700438 41828 700498
rect 41892 700496 41939 700500
rect 41934 700440 41939 700496
rect 41822 700436 41828 700438
rect 41892 700436 41939 700440
rect 41873 700435 41939 700436
rect 64646 700314 64706 700846
rect 61377 699682 61443 699685
rect 61377 699680 64706 699682
rect 61377 699624 61382 699680
rect 61438 699624 64706 699680
rect 61377 699622 64706 699624
rect 61377 699619 61443 699622
rect 64646 699132 64706 699622
rect 667657 698322 667723 698325
rect 675109 698322 675175 698325
rect 667657 698320 675175 698322
rect 667657 698264 667662 698320
rect 667718 698264 675114 698320
rect 675170 698264 675175 698320
rect 667657 698262 675175 698264
rect 667657 698259 667723 698262
rect 675109 698259 675175 698262
rect 62205 698050 62271 698053
rect 62205 698048 64706 698050
rect 62205 697992 62210 698048
rect 62266 697992 64706 698048
rect 62205 697990 64706 697992
rect 62205 697987 62271 697990
rect 64646 697950 64706 697990
rect 673269 696962 673335 696965
rect 675109 696962 675175 696965
rect 673269 696960 675175 696962
rect 673269 696904 673274 696960
rect 673330 696904 675114 696960
rect 675170 696904 675175 696960
rect 673269 696902 675175 696904
rect 673269 696899 673335 696902
rect 675109 696899 675175 696902
rect 675477 696828 675543 696829
rect 675477 696824 675524 696828
rect 675588 696826 675594 696828
rect 675477 696768 675482 696824
rect 675477 696764 675524 696768
rect 675588 696766 675634 696826
rect 675588 696764 675594 696766
rect 675477 696763 675543 696764
rect 670877 695874 670943 695877
rect 675109 695874 675175 695877
rect 670877 695872 675175 695874
rect 670877 695816 670882 695872
rect 670938 695816 675114 695872
rect 675170 695816 675175 695872
rect 670877 695814 675175 695816
rect 670877 695811 670943 695814
rect 675109 695811 675175 695814
rect 674414 694588 674420 694652
rect 674484 694650 674490 694652
rect 675109 694650 675175 694653
rect 674484 694648 675175 694650
rect 674484 694592 675114 694648
rect 675170 694592 675175 694648
rect 674484 694590 675175 694592
rect 674484 694588 674490 694590
rect 675109 694587 675175 694590
rect 673729 692882 673795 692885
rect 675109 692882 675175 692885
rect 673729 692880 675175 692882
rect 673729 692824 673734 692880
rect 673790 692824 675114 692880
rect 675170 692824 675175 692880
rect 673729 692822 675175 692824
rect 673729 692819 673795 692822
rect 675109 692819 675175 692822
rect 673729 690162 673795 690165
rect 674925 690162 674991 690165
rect 673729 690160 674991 690162
rect 673729 690104 673734 690160
rect 673790 690104 674930 690160
rect 674986 690104 674991 690160
rect 673729 690102 674991 690104
rect 673729 690099 673795 690102
rect 674925 690099 674991 690102
rect 649950 689482 650010 689980
rect 674097 689890 674163 689893
rect 675109 689890 675175 689893
rect 674097 689888 675175 689890
rect 674097 689832 674102 689888
rect 674158 689832 675114 689888
rect 675170 689832 675175 689888
rect 674097 689830 675175 689832
rect 674097 689827 674163 689830
rect 675109 689827 675175 689830
rect 651465 689482 651531 689485
rect 649950 689480 651531 689482
rect 649950 689424 651470 689480
rect 651526 689424 651531 689480
rect 649950 689422 651531 689424
rect 651465 689419 651531 689422
rect 669037 689482 669103 689485
rect 675109 689482 675175 689485
rect 669037 689480 675175 689482
rect 669037 689424 669042 689480
rect 669098 689424 675114 689480
rect 675170 689424 675175 689480
rect 669037 689422 675175 689424
rect 669037 689419 669103 689422
rect 675109 689419 675175 689422
rect 649980 688802 650562 688828
rect 651649 688802 651715 688805
rect 649980 688800 651715 688802
rect 649980 688768 651654 688800
rect 650502 688744 651654 688768
rect 651710 688744 651715 688800
rect 650502 688742 651715 688744
rect 651649 688739 651715 688742
rect 673729 688802 673795 688805
rect 674925 688802 674991 688805
rect 673729 688800 674991 688802
rect 673729 688744 673734 688800
rect 673790 688744 674930 688800
rect 674986 688744 674991 688800
rect 673729 688742 674991 688744
rect 673729 688739 673795 688742
rect 674925 688739 674991 688742
rect 35433 688394 35499 688397
rect 35390 688392 35499 688394
rect 35390 688336 35438 688392
rect 35494 688336 35499 688392
rect 35390 688331 35499 688336
rect 35390 688092 35450 688331
rect 673729 688122 673795 688125
rect 674281 688122 674347 688125
rect 673729 688120 674347 688122
rect 673729 688064 673734 688120
rect 673790 688064 674286 688120
rect 674342 688064 674347 688120
rect 673729 688062 674347 688064
rect 673729 688059 673795 688062
rect 674281 688059 674347 688062
rect 668209 687850 668275 687853
rect 675109 687850 675175 687853
rect 668209 687848 675175 687850
rect 668209 687792 668214 687848
rect 668270 687792 675114 687848
rect 675170 687792 675175 687848
rect 668209 687790 675175 687792
rect 668209 687787 668275 687790
rect 675109 687787 675175 687790
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 41689 687578 41755 687581
rect 45461 687578 45527 687581
rect 41689 687576 45527 687578
rect 41689 687520 41694 687576
rect 41750 687520 45466 687576
rect 45522 687520 45527 687576
rect 41689 687518 45527 687520
rect 41689 687515 41755 687518
rect 45461 687515 45527 687518
rect 649950 687442 650010 687616
rect 651465 687442 651531 687445
rect 649950 687440 651531 687442
rect 649950 687384 651470 687440
rect 651526 687384 651531 687440
rect 649950 687382 651531 687384
rect 651465 687379 651531 687382
rect 35617 687306 35683 687309
rect 35604 687304 35683 687306
rect 35604 687248 35622 687304
rect 35678 687248 35683 687304
rect 35604 687246 35683 687248
rect 35617 687243 35683 687246
rect 41689 687170 41755 687173
rect 46197 687170 46263 687173
rect 41689 687168 46263 687170
rect 41689 687112 41694 687168
rect 41750 687112 46202 687168
rect 46258 687112 46263 687168
rect 41689 687110 46263 687112
rect 41689 687107 41755 687110
rect 46197 687107 46263 687110
rect 35433 686898 35499 686901
rect 35420 686896 35499 686898
rect 35420 686840 35438 686896
rect 35494 686840 35499 686896
rect 35420 686838 35499 686840
rect 35433 686835 35499 686838
rect 651465 686762 651531 686765
rect 649950 686760 651531 686762
rect 649950 686704 651470 686760
rect 651526 686704 651531 686760
rect 649950 686702 651531 686704
rect 35801 686490 35867 686493
rect 35788 686488 35867 686490
rect 35788 686432 35806 686488
rect 35862 686432 35867 686488
rect 649950 686434 650010 686702
rect 651465 686699 651531 686702
rect 35788 686430 35867 686432
rect 35801 686427 35867 686430
rect 673085 686218 673151 686221
rect 675109 686218 675175 686221
rect 673085 686216 675175 686218
rect 673085 686160 673090 686216
rect 673146 686160 675114 686216
rect 675170 686160 675175 686216
rect 673085 686158 675175 686160
rect 673085 686155 673151 686158
rect 675109 686155 675175 686158
rect 35801 686082 35867 686085
rect 35788 686080 35867 686082
rect 35788 686024 35806 686080
rect 35862 686024 35867 686080
rect 35788 686022 35867 686024
rect 35801 686019 35867 686022
rect 669773 685810 669839 685813
rect 674925 685810 674991 685813
rect 669773 685808 674991 685810
rect 669773 685752 669778 685808
rect 669834 685752 674930 685808
rect 674986 685752 674991 685808
rect 669773 685750 674991 685752
rect 669773 685747 669839 685750
rect 674925 685747 674991 685750
rect 35801 685674 35867 685677
rect 35788 685672 35867 685674
rect 35788 685616 35806 685672
rect 35862 685616 35867 685672
rect 35788 685614 35867 685616
rect 35801 685611 35867 685614
rect 670601 685538 670667 685541
rect 675109 685538 675175 685541
rect 670601 685536 675175 685538
rect 670601 685480 670606 685536
rect 670662 685480 675114 685536
rect 675170 685480 675175 685536
rect 670601 685478 675175 685480
rect 670601 685475 670667 685478
rect 675109 685475 675175 685478
rect 35617 685266 35683 685269
rect 651465 685266 651531 685269
rect 35604 685264 35683 685266
rect 35604 685208 35622 685264
rect 35678 685208 35683 685264
rect 35604 685206 35683 685208
rect 649950 685264 651531 685266
rect 649950 685208 651470 685264
rect 651526 685208 651531 685264
rect 649950 685206 651531 685208
rect 35617 685203 35683 685206
rect 651465 685203 651531 685206
rect 35801 684858 35867 684861
rect 35788 684856 35867 684858
rect 35788 684800 35806 684856
rect 35862 684800 35867 684856
rect 35788 684798 35867 684800
rect 35801 684795 35867 684798
rect 41689 684722 41755 684725
rect 43069 684722 43135 684725
rect 41689 684720 43135 684722
rect 41689 684664 41694 684720
rect 41750 684664 43074 684720
rect 43130 684664 43135 684720
rect 41689 684662 43135 684664
rect 41689 684659 41755 684662
rect 43069 684659 43135 684662
rect 35617 684450 35683 684453
rect 652569 684450 652635 684453
rect 35604 684448 35683 684450
rect 35604 684392 35622 684448
rect 35678 684392 35683 684448
rect 35604 684390 35683 684392
rect 35617 684387 35683 684390
rect 649950 684448 652635 684450
rect 649950 684392 652574 684448
rect 652630 684392 652635 684448
rect 649950 684390 652635 684392
rect 649950 684070 650010 684390
rect 652569 684387 652635 684390
rect 35433 684042 35499 684045
rect 35420 684040 35499 684042
rect 35420 683984 35438 684040
rect 35494 683984 35499 684040
rect 35420 683982 35499 683984
rect 35433 683979 35499 683982
rect 675109 684042 675175 684045
rect 675518 684042 675524 684044
rect 675109 684040 675524 684042
rect 675109 683984 675114 684040
rect 675170 683984 675524 684040
rect 675109 683982 675524 683984
rect 675109 683979 675175 683982
rect 675518 683980 675524 683982
rect 675588 683980 675594 684044
rect 41689 683906 41755 683909
rect 43437 683906 43503 683909
rect 41689 683904 43503 683906
rect 41689 683848 41694 683904
rect 41750 683848 43442 683904
rect 43498 683848 43503 683904
rect 41689 683846 43503 683848
rect 41689 683843 41755 683846
rect 43437 683843 43503 683846
rect 675293 683772 675359 683773
rect 675293 683770 675340 683772
rect 675248 683768 675340 683770
rect 675248 683712 675298 683768
rect 675248 683710 675340 683712
rect 675293 683708 675340 683710
rect 675404 683708 675410 683772
rect 675293 683707 675359 683708
rect 42006 683634 42012 683636
rect 41492 683574 42012 683634
rect 42006 683572 42012 683574
rect 42076 683572 42082 683636
rect 35801 683226 35867 683229
rect 35788 683224 35867 683226
rect 35788 683168 35806 683224
rect 35862 683168 35867 683224
rect 35788 683166 35867 683168
rect 35801 683163 35867 683166
rect 41689 683090 41755 683093
rect 45093 683090 45159 683093
rect 41689 683088 45159 683090
rect 41689 683032 41694 683088
rect 41750 683032 45098 683088
rect 45154 683032 45159 683088
rect 41689 683030 45159 683032
rect 41689 683027 41755 683030
rect 45093 683027 45159 683030
rect 35617 682818 35683 682821
rect 35604 682816 35683 682818
rect 35604 682760 35622 682816
rect 35678 682760 35683 682816
rect 35604 682758 35683 682760
rect 35617 682755 35683 682758
rect 674230 682620 674236 682684
rect 674300 682682 674306 682684
rect 684125 682682 684191 682685
rect 674300 682680 684191 682682
rect 674300 682624 684130 682680
rect 684186 682624 684191 682680
rect 674300 682622 684191 682624
rect 674300 682620 674306 682622
rect 684125 682619 684191 682622
rect 35801 682410 35867 682413
rect 35788 682408 35867 682410
rect 35788 682352 35806 682408
rect 35862 682352 35867 682408
rect 35788 682350 35867 682352
rect 35801 682347 35867 682350
rect 673453 682410 673519 682413
rect 674833 682410 674899 682413
rect 673453 682408 674899 682410
rect 673453 682352 673458 682408
rect 673514 682352 674838 682408
rect 674894 682352 674899 682408
rect 673453 682350 674899 682352
rect 673453 682347 673519 682350
rect 674833 682347 674899 682350
rect 35157 682002 35223 682005
rect 673545 682002 673611 682005
rect 675477 682002 675543 682005
rect 35157 682000 35236 682002
rect 35157 681944 35162 682000
rect 35218 681944 35236 682000
rect 35157 681942 35236 681944
rect 673545 682000 675543 682002
rect 673545 681944 673550 682000
rect 673606 681944 675482 682000
rect 675538 681944 675543 682000
rect 673545 681942 675543 681944
rect 35157 681939 35223 681942
rect 673545 681939 673611 681942
rect 675477 681939 675543 681942
rect 33041 681594 33107 681597
rect 33028 681592 33107 681594
rect 33028 681536 33046 681592
rect 33102 681536 33107 681592
rect 33028 681534 33107 681536
rect 33041 681531 33107 681534
rect 41689 681458 41755 681461
rect 42190 681458 42196 681460
rect 41689 681456 42196 681458
rect 41689 681400 41694 681456
rect 41750 681400 42196 681456
rect 41689 681398 42196 681400
rect 41689 681395 41755 681398
rect 42190 681396 42196 681398
rect 42260 681396 42266 681460
rect 33777 681186 33843 681189
rect 33764 681184 33843 681186
rect 33764 681128 33782 681184
rect 33838 681128 33843 681184
rect 33764 681126 33843 681128
rect 33777 681123 33843 681126
rect 41689 681050 41755 681053
rect 42701 681050 42767 681053
rect 41689 681048 42767 681050
rect 41689 680992 41694 681048
rect 41750 680992 42706 681048
rect 42762 680992 42767 681048
rect 41689 680990 42767 680992
rect 41689 680987 41755 680990
rect 42701 680987 42767 680990
rect 31017 680778 31083 680781
rect 31004 680776 31083 680778
rect 31004 680720 31022 680776
rect 31078 680720 31083 680776
rect 31004 680718 31083 680720
rect 31017 680715 31083 680718
rect 35801 680370 35867 680373
rect 35788 680368 35867 680370
rect 35788 680312 35806 680368
rect 35862 680312 35867 680368
rect 35788 680310 35867 680312
rect 35801 680307 35867 680310
rect 41689 680234 41755 680237
rect 44449 680234 44515 680237
rect 41689 680232 44515 680234
rect 41689 680176 41694 680232
rect 41750 680176 44454 680232
rect 44510 680176 44515 680232
rect 41689 680174 44515 680176
rect 41689 680171 41755 680174
rect 44449 680171 44515 680174
rect 35801 679962 35867 679965
rect 35788 679960 35867 679962
rect 35788 679904 35806 679960
rect 35862 679904 35867 679960
rect 35788 679902 35867 679904
rect 35801 679899 35867 679902
rect 35617 679554 35683 679557
rect 35604 679552 35683 679554
rect 35604 679496 35622 679552
rect 35678 679496 35683 679552
rect 35604 679494 35683 679496
rect 35617 679491 35683 679494
rect 41689 679418 41755 679421
rect 44265 679418 44331 679421
rect 41689 679416 44331 679418
rect 41689 679360 41694 679416
rect 41750 679360 44270 679416
rect 44326 679360 44331 679416
rect 41689 679358 44331 679360
rect 41689 679355 41755 679358
rect 44265 679355 44331 679358
rect 35801 679146 35867 679149
rect 35788 679144 35867 679146
rect 35788 679088 35806 679144
rect 35862 679088 35867 679144
rect 35788 679086 35867 679088
rect 35801 679083 35867 679086
rect 41689 679010 41755 679013
rect 44725 679010 44791 679013
rect 41689 679008 44791 679010
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 41689 678952 41694 679008
rect 41750 678952 44730 679008
rect 44786 678952 44791 679008
rect 41689 678950 44791 678952
rect 41689 678947 41755 678950
rect 44725 678947 44791 678950
rect 40542 678708 40602 678928
rect 41689 678602 41755 678605
rect 43805 678602 43871 678605
rect 41689 678600 43871 678602
rect 41689 678544 41694 678600
rect 41750 678544 43810 678600
rect 43866 678544 43871 678600
rect 41689 678542 43871 678544
rect 41689 678539 41755 678542
rect 43805 678539 43871 678542
rect 41822 678330 41828 678332
rect 41492 678270 41828 678330
rect 41822 678268 41828 678270
rect 41892 678268 41898 678332
rect 43437 677922 43503 677925
rect 41492 677920 43503 677922
rect 41492 677864 43442 677920
rect 43498 677864 43503 677920
rect 41492 677862 43503 677864
rect 43437 677859 43503 677862
rect 43989 677106 44055 677109
rect 41492 677104 44055 677106
rect 41492 677048 43994 677104
rect 44050 677048 44055 677104
rect 41492 677046 44055 677048
rect 43989 677043 44055 677046
rect 675109 676426 675175 676429
rect 676070 676426 676076 676428
rect 675109 676424 676076 676426
rect 675109 676368 675114 676424
rect 675170 676368 676076 676424
rect 675109 676366 676076 676368
rect 675109 676363 675175 676366
rect 676070 676364 676076 676366
rect 676140 676364 676146 676428
rect 33777 672754 33843 672757
rect 41822 672754 41828 672756
rect 33777 672752 41828 672754
rect 33777 672696 33782 672752
rect 33838 672696 41828 672752
rect 33777 672694 41828 672696
rect 33777 672691 33843 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 42241 672620 42307 672621
rect 42190 672618 42196 672620
rect 42150 672558 42196 672618
rect 42260 672616 42307 672620
rect 42302 672560 42307 672616
rect 42190 672556 42196 672558
rect 42260 672556 42307 672560
rect 42241 672555 42307 672556
rect 673545 671394 673611 671397
rect 673545 671392 676292 671394
rect 673545 671336 673550 671392
rect 673606 671336 676292 671392
rect 673545 671334 676292 671336
rect 673545 671331 673611 671334
rect 673545 670986 673611 670989
rect 673545 670984 676292 670986
rect 673545 670928 673550 670984
rect 673606 670928 676292 670984
rect 673545 670926 676292 670928
rect 673545 670923 673611 670926
rect 673545 670578 673611 670581
rect 673545 670576 676292 670578
rect 673545 670520 673550 670576
rect 673606 670520 676292 670576
rect 673545 670518 676292 670520
rect 673545 670515 673611 670518
rect 672441 670034 672507 670037
rect 676262 670034 676322 670140
rect 672441 670032 676322 670034
rect 672441 669976 672446 670032
rect 672502 669976 676322 670032
rect 672441 669974 676322 669976
rect 672441 669971 672507 669974
rect 673545 669762 673611 669765
rect 673545 669760 676292 669762
rect 673545 669704 673550 669760
rect 673606 669704 676292 669760
rect 673545 669702 676292 669704
rect 673545 669699 673611 669702
rect 672625 669490 672691 669493
rect 672625 669488 676322 669490
rect 672625 669432 672630 669488
rect 672686 669432 676322 669488
rect 672625 669430 676322 669432
rect 672625 669427 672691 669430
rect 676262 669324 676322 669430
rect 673545 668946 673611 668949
rect 673545 668944 676292 668946
rect 673545 668888 673550 668944
rect 673606 668888 676292 668944
rect 673545 668886 676292 668888
rect 673545 668883 673611 668886
rect 41965 668538 42031 668541
rect 42190 668538 42196 668540
rect 41965 668536 42196 668538
rect 41965 668480 41970 668536
rect 42026 668480 42196 668536
rect 41965 668478 42196 668480
rect 41965 668475 42031 668478
rect 42190 668476 42196 668478
rect 42260 668476 42266 668540
rect 673545 668538 673611 668541
rect 673545 668536 676292 668538
rect 673545 668480 673550 668536
rect 673606 668480 676292 668536
rect 673545 668478 676292 668480
rect 673545 668475 673611 668478
rect 673545 668130 673611 668133
rect 673545 668128 676292 668130
rect 673545 668072 673550 668128
rect 673606 668072 676292 668128
rect 673545 668070 676292 668072
rect 673545 668067 673611 668070
rect 42057 667722 42123 667725
rect 44081 667722 44147 667725
rect 42057 667720 44147 667722
rect 42057 667664 42062 667720
rect 42118 667664 44086 667720
rect 44142 667664 44147 667720
rect 42057 667662 44147 667664
rect 42057 667659 42123 667662
rect 44081 667659 44147 667662
rect 673545 667722 673611 667725
rect 673545 667720 676292 667722
rect 673545 667664 673550 667720
rect 673606 667664 676292 667720
rect 673545 667662 676292 667664
rect 673545 667659 673611 667662
rect 676029 667314 676095 667317
rect 676029 667312 676292 667314
rect 676029 667256 676034 667312
rect 676090 667256 676292 667312
rect 676029 667254 676292 667256
rect 676029 667251 676095 667254
rect 42057 667178 42123 667181
rect 44725 667178 44791 667181
rect 42057 667176 44791 667178
rect 42057 667120 42062 667176
rect 42118 667120 44730 667176
rect 44786 667120 44791 667176
rect 42057 667118 44791 667120
rect 42057 667115 42123 667118
rect 44725 667115 44791 667118
rect 673545 666906 673611 666909
rect 673545 666904 676292 666906
rect 673545 666848 673550 666904
rect 673606 666848 676292 666904
rect 673545 666846 676292 666848
rect 673545 666843 673611 666846
rect 42057 666634 42123 666637
rect 44265 666634 44331 666637
rect 42057 666632 44331 666634
rect 42057 666576 42062 666632
rect 42118 666576 44270 666632
rect 44326 666576 44331 666632
rect 42057 666574 44331 666576
rect 42057 666571 42123 666574
rect 44265 666571 44331 666574
rect 673545 666634 673611 666637
rect 674833 666634 674899 666637
rect 673545 666632 674899 666634
rect 673545 666576 673550 666632
rect 673606 666576 674838 666632
rect 674894 666576 674899 666632
rect 673545 666574 674899 666576
rect 673545 666571 673611 666574
rect 674833 666571 674899 666574
rect 675293 666498 675359 666501
rect 675293 666496 676292 666498
rect 675293 666440 675298 666496
rect 675354 666440 676292 666496
rect 675293 666438 676292 666440
rect 675293 666435 675359 666438
rect 684125 666226 684191 666229
rect 684125 666224 684234 666226
rect 684125 666168 684130 666224
rect 684186 666168 684234 666224
rect 684125 666163 684234 666168
rect 684174 666060 684234 666163
rect 676806 665756 676812 665820
rect 676876 665756 676882 665820
rect 676814 665652 676874 665756
rect 673545 665274 673611 665277
rect 673545 665272 676292 665274
rect 673545 665216 673550 665272
rect 673606 665216 676292 665272
rect 673545 665214 676292 665216
rect 673545 665211 673611 665214
rect 40718 665076 40724 665140
rect 40788 665138 40794 665140
rect 41781 665138 41847 665141
rect 40788 665136 41847 665138
rect 40788 665080 41786 665136
rect 41842 665080 41847 665136
rect 40788 665078 41847 665080
rect 40788 665076 40794 665078
rect 41781 665075 41847 665078
rect 676029 664866 676095 664869
rect 676029 664864 676292 664866
rect 676029 664808 676034 664864
rect 676090 664808 676292 664864
rect 676029 664806 676292 664808
rect 676029 664803 676095 664806
rect 673545 664458 673611 664461
rect 673545 664456 676292 664458
rect 673545 664400 673550 664456
rect 673606 664400 676292 664456
rect 673545 664398 676292 664400
rect 673545 664395 673611 664398
rect 40534 663988 40540 664052
rect 40604 664050 40610 664052
rect 41781 664050 41847 664053
rect 40604 664048 41847 664050
rect 40604 663992 41786 664048
rect 41842 663992 41847 664048
rect 40604 663990 41847 663992
rect 40604 663988 40610 663990
rect 41781 663987 41847 663990
rect 672257 664050 672323 664053
rect 672257 664048 676292 664050
rect 672257 663992 672262 664048
rect 672318 663992 676292 664048
rect 672257 663990 676292 663992
rect 672257 663987 672323 663990
rect 673545 663778 673611 663781
rect 674833 663778 674899 663781
rect 673545 663776 674899 663778
rect 673545 663720 673550 663776
rect 673606 663720 674838 663776
rect 674894 663720 674899 663776
rect 673545 663718 674899 663720
rect 673545 663715 673611 663718
rect 674833 663715 674899 663718
rect 683205 663778 683271 663781
rect 683205 663776 683314 663778
rect 683205 663720 683210 663776
rect 683266 663720 683314 663776
rect 683205 663715 683314 663720
rect 683254 663612 683314 663715
rect 672901 662962 672967 662965
rect 676262 662962 676322 663204
rect 683481 662962 683547 662965
rect 672901 662960 676322 662962
rect 672901 662904 672906 662960
rect 672962 662904 676322 662960
rect 672901 662902 676322 662904
rect 683438 662960 683547 662962
rect 683438 662904 683486 662960
rect 683542 662904 683547 662960
rect 672901 662899 672967 662902
rect 683438 662899 683547 662904
rect 683438 662796 683498 662899
rect 674598 662356 674604 662420
rect 674668 662418 674674 662420
rect 674668 662358 676292 662418
rect 674668 662356 674674 662358
rect 673913 662010 673979 662013
rect 673913 662008 676292 662010
rect 673913 661952 673918 662008
rect 673974 661952 676292 662008
rect 673913 661950 676292 661952
rect 673913 661947 673979 661950
rect 674005 661602 674071 661605
rect 674005 661600 676292 661602
rect 674005 661544 674010 661600
rect 674066 661544 676292 661600
rect 674005 661542 676292 661544
rect 674005 661539 674071 661542
rect 674005 661194 674071 661197
rect 674005 661192 676292 661194
rect 674005 661136 674010 661192
rect 674066 661136 676292 661192
rect 674005 661134 676292 661136
rect 674005 661131 674071 661134
rect 62113 660922 62179 660925
rect 62113 660920 64706 660922
rect 62113 660864 62118 660920
rect 62174 660864 64706 660920
rect 62113 660862 64706 660864
rect 62113 660859 62179 660862
rect 64646 660638 64706 660862
rect 674005 660242 674071 660245
rect 674833 660242 674899 660245
rect 674005 660240 674899 660242
rect 674005 660184 674010 660240
rect 674066 660184 674838 660240
rect 674894 660184 674899 660240
rect 674005 660182 674899 660184
rect 674005 660179 674071 660182
rect 674833 660179 674899 660182
rect 683070 660109 683130 660756
rect 683070 660104 683179 660109
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660046 683179 660048
rect 683113 660043 683179 660046
rect 674005 659970 674071 659973
rect 674005 659968 676292 659970
rect 674005 659912 674010 659968
rect 674066 659912 676292 659968
rect 674005 659910 676292 659912
rect 674005 659907 674071 659910
rect 61377 659562 61443 659565
rect 61377 659560 64706 659562
rect 61377 659504 61382 659560
rect 61438 659504 64706 659560
rect 61377 659502 64706 659504
rect 61377 659499 61443 659502
rect 64646 659456 64706 659502
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42517 658610 42583 658613
rect 41708 658608 42583 658610
rect 41708 658552 42522 658608
rect 42578 658552 42583 658608
rect 41708 658550 42583 658552
rect 41708 658548 41714 658550
rect 42517 658547 42583 658550
rect 41781 658340 41847 658341
rect 41781 658336 41828 658340
rect 41892 658338 41898 658340
rect 62113 658338 62179 658341
rect 41781 658280 41786 658336
rect 41781 658276 41828 658280
rect 41892 658278 41938 658338
rect 62113 658336 64706 658338
rect 62113 658280 62118 658336
rect 62174 658280 64706 658336
rect 62113 658278 64706 658280
rect 41892 658276 41898 658278
rect 41781 658275 41847 658276
rect 62113 658275 62179 658278
rect 64646 658274 64706 658278
rect 62941 657658 63007 657661
rect 62941 657656 64706 657658
rect 62941 657600 62946 657656
rect 63002 657600 64706 657656
rect 62941 657598 64706 657600
rect 62941 657595 63007 657598
rect 41454 657188 41460 657252
rect 41524 657250 41530 657252
rect 41781 657250 41847 657253
rect 41524 657248 41847 657250
rect 41524 657192 41786 657248
rect 41842 657192 41847 657248
rect 41524 657190 41847 657192
rect 41524 657188 41530 657190
rect 41781 657187 41847 657190
rect 64646 657092 64706 657598
rect 62113 656570 62179 656573
rect 62113 656568 64706 656570
rect 62113 656512 62118 656568
rect 62174 656512 64706 656568
rect 62113 656510 64706 656512
rect 62113 656507 62179 656510
rect 64646 655910 64706 656510
rect 674005 655618 674071 655621
rect 675109 655618 675175 655621
rect 674005 655616 675175 655618
rect 674005 655560 674010 655616
rect 674066 655560 675114 655616
rect 675170 655560 675175 655616
rect 674005 655558 675175 655560
rect 674005 655555 674071 655558
rect 675109 655555 675175 655558
rect 62113 655346 62179 655349
rect 62113 655344 64706 655346
rect 62113 655288 62118 655344
rect 62174 655288 64706 655344
rect 62113 655286 64706 655288
rect 62113 655283 62179 655286
rect 64646 654728 64706 655286
rect 674230 652836 674236 652900
rect 674300 652898 674306 652900
rect 675385 652898 675451 652901
rect 674300 652896 675451 652898
rect 674300 652840 675390 652896
rect 675446 652840 675451 652896
rect 674300 652838 675451 652840
rect 674300 652836 674306 652838
rect 675385 652835 675451 652838
rect 671981 652490 672047 652493
rect 675109 652490 675175 652493
rect 671981 652488 675175 652490
rect 671981 652432 671986 652488
rect 672042 652432 675114 652488
rect 675170 652432 675175 652488
rect 671981 652430 675175 652432
rect 671981 652427 672047 652430
rect 675109 652427 675175 652430
rect 672809 649226 672875 649229
rect 675385 649226 675451 649229
rect 672809 649224 675451 649226
rect 672809 649168 672814 649224
rect 672870 649168 675390 649224
rect 675446 649168 675451 649224
rect 672809 649166 675451 649168
rect 672809 649163 672875 649166
rect 675385 649163 675451 649166
rect 672993 648818 673059 648821
rect 675109 648818 675175 648821
rect 672993 648816 675175 648818
rect 672993 648760 672998 648816
rect 673054 648760 675114 648816
rect 675170 648760 675175 648816
rect 672993 648758 675175 648760
rect 672993 648755 673059 648758
rect 675109 648755 675175 648758
rect 671705 647866 671771 647869
rect 675385 647866 675451 647869
rect 671705 647864 675451 647866
rect 671705 647808 671710 647864
rect 671766 647808 675390 647864
rect 675446 647808 675451 647864
rect 671705 647806 675451 647808
rect 671705 647803 671771 647806
rect 675385 647803 675451 647806
rect 667473 645826 667539 645829
rect 675109 645826 675175 645829
rect 667473 645824 675175 645826
rect 667473 645768 667478 645824
rect 667534 645768 675114 645824
rect 675170 645768 675175 645824
rect 667473 645766 675175 645768
rect 667473 645763 667539 645766
rect 675109 645763 675175 645766
rect 671245 645554 671311 645557
rect 675518 645554 675524 645556
rect 671245 645552 675524 645554
rect 671245 645496 671250 645552
rect 671306 645496 675524 645552
rect 671245 645494 675524 645496
rect 671245 645491 671311 645494
rect 675518 645492 675524 645494
rect 675588 645492 675594 645556
rect 35758 644741 35818 644912
rect 35758 644736 35867 644741
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644678 35867 644680
rect 35801 644675 35867 644678
rect 674189 644602 674255 644605
rect 675293 644602 675359 644605
rect 674189 644600 675359 644602
rect 674189 644544 674194 644600
rect 674250 644544 675298 644600
rect 675354 644544 675359 644600
rect 674189 644542 675359 644544
rect 674189 644539 674255 644542
rect 675293 644539 675359 644542
rect 38518 644333 38578 644504
rect 38518 644328 38627 644333
rect 38518 644272 38566 644328
rect 38622 644272 38627 644328
rect 38518 644270 38627 644272
rect 38561 644267 38627 644270
rect 669589 644330 669655 644333
rect 675385 644330 675451 644333
rect 669589 644328 675451 644330
rect 669589 644272 669594 644328
rect 669650 644272 675390 644328
rect 675446 644272 675451 644328
rect 669589 644270 675451 644272
rect 669589 644267 669655 644270
rect 675385 644267 675451 644270
rect 35390 643925 35450 644096
rect 35341 643920 35450 643925
rect 35341 643864 35346 643920
rect 35402 643864 35450 643920
rect 35341 643862 35450 643864
rect 35341 643859 35407 643862
rect 35574 643517 35634 643688
rect 675569 643652 675635 643653
rect 675518 643588 675524 643652
rect 675588 643650 675635 643652
rect 675588 643648 675680 643650
rect 675630 643592 675680 643648
rect 675588 643590 675680 643592
rect 675588 643588 675635 643590
rect 675569 643587 675635 643588
rect 35525 643512 35634 643517
rect 35801 643514 35867 643517
rect 35525 643456 35530 643512
rect 35586 643456 35634 643512
rect 35525 643454 35634 643456
rect 35758 643512 35867 643514
rect 35758 643456 35806 643512
rect 35862 643456 35867 643512
rect 35525 643451 35591 643454
rect 35758 643451 35867 643456
rect 35758 643280 35818 643451
rect 649950 643242 650010 643558
rect 673545 643514 673611 643517
rect 675293 643514 675359 643517
rect 673545 643512 675359 643514
rect 673545 643456 673550 643512
rect 673606 643456 675298 643512
rect 675354 643456 675359 643512
rect 673545 643454 675359 643456
rect 673545 643451 673611 643454
rect 675293 643451 675359 643454
rect 651465 643242 651531 643245
rect 649950 643240 651531 643242
rect 649950 643184 651470 643240
rect 651526 643184 651531 643240
rect 649950 643182 651531 643184
rect 651465 643179 651531 643182
rect 35390 642701 35450 642872
rect 35390 642696 35499 642701
rect 35801 642698 35867 642701
rect 35390 642640 35438 642696
rect 35494 642640 35499 642696
rect 35390 642638 35499 642640
rect 35433 642635 35499 642638
rect 35758 642696 35867 642698
rect 35758 642640 35806 642696
rect 35862 642640 35867 642696
rect 35758 642635 35867 642640
rect 35758 642464 35818 642635
rect 35617 642290 35683 642293
rect 35574 642288 35683 642290
rect 35574 642232 35622 642288
rect 35678 642232 35683 642288
rect 35574 642227 35683 642232
rect 35574 642056 35634 642227
rect 649950 641882 650010 642376
rect 652017 641882 652083 641885
rect 649950 641880 652083 641882
rect 649950 641824 652022 641880
rect 652078 641824 652083 641880
rect 649950 641822 652083 641824
rect 652017 641819 652083 641822
rect 673453 641746 673519 641749
rect 675293 641746 675359 641749
rect 673453 641744 675359 641746
rect 673453 641688 673458 641744
rect 673514 641688 675298 641744
rect 675354 641688 675359 641744
rect 673453 641686 675359 641688
rect 673453 641683 673519 641686
rect 675293 641683 675359 641686
rect 35758 641477 35818 641648
rect 35758 641472 35867 641477
rect 35758 641416 35806 641472
rect 35862 641416 35867 641472
rect 35758 641414 35867 641416
rect 35801 641411 35867 641414
rect 671245 641474 671311 641477
rect 675201 641474 675267 641477
rect 671245 641472 675267 641474
rect 671245 641416 671250 641472
rect 671306 641416 675206 641472
rect 675262 641416 675267 641472
rect 671245 641414 675267 641416
rect 671245 641411 671311 641414
rect 675201 641411 675267 641414
rect 35574 641069 35634 641240
rect 35574 641064 35683 641069
rect 35574 641008 35622 641064
rect 35678 641008 35683 641064
rect 35574 641006 35683 641008
rect 35617 641003 35683 641006
rect 41137 641066 41203 641069
rect 44541 641066 44607 641069
rect 41137 641064 44607 641066
rect 41137 641008 41142 641064
rect 41198 641008 44546 641064
rect 44602 641008 44607 641064
rect 41137 641006 44607 641008
rect 41137 641003 41203 641006
rect 44541 641003 44607 641006
rect 35758 640661 35818 640832
rect 649950 640794 650010 641194
rect 651465 640794 651531 640797
rect 649950 640792 651531 640794
rect 649950 640736 651470 640792
rect 651526 640736 651531 640792
rect 649950 640734 651531 640736
rect 651465 640731 651531 640734
rect 35758 640656 35867 640661
rect 35758 640600 35806 640656
rect 35862 640600 35867 640656
rect 35758 640598 35867 640600
rect 35801 640595 35867 640598
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 40861 640250 40927 640253
rect 45093 640250 45159 640253
rect 40861 640248 45159 640250
rect 40861 640192 40866 640248
rect 40922 640192 45098 640248
rect 45154 640192 45159 640248
rect 40861 640190 45159 640192
rect 40861 640187 40927 640190
rect 45093 640187 45159 640190
rect 651373 640114 651439 640117
rect 649950 640112 651439 640114
rect 649950 640056 651378 640112
rect 651434 640056 651439 640112
rect 649950 640054 651439 640056
rect 34470 639845 34530 640016
rect 649950 640012 650010 640054
rect 651373 640051 651439 640054
rect 34421 639840 34530 639845
rect 34421 639784 34426 639840
rect 34482 639784 34530 639840
rect 34421 639782 34530 639784
rect 39389 639842 39455 639845
rect 44357 639842 44423 639845
rect 39389 639840 44423 639842
rect 39389 639784 39394 639840
rect 39450 639784 44362 639840
rect 44418 639784 44423 639840
rect 39389 639782 44423 639784
rect 34421 639779 34487 639782
rect 39389 639779 39455 639782
rect 44357 639779 44423 639782
rect 35574 639437 35634 639608
rect 35525 639432 35634 639437
rect 35801 639434 35867 639437
rect 35525 639376 35530 639432
rect 35586 639376 35634 639432
rect 35525 639374 35634 639376
rect 35758 639432 35867 639434
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35525 639371 35591 639374
rect 35758 639371 35867 639376
rect 35758 639200 35818 639371
rect 35574 638621 35634 638792
rect 35574 638616 35683 638621
rect 35574 638560 35622 638616
rect 35678 638560 35683 638616
rect 35574 638558 35683 638560
rect 649766 638618 649826 638830
rect 651465 638618 651531 638621
rect 649766 638616 651531 638618
rect 649766 638560 651470 638616
rect 651526 638560 651531 638616
rect 649766 638558 651531 638560
rect 35617 638555 35683 638558
rect 651465 638555 651531 638558
rect 671337 638618 671403 638621
rect 675477 638618 675543 638621
rect 671337 638616 675543 638618
rect 671337 638560 671342 638616
rect 671398 638560 675482 638616
rect 675538 638560 675543 638616
rect 671337 638558 675543 638560
rect 671337 638555 671403 638558
rect 675477 638555 675543 638558
rect 35758 638213 35818 638384
rect 35758 638208 35867 638213
rect 651649 638210 651715 638213
rect 35758 638152 35806 638208
rect 35862 638152 35867 638208
rect 35758 638150 35867 638152
rect 35801 638147 35867 638150
rect 649950 638208 651715 638210
rect 649950 638152 651654 638208
rect 651710 638152 651715 638208
rect 649950 638150 651715 638152
rect 32446 637805 32506 637976
rect 32397 637800 32506 637805
rect 32397 637744 32402 637800
rect 32458 637744 32506 637800
rect 32397 637742 32506 637744
rect 32397 637739 32463 637742
rect 649950 637648 650010 638150
rect 651649 638147 651715 638150
rect 35206 637397 35266 637568
rect 676070 637468 676076 637532
rect 676140 637530 676146 637532
rect 680997 637530 681063 637533
rect 676140 637528 681063 637530
rect 676140 637472 681002 637528
rect 681058 637472 681063 637528
rect 676140 637470 681063 637472
rect 676140 637468 676146 637470
rect 680997 637467 681063 637470
rect 35157 637392 35266 637397
rect 35157 637336 35162 637392
rect 35218 637336 35266 637392
rect 35157 637334 35266 637336
rect 35157 637331 35223 637334
rect 35758 636989 35818 637160
rect 35758 636984 35867 636989
rect 35758 636928 35806 636984
rect 35862 636928 35867 636984
rect 35758 636926 35867 636928
rect 35801 636923 35867 636926
rect 35574 636581 35634 636752
rect 35525 636576 35634 636581
rect 35801 636578 35867 636581
rect 35525 636520 35530 636576
rect 35586 636520 35634 636576
rect 35525 636518 35634 636520
rect 35758 636576 35867 636578
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35525 636515 35591 636518
rect 35758 636515 35867 636520
rect 40033 636578 40099 636581
rect 43805 636578 43871 636581
rect 40033 636576 43871 636578
rect 40033 636520 40038 636576
rect 40094 636520 43810 636576
rect 43866 636520 43871 636576
rect 40033 636518 43871 636520
rect 40033 636515 40099 636518
rect 43805 636515 43871 636518
rect 35758 636344 35818 636515
rect 39113 636170 39179 636173
rect 44173 636170 44239 636173
rect 39113 636168 44239 636170
rect 39113 636112 39118 636168
rect 39174 636112 44178 636168
rect 44234 636112 44239 636168
rect 39113 636110 44239 636112
rect 39113 636107 39179 636110
rect 44173 636107 44239 636110
rect 35758 635765 35818 635936
rect 35758 635760 35867 635765
rect 35758 635704 35806 635760
rect 35862 635704 35867 635760
rect 35758 635702 35867 635704
rect 35801 635699 35867 635702
rect 39573 635762 39639 635765
rect 43989 635762 44055 635765
rect 39573 635760 44055 635762
rect 39573 635704 39578 635760
rect 39634 635704 43994 635760
rect 44050 635704 44055 635760
rect 39573 635702 44055 635704
rect 39573 635699 39639 635702
rect 43989 635699 44055 635702
rect 40542 635356 40602 635528
rect 40534 635292 40540 635356
rect 40604 635292 40610 635356
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 35758 634541 35818 634712
rect 35758 634536 35867 634541
rect 35758 634480 35806 634536
rect 35862 634480 35867 634536
rect 35758 634478 35867 634480
rect 35801 634475 35867 634478
rect 40125 634130 40191 634133
rect 43069 634130 43135 634133
rect 40125 634128 43135 634130
rect 40125 634072 40130 634128
rect 40186 634072 43074 634128
rect 43130 634072 43135 634128
rect 40125 634070 43135 634072
rect 40125 634067 40191 634070
rect 43069 634067 43135 634070
rect 35758 633725 35818 633896
rect 35758 633720 35867 633725
rect 35758 633664 35806 633720
rect 35862 633664 35867 633720
rect 35758 633662 35867 633664
rect 35801 633659 35867 633662
rect 41597 633314 41663 633317
rect 42057 633314 42123 633317
rect 41597 633312 42123 633314
rect 41597 633256 41602 633312
rect 41658 633256 42062 633312
rect 42118 633256 42123 633312
rect 41597 633254 42123 633256
rect 41597 633251 41663 633254
rect 42057 633251 42123 633254
rect 40585 632906 40651 632909
rect 42609 632906 42675 632909
rect 40585 632904 42675 632906
rect 40585 632848 40590 632904
rect 40646 632848 42614 632904
rect 42670 632848 42675 632904
rect 40585 632846 42675 632848
rect 40585 632843 40651 632846
rect 42609 632843 42675 632846
rect 675150 631348 675156 631412
rect 675220 631410 675226 631412
rect 675477 631410 675543 631413
rect 675220 631408 675543 631410
rect 675220 631352 675482 631408
rect 675538 631352 675543 631408
rect 675220 631350 675543 631352
rect 675220 631348 675226 631350
rect 675477 631347 675543 631350
rect 675661 631410 675727 631413
rect 676070 631410 676076 631412
rect 675661 631408 676076 631410
rect 675661 631352 675666 631408
rect 675722 631352 676076 631408
rect 675661 631350 676076 631352
rect 675661 631347 675727 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 40033 630866 40099 630869
rect 43621 630866 43687 630869
rect 40033 630864 43687 630866
rect 40033 630808 40038 630864
rect 40094 630808 43626 630864
rect 43682 630808 43687 630864
rect 40033 630806 43687 630808
rect 40033 630803 40099 630806
rect 43621 630803 43687 630806
rect 32397 629914 32463 629917
rect 41638 629914 41644 629916
rect 32397 629912 41644 629914
rect 32397 629856 32402 629912
rect 32458 629856 41644 629912
rect 32397 629854 41644 629856
rect 32397 629851 32463 629854
rect 41638 629852 41644 629854
rect 41708 629852 41714 629916
rect 39297 629234 39363 629237
rect 41822 629234 41828 629236
rect 39297 629232 41828 629234
rect 39297 629176 39302 629232
rect 39358 629176 41828 629232
rect 39297 629174 41828 629176
rect 39297 629171 39363 629174
rect 41822 629172 41828 629174
rect 41892 629172 41898 629236
rect 39389 628690 39455 628693
rect 42609 628690 42675 628693
rect 39389 628688 42675 628690
rect 39389 628632 39394 628688
rect 39450 628632 42614 628688
rect 42670 628632 42675 628688
rect 39389 628630 42675 628632
rect 39389 628627 39455 628630
rect 42609 628627 42675 628630
rect 41781 627464 41847 627469
rect 41781 627408 41786 627464
rect 41842 627408 41847 627464
rect 41781 627403 41847 627408
rect 41784 627197 41844 627403
rect 41781 627192 41847 627197
rect 41781 627136 41786 627192
rect 41842 627136 41847 627192
rect 41781 627131 41847 627136
rect 673269 626106 673335 626109
rect 676262 626106 676322 626348
rect 673269 626104 676322 626106
rect 673269 626048 673274 626104
rect 673330 626048 676322 626104
rect 673269 626046 676322 626048
rect 673269 626043 673335 626046
rect 676262 625701 676322 625940
rect 676213 625696 676322 625701
rect 676213 625640 676218 625696
rect 676274 625640 676322 625696
rect 676213 625638 676322 625640
rect 676213 625635 676279 625638
rect 676262 625460 676322 625532
rect 673269 625426 673335 625429
rect 676078 625426 676322 625460
rect 673269 625424 676322 625426
rect 673269 625368 673274 625424
rect 673330 625400 676322 625424
rect 673330 625368 676138 625400
rect 673269 625366 676138 625368
rect 673269 625363 673335 625366
rect 673269 625154 673335 625157
rect 674281 625154 674347 625157
rect 673269 625152 674347 625154
rect 673269 625096 673274 625152
rect 673330 625096 674286 625152
rect 674342 625096 674347 625152
rect 673269 625094 674347 625096
rect 673269 625091 673335 625094
rect 674281 625091 674347 625094
rect 676262 624882 676322 625124
rect 674422 624822 676322 624882
rect 42149 624610 42215 624613
rect 44173 624610 44239 624613
rect 42149 624608 44239 624610
rect 42149 624552 42154 624608
rect 42210 624552 44178 624608
rect 44234 624552 44239 624608
rect 42149 624550 44239 624552
rect 42149 624547 42215 624550
rect 44173 624547 44239 624550
rect 672625 624474 672691 624477
rect 674422 624474 674482 624822
rect 676262 624477 676322 624716
rect 672625 624472 674482 624474
rect 672625 624416 672630 624472
rect 672686 624416 674482 624472
rect 672625 624414 674482 624416
rect 676213 624472 676322 624477
rect 676213 624416 676218 624472
rect 676274 624416 676322 624472
rect 676213 624414 676322 624416
rect 672625 624411 672691 624414
rect 676213 624411 676279 624414
rect 676262 624236 676322 624308
rect 671429 624202 671495 624205
rect 676078 624202 676322 624236
rect 671429 624200 676322 624202
rect 671429 624144 671434 624200
rect 671490 624176 676322 624200
rect 671490 624144 676138 624176
rect 671429 624142 676138 624144
rect 671429 624139 671495 624142
rect 674005 623930 674071 623933
rect 674005 623928 676292 623930
rect 674005 623872 674010 623928
rect 674066 623872 676292 623928
rect 674005 623870 676292 623872
rect 674005 623867 674071 623870
rect 672625 623794 672691 623797
rect 673318 623794 673562 623828
rect 672625 623792 673562 623794
rect 672625 623736 672630 623792
rect 672686 623768 673562 623792
rect 672686 623736 673378 623768
rect 672625 623734 673378 623736
rect 672625 623731 672691 623734
rect 673502 623658 673562 623768
rect 674281 623658 674347 623661
rect 673502 623656 674347 623658
rect 673502 623600 674286 623656
rect 674342 623600 674347 623656
rect 673502 623598 674347 623600
rect 674281 623595 674347 623598
rect 672625 623250 672691 623253
rect 676262 623250 676322 623492
rect 672625 623248 676322 623250
rect 672625 623192 672630 623248
rect 672686 623192 676322 623248
rect 672625 623190 676322 623192
rect 672625 623187 672691 623190
rect 676446 622845 676506 623084
rect 676397 622840 676506 622845
rect 676397 622784 676402 622840
rect 676458 622784 676506 622840
rect 676397 622782 676506 622784
rect 676397 622779 676463 622782
rect 676029 622706 676095 622709
rect 676029 622704 676292 622706
rect 676029 622648 676034 622704
rect 676090 622648 676292 622704
rect 676029 622646 676292 622648
rect 676029 622643 676095 622646
rect 672625 622434 672691 622437
rect 674281 622434 674347 622437
rect 672625 622432 674347 622434
rect 672625 622376 672630 622432
rect 672686 622376 674286 622432
rect 674342 622376 674347 622432
rect 672625 622374 674347 622376
rect 672625 622371 672691 622374
rect 674281 622371 674347 622374
rect 40718 621964 40724 622028
rect 40788 622026 40794 622028
rect 41781 622026 41847 622029
rect 40788 622024 41847 622026
rect 40788 621968 41786 622024
rect 41842 621968 41847 622024
rect 40788 621966 41847 621968
rect 40788 621964 40794 621966
rect 41781 621963 41847 621966
rect 42149 622026 42215 622029
rect 44173 622026 44239 622029
rect 676262 622026 676322 622268
rect 42149 622024 44239 622026
rect 42149 621968 42154 622024
rect 42210 621968 44178 622024
rect 44234 621968 44239 622024
rect 42149 621966 44239 621968
rect 42149 621963 42215 621966
rect 44173 621963 44239 621966
rect 674606 621966 676322 622026
rect 680997 622026 681063 622029
rect 680997 622024 681106 622026
rect 680997 621968 681002 622024
rect 681058 621968 681106 622024
rect 674606 621346 674666 621966
rect 680997 621963 681106 621968
rect 681046 621860 681106 621963
rect 676029 621482 676095 621485
rect 676029 621480 676292 621482
rect 676029 621424 676034 621480
rect 676090 621424 676292 621480
rect 676029 621422 676292 621424
rect 676029 621419 676095 621422
rect 673686 621286 674666 621346
rect 673269 621210 673335 621213
rect 673686 621210 673746 621286
rect 673269 621208 673746 621210
rect 673269 621152 673274 621208
rect 673330 621152 673746 621208
rect 673269 621150 673746 621152
rect 673269 621147 673335 621150
rect 674005 621074 674071 621077
rect 674005 621072 676292 621074
rect 674005 621016 674010 621072
rect 674066 621016 676292 621072
rect 674005 621014 676292 621016
rect 674005 621011 674071 621014
rect 40534 620740 40540 620804
rect 40604 620802 40610 620804
rect 41781 620802 41847 620805
rect 40604 620800 41847 620802
rect 40604 620744 41786 620800
rect 41842 620744 41847 620800
rect 40604 620742 41847 620744
rect 40604 620740 40610 620742
rect 41781 620739 41847 620742
rect 676213 620802 676279 620805
rect 676213 620800 676322 620802
rect 676213 620744 676218 620800
rect 676274 620744 676322 620800
rect 676213 620739 676322 620744
rect 676262 620636 676322 620739
rect 676262 619989 676322 620228
rect 676213 619984 676322 619989
rect 676489 619986 676555 619989
rect 676213 619928 676218 619984
rect 676274 619928 676322 619984
rect 676213 619926 676322 619928
rect 676446 619984 676555 619986
rect 676446 619928 676494 619984
rect 676550 619928 676555 619984
rect 676213 619923 676279 619926
rect 676446 619923 676555 619928
rect 676446 619820 676506 619923
rect 676213 619578 676279 619581
rect 676213 619576 676322 619578
rect 676213 619520 676218 619576
rect 676274 619520 676322 619576
rect 676213 619515 676322 619520
rect 676262 619412 676322 619515
rect 674414 618972 674420 619036
rect 674484 619034 674490 619036
rect 674484 618974 676292 619034
rect 674484 618972 674490 618974
rect 683205 618762 683271 618765
rect 683205 618760 683314 618762
rect 683205 618704 683210 618760
rect 683266 618704 683314 618760
rect 683205 618699 683314 618704
rect 683254 618596 683314 618699
rect 673269 618218 673335 618221
rect 673269 618216 676292 618218
rect 673269 618160 673274 618216
rect 673330 618160 676292 618216
rect 673269 618158 676292 618160
rect 673269 618155 673335 618158
rect 63125 618082 63191 618085
rect 63125 618080 64706 618082
rect 63125 618024 63130 618080
rect 63186 618024 64706 618080
rect 63125 618022 64706 618024
rect 63125 618019 63191 618022
rect 64646 617416 64706 618022
rect 676029 617810 676095 617813
rect 676029 617808 676292 617810
rect 676029 617752 676034 617808
rect 676090 617752 676292 617808
rect 676029 617750 676292 617752
rect 676029 617747 676095 617750
rect 673729 617402 673795 617405
rect 673729 617400 676292 617402
rect 673729 617344 673734 617400
rect 673790 617344 676292 617400
rect 673729 617342 676292 617344
rect 673729 617339 673795 617342
rect 675293 617130 675359 617133
rect 676806 617130 676812 617132
rect 675293 617128 676812 617130
rect 675293 617072 675298 617128
rect 675354 617072 676812 617128
rect 675293 617070 676812 617072
rect 675293 617067 675359 617070
rect 676806 617068 676812 617070
rect 676876 617068 676882 617132
rect 683573 617130 683639 617133
rect 683573 617128 683682 617130
rect 683573 617072 683578 617128
rect 683634 617072 683682 617128
rect 683573 617067 683682 617072
rect 683622 616964 683682 617067
rect 683389 616722 683455 616725
rect 683389 616720 683498 616722
rect 683389 616664 683394 616720
rect 683450 616664 683498 616720
rect 683389 616659 683498 616664
rect 62113 616586 62179 616589
rect 62113 616584 64706 616586
rect 62113 616528 62118 616584
rect 62174 616528 64706 616584
rect 683438 616556 683498 616659
rect 62113 616526 64706 616528
rect 62113 616523 62179 616526
rect 64646 616234 64706 616526
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 41454 615708 41460 615772
rect 41524 615770 41530 615772
rect 42333 615770 42399 615773
rect 41524 615768 42399 615770
rect 41524 615712 42338 615768
rect 42394 615712 42399 615768
rect 41524 615710 42399 615712
rect 41524 615708 41530 615710
rect 42333 615707 42399 615710
rect 683070 615501 683130 615740
rect 41822 615436 41828 615500
rect 41892 615498 41898 615500
rect 42609 615498 42675 615501
rect 41892 615496 42675 615498
rect 41892 615440 42614 615496
rect 42670 615440 42675 615496
rect 41892 615438 42675 615440
rect 41892 615436 41898 615438
rect 42609 615435 42675 615438
rect 683070 615498 683179 615501
rect 683070 615496 683260 615498
rect 683070 615440 683118 615496
rect 683174 615440 683260 615496
rect 683070 615438 683260 615440
rect 683070 615435 683179 615438
rect 683070 615332 683130 615435
rect 62113 614682 62179 614685
rect 64646 614682 64706 615052
rect 674005 614954 674071 614957
rect 674005 614952 676292 614954
rect 674005 614896 674010 614952
rect 674066 614896 676292 614952
rect 674005 614894 676292 614896
rect 674005 614891 674071 614894
rect 62113 614680 64706 614682
rect 62113 614624 62118 614680
rect 62174 614624 64706 614680
rect 62113 614622 64706 614624
rect 62113 614619 62179 614622
rect 42885 614274 42951 614277
rect 44081 614274 44147 614277
rect 42885 614272 44147 614274
rect 42885 614216 42890 614272
rect 42946 614216 44086 614272
rect 44142 614216 44147 614272
rect 42885 614214 44147 614216
rect 42885 614211 42951 614214
rect 44081 614211 44147 614214
rect 61377 613866 61443 613869
rect 64646 613866 64706 613870
rect 61377 613864 64706 613866
rect 61377 613808 61382 613864
rect 61438 613808 64706 613864
rect 61377 613806 64706 613808
rect 61377 613803 61443 613806
rect 41873 613460 41939 613461
rect 41822 613458 41828 613460
rect 41782 613398 41828 613458
rect 41892 613456 41939 613460
rect 41934 613400 41939 613456
rect 41822 613396 41828 613398
rect 41892 613396 41939 613400
rect 41873 613395 41939 613396
rect 62113 612642 62179 612645
rect 64646 612642 64706 612688
rect 62113 612640 64706 612642
rect 62113 612584 62118 612640
rect 62174 612584 64706 612640
rect 62113 612582 64706 612584
rect 62113 612579 62179 612582
rect 40534 612308 40540 612372
rect 40604 612370 40610 612372
rect 42241 612370 42307 612373
rect 40604 612368 42307 612370
rect 40604 612312 42246 612368
rect 42302 612312 42307 612368
rect 40604 612310 42307 612312
rect 40604 612308 40610 612310
rect 42241 612307 42307 612310
rect 62941 612098 63007 612101
rect 62941 612096 64706 612098
rect 62941 612040 62946 612096
rect 63002 612040 64706 612096
rect 62941 612038 64706 612040
rect 62941 612035 63007 612038
rect 43759 611826 43825 611829
rect 43759 611824 51090 611826
rect 43759 611768 43764 611824
rect 43820 611768 51090 611824
rect 43759 611766 51090 611768
rect 43759 611763 43825 611766
rect 51030 611690 51090 611766
rect 55857 611690 55923 611693
rect 51030 611688 55923 611690
rect 51030 611632 55862 611688
rect 55918 611632 55923 611688
rect 51030 611630 55923 611632
rect 55857 611627 55923 611630
rect 64646 611506 64706 612038
rect 43989 611418 44055 611421
rect 64137 611418 64203 611421
rect 43989 611416 64203 611418
rect 43989 611360 43994 611416
rect 44050 611360 64142 611416
rect 64198 611360 64203 611416
rect 43989 611358 64203 611360
rect 43989 611355 44055 611358
rect 64137 611355 64203 611358
rect 43437 611146 43503 611149
rect 44725 611146 44791 611149
rect 43437 611144 44791 611146
rect 43437 611088 43442 611144
rect 43498 611088 44730 611144
rect 44786 611088 44791 611144
rect 43437 611086 44791 611088
rect 43437 611083 43503 611086
rect 44725 611083 44791 611086
rect 43621 610738 43687 610741
rect 44725 610738 44791 610741
rect 43621 610736 44791 610738
rect 43621 610680 43626 610736
rect 43682 610680 44730 610736
rect 44786 610680 44791 610736
rect 43621 610678 44791 610680
rect 43621 610675 43687 610678
rect 44725 610675 44791 610678
rect 670969 607746 671035 607749
rect 675477 607746 675543 607749
rect 670969 607744 675543 607746
rect 670969 607688 670974 607744
rect 671030 607688 675482 607744
rect 675538 607688 675543 607744
rect 670969 607686 675543 607688
rect 670969 607683 671035 607686
rect 675477 607683 675543 607686
rect 673269 607338 673335 607341
rect 675293 607338 675359 607341
rect 673269 607336 675359 607338
rect 673269 607280 673274 607336
rect 673330 607280 675298 607336
rect 675354 607280 675359 607336
rect 673269 607278 675359 607280
rect 673269 607275 673335 607278
rect 675293 607275 675359 607278
rect 672349 604482 672415 604485
rect 675109 604482 675175 604485
rect 672349 604480 675175 604482
rect 672349 604424 672354 604480
rect 672410 604424 675114 604480
rect 675170 604424 675175 604480
rect 672349 604422 675175 604424
rect 672349 604419 672415 604422
rect 675109 604419 675175 604422
rect 674414 602924 674420 602988
rect 674484 602986 674490 602988
rect 675109 602986 675175 602989
rect 674484 602984 675175 602986
rect 674484 602928 675114 602984
rect 675170 602928 675175 602984
rect 674484 602926 675175 602928
rect 674484 602924 674490 602926
rect 675109 602923 675175 602926
rect 40309 602034 40375 602037
rect 40534 602034 40540 602036
rect 40309 602032 40540 602034
rect 40309 601976 40314 602032
rect 40370 601976 40540 602032
rect 40309 601974 40540 601976
rect 40309 601971 40375 601974
rect 40534 601972 40540 601974
rect 40604 601972 40610 602036
rect 35801 601762 35867 601765
rect 35788 601760 35867 601762
rect 35788 601704 35806 601760
rect 35862 601704 35867 601760
rect 35788 601702 35867 601704
rect 35801 601699 35867 601702
rect 39941 601354 40007 601357
rect 39941 601352 40020 601354
rect 39941 601296 39946 601352
rect 40002 601296 40020 601352
rect 39941 601294 40020 601296
rect 39941 601291 40007 601294
rect 40125 600946 40191 600949
rect 667289 600946 667355 600949
rect 675385 600946 675451 600949
rect 40125 600944 40204 600946
rect 40125 600888 40130 600944
rect 40186 600888 40204 600944
rect 40125 600886 40204 600888
rect 667289 600944 675451 600946
rect 667289 600888 667294 600944
rect 667350 600888 675390 600944
rect 675446 600888 675451 600944
rect 667289 600886 675451 600888
rect 40125 600883 40191 600886
rect 667289 600883 667355 600886
rect 675385 600883 675451 600886
rect 44541 600538 44607 600541
rect 41492 600536 44607 600538
rect 41492 600480 44546 600536
rect 44602 600480 44607 600536
rect 41492 600478 44607 600480
rect 44541 600475 44607 600478
rect 44633 600130 44699 600133
rect 41492 600128 44699 600130
rect 41492 600072 44638 600128
rect 44694 600072 44699 600128
rect 41492 600070 44699 600072
rect 44633 600067 44699 600070
rect 44449 599722 44515 599725
rect 41492 599720 44515 599722
rect 41492 599664 44454 599720
rect 44510 599664 44515 599720
rect 41492 599662 44515 599664
rect 44449 599659 44515 599662
rect 44909 599314 44975 599317
rect 41492 599312 44975 599314
rect 41492 599256 44914 599312
rect 44970 599256 44975 599312
rect 41492 599254 44975 599256
rect 44909 599251 44975 599254
rect 674189 599042 674255 599045
rect 675477 599042 675543 599045
rect 674189 599040 675543 599042
rect 674189 598984 674194 599040
rect 674250 598984 675482 599040
rect 675538 598984 675543 599040
rect 674189 598982 675543 598984
rect 674189 598979 674255 598982
rect 675477 598979 675543 598982
rect 45093 598906 45159 598909
rect 41492 598904 45159 598906
rect 41492 598848 45098 598904
rect 45154 598848 45159 598904
rect 41492 598846 45159 598848
rect 45093 598843 45159 598846
rect 673913 598634 673979 598637
rect 675477 598634 675543 598637
rect 673913 598632 675543 598634
rect 673913 598576 673918 598632
rect 673974 598576 675482 598632
rect 675538 598576 675543 598632
rect 673913 598574 675543 598576
rect 673913 598571 673979 598574
rect 675477 598571 675543 598574
rect 43110 598498 43116 598500
rect 41492 598438 43116 598498
rect 43110 598436 43116 598438
rect 43180 598436 43186 598500
rect 45277 598090 45343 598093
rect 41492 598088 45343 598090
rect 41492 598032 45282 598088
rect 45338 598032 45343 598088
rect 41492 598030 45343 598032
rect 45277 598027 45343 598030
rect 649950 597954 650010 598336
rect 651465 597954 651531 597957
rect 649950 597952 651531 597954
rect 649950 597896 651470 597952
rect 651526 597896 651531 597952
rect 649950 597894 651531 597896
rect 651465 597891 651531 597894
rect 42885 597682 42951 597685
rect 41492 597680 42951 597682
rect 41492 597624 42890 597680
rect 42946 597624 42951 597680
rect 41492 597622 42951 597624
rect 42885 597619 42951 597622
rect 672533 597410 672599 597413
rect 675477 597410 675543 597413
rect 672533 597408 675543 597410
rect 672533 597352 672538 597408
rect 672594 597352 675482 597408
rect 675538 597352 675543 597408
rect 672533 597350 675543 597352
rect 672533 597347 672599 597350
rect 675477 597347 675543 597350
rect 42006 597274 42012 597276
rect 41492 597214 42012 597274
rect 42006 597212 42012 597214
rect 42076 597212 42082 597276
rect 43069 597004 43135 597005
rect 43069 597000 43116 597004
rect 43180 597002 43186 597004
rect 43069 596944 43074 597000
rect 43069 596940 43116 596944
rect 43180 596942 43226 597002
rect 43180 596940 43186 596942
rect 43069 596939 43135 596940
rect 40953 596866 41019 596869
rect 40940 596864 41019 596866
rect 40940 596808 40958 596864
rect 41014 596808 41019 596864
rect 40940 596806 41019 596808
rect 40953 596803 41019 596806
rect 649950 596730 650010 597154
rect 651465 596730 651531 596733
rect 649950 596728 651531 596730
rect 649950 596672 651470 596728
rect 651526 596672 651531 596728
rect 649950 596670 651531 596672
rect 651465 596667 651531 596670
rect 41137 596458 41203 596461
rect 41124 596456 41203 596458
rect 41124 596400 41142 596456
rect 41198 596400 41203 596456
rect 41124 596398 41203 596400
rect 41137 596395 41203 596398
rect 41278 595815 41338 596020
rect 35157 595812 35223 595815
rect 35157 595810 35266 595812
rect 35157 595754 35162 595810
rect 35218 595754 35266 595810
rect 35157 595749 35266 595754
rect 41278 595810 41387 595815
rect 41278 595754 41326 595810
rect 41382 595754 41387 595810
rect 41278 595752 41387 595754
rect 41321 595749 41387 595752
rect 41689 595778 41755 595781
rect 63309 595778 63375 595781
rect 41689 595776 63375 595778
rect 35206 595612 35266 595749
rect 41689 595720 41694 595776
rect 41750 595720 63314 595776
rect 63370 595720 63375 595776
rect 41689 595718 63375 595720
rect 41689 595715 41755 595718
rect 63309 595715 63375 595718
rect 649950 595370 650010 595972
rect 651465 595370 651531 595373
rect 649950 595368 651531 595370
rect 649950 595312 651470 595368
rect 651526 595312 651531 595368
rect 649950 595310 651531 595312
rect 651465 595307 651531 595310
rect 674966 595308 674972 595372
rect 675036 595370 675042 595372
rect 675385 595370 675451 595373
rect 675036 595368 675451 595370
rect 675036 595312 675390 595368
rect 675446 595312 675451 595368
rect 675036 595310 675451 595312
rect 675036 595308 675042 595310
rect 675385 595307 675451 595310
rect 33041 595234 33107 595237
rect 33028 595232 33107 595234
rect 33028 595176 33046 595232
rect 33102 595176 33107 595232
rect 33028 595174 33107 595176
rect 33041 595171 33107 595174
rect 651649 595098 651715 595101
rect 649950 595096 651715 595098
rect 649950 595040 651654 595096
rect 651710 595040 651715 595096
rect 649950 595038 651715 595040
rect 37966 594591 38026 594796
rect 649950 594790 650010 595038
rect 651649 595035 651715 595038
rect 668761 594826 668827 594829
rect 675201 594826 675267 594829
rect 668761 594824 675267 594826
rect 668761 594768 668766 594824
rect 668822 594768 675206 594824
rect 675262 594768 675267 594824
rect 668761 594766 675267 594768
rect 668761 594763 668827 594766
rect 675201 594763 675267 594766
rect 37917 594586 38026 594591
rect 37917 594530 37922 594586
rect 37978 594530 38026 594586
rect 37917 594528 38026 594530
rect 41689 594554 41755 594557
rect 673453 594554 673519 594557
rect 675201 594554 675267 594557
rect 41689 594552 51090 594554
rect 37917 594525 37983 594528
rect 41689 594496 41694 594552
rect 41750 594496 51090 594552
rect 41689 594494 51090 594496
rect 41689 594491 41755 594494
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 51030 594146 51090 594494
rect 673453 594552 675267 594554
rect 673453 594496 673458 594552
rect 673514 594496 675206 594552
rect 675262 594496 675267 594552
rect 673453 594494 675267 594496
rect 673453 594491 673519 594494
rect 675201 594491 675267 594494
rect 63125 594146 63191 594149
rect 651465 594146 651531 594149
rect 51030 594144 63191 594146
rect 51030 594088 63130 594144
rect 63186 594088 63191 594144
rect 51030 594086 63191 594088
rect 63125 594083 63191 594086
rect 649950 594144 651531 594146
rect 649950 594088 651470 594144
rect 651526 594088 651531 594144
rect 649950 594086 651531 594088
rect 41822 594010 41828 594012
rect 41492 593950 41828 594010
rect 41822 593948 41828 593950
rect 41892 593948 41898 594012
rect 649950 593608 650010 594086
rect 651465 594083 651531 594086
rect 33777 593602 33843 593605
rect 33764 593600 33843 593602
rect 33764 593544 33782 593600
rect 33838 593544 33843 593600
rect 33764 593542 33843 593544
rect 33777 593539 33843 593542
rect 668945 593466 669011 593469
rect 675385 593466 675451 593469
rect 668945 593464 675451 593466
rect 668945 593408 668950 593464
rect 669006 593408 675390 593464
rect 675446 593408 675451 593464
rect 668945 593406 675451 593408
rect 668945 593403 669011 593406
rect 675385 593403 675451 593406
rect 44357 593194 44423 593197
rect 41492 593192 44423 593194
rect 41492 593136 44362 593192
rect 44418 593136 44423 593192
rect 41492 593134 44423 593136
rect 44357 593131 44423 593134
rect 675150 593132 675156 593196
rect 675220 593194 675226 593196
rect 675477 593194 675543 593197
rect 675220 593192 675543 593194
rect 675220 593136 675482 593192
rect 675538 593136 675543 593192
rect 675220 593134 675543 593136
rect 675220 593132 675226 593134
rect 675477 593131 675543 593134
rect 651465 592922 651531 592925
rect 649950 592920 651531 592922
rect 649950 592864 651470 592920
rect 651526 592864 651531 592920
rect 649950 592862 651531 592864
rect 40726 592550 40786 592756
rect 40718 592486 40724 592550
rect 40788 592486 40794 592550
rect 649950 592426 650010 592862
rect 651465 592859 651531 592862
rect 41822 592378 41828 592380
rect 41492 592318 41828 592378
rect 41822 592316 41828 592318
rect 41892 592316 41898 592380
rect 41689 592106 41755 592109
rect 42190 592106 42196 592108
rect 41689 592104 42196 592106
rect 41689 592048 41694 592104
rect 41750 592048 42196 592104
rect 41689 592046 42196 592048
rect 41689 592043 41755 592046
rect 42190 592044 42196 592046
rect 42260 592044 42266 592108
rect 35617 591970 35683 591973
rect 35604 591968 35683 591970
rect 35604 591912 35622 591968
rect 35678 591912 35683 591968
rect 35604 591910 35683 591912
rect 35617 591907 35683 591910
rect 676070 591636 676076 591700
rect 676140 591698 676146 591700
rect 680997 591698 681063 591701
rect 676140 591696 681063 591698
rect 676140 591640 681002 591696
rect 681058 591640 681063 591696
rect 676140 591638 681063 591640
rect 676140 591636 676146 591638
rect 680997 591635 681063 591638
rect 35801 591562 35867 591565
rect 35788 591560 35867 591562
rect 35788 591504 35806 591560
rect 35862 591504 35867 591560
rect 35788 591502 35867 591504
rect 35801 591499 35867 591502
rect 674230 591228 674236 591292
rect 674300 591290 674306 591292
rect 684217 591290 684283 591293
rect 674300 591288 684283 591290
rect 674300 591232 684222 591288
rect 684278 591232 684283 591288
rect 674300 591230 684283 591232
rect 674300 591228 674306 591230
rect 684217 591227 684283 591230
rect 41462 590746 41522 591124
rect 62941 590746 63007 590749
rect 41462 590744 63007 590746
rect 41462 590716 62946 590744
rect 41492 590688 62946 590716
rect 63002 590688 63007 590744
rect 41492 590686 63007 590688
rect 62941 590683 63007 590686
rect 41689 590474 41755 590477
rect 43253 590474 43319 590477
rect 674925 590476 674991 590477
rect 674925 590474 674972 590476
rect 41689 590472 43319 590474
rect 41689 590416 41694 590472
rect 41750 590416 43258 590472
rect 43314 590416 43319 590472
rect 41689 590414 43319 590416
rect 674880 590472 674972 590474
rect 674880 590416 674930 590472
rect 674880 590414 674972 590416
rect 41689 590411 41755 590414
rect 43253 590411 43319 590414
rect 674925 590412 674972 590414
rect 675036 590412 675042 590476
rect 674925 590411 674991 590412
rect 62481 590066 62547 590069
rect 51030 590064 62547 590066
rect 51030 590008 62486 590064
rect 62542 590008 62547 590064
rect 51030 590006 62547 590008
rect 36537 589658 36603 589661
rect 51030 589658 51090 590006
rect 62481 590003 62547 590006
rect 36537 589656 51090 589658
rect 36537 589600 36542 589656
rect 36598 589600 51090 589656
rect 36537 589598 51090 589600
rect 36537 589595 36603 589598
rect 39757 589386 39823 589389
rect 43437 589386 43503 589389
rect 39757 589384 43503 589386
rect 39757 589328 39762 589384
rect 39818 589328 43442 589384
rect 43498 589328 43503 589384
rect 39757 589326 43503 589328
rect 39757 589323 39823 589326
rect 43437 589323 43503 589326
rect 675201 586258 675267 586261
rect 676070 586258 676076 586260
rect 675201 586256 676076 586258
rect 675201 586200 675206 586256
rect 675262 586200 676076 586256
rect 675201 586198 676076 586200
rect 675201 586195 675267 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 40585 585986 40651 585989
rect 42425 585986 42491 585989
rect 40585 585984 42491 585986
rect 40585 585928 40590 585984
rect 40646 585928 42430 585984
rect 42486 585928 42491 585984
rect 40585 585926 42491 585928
rect 40585 585923 40651 585926
rect 42425 585923 42491 585926
rect 40401 585714 40467 585717
rect 62062 585714 62068 585716
rect 40401 585712 62068 585714
rect 40401 585656 40406 585712
rect 40462 585656 62068 585712
rect 40401 585654 62068 585656
rect 40401 585651 40467 585654
rect 62062 585652 62068 585654
rect 62132 585652 62138 585716
rect 37917 585170 37983 585173
rect 41822 585170 41828 585172
rect 37917 585168 41828 585170
rect 37917 585112 37922 585168
rect 37978 585112 41828 585168
rect 37917 585110 41828 585112
rect 37917 585107 37983 585110
rect 41822 585108 41828 585110
rect 41892 585108 41898 585172
rect 39849 584626 39915 584629
rect 40350 584626 40356 584628
rect 39849 584624 40356 584626
rect 39849 584568 39854 584624
rect 39910 584568 40356 584624
rect 39849 584566 40356 584568
rect 39849 584563 39915 584566
rect 40350 584564 40356 584566
rect 40420 584564 40426 584628
rect 673545 581362 673611 581365
rect 674465 581362 674531 581365
rect 673545 581360 674531 581362
rect 673545 581304 673550 581360
rect 673606 581304 674470 581360
rect 674526 581304 674531 581360
rect 673545 581302 674531 581304
rect 673545 581299 673611 581302
rect 674465 581299 674531 581302
rect 674005 581090 674071 581093
rect 674005 581088 676292 581090
rect 674005 581032 674010 581088
rect 674066 581032 676292 581088
rect 674005 581030 676292 581032
rect 674005 581027 674071 581030
rect 673545 580682 673611 580685
rect 673545 580680 676292 580682
rect 673545 580624 673550 580680
rect 673606 580624 676292 580680
rect 673545 580622 676292 580624
rect 673545 580619 673611 580622
rect 40350 580212 40356 580276
rect 40420 580274 40426 580276
rect 41781 580274 41847 580277
rect 40420 580272 41847 580274
rect 40420 580216 41786 580272
rect 41842 580216 41847 580272
rect 40420 580214 41847 580216
rect 40420 580212 40426 580214
rect 41781 580211 41847 580214
rect 42241 580274 42307 580277
rect 45093 580274 45159 580277
rect 42241 580272 45159 580274
rect 42241 580216 42246 580272
rect 42302 580216 45098 580272
rect 45154 580216 45159 580272
rect 42241 580214 45159 580216
rect 42241 580211 42307 580214
rect 45093 580211 45159 580214
rect 674005 580274 674071 580277
rect 674005 580272 676292 580274
rect 674005 580216 674010 580272
rect 674066 580216 676292 580272
rect 674005 580214 676292 580216
rect 674005 580211 674071 580214
rect 674005 579866 674071 579869
rect 674005 579864 676292 579866
rect 674005 579808 674010 579864
rect 674066 579808 676292 579864
rect 674005 579806 676292 579808
rect 674005 579803 674071 579806
rect 44357 579730 44423 579733
rect 42198 579728 44423 579730
rect 42198 579672 44362 579728
rect 44418 579672 44423 579728
rect 42198 579670 44423 579672
rect 41965 578914 42031 578917
rect 41965 578912 42074 578914
rect 41965 578856 41970 578912
rect 42026 578856 42074 578912
rect 41965 578851 42074 578856
rect 42014 578234 42074 578851
rect 42198 578509 42258 579670
rect 44357 579667 44423 579670
rect 674005 579458 674071 579461
rect 674005 579456 676292 579458
rect 674005 579400 674010 579456
rect 674066 579400 676292 579456
rect 674005 579398 676292 579400
rect 674005 579395 674071 579398
rect 674005 579050 674071 579053
rect 674005 579048 676292 579050
rect 674005 578992 674010 579048
rect 674066 578992 676292 579048
rect 674005 578990 676292 578992
rect 674005 578987 674071 578990
rect 674005 578642 674071 578645
rect 674005 578640 676292 578642
rect 674005 578584 674010 578640
rect 674066 578584 676292 578640
rect 674005 578582 676292 578584
rect 674005 578579 674071 578582
rect 42198 578504 42307 578509
rect 42198 578448 42246 578504
rect 42302 578448 42307 578504
rect 42198 578446 42307 578448
rect 42241 578443 42307 578446
rect 46933 578234 46999 578237
rect 42014 578232 46999 578234
rect 42014 578176 46938 578232
rect 46994 578176 46999 578232
rect 42014 578174 46999 578176
rect 46933 578171 46999 578174
rect 674005 578234 674071 578237
rect 674005 578232 676292 578234
rect 674005 578176 674010 578232
rect 674066 578176 676292 578232
rect 674005 578174 676292 578176
rect 674005 578171 674071 578174
rect 40902 577764 40908 577828
rect 40972 577826 40978 577828
rect 41781 577826 41847 577829
rect 40972 577824 41847 577826
rect 40972 577768 41786 577824
rect 41842 577768 41847 577824
rect 40972 577766 41847 577768
rect 40972 577764 40978 577766
rect 41781 577763 41847 577766
rect 674005 577826 674071 577829
rect 674005 577824 676292 577826
rect 674005 577768 674010 577824
rect 674066 577768 676292 577824
rect 674005 577766 676292 577768
rect 674005 577763 674071 577766
rect 674005 577418 674071 577421
rect 674005 577416 676292 577418
rect 674005 577360 674010 577416
rect 674066 577360 676292 577416
rect 674005 577358 676292 577360
rect 674005 577355 674071 577358
rect 674005 577010 674071 577013
rect 674005 577008 676292 577010
rect 674005 576952 674010 577008
rect 674066 576952 676292 577008
rect 674005 576950 676292 576952
rect 674005 576947 674071 576950
rect 676806 576812 676812 576876
rect 676876 576812 676882 576876
rect 676814 576572 676874 576812
rect 682377 576466 682443 576469
rect 682334 576464 682443 576466
rect 682334 576408 682382 576464
rect 682438 576408 682443 576464
rect 682334 576403 682443 576408
rect 682334 576164 682394 576403
rect 684217 576058 684283 576061
rect 684174 576056 684283 576058
rect 684174 576000 684222 576056
rect 684278 576000 684283 576056
rect 684174 575995 684283 576000
rect 40718 575860 40724 575924
rect 40788 575922 40794 575924
rect 42241 575922 42307 575925
rect 40788 575920 42307 575922
rect 40788 575864 42246 575920
rect 42302 575864 42307 575920
rect 40788 575862 42307 575864
rect 40788 575860 40794 575862
rect 42241 575859 42307 575862
rect 684174 575756 684234 575995
rect 680997 575650 681063 575653
rect 680997 575648 681106 575650
rect 680997 575592 681002 575648
rect 681058 575592 681106 575648
rect 680997 575587 681106 575592
rect 40534 575452 40540 575516
rect 40604 575514 40610 575516
rect 42006 575514 42012 575516
rect 40604 575454 42012 575514
rect 40604 575452 40610 575454
rect 42006 575452 42012 575454
rect 42076 575452 42082 575516
rect 681046 575348 681106 575587
rect 674005 574970 674071 574973
rect 674005 574968 676292 574970
rect 674005 574912 674010 574968
rect 674066 574912 676292 574968
rect 674005 574910 676292 574912
rect 674005 574907 674071 574910
rect 62113 574834 62179 574837
rect 62113 574832 64706 574834
rect 62113 574776 62118 574832
rect 62174 574776 64706 574832
rect 62113 574774 64706 574776
rect 62113 574771 62179 574774
rect 64646 574194 64706 574774
rect 673545 574562 673611 574565
rect 673545 574560 676292 574562
rect 673545 574504 673550 574560
rect 673606 574504 676292 574560
rect 673545 574502 676292 574504
rect 673545 574499 673611 574502
rect 673545 574154 673611 574157
rect 673545 574152 676292 574154
rect 673545 574096 673550 574152
rect 673606 574096 676292 574152
rect 673545 574094 676292 574096
rect 673545 574091 673611 574094
rect 41965 573884 42031 573885
rect 41965 573880 42012 573884
rect 42076 573882 42082 573884
rect 41965 573824 41970 573880
rect 41965 573820 42012 573824
rect 42076 573822 42122 573882
rect 42076 573820 42082 573822
rect 41965 573819 42031 573820
rect 672809 573746 672875 573749
rect 672809 573744 676292 573746
rect 672809 573688 672814 573744
rect 672870 573688 676292 573744
rect 672809 573686 676292 573688
rect 672809 573683 672875 573686
rect 62113 573610 62179 573613
rect 62113 573608 64706 573610
rect 62113 573552 62118 573608
rect 62174 573552 64706 573608
rect 62113 573550 64706 573552
rect 62113 573547 62179 573550
rect 41454 573276 41460 573340
rect 41524 573338 41530 573340
rect 42609 573338 42675 573341
rect 41524 573336 42675 573338
rect 41524 573280 42614 573336
rect 42670 573280 42675 573336
rect 41524 573278 42675 573280
rect 41524 573276 41530 573278
rect 42609 573275 42675 573278
rect 64646 573012 64706 573550
rect 672993 573338 673059 573341
rect 672993 573336 676292 573338
rect 672993 573280 672998 573336
rect 673054 573280 676292 573336
rect 672993 573278 676292 573280
rect 672993 573275 673059 573278
rect 683389 573202 683455 573205
rect 683389 573200 683498 573202
rect 683389 573144 683394 573200
rect 683450 573144 683498 573200
rect 683389 573139 683498 573144
rect 683438 572900 683498 573139
rect 674005 572522 674071 572525
rect 674005 572520 676292 572522
rect 674005 572464 674010 572520
rect 674066 572464 676292 572520
rect 674005 572462 676292 572464
rect 674005 572459 674071 572462
rect 674005 572114 674071 572117
rect 674005 572112 676292 572114
rect 674005 572056 674010 572112
rect 674066 572056 676292 572112
rect 674005 572054 676292 572056
rect 674005 572051 674071 572054
rect 684033 571978 684099 571981
rect 683990 571976 684099 571978
rect 683990 571920 684038 571976
rect 684094 571920 684099 571976
rect 683990 571915 684099 571920
rect 41638 571508 41644 571572
rect 41708 571570 41714 571572
rect 42057 571570 42123 571573
rect 41708 571568 42123 571570
rect 41708 571512 42062 571568
rect 42118 571512 42123 571568
rect 41708 571510 42123 571512
rect 41708 571508 41714 571510
rect 42057 571507 42123 571510
rect 42425 571434 42491 571437
rect 64646 571434 64706 571830
rect 683990 571676 684050 571915
rect 676213 571570 676279 571573
rect 676213 571568 676322 571570
rect 676213 571512 676218 571568
rect 676274 571512 676322 571568
rect 676213 571507 676322 571512
rect 42425 571432 64706 571434
rect 42425 571376 42430 571432
rect 42486 571376 64706 571432
rect 42425 571374 64706 571376
rect 42425 571371 42491 571374
rect 676262 571268 676322 571507
rect 63309 571162 63375 571165
rect 63309 571160 64706 571162
rect 63309 571104 63314 571160
rect 63370 571104 64706 571160
rect 63309 571102 64706 571104
rect 63309 571099 63375 571102
rect 64646 570648 64706 571102
rect 674005 570890 674071 570893
rect 674005 570888 676292 570890
rect 674005 570832 674010 570888
rect 674066 570832 676292 570888
rect 674005 570830 676292 570832
rect 674005 570827 674071 570830
rect 673545 570482 673611 570485
rect 674833 570482 674899 570485
rect 673545 570480 674899 570482
rect 673545 570424 673550 570480
rect 673606 570424 674838 570480
rect 674894 570424 674899 570480
rect 673545 570422 674899 570424
rect 673545 570419 673611 570422
rect 674833 570419 674899 570422
rect 682886 570346 682946 570452
rect 683113 570346 683179 570349
rect 682886 570344 683179 570346
rect 682886 570288 683118 570344
rect 683174 570288 683179 570344
rect 682886 570286 683179 570288
rect 41781 570212 41847 570213
rect 41781 570208 41828 570212
rect 41892 570210 41898 570212
rect 41781 570152 41786 570208
rect 41781 570148 41828 570152
rect 41892 570150 41938 570210
rect 41892 570148 41898 570150
rect 41781 570147 41847 570148
rect 682886 570044 682946 570286
rect 683113 570283 683179 570286
rect 62481 569938 62547 569941
rect 62481 569936 64706 569938
rect 62481 569880 62486 569936
rect 62542 569880 64706 569936
rect 62481 569878 64706 569880
rect 62481 569875 62547 569878
rect 64646 569466 64706 569878
rect 674005 569666 674071 569669
rect 674005 569664 676292 569666
rect 674005 569608 674010 569664
rect 674066 569608 676292 569664
rect 674005 569606 676292 569608
rect 674005 569603 674071 569606
rect 63125 568578 63191 568581
rect 63125 568576 64706 568578
rect 63125 568520 63130 568576
rect 63186 568520 64706 568576
rect 63125 568518 64706 568520
rect 63125 568515 63191 568518
rect 64646 568284 64706 568518
rect 673545 565858 673611 565861
rect 675385 565858 675451 565861
rect 673545 565856 675451 565858
rect 673545 565800 673550 565856
rect 673606 565800 675390 565856
rect 675446 565800 675451 565856
rect 673545 565798 675451 565800
rect 673545 565795 673611 565798
rect 675385 565795 675451 565798
rect 673545 564498 673611 564501
rect 675109 564498 675175 564501
rect 673545 564496 675175 564498
rect 673545 564440 673550 564496
rect 673606 564440 675114 564496
rect 675170 564440 675175 564496
rect 673545 564438 675175 564440
rect 673545 564435 673611 564438
rect 675109 564435 675175 564438
rect 668577 562322 668643 562325
rect 675109 562322 675175 562325
rect 668577 562320 675175 562322
rect 668577 562264 668582 562320
rect 668638 562264 675114 562320
rect 675170 562264 675175 562320
rect 668577 562262 675175 562264
rect 668577 562259 668643 562262
rect 675109 562259 675175 562262
rect 675385 561916 675451 561917
rect 675334 561914 675340 561916
rect 675294 561854 675340 561914
rect 675404 561912 675451 561916
rect 675446 561856 675451 561912
rect 675334 561852 675340 561854
rect 675404 561852 675451 561856
rect 675385 561851 675451 561852
rect 673085 560146 673151 560149
rect 673085 560144 675586 560146
rect 673085 560088 673090 560144
rect 673146 560088 675586 560144
rect 673085 560086 675586 560088
rect 673085 560083 673151 560086
rect 671797 559738 671863 559741
rect 675293 559738 675359 559741
rect 671797 559736 675359 559738
rect 671797 559680 671802 559736
rect 671858 559680 675298 559736
rect 675354 559680 675359 559736
rect 671797 559678 675359 559680
rect 671797 559675 671863 559678
rect 675293 559675 675359 559678
rect 675526 559469 675586 560086
rect 675477 559464 675586 559469
rect 675477 559408 675482 559464
rect 675538 559408 675586 559464
rect 675477 559406 675586 559408
rect 675477 559403 675543 559406
rect 41270 559268 41276 559332
rect 41340 559330 41346 559332
rect 44633 559330 44699 559333
rect 41340 559328 44699 559330
rect 41340 559272 44638 559328
rect 44694 559272 44699 559328
rect 41340 559270 44699 559272
rect 41340 559268 41346 559270
rect 44633 559267 44699 559270
rect 39849 559058 39915 559061
rect 42793 559058 42859 559061
rect 39849 559056 42859 559058
rect 39849 559000 39854 559056
rect 39910 559000 42798 559056
rect 42854 559000 42859 559056
rect 39849 558998 42859 559000
rect 39849 558995 39915 558998
rect 42793 558995 42859 558998
rect 40493 558786 40559 558789
rect 43069 558786 43135 558789
rect 40493 558784 43135 558786
rect 40493 558728 40498 558784
rect 40554 558728 43074 558784
rect 43130 558728 43135 558784
rect 40493 558726 43135 558728
rect 40493 558723 40559 558726
rect 43069 558723 43135 558726
rect 47577 558514 47643 558517
rect 41492 558512 47643 558514
rect 41492 558456 47582 558512
rect 47638 558456 47643 558512
rect 41492 558454 47643 558456
rect 47577 558451 47643 558454
rect 674097 558378 674163 558381
rect 675477 558378 675543 558381
rect 674097 558376 675543 558378
rect 674097 558320 674102 558376
rect 674158 558320 675482 558376
rect 675538 558320 675543 558376
rect 674097 558318 675543 558320
rect 674097 558315 674163 558318
rect 675477 558315 675543 558318
rect 35801 558106 35867 558109
rect 35788 558104 35867 558106
rect 35788 558048 35806 558104
rect 35862 558048 35867 558104
rect 35788 558046 35867 558048
rect 35801 558043 35867 558046
rect 38518 557550 38578 557668
rect 38702 557638 48330 557698
rect 38702 557550 38762 557638
rect 38518 557490 38762 557550
rect 41270 557488 41276 557552
rect 41340 557488 41346 557552
rect 41278 557260 41338 557488
rect 48270 557426 48330 557638
rect 675293 557562 675359 557565
rect 676254 557562 676260 557564
rect 675293 557560 676260 557562
rect 675293 557504 675298 557560
rect 675354 557504 676260 557560
rect 675293 557502 676260 557504
rect 675293 557499 675359 557502
rect 676254 557500 676260 557502
rect 676324 557500 676330 557564
rect 48270 557366 51090 557426
rect 44541 556882 44607 556885
rect 41492 556880 44607 556882
rect 41492 556824 44546 556880
rect 44602 556824 44607 556880
rect 41492 556822 44607 556824
rect 44541 556819 44607 556822
rect 51030 556746 51090 557366
rect 62481 556746 62547 556749
rect 51030 556744 62547 556746
rect 51030 556688 62486 556744
rect 62542 556688 62547 556744
rect 51030 556686 62547 556688
rect 62481 556683 62547 556686
rect 44909 556474 44975 556477
rect 41492 556472 44975 556474
rect 41492 556416 44914 556472
rect 44970 556416 44975 556472
rect 41492 556414 44975 556416
rect 44909 556411 44975 556414
rect 45001 556066 45067 556069
rect 41492 556064 45067 556066
rect 41492 556008 45006 556064
rect 45062 556008 45067 556064
rect 41492 556006 45067 556008
rect 45001 556003 45067 556006
rect 35801 555658 35867 555661
rect 35788 555656 35867 555658
rect 35788 555600 35806 555656
rect 35862 555600 35867 555656
rect 35788 555598 35867 555600
rect 35801 555595 35867 555598
rect 44357 555250 44423 555253
rect 41492 555248 44423 555250
rect 41492 555192 44362 555248
rect 44418 555192 44423 555248
rect 41492 555190 44423 555192
rect 44357 555187 44423 555190
rect 672901 555250 672967 555253
rect 675385 555250 675451 555253
rect 672901 555248 675451 555250
rect 672901 555192 672906 555248
rect 672962 555192 675390 555248
rect 675446 555192 675451 555248
rect 672901 555190 675451 555192
rect 672901 555187 672967 555190
rect 675385 555187 675451 555190
rect 35801 554842 35867 554845
rect 35788 554840 35867 554842
rect 35788 554784 35806 554840
rect 35862 554784 35867 554840
rect 35788 554782 35867 554784
rect 35801 554779 35867 554782
rect 673545 554842 673611 554845
rect 675293 554842 675359 554845
rect 673545 554840 675359 554842
rect 673545 554784 673550 554840
rect 673606 554784 675298 554840
rect 675354 554784 675359 554840
rect 673545 554782 675359 554784
rect 673545 554779 673611 554782
rect 675293 554779 675359 554782
rect 35617 554434 35683 554437
rect 35604 554432 35683 554434
rect 35604 554376 35622 554432
rect 35678 554376 35683 554432
rect 35604 554374 35683 554376
rect 35617 554371 35683 554374
rect 41822 554026 41828 554028
rect 41492 553966 41828 554026
rect 41822 553964 41828 553966
rect 41892 553964 41898 554028
rect 35801 553618 35867 553621
rect 35788 553616 35867 553618
rect 35788 553560 35806 553616
rect 35862 553560 35867 553616
rect 35788 553558 35867 553560
rect 35801 553555 35867 553558
rect 649950 553482 650010 553914
rect 675753 553890 675819 553893
rect 676806 553890 676812 553892
rect 675753 553888 676812 553890
rect 675753 553832 675758 553888
rect 675814 553832 676812 553888
rect 675753 553830 676812 553832
rect 675753 553827 675819 553830
rect 676806 553828 676812 553830
rect 676876 553828 676882 553892
rect 651465 553482 651531 553485
rect 675569 553482 675635 553485
rect 649950 553480 651531 553482
rect 649950 553424 651470 553480
rect 651526 553424 651531 553480
rect 649950 553422 651531 553424
rect 651465 553419 651531 553422
rect 675526 553480 675635 553482
rect 675526 553424 675574 553480
rect 675630 553424 675635 553480
rect 675526 553419 675635 553424
rect 37917 553410 37983 553413
rect 37917 553408 38026 553410
rect 37917 553352 37922 553408
rect 37978 553352 38026 553408
rect 37917 553347 38026 553352
rect 37966 553180 38026 553347
rect 673545 553210 673611 553213
rect 675526 553210 675586 553419
rect 673545 553208 675586 553210
rect 673545 553152 673550 553208
rect 673606 553152 675586 553208
rect 673545 553150 675586 553152
rect 673545 553147 673611 553150
rect 41689 553074 41755 553077
rect 43161 553074 43227 553077
rect 41689 553072 43227 553074
rect 41689 553016 41694 553072
rect 41750 553016 43166 553072
rect 43222 553016 43227 553072
rect 41689 553014 43227 553016
rect 41689 553011 41755 553014
rect 43161 553011 43227 553014
rect 41822 552802 41828 552804
rect 41492 552742 41828 552802
rect 41822 552740 41828 552742
rect 41892 552740 41898 552804
rect 41321 552394 41387 552397
rect 41308 552392 41387 552394
rect 41308 552336 41326 552392
rect 41382 552336 41387 552392
rect 41308 552334 41387 552336
rect 41321 552331 41387 552334
rect 649950 552122 650010 552732
rect 651649 552122 651715 552125
rect 649950 552120 651715 552122
rect 649950 552064 651654 552120
rect 651710 552064 651715 552120
rect 649950 552062 651715 552064
rect 651649 552059 651715 552062
rect 674465 552122 674531 552125
rect 675385 552122 675451 552125
rect 674465 552120 675451 552122
rect 674465 552064 674470 552120
rect 674526 552064 675390 552120
rect 675446 552064 675451 552120
rect 674465 552062 675451 552064
rect 674465 552059 674531 552062
rect 675385 552059 675451 552062
rect 29637 551986 29703 551989
rect 29637 551984 29716 551986
rect 29637 551928 29642 551984
rect 29698 551928 29716 551984
rect 29637 551926 29716 551928
rect 29637 551923 29703 551926
rect 41689 551850 41755 551853
rect 43989 551850 44055 551853
rect 41689 551848 44055 551850
rect 41689 551792 41694 551848
rect 41750 551792 43994 551848
rect 44050 551792 44055 551848
rect 41689 551790 44055 551792
rect 41689 551787 41755 551790
rect 43989 551787 44055 551790
rect 45185 551578 45251 551581
rect 41492 551576 45251 551578
rect 41492 551520 45190 551576
rect 45246 551520 45251 551576
rect 670417 551578 670483 551581
rect 675385 551578 675451 551581
rect 670417 551576 675451 551578
rect 41492 551518 45251 551520
rect 45185 551515 45251 551518
rect 41137 551170 41203 551173
rect 41124 551168 41203 551170
rect 41124 551112 41142 551168
rect 41198 551112 41203 551168
rect 41124 551110 41203 551112
rect 649950 551170 650010 551550
rect 670417 551520 670422 551576
rect 670478 551520 675390 551576
rect 675446 551520 675451 551576
rect 670417 551518 675451 551520
rect 670417 551515 670483 551518
rect 675385 551515 675451 551518
rect 651465 551170 651531 551173
rect 649950 551168 651531 551170
rect 649950 551112 651470 551168
rect 651526 551112 651531 551168
rect 649950 551110 651531 551112
rect 41137 551107 41203 551110
rect 651465 551107 651531 551110
rect 43805 550762 43871 550765
rect 41492 550760 43871 550762
rect 41492 550704 43810 550760
rect 43866 550704 43871 550760
rect 41492 550702 43871 550704
rect 43805 550699 43871 550702
rect 45369 550490 45435 550493
rect 41784 550488 45435 550490
rect 41784 550432 45374 550488
rect 45430 550432 45435 550488
rect 41784 550430 45435 550432
rect 41784 550354 41844 550430
rect 45369 550427 45435 550430
rect 41492 550294 41844 550354
rect 649950 550354 650010 550368
rect 651373 550354 651439 550357
rect 649950 550352 651439 550354
rect 649950 550296 651378 550352
rect 651434 550296 651439 550352
rect 649950 550294 651439 550296
rect 651373 550291 651439 550294
rect 42057 550218 42123 550221
rect 63309 550218 63375 550221
rect 42057 550216 63375 550218
rect 42057 550160 42062 550216
rect 42118 550160 63314 550216
rect 63370 550160 63375 550216
rect 42057 550158 63375 550160
rect 42057 550155 42123 550158
rect 63309 550155 63375 550158
rect 41781 549946 41847 549949
rect 41492 549944 41847 549946
rect 41492 549888 41786 549944
rect 41842 549888 41847 549944
rect 41492 549886 41847 549888
rect 41781 549883 41847 549886
rect 670417 549674 670483 549677
rect 675477 549674 675543 549677
rect 670417 549672 675543 549674
rect 670417 549616 670422 549672
rect 670478 549616 675482 549672
rect 675538 549616 675543 549672
rect 670417 549614 675543 549616
rect 670417 549611 670483 549614
rect 675477 549611 675543 549614
rect 40493 549538 40559 549541
rect 40493 549536 40572 549538
rect 40493 549480 40498 549536
rect 40554 549480 40572 549536
rect 40493 549478 40572 549480
rect 40493 549475 40559 549478
rect 651465 549266 651531 549269
rect 649950 549264 651531 549266
rect 649950 549208 651470 549264
rect 651526 549208 651531 549264
rect 649950 549206 651531 549208
rect 649950 549186 650010 549206
rect 651465 549203 651531 549206
rect 42793 549130 42859 549133
rect 41492 549128 42859 549130
rect 41492 549072 42798 549128
rect 42854 549072 42859 549128
rect 41492 549070 42859 549072
rect 42793 549067 42859 549070
rect 44173 548722 44239 548725
rect 41492 548720 44239 548722
rect 41492 548664 44178 548720
rect 44234 548664 44239 548720
rect 41492 548662 44239 548664
rect 44173 548659 44239 548662
rect 651465 548450 651531 548453
rect 649950 548448 651531 548450
rect 649950 548392 651470 548448
rect 651526 548392 651531 548448
rect 649950 548390 651531 548392
rect 41321 548314 41387 548317
rect 41308 548312 41387 548314
rect 41308 548256 41326 548312
rect 41382 548256 41387 548312
rect 41308 548254 41387 548256
rect 41321 548251 41387 548254
rect 649950 548004 650010 548390
rect 651465 548387 651531 548390
rect 675753 548314 675819 548317
rect 676990 548314 676996 548316
rect 675753 548312 676996 548314
rect 675753 548256 675758 548312
rect 675814 548256 676996 548312
rect 675753 548254 676996 548256
rect 675753 548251 675819 548254
rect 676990 548252 676996 548254
rect 677060 548252 677066 548316
rect 41689 547770 41755 547773
rect 43621 547770 43687 547773
rect 41689 547768 43687 547770
rect 41689 547712 41694 547768
rect 41750 547712 43626 547768
rect 43682 547712 43687 547768
rect 41689 547710 43687 547712
rect 41689 547707 41755 547710
rect 43621 547707 43687 547710
rect 676254 547572 676260 547636
rect 676324 547634 676330 547636
rect 677409 547634 677475 547637
rect 676324 547632 677475 547634
rect 676324 547576 677414 547632
rect 677470 547576 677475 547632
rect 676324 547574 677475 547576
rect 676324 547572 676330 547574
rect 677409 547571 677475 547574
rect 39205 547498 39271 547501
rect 39205 547496 39284 547498
rect 39205 547440 39210 547496
rect 39266 547440 39284 547496
rect 39205 547438 39284 547440
rect 39205 547435 39271 547438
rect 673913 547362 673979 547365
rect 675569 547362 675635 547365
rect 673913 547360 675635 547362
rect 673913 547304 673918 547360
rect 673974 547304 675574 547360
rect 675630 547304 675635 547360
rect 673913 547302 675635 547304
rect 673913 547299 673979 547302
rect 675569 547299 675635 547302
rect 674414 547028 674420 547092
rect 674484 547090 674490 547092
rect 683389 547090 683455 547093
rect 674484 547088 683455 547090
rect 674484 547032 683394 547088
rect 683450 547032 683455 547088
rect 674484 547030 683455 547032
rect 674484 547028 674490 547030
rect 683389 547027 683455 547030
rect 676070 546756 676076 546820
rect 676140 546818 676146 546820
rect 680997 546818 681063 546821
rect 676140 546816 681063 546818
rect 676140 546760 681002 546816
rect 681058 546760 681063 546816
rect 676140 546758 681063 546760
rect 676140 546756 676146 546758
rect 680997 546755 681063 546758
rect 674925 545730 674991 545733
rect 675334 545730 675340 545732
rect 674925 545728 675340 545730
rect 674925 545672 674930 545728
rect 674986 545672 675340 545728
rect 674925 545670 675340 545672
rect 674925 545667 674991 545670
rect 675334 545668 675340 545670
rect 675404 545668 675410 545732
rect 40718 545532 40724 545596
rect 40788 545594 40794 545596
rect 41505 545594 41571 545597
rect 40788 545592 41571 545594
rect 40788 545536 41510 545592
rect 41566 545536 41571 545592
rect 40788 545534 41571 545536
rect 40788 545532 40794 545534
rect 41505 545531 41571 545534
rect 40493 545324 40559 545325
rect 40493 545320 40540 545324
rect 40604 545322 40610 545324
rect 40493 545264 40498 545320
rect 40493 545260 40540 545264
rect 40604 545262 40650 545322
rect 40604 545260 40610 545262
rect 40493 545259 40559 545260
rect 39205 543690 39271 543693
rect 44766 543690 44772 543692
rect 39205 543688 44772 543690
rect 39205 543632 39210 543688
rect 39266 543632 44772 543688
rect 39205 543630 44772 543632
rect 39205 543627 39271 543630
rect 44766 543628 44772 543630
rect 44836 543628 44842 543692
rect 37917 542330 37983 542333
rect 41822 542330 41828 542332
rect 37917 542328 41828 542330
rect 37917 542272 37922 542328
rect 37978 542272 41828 542328
rect 37917 542270 41828 542272
rect 37917 542267 37983 542270
rect 41822 542268 41828 542270
rect 41892 542268 41898 542332
rect 42609 539610 42675 539613
rect 45369 539610 45435 539613
rect 42609 539608 45435 539610
rect 42609 539552 42614 539608
rect 42670 539552 45374 539608
rect 45430 539552 45435 539608
rect 42609 539550 45435 539552
rect 42609 539547 42675 539550
rect 45369 539547 45435 539550
rect 42425 538250 42491 538253
rect 51717 538250 51783 538253
rect 42425 538248 51783 538250
rect 42425 538192 42430 538248
rect 42486 538192 51722 538248
rect 51778 538192 51783 538248
rect 42425 538190 51783 538192
rect 42425 538187 42491 538190
rect 51717 538187 51783 538190
rect 42057 537434 42123 537437
rect 44725 537434 44791 537437
rect 42057 537432 44791 537434
rect 42057 537376 42062 537432
rect 42118 537376 44730 537432
rect 44786 537376 44791 537432
rect 42057 537374 44791 537376
rect 42057 537371 42123 537374
rect 44725 537371 44791 537374
rect 42057 537026 42123 537029
rect 42609 537026 42675 537029
rect 42057 537024 42675 537026
rect 42057 536968 42062 537024
rect 42118 536968 42614 537024
rect 42670 536968 42675 537024
rect 42057 536966 42675 536968
rect 42057 536963 42123 536966
rect 42609 536963 42675 536966
rect 44173 536890 44239 536893
rect 42750 536888 44239 536890
rect 42750 536832 44178 536888
rect 44234 536832 44239 536888
rect 42750 536830 44239 536832
rect 42750 536757 42810 536830
rect 44173 536827 44239 536830
rect 42701 536752 42810 536757
rect 42701 536696 42706 536752
rect 42762 536696 42810 536752
rect 42701 536694 42810 536696
rect 42701 536691 42767 536694
rect 676262 535941 676322 536112
rect 676213 535936 676322 535941
rect 676213 535880 676218 535936
rect 676274 535880 676322 535936
rect 676213 535878 676322 535880
rect 676213 535875 676279 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 42057 535666 42123 535669
rect 42701 535666 42767 535669
rect 42057 535664 42767 535666
rect 42057 535608 42062 535664
rect 42118 535608 42706 535664
rect 42762 535608 42767 535664
rect 42057 535606 42767 535608
rect 42057 535603 42123 535606
rect 42701 535603 42767 535606
rect 40718 535196 40724 535260
rect 40788 535258 40794 535260
rect 41781 535258 41847 535261
rect 40788 535256 41847 535258
rect 40788 535200 41786 535256
rect 41842 535200 41847 535256
rect 40788 535198 41847 535200
rect 40788 535196 40794 535198
rect 41781 535195 41847 535198
rect 676262 535125 676322 535296
rect 676213 535120 676322 535125
rect 676213 535064 676218 535120
rect 676274 535064 676322 535120
rect 676213 535062 676322 535064
rect 676213 535059 676279 535062
rect 676029 534918 676095 534921
rect 676029 534916 676292 534918
rect 676029 534860 676034 534916
rect 676090 534860 676292 534916
rect 676029 534858 676292 534860
rect 676029 534855 676095 534858
rect 676029 534510 676095 534513
rect 676029 534508 676292 534510
rect 676029 534452 676034 534508
rect 676090 534452 676292 534508
rect 676029 534450 676292 534452
rect 676029 534447 676095 534450
rect 676029 534102 676095 534105
rect 676029 534100 676292 534102
rect 676029 534044 676034 534100
rect 676090 534044 676292 534100
rect 676029 534042 676292 534044
rect 676029 534039 676095 534042
rect 42425 533898 42491 533901
rect 43989 533898 44055 533901
rect 42425 533896 44055 533898
rect 42425 533840 42430 533896
rect 42486 533840 43994 533896
rect 44050 533840 44055 533896
rect 42425 533838 44055 533840
rect 42425 533835 42491 533838
rect 43989 533835 44055 533838
rect 42701 533626 42767 533629
rect 43805 533626 43871 533629
rect 42701 533624 43871 533626
rect 42701 533568 42706 533624
rect 42762 533568 43810 533624
rect 43866 533568 43871 533624
rect 42701 533566 43871 533568
rect 42701 533563 42767 533566
rect 43805 533563 43871 533566
rect 676446 533493 676506 533664
rect 676397 533488 676506 533493
rect 676397 533432 676402 533488
rect 676458 533432 676506 533488
rect 676397 533430 676506 533432
rect 676397 533427 676463 533430
rect 40534 533292 40540 533356
rect 40604 533354 40610 533356
rect 42241 533354 42307 533357
rect 40604 533352 42307 533354
rect 40604 533296 42246 533352
rect 42302 533296 42307 533352
rect 40604 533294 42307 533296
rect 40604 533292 40610 533294
rect 42241 533291 42307 533294
rect 676029 533286 676095 533289
rect 676029 533284 676292 533286
rect 676029 533228 676034 533284
rect 676090 533228 676292 533284
rect 676029 533226 676292 533228
rect 676029 533223 676095 533226
rect 676213 533082 676279 533085
rect 676213 533080 676322 533082
rect 676213 533024 676218 533080
rect 676274 533024 676322 533080
rect 676213 533019 676322 533024
rect 676262 532848 676322 533019
rect 41638 532612 41644 532676
rect 41708 532674 41714 532676
rect 42517 532674 42583 532677
rect 41708 532672 42583 532674
rect 41708 532616 42522 532672
rect 42578 532616 42583 532672
rect 41708 532614 42583 532616
rect 41708 532612 41714 532614
rect 42517 532611 42583 532614
rect 676262 532269 676322 532440
rect 676213 532264 676322 532269
rect 676213 532208 676218 532264
rect 676274 532208 676322 532264
rect 676213 532206 676322 532208
rect 676213 532203 676279 532206
rect 676029 532062 676095 532065
rect 676029 532060 676292 532062
rect 676029 532004 676034 532060
rect 676090 532004 676292 532060
rect 676029 532002 676292 532004
rect 676029 531999 676095 532002
rect 676397 531858 676463 531861
rect 676397 531856 676506 531858
rect 676397 531800 676402 531856
rect 676458 531800 676506 531856
rect 676397 531795 676506 531800
rect 676446 531624 676506 531795
rect 682377 531450 682443 531453
rect 682334 531448 682443 531450
rect 682334 531392 682382 531448
rect 682438 531392 682443 531448
rect 682334 531387 682443 531392
rect 682334 531216 682394 531387
rect 62113 531178 62179 531181
rect 62113 531176 64706 531178
rect 62113 531120 62118 531176
rect 62174 531120 64706 531176
rect 62113 531118 64706 531120
rect 62113 531115 62179 531118
rect 62297 530634 62363 530637
rect 676262 530634 676322 530808
rect 62297 530632 64706 530634
rect 62297 530576 62302 530632
rect 62358 530576 64706 530632
rect 62297 530574 64706 530576
rect 62297 530571 62363 530574
rect 41454 530028 41460 530092
rect 41524 530090 41530 530092
rect 42609 530090 42675 530093
rect 41524 530088 42675 530090
rect 41524 530032 42614 530088
rect 42670 530032 42675 530088
rect 41524 530030 42675 530032
rect 41524 530028 41530 530030
rect 42609 530027 42675 530030
rect 64646 529990 64706 530574
rect 675710 530574 676322 530634
rect 680997 530634 681063 530637
rect 680997 530632 681106 530634
rect 680997 530576 681002 530632
rect 681058 530576 681106 530632
rect 673269 530090 673335 530093
rect 675710 530090 675770 530574
rect 680997 530571 681106 530576
rect 681046 530400 681106 530571
rect 673269 530088 675770 530090
rect 673269 530032 673274 530088
rect 673330 530032 675770 530088
rect 673269 530030 675770 530032
rect 673269 530027 673335 530030
rect 676029 530022 676095 530025
rect 676029 530020 676292 530022
rect 676029 529964 676034 530020
rect 676090 529964 676292 530020
rect 676029 529962 676292 529964
rect 676029 529959 676095 529962
rect 676262 529413 676322 529584
rect 676213 529408 676322 529413
rect 676213 529352 676218 529408
rect 676274 529352 676322 529408
rect 676213 529350 676322 529352
rect 676213 529347 676279 529350
rect 676262 529005 676322 529176
rect 42701 529002 42767 529005
rect 45185 529002 45251 529005
rect 42701 529000 45251 529002
rect 42701 528944 42706 529000
rect 42762 528944 45190 529000
rect 45246 528944 45251 529000
rect 42701 528942 45251 528944
rect 42701 528939 42767 528942
rect 45185 528939 45251 528942
rect 676213 529000 676322 529005
rect 676213 528944 676218 529000
rect 676274 528944 676322 529000
rect 676213 528942 676322 528944
rect 676213 528939 676279 528942
rect 41822 528668 41828 528732
rect 41892 528730 41898 528732
rect 42701 528730 42767 528733
rect 41892 528728 42767 528730
rect 41892 528672 42706 528728
rect 42762 528672 42767 528728
rect 41892 528670 42767 528672
rect 41892 528668 41898 528670
rect 42701 528667 42767 528670
rect 62113 528594 62179 528597
rect 64646 528594 64706 528808
rect 676029 528798 676095 528801
rect 676029 528796 676292 528798
rect 676029 528740 676034 528796
rect 676090 528740 676292 528796
rect 676029 528738 676292 528740
rect 676029 528735 676095 528738
rect 62113 528592 64706 528594
rect 62113 528536 62118 528592
rect 62174 528536 64706 528592
rect 62113 528534 64706 528536
rect 683573 528594 683639 528597
rect 683573 528592 683682 528594
rect 683573 528536 683578 528592
rect 683634 528536 683682 528592
rect 62113 528531 62179 528534
rect 683573 528531 683682 528536
rect 683622 528360 683682 528531
rect 62481 528050 62547 528053
rect 62481 528048 64706 528050
rect 62481 527992 62486 528048
rect 62542 527992 64706 528048
rect 62481 527990 64706 527992
rect 62481 527987 62547 527990
rect 64646 527626 64706 527990
rect 673361 527778 673427 527781
rect 676262 527778 676322 527952
rect 673361 527776 676322 527778
rect 673361 527720 673366 527776
rect 673422 527720 676322 527776
rect 673361 527718 676322 527720
rect 683205 527778 683271 527781
rect 683205 527776 683314 527778
rect 683205 527720 683210 527776
rect 683266 527720 683314 527776
rect 673361 527715 673427 527718
rect 683205 527715 683314 527720
rect 683254 527544 683314 527715
rect 683389 527370 683455 527373
rect 683389 527368 683498 527370
rect 683389 527312 683394 527368
rect 683450 527312 683498 527368
rect 683389 527307 683498 527312
rect 42885 527234 42951 527237
rect 44817 527234 44883 527237
rect 42885 527232 44883 527234
rect 42885 527176 42890 527232
rect 42946 527176 44822 527232
rect 44878 527176 44883 527232
rect 42885 527174 44883 527176
rect 42885 527171 42951 527174
rect 44817 527171 44883 527174
rect 683438 527136 683498 527307
rect 62113 527098 62179 527101
rect 62113 527096 64706 527098
rect 62113 527040 62118 527096
rect 62174 527040 64706 527096
rect 62113 527038 64706 527040
rect 62113 527035 62179 527038
rect 64646 526444 64706 527038
rect 676029 526758 676095 526761
rect 676029 526756 676292 526758
rect 676029 526700 676034 526756
rect 676090 526700 676292 526756
rect 676029 526698 676292 526700
rect 676029 526695 676095 526698
rect 676029 526350 676095 526353
rect 676029 526348 676292 526350
rect 676029 526292 676034 526348
rect 676090 526292 676292 526348
rect 676029 526290 676292 526292
rect 676029 526287 676095 526290
rect 677918 525741 677978 525912
rect 63309 525738 63375 525741
rect 63309 525736 64706 525738
rect 63309 525680 63314 525736
rect 63370 525680 64706 525736
rect 63309 525678 64706 525680
rect 63309 525675 63375 525678
rect 64646 525262 64706 525678
rect 677869 525736 677978 525741
rect 677869 525680 677874 525736
rect 677930 525680 677978 525736
rect 677869 525678 677978 525680
rect 677869 525675 677935 525678
rect 683070 524925 683130 525504
rect 683070 524920 683179 524925
rect 683070 524864 683118 524920
rect 683174 524864 683179 524920
rect 683070 524862 683179 524864
rect 683113 524859 683179 524862
rect 679022 524517 679082 524688
rect 678973 524512 679082 524517
rect 678973 524456 678978 524512
rect 679034 524456 679082 524512
rect 678973 524454 679082 524456
rect 678973 524451 679039 524454
rect 676990 503644 676996 503708
rect 677060 503706 677066 503708
rect 683389 503706 683455 503709
rect 677060 503704 683455 503706
rect 677060 503648 683394 503704
rect 683450 503648 683455 503704
rect 677060 503646 683455 503648
rect 677060 503644 677066 503646
rect 683389 503643 683455 503646
rect 676806 500924 676812 500988
rect 676876 500986 676882 500988
rect 683205 500986 683271 500989
rect 676876 500984 683271 500986
rect 676876 500928 683210 500984
rect 683266 500928 683271 500984
rect 676876 500926 683271 500928
rect 676876 500924 676882 500926
rect 683205 500923 683271 500926
rect 673821 492146 673887 492149
rect 673821 492144 676292 492146
rect 673821 492088 673826 492144
rect 673882 492088 676292 492144
rect 673821 492086 676292 492088
rect 673821 492083 673887 492086
rect 676029 491738 676095 491741
rect 676029 491736 676292 491738
rect 676029 491680 676034 491736
rect 676090 491680 676292 491736
rect 676029 491678 676292 491680
rect 676029 491675 676095 491678
rect 674005 491330 674071 491333
rect 674005 491328 676292 491330
rect 674005 491272 674010 491328
rect 674066 491272 676292 491328
rect 674005 491270 676292 491272
rect 674005 491267 674071 491270
rect 674005 490922 674071 490925
rect 674005 490920 676292 490922
rect 674005 490864 674010 490920
rect 674066 490864 676292 490920
rect 674005 490862 676292 490864
rect 674005 490859 674071 490862
rect 673361 490514 673427 490517
rect 673361 490512 676292 490514
rect 673361 490456 673366 490512
rect 673422 490456 676292 490512
rect 673361 490454 676292 490456
rect 673361 490451 673427 490454
rect 672717 490106 672783 490109
rect 672717 490104 676292 490106
rect 672717 490048 672722 490104
rect 672778 490048 676292 490104
rect 672717 490046 676292 490048
rect 672717 490043 672783 490046
rect 44766 489908 44772 489972
rect 44836 489970 44842 489972
rect 47577 489970 47643 489973
rect 44836 489968 47643 489970
rect 44836 489912 47582 489968
rect 47638 489912 47643 489968
rect 44836 489910 47643 489912
rect 44836 489908 44842 489910
rect 47577 489907 47643 489910
rect 674005 489698 674071 489701
rect 674005 489696 676292 489698
rect 674005 489640 674010 489696
rect 674066 489640 676292 489696
rect 674005 489638 676292 489640
rect 674005 489635 674071 489638
rect 674005 489290 674071 489293
rect 674005 489288 676292 489290
rect 674005 489232 674010 489288
rect 674066 489232 676292 489288
rect 674005 489230 676292 489232
rect 674005 489227 674071 489230
rect 676024 488820 676030 488884
rect 676094 488882 676100 488884
rect 676094 488822 676292 488882
rect 676094 488820 676100 488822
rect 674005 488474 674071 488477
rect 674005 488472 676292 488474
rect 674005 488416 674010 488472
rect 674066 488416 676292 488472
rect 674005 488414 676292 488416
rect 674005 488411 674071 488414
rect 676170 488006 676292 488066
rect 675886 487868 675892 487932
rect 675956 487930 675962 487932
rect 676170 487930 676230 488006
rect 675956 487870 676230 487930
rect 675956 487868 675962 487870
rect 681181 487658 681247 487661
rect 681181 487656 681260 487658
rect 681181 487600 681186 487656
rect 681242 487600 681260 487656
rect 681181 487598 681260 487600
rect 681181 487595 681247 487598
rect 679617 487250 679683 487253
rect 679604 487248 679683 487250
rect 679604 487192 679622 487248
rect 679678 487192 679683 487248
rect 679604 487190 679683 487192
rect 679617 487187 679683 487190
rect 676029 486842 676095 486845
rect 676029 486840 676292 486842
rect 676029 486784 676034 486840
rect 676090 486784 676292 486840
rect 676029 486782 676292 486784
rect 676029 486779 676095 486782
rect 680997 486434 681063 486437
rect 680997 486432 681076 486434
rect 680997 486376 681002 486432
rect 681058 486376 681076 486432
rect 680997 486374 681076 486376
rect 680997 486371 681063 486374
rect 672901 486026 672967 486029
rect 672901 486024 676292 486026
rect 672901 485968 672906 486024
rect 672962 485968 676292 486024
rect 672901 485966 676292 485968
rect 672901 485963 672967 485966
rect 683389 485618 683455 485621
rect 683389 485616 683468 485618
rect 683389 485560 683394 485616
rect 683450 485560 683468 485616
rect 683389 485558 683468 485560
rect 683389 485555 683455 485558
rect 676029 485210 676095 485213
rect 676029 485208 676292 485210
rect 676029 485152 676034 485208
rect 676090 485152 676292 485208
rect 676029 485150 676292 485152
rect 676029 485147 676095 485150
rect 673085 484802 673151 484805
rect 673085 484800 676292 484802
rect 673085 484744 673090 484800
rect 673146 484744 676292 484800
rect 673085 484742 676292 484744
rect 673085 484739 673151 484742
rect 674649 484394 674715 484397
rect 674649 484392 676292 484394
rect 674649 484336 674654 484392
rect 674710 484336 676292 484392
rect 674649 484334 676292 484336
rect 674649 484331 674715 484334
rect 676029 483986 676095 483989
rect 676029 483984 676292 483986
rect 676029 483928 676034 483984
rect 676090 483928 676292 483984
rect 676029 483926 676292 483928
rect 676029 483923 676095 483926
rect 683205 483578 683271 483581
rect 683205 483576 683284 483578
rect 683205 483520 683210 483576
rect 683266 483520 683284 483576
rect 683205 483518 683284 483520
rect 683205 483515 683271 483518
rect 674005 483170 674071 483173
rect 674005 483168 676292 483170
rect 674005 483112 674010 483168
rect 674066 483112 676292 483168
rect 674005 483110 676292 483112
rect 674005 483107 674071 483110
rect 676029 482762 676095 482765
rect 676029 482760 676292 482762
rect 676029 482704 676034 482760
rect 676090 482704 676292 482760
rect 676029 482702 676292 482704
rect 676029 482699 676095 482702
rect 673545 482354 673611 482357
rect 673545 482352 676292 482354
rect 673545 482296 673550 482352
rect 673606 482296 676292 482352
rect 673545 482294 676292 482296
rect 673545 482291 673611 482294
rect 680353 481946 680419 481949
rect 680340 481944 680419 481946
rect 680340 481888 680358 481944
rect 680414 481888 680419 481944
rect 680340 481886 680419 481888
rect 680353 481883 680419 481886
rect 677182 481130 677242 481508
rect 683113 481130 683179 481133
rect 677182 481128 683179 481130
rect 677182 481100 683118 481128
rect 677212 481072 683118 481100
rect 683174 481072 683179 481128
rect 677212 481070 683179 481072
rect 683113 481067 683179 481070
rect 675845 480722 675911 480725
rect 675845 480720 676292 480722
rect 675845 480664 675850 480720
rect 675906 480664 676292 480720
rect 675845 480662 676292 480664
rect 675845 480659 675911 480662
rect 669773 455426 669839 455429
rect 673269 455426 673335 455429
rect 669773 455424 673335 455426
rect 669773 455368 669778 455424
rect 669834 455368 673274 455424
rect 673330 455368 673335 455424
rect 669773 455366 673335 455368
rect 669773 455363 669839 455366
rect 673269 455363 673335 455366
rect 673381 455290 673447 455293
rect 673862 455290 673868 455292
rect 673381 455288 673868 455290
rect 673381 455232 673386 455288
rect 673442 455232 673868 455288
rect 673381 455230 673868 455232
rect 673381 455227 673447 455230
rect 673862 455228 673868 455230
rect 673932 455228 673938 455292
rect 670601 455154 670667 455157
rect 673269 455154 673335 455157
rect 670601 455152 673335 455154
rect 670601 455096 670606 455152
rect 670662 455096 673274 455152
rect 673330 455096 673335 455152
rect 670601 455094 673335 455096
rect 670601 455091 670667 455094
rect 673269 455091 673335 455094
rect 672809 454882 672875 454885
rect 674281 454882 674347 454885
rect 672809 454880 674347 454882
rect 672809 454824 672814 454880
rect 672870 454824 674286 454880
rect 674342 454824 674347 454880
rect 672809 454822 674347 454824
rect 672809 454819 672875 454822
rect 674281 454819 674347 454822
rect 673039 454610 673105 454613
rect 674281 454610 674347 454613
rect 673039 454608 674347 454610
rect 673039 454552 673044 454608
rect 673100 454552 674286 454608
rect 674342 454552 674347 454608
rect 673039 454550 674347 454552
rect 673039 454547 673105 454550
rect 674281 454547 674347 454550
rect 672947 454338 673013 454341
rect 674281 454338 674347 454341
rect 672947 454336 674347 454338
rect 672947 454280 672952 454336
rect 673008 454280 674286 454336
rect 674342 454280 674347 454336
rect 672947 454278 674347 454280
rect 672947 454275 673013 454278
rect 674281 454275 674347 454278
rect 672257 453930 672323 453933
rect 674281 453930 674347 453933
rect 672257 453928 674347 453930
rect 672257 453872 672262 453928
rect 672318 453872 674286 453928
rect 674342 453872 674347 453928
rect 672257 453870 674347 453872
rect 672257 453867 672323 453870
rect 674281 453867 674347 453870
rect 44817 430946 44883 430949
rect 41492 430944 44883 430946
rect 41492 430888 44822 430944
rect 44878 430888 44883 430944
rect 41492 430886 44883 430888
rect 44817 430883 44883 430886
rect 47761 430538 47827 430541
rect 41492 430536 47827 430538
rect 41492 430480 47766 430536
rect 47822 430480 47827 430536
rect 41492 430478 47827 430480
rect 47761 430475 47827 430478
rect 35801 430130 35867 430133
rect 35788 430128 35867 430130
rect 35788 430072 35806 430128
rect 35862 430072 35867 430128
rect 35788 430070 35867 430072
rect 35801 430067 35867 430070
rect 44541 429722 44607 429725
rect 41492 429720 44607 429722
rect 41492 429664 44546 429720
rect 44602 429664 44607 429720
rect 41492 429662 44607 429664
rect 44541 429659 44607 429662
rect 44633 429314 44699 429317
rect 41492 429312 44699 429314
rect 41492 429256 44638 429312
rect 44694 429256 44699 429312
rect 41492 429254 44699 429256
rect 44633 429251 44699 429254
rect 45001 428906 45067 428909
rect 41492 428904 45067 428906
rect 41492 428848 45006 428904
rect 45062 428848 45067 428904
rect 41492 428846 45067 428848
rect 45001 428843 45067 428846
rect 35801 428498 35867 428501
rect 35788 428496 35867 428498
rect 35788 428440 35806 428496
rect 35862 428440 35867 428496
rect 35788 428438 35867 428440
rect 35801 428435 35867 428438
rect 44357 428090 44423 428093
rect 41492 428088 44423 428090
rect 41492 428032 44362 428088
rect 44418 428032 44423 428088
rect 41492 428030 44423 428032
rect 44357 428027 44423 428030
rect 44449 427682 44515 427685
rect 41492 427680 44515 427682
rect 41492 427624 44454 427680
rect 44510 427624 44515 427680
rect 41492 427622 44515 427624
rect 44449 427619 44515 427622
rect 43161 427410 43227 427413
rect 41784 427408 43227 427410
rect 41784 427352 43166 427408
rect 43222 427352 43227 427408
rect 41784 427350 43227 427352
rect 41784 427274 41844 427350
rect 43161 427347 43227 427350
rect 41492 427214 41844 427274
rect 42149 427138 42215 427141
rect 62481 427138 62547 427141
rect 42149 427136 62547 427138
rect 42149 427080 42154 427136
rect 42210 427080 62486 427136
rect 62542 427080 62547 427136
rect 42149 427078 62547 427080
rect 42149 427075 42215 427078
rect 62481 427075 62547 427078
rect 44265 426866 44331 426869
rect 41492 426864 44331 426866
rect 41492 426808 44270 426864
rect 44326 426808 44331 426864
rect 41492 426806 44331 426808
rect 44265 426803 44331 426806
rect 41965 426594 42031 426597
rect 42885 426594 42951 426597
rect 41965 426592 42951 426594
rect 41965 426536 41970 426592
rect 42026 426536 42890 426592
rect 42946 426536 42951 426592
rect 41965 426534 42951 426536
rect 41965 426531 42031 426534
rect 42885 426531 42951 426534
rect 40953 426458 41019 426461
rect 40940 426456 41019 426458
rect 40940 426400 40958 426456
rect 41014 426400 41019 426456
rect 40940 426398 41019 426400
rect 40953 426395 41019 426398
rect 41137 426050 41203 426053
rect 41124 426048 41203 426050
rect 41124 425992 41142 426048
rect 41198 425992 41203 426048
rect 41124 425990 41203 425992
rect 41137 425987 41203 425990
rect 39297 425642 39363 425645
rect 39284 425640 39363 425642
rect 39284 425584 39302 425640
rect 39358 425584 39363 425640
rect 39284 425582 39363 425584
rect 39297 425579 39363 425582
rect 43069 425234 43135 425237
rect 41492 425232 43135 425234
rect 41492 425176 43074 425232
rect 43130 425176 43135 425232
rect 41492 425174 43135 425176
rect 43069 425171 43135 425174
rect 32765 424826 32831 424829
rect 32765 424824 32844 424826
rect 32765 424768 32770 424824
rect 32826 424768 32844 424824
rect 32765 424766 32844 424768
rect 32765 424763 32831 424766
rect 34513 424418 34579 424421
rect 34500 424416 34579 424418
rect 34500 424360 34518 424416
rect 34574 424360 34579 424416
rect 34500 424358 34579 424360
rect 34513 424355 34579 424358
rect 33777 424010 33843 424013
rect 33764 424008 33843 424010
rect 33764 423952 33782 424008
rect 33838 423952 33843 424008
rect 33764 423950 33843 423952
rect 33777 423947 33843 423950
rect 41776 423602 41782 423604
rect 41492 423542 41782 423602
rect 41776 423540 41782 423542
rect 41846 423540 41852 423604
rect 45093 423194 45159 423197
rect 41492 423192 45159 423194
rect 41492 423136 45098 423192
rect 45154 423136 45159 423192
rect 41492 423134 45159 423136
rect 45093 423131 45159 423134
rect 43805 422786 43871 422789
rect 41492 422784 43871 422786
rect 41492 422728 43810 422784
rect 43866 422728 43871 422784
rect 41492 422726 43871 422728
rect 43805 422723 43871 422726
rect 41781 422378 41847 422381
rect 41492 422376 41847 422378
rect 41492 422320 41786 422376
rect 41842 422320 41847 422376
rect 41492 422318 41847 422320
rect 41781 422315 41847 422318
rect 42006 421970 42012 421972
rect 41492 421910 42012 421970
rect 42006 421908 42012 421910
rect 42076 421908 42082 421972
rect 42149 421562 42215 421565
rect 41492 421560 42215 421562
rect 41492 421504 42154 421560
rect 42210 421504 42215 421560
rect 41492 421502 42215 421504
rect 42149 421499 42215 421502
rect 43989 421154 44055 421157
rect 41492 421152 44055 421154
rect 41492 421096 43994 421152
rect 44050 421096 44055 421152
rect 41492 421094 44055 421096
rect 43989 421091 44055 421094
rect 45461 420746 45527 420749
rect 41492 420744 45527 420746
rect 41492 420688 45466 420744
rect 45522 420688 45527 420744
rect 41492 420686 45527 420688
rect 45461 420683 45527 420686
rect 41321 419930 41387 419933
rect 41308 419928 41387 419930
rect 41308 419872 41326 419928
rect 41382 419872 41387 419928
rect 41308 419870 41387 419872
rect 41321 419867 41387 419870
rect 41321 418842 41387 418845
rect 49325 418842 49391 418845
rect 41321 418840 49391 418842
rect 41321 418784 41326 418840
rect 41382 418784 49330 418840
rect 49386 418784 49391 418840
rect 41321 418782 49391 418784
rect 41321 418779 41387 418782
rect 49325 418779 49391 418782
rect 40902 418508 40908 418572
rect 40972 418570 40978 418572
rect 41781 418570 41847 418573
rect 40972 418568 41847 418570
rect 40972 418512 41786 418568
rect 41842 418512 41847 418568
rect 40972 418510 41847 418512
rect 40972 418508 40978 418510
rect 41781 418507 41847 418510
rect 40534 418236 40540 418300
rect 40604 418298 40610 418300
rect 42149 418298 42215 418301
rect 40604 418296 42215 418298
rect 40604 418240 42154 418296
rect 42210 418240 42215 418296
rect 40604 418238 42215 418240
rect 40604 418236 40610 418238
rect 42149 418235 42215 418238
rect 40718 417964 40724 418028
rect 40788 418026 40794 418028
rect 42006 418026 42012 418028
rect 40788 417966 42012 418026
rect 40788 417964 40794 417966
rect 42006 417964 42012 417966
rect 42076 417964 42082 418028
rect 40953 417754 41019 417757
rect 41454 417754 41460 417756
rect 40953 417752 41460 417754
rect 40953 417696 40958 417752
rect 41014 417696 41460 417752
rect 40953 417694 41460 417696
rect 40953 417691 41019 417694
rect 41454 417692 41460 417694
rect 41524 417692 41530 417756
rect 41822 417692 41828 417756
rect 41892 417754 41898 417756
rect 42977 417754 43043 417757
rect 41892 417752 43043 417754
rect 41892 417696 42982 417752
rect 43038 417696 43043 417752
rect 41892 417694 43043 417696
rect 41892 417692 41898 417694
rect 42977 417691 43043 417694
rect 39297 415306 39363 415309
rect 42006 415306 42012 415308
rect 39297 415304 42012 415306
rect 39297 415248 39302 415304
rect 39358 415248 42012 415304
rect 39297 415246 42012 415248
rect 39297 415243 39363 415246
rect 42006 415244 42012 415246
rect 42076 415244 42082 415308
rect 33777 414626 33843 414629
rect 41822 414626 41828 414628
rect 33777 414624 41828 414626
rect 33777 414568 33782 414624
rect 33838 414568 41828 414624
rect 33777 414566 41828 414568
rect 33777 414563 33843 414566
rect 41822 414564 41828 414566
rect 41892 414564 41898 414628
rect 41781 413538 41847 413541
rect 41781 413536 41890 413538
rect 41781 413480 41786 413536
rect 41842 413480 41890 413536
rect 41781 413475 41890 413480
rect 41830 413133 41890 413475
rect 41781 413128 41890 413133
rect 41781 413072 41786 413128
rect 41842 413072 41890 413128
rect 41781 413070 41890 413072
rect 41781 413067 41847 413070
rect 42241 409866 42307 409869
rect 43805 409866 43871 409869
rect 42241 409864 43871 409866
rect 42241 409808 42246 409864
rect 42302 409808 43810 409864
rect 43866 409808 43871 409864
rect 42241 409806 43871 409808
rect 42241 409803 42307 409806
rect 43805 409803 43871 409806
rect 42057 408098 42123 408101
rect 43989 408098 44055 408101
rect 42057 408096 44055 408098
rect 42057 408040 42062 408096
rect 42118 408040 43994 408096
rect 44050 408040 44055 408096
rect 42057 408038 44055 408040
rect 42057 408035 42123 408038
rect 43989 408035 44055 408038
rect 42425 407282 42491 407285
rect 45277 407282 45343 407285
rect 42425 407280 45343 407282
rect 42425 407224 42430 407280
rect 42486 407224 45282 407280
rect 45338 407224 45343 407280
rect 42425 407222 45343 407224
rect 42425 407219 42491 407222
rect 45277 407219 45343 407222
rect 40902 406948 40908 407012
rect 40972 407010 40978 407012
rect 41781 407010 41847 407013
rect 40972 407008 41847 407010
rect 40972 406952 41786 407008
rect 41842 406952 41847 407008
rect 40972 406950 41847 406952
rect 40972 406948 40978 406950
rect 41781 406947 41847 406950
rect 40534 406676 40540 406740
rect 40604 406738 40610 406740
rect 41781 406738 41847 406741
rect 40604 406736 41847 406738
rect 40604 406680 41786 406736
rect 41842 406680 41847 406736
rect 40604 406678 41847 406680
rect 40604 406676 40610 406678
rect 41781 406675 41847 406678
rect 42425 404970 42491 404973
rect 51441 404970 51507 404973
rect 42425 404968 51507 404970
rect 42425 404912 42430 404968
rect 42486 404912 51446 404968
rect 51502 404912 51507 404968
rect 42425 404910 51507 404912
rect 42425 404907 42491 404910
rect 51441 404907 51507 404910
rect 40718 404500 40724 404564
rect 40788 404562 40794 404564
rect 42241 404562 42307 404565
rect 40788 404560 42307 404562
rect 40788 404504 42246 404560
rect 42302 404504 42307 404560
rect 40788 404502 42307 404504
rect 40788 404500 40794 404502
rect 42241 404499 42307 404502
rect 62113 404154 62179 404157
rect 62113 404152 64706 404154
rect 62113 404096 62118 404152
rect 62174 404096 64706 404152
rect 62113 404094 64706 404096
rect 62113 404091 62179 404094
rect 64646 403550 64706 404094
rect 676262 403746 676322 403852
rect 663750 403686 676322 403746
rect 657537 403338 657603 403341
rect 663750 403338 663810 403686
rect 676262 403341 676322 403444
rect 657537 403336 663810 403338
rect 657537 403280 657542 403336
rect 657598 403280 663810 403336
rect 657537 403278 663810 403280
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 657537 403275 657603 403278
rect 676213 403275 676279 403278
rect 676630 402933 676690 403036
rect 42333 402930 42399 402933
rect 45093 402930 45159 402933
rect 42333 402928 45159 402930
rect 42333 402872 42338 402928
rect 42394 402872 45098 402928
rect 45154 402872 45159 402928
rect 42333 402870 45159 402872
rect 42333 402867 42399 402870
rect 45093 402867 45159 402870
rect 676581 402928 676690 402933
rect 676581 402872 676586 402928
rect 676642 402872 676690 402928
rect 676581 402870 676690 402872
rect 676581 402867 676647 402870
rect 62113 402658 62179 402661
rect 62113 402656 64706 402658
rect 62113 402600 62118 402656
rect 62174 402600 64706 402656
rect 62113 402598 64706 402600
rect 62113 402595 62179 402598
rect 64646 402368 64706 402598
rect 672625 402522 672691 402525
rect 676262 402522 676322 402628
rect 672625 402520 676322 402522
rect 672625 402464 672630 402520
rect 672686 402464 676322 402520
rect 672625 402462 676322 402464
rect 672625 402459 672691 402462
rect 674833 402250 674899 402253
rect 674833 402248 676292 402250
rect 674833 402192 674838 402248
rect 674894 402192 676292 402248
rect 674833 402190 676292 402192
rect 674833 402187 674899 402190
rect 672441 401978 672507 401981
rect 672441 401976 676322 401978
rect 672441 401920 672446 401976
rect 672502 401920 676322 401976
rect 672441 401918 676322 401920
rect 672441 401915 672507 401918
rect 676262 401812 676322 401918
rect 673177 401706 673243 401709
rect 674833 401706 674899 401709
rect 673177 401704 674899 401706
rect 673177 401648 673182 401704
rect 673238 401648 674838 401704
rect 674894 401648 674899 401704
rect 673177 401646 674899 401648
rect 673177 401643 673243 401646
rect 674833 401643 674899 401646
rect 673913 401434 673979 401437
rect 673913 401432 676292 401434
rect 673913 401376 673918 401432
rect 673974 401376 676292 401432
rect 673913 401374 676292 401376
rect 673913 401371 673979 401374
rect 677174 401236 677180 401300
rect 677244 401236 677250 401300
rect 62113 400618 62179 400621
rect 64646 400618 64706 401186
rect 677182 400996 677242 401236
rect 652017 400890 652083 400893
rect 676581 400890 676647 400893
rect 652017 400888 676647 400890
rect 652017 400832 652022 400888
rect 652078 400832 676586 400888
rect 676642 400832 676647 400888
rect 652017 400830 676647 400832
rect 652017 400827 652083 400830
rect 676581 400827 676647 400830
rect 62113 400616 64706 400618
rect 62113 400560 62118 400616
rect 62174 400560 64706 400616
rect 62113 400558 64706 400560
rect 62113 400555 62179 400558
rect 673361 400482 673427 400485
rect 676262 400482 676322 400588
rect 673361 400480 676322 400482
rect 673361 400424 673366 400480
rect 673422 400424 676322 400480
rect 673361 400422 676322 400424
rect 673361 400419 673427 400422
rect 676806 400420 676812 400484
rect 676876 400420 676882 400484
rect 62481 400210 62547 400213
rect 62481 400208 64706 400210
rect 62481 400152 62486 400208
rect 62542 400152 64706 400208
rect 676814 400180 676874 400420
rect 62481 400150 64706 400152
rect 62481 400147 62547 400150
rect 41454 400012 41460 400076
rect 41524 400074 41530 400076
rect 41781 400074 41847 400077
rect 41524 400072 41847 400074
rect 41524 400016 41786 400072
rect 41842 400016 41847 400072
rect 41524 400014 41847 400016
rect 41524 400012 41530 400014
rect 41781 400011 41847 400014
rect 64646 400004 64706 400150
rect 672809 399666 672875 399669
rect 676262 399666 676322 399772
rect 672809 399664 676322 399666
rect 672809 399608 672814 399664
rect 672870 399608 676322 399664
rect 672809 399606 676322 399608
rect 672809 399603 672875 399606
rect 41781 399396 41847 399397
rect 41781 399392 41828 399396
rect 41892 399394 41898 399396
rect 62113 399394 62179 399397
rect 676029 399394 676095 399397
rect 41781 399336 41786 399392
rect 41781 399332 41828 399336
rect 41892 399334 41938 399394
rect 62113 399392 64706 399394
rect 62113 399336 62118 399392
rect 62174 399336 64706 399392
rect 62113 399334 64706 399336
rect 41892 399332 41898 399334
rect 41781 399331 41847 399332
rect 62113 399331 62179 399334
rect 41965 398852 42031 398853
rect 41965 398848 42012 398852
rect 42076 398850 42082 398852
rect 41965 398792 41970 398848
rect 41965 398788 42012 398792
rect 42076 398790 42122 398850
rect 64646 398822 64706 399334
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 42076 398788 42082 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 41965 398787 42031 398788
rect 679574 398445 679634 398548
rect 679574 398440 679683 398445
rect 679574 398384 679622 398440
rect 679678 398384 679683 398440
rect 679574 398382 679683 398384
rect 679617 398379 679683 398382
rect 62113 398306 62179 398309
rect 62113 398304 64706 398306
rect 62113 398248 62118 398304
rect 62174 398248 64706 398304
rect 62113 398246 64706 398248
rect 62113 398243 62179 398246
rect 64646 397640 64706 398246
rect 676262 398037 676322 398140
rect 676213 398032 676322 398037
rect 676213 397976 676218 398032
rect 676274 397976 676322 398032
rect 676213 397974 676322 397976
rect 676213 397971 676279 397974
rect 678286 397629 678346 397732
rect 678237 397624 678346 397629
rect 678237 397568 678242 397624
rect 678298 397568 678346 397624
rect 678237 397566 678346 397568
rect 678237 397563 678303 397566
rect 674741 397354 674807 397357
rect 674741 397352 676292 397354
rect 674741 397296 674746 397352
rect 674802 397296 676292 397352
rect 674741 397294 676292 397296
rect 674741 397291 674807 397294
rect 676262 396812 676322 396916
rect 676254 396748 676260 396812
rect 676324 396748 676330 396812
rect 652201 396674 652267 396677
rect 674557 396674 674623 396677
rect 652201 396672 674623 396674
rect 652201 396616 652206 396672
rect 652262 396616 674562 396672
rect 674618 396616 674623 396672
rect 652201 396614 674623 396616
rect 652201 396611 652267 396614
rect 674557 396611 674623 396614
rect 676446 396404 676506 396508
rect 676438 396340 676444 396404
rect 676508 396340 676514 396404
rect 676029 396130 676095 396133
rect 676029 396128 676292 396130
rect 676029 396072 676034 396128
rect 676090 396072 676292 396128
rect 676029 396070 676292 396072
rect 676029 396067 676095 396070
rect 42149 395722 42215 395725
rect 51073 395722 51139 395725
rect 42149 395720 51139 395722
rect 42149 395664 42154 395720
rect 42210 395664 51078 395720
rect 51134 395664 51139 395720
rect 42149 395662 51139 395664
rect 42149 395659 42215 395662
rect 51073 395659 51139 395662
rect 673729 395722 673795 395725
rect 673729 395720 676292 395722
rect 673729 395664 673734 395720
rect 673790 395664 676292 395720
rect 673729 395662 676292 395664
rect 673729 395659 673795 395662
rect 676630 395180 676690 395284
rect 676622 395116 676628 395180
rect 676692 395116 676698 395180
rect 672993 395042 673059 395045
rect 672993 395040 676322 395042
rect 672993 394984 672998 395040
rect 673054 394984 676322 395040
rect 672993 394982 676322 394984
rect 672993 394979 673059 394982
rect 676262 394876 676322 394982
rect 676262 394365 676322 394468
rect 676213 394360 676322 394365
rect 676213 394304 676218 394360
rect 676274 394304 676322 394360
rect 676213 394302 676322 394304
rect 676213 394299 676279 394302
rect 672625 393954 672691 393957
rect 676262 393954 676322 394060
rect 672625 393952 676322 393954
rect 672625 393896 672630 393952
rect 672686 393896 676322 393952
rect 672625 393894 676322 393896
rect 672625 393891 672691 393894
rect 671889 393682 671955 393685
rect 671889 393680 676292 393682
rect 671889 393624 671894 393680
rect 671950 393624 676292 393680
rect 671889 393622 676292 393624
rect 671889 393619 671955 393622
rect 675886 392804 675892 392868
rect 675956 392866 675962 392868
rect 676262 392866 676322 393244
rect 675956 392836 676322 392866
rect 675956 392806 676292 392836
rect 675956 392804 675962 392806
rect 670509 392594 670575 392597
rect 670509 392592 676322 392594
rect 670509 392536 670514 392592
rect 670570 392536 676322 392592
rect 670509 392534 676322 392536
rect 670509 392531 670575 392534
rect 676262 392428 676322 392534
rect 47761 387698 47827 387701
rect 41492 387696 47827 387698
rect 41492 387640 47766 387696
rect 47822 387640 47827 387696
rect 41492 387638 47827 387640
rect 47761 387635 47827 387638
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 678237 387698 678303 387701
rect 675772 387696 678303 387698
rect 675772 387640 678242 387696
rect 678298 387640 678303 387696
rect 675772 387638 678303 387640
rect 675772 387636 675778 387638
rect 678237 387635 678303 387638
rect 41278 387157 41338 387260
rect 41278 387152 41387 387157
rect 41278 387096 41326 387152
rect 41382 387096 41387 387152
rect 41278 387094 41387 387096
rect 41321 387091 41387 387094
rect 41094 386749 41154 386852
rect 41094 386744 41203 386749
rect 41094 386688 41142 386744
rect 41198 386688 41203 386744
rect 41094 386686 41203 386688
rect 41137 386683 41203 386686
rect 44633 386474 44699 386477
rect 41492 386472 44699 386474
rect 41492 386416 44638 386472
rect 44694 386416 44699 386472
rect 41492 386414 44699 386416
rect 44633 386411 44699 386414
rect 40910 385933 40970 386036
rect 40910 385928 41019 385933
rect 40910 385872 40958 385928
rect 41014 385872 41019 385928
rect 40910 385870 41019 385872
rect 40953 385867 41019 385870
rect 41137 385930 41203 385933
rect 62481 385930 62547 385933
rect 41137 385928 62547 385930
rect 41137 385872 41142 385928
rect 41198 385872 62486 385928
rect 62542 385872 62547 385928
rect 41137 385870 62547 385872
rect 41137 385867 41203 385870
rect 62481 385867 62547 385870
rect 42793 385658 42859 385661
rect 41492 385656 42859 385658
rect 41492 385600 42798 385656
rect 42854 385600 42859 385656
rect 41492 385598 42859 385600
rect 42793 385595 42859 385598
rect 43253 385250 43319 385253
rect 41492 385248 43319 385250
rect 41492 385192 43258 385248
rect 43314 385192 43319 385248
rect 41492 385190 43319 385192
rect 43253 385187 43319 385190
rect 675753 384978 675819 384981
rect 676254 384978 676260 384980
rect 675753 384976 676260 384978
rect 675753 384920 675758 384976
rect 675814 384920 676260 384976
rect 675753 384918 676260 384920
rect 675753 384915 675819 384918
rect 676254 384916 676260 384918
rect 676324 384916 676330 384980
rect 44449 384842 44515 384845
rect 41492 384840 44515 384842
rect 41492 384784 44454 384840
rect 44510 384784 44515 384840
rect 41492 384782 44515 384784
rect 44449 384779 44515 384782
rect 45093 384434 45159 384437
rect 41492 384432 45159 384434
rect 41492 384376 45098 384432
rect 45154 384376 45159 384432
rect 41492 384374 45159 384376
rect 45093 384371 45159 384374
rect 44265 384026 44331 384029
rect 41492 384024 44331 384026
rect 41492 383968 44270 384024
rect 44326 383968 44331 384024
rect 41492 383966 44331 383968
rect 44265 383963 44331 383966
rect 45277 383618 45343 383621
rect 41492 383616 45343 383618
rect 41492 383560 45282 383616
rect 45338 383560 45343 383616
rect 41492 383558 45343 383560
rect 45277 383555 45343 383558
rect 41094 383077 41154 383180
rect 41094 383072 41203 383077
rect 41094 383016 41142 383072
rect 41198 383016 41203 383072
rect 41094 383014 41203 383016
rect 41137 383011 41203 383014
rect 654777 382938 654843 382941
rect 675109 382938 675175 382941
rect 654777 382936 675175 382938
rect 654777 382880 654782 382936
rect 654838 382880 675114 382936
rect 675170 382880 675175 382936
rect 654777 382878 675175 382880
rect 654777 382875 654843 382878
rect 675109 382875 675175 382878
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 39990 382261 40050 382364
rect 39990 382256 40099 382261
rect 39990 382200 40038 382256
rect 40094 382200 40099 382256
rect 39990 382198 40099 382200
rect 40033 382195 40099 382198
rect 40953 382258 41019 382261
rect 44909 382258 44975 382261
rect 40953 382256 44975 382258
rect 40953 382200 40958 382256
rect 41014 382200 44914 382256
rect 44970 382200 44975 382256
rect 40953 382198 44975 382200
rect 40953 382195 41019 382198
rect 44909 382195 44975 382198
rect 675753 382258 675819 382261
rect 676438 382258 676444 382260
rect 675753 382256 676444 382258
rect 675753 382200 675758 382256
rect 675814 382200 676444 382256
rect 675753 382198 676444 382200
rect 675753 382195 675819 382198
rect 676438 382196 676444 382198
rect 676508 382196 676514 382260
rect 35390 381853 35450 381956
rect 35390 381848 35499 381853
rect 35390 381792 35438 381848
rect 35494 381792 35499 381848
rect 35390 381790 35499 381792
rect 35433 381787 35499 381790
rect 41137 381850 41203 381853
rect 41454 381850 41460 381852
rect 41137 381848 41460 381850
rect 41137 381792 41142 381848
rect 41198 381792 41460 381848
rect 41137 381790 41460 381792
rect 41137 381787 41203 381790
rect 41454 381788 41460 381790
rect 41524 381788 41530 381852
rect 41873 381578 41939 381581
rect 63309 381578 63375 381581
rect 41873 381576 63375 381578
rect 39254 381445 39314 381548
rect 41873 381520 41878 381576
rect 41934 381520 63314 381576
rect 63370 381520 63375 381576
rect 41873 381518 63375 381520
rect 41873 381515 41939 381518
rect 63309 381515 63375 381518
rect 39254 381440 39363 381445
rect 39254 381384 39302 381440
rect 39358 381384 39363 381440
rect 39254 381382 39363 381384
rect 39297 381379 39363 381382
rect 33918 381037 33978 381140
rect 33918 381032 34027 381037
rect 33918 380976 33966 381032
rect 34022 380976 34027 381032
rect 33918 380974 34027 380976
rect 33961 380971 34027 380974
rect 672993 381034 673059 381037
rect 675385 381034 675451 381037
rect 672993 381032 675451 381034
rect 672993 380976 672998 381032
rect 673054 380976 675390 381032
rect 675446 380976 675451 381032
rect 672993 380974 675451 380976
rect 672993 380971 673059 380974
rect 675385 380971 675451 380974
rect 42885 380762 42951 380765
rect 41492 380760 42951 380762
rect 41492 380704 42890 380760
rect 42946 380704 42951 380760
rect 41492 380702 42951 380704
rect 42885 380699 42951 380702
rect 44633 380354 44699 380357
rect 41492 380352 44699 380354
rect 41492 380296 44638 380352
rect 44694 380296 44699 380352
rect 41492 380294 44699 380296
rect 44633 380291 44699 380294
rect 41278 379813 41338 379916
rect 41278 379808 41387 379813
rect 41278 379752 41326 379808
rect 41382 379752 41387 379808
rect 41278 379750 41387 379752
rect 41321 379747 41387 379750
rect 41505 379810 41571 379813
rect 43805 379810 43871 379813
rect 41505 379808 43871 379810
rect 41505 379752 41510 379808
rect 41566 379752 43810 379808
rect 43866 379752 43871 379808
rect 41505 379750 43871 379752
rect 41505 379747 41571 379750
rect 43805 379747 43871 379750
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 40033 379402 40099 379405
rect 41638 379402 41644 379404
rect 40033 379400 41644 379402
rect 40033 379344 40038 379400
rect 40094 379344 41644 379400
rect 40033 379342 41644 379344
rect 40033 379339 40099 379342
rect 41638 379340 41644 379342
rect 41708 379340 41714 379404
rect 40726 378996 40786 379100
rect 40718 378932 40724 378996
rect 40788 378932 40794 378996
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 35758 378181 35818 378284
rect 35758 378176 35867 378181
rect 35758 378120 35806 378176
rect 35862 378120 35867 378176
rect 35758 378118 35867 378120
rect 35801 378115 35867 378118
rect 41689 378178 41755 378181
rect 43989 378178 44055 378181
rect 41689 378176 44055 378178
rect 41689 378120 41694 378176
rect 41750 378120 43994 378176
rect 44050 378120 44055 378176
rect 41689 378118 44055 378120
rect 41689 378115 41755 378118
rect 43989 378115 44055 378118
rect 40910 377772 40970 377876
rect 40902 377708 40908 377772
rect 40972 377708 40978 377772
rect 44265 377498 44331 377501
rect 41492 377496 44331 377498
rect 41492 377440 44270 377496
rect 44326 377440 44331 377496
rect 41492 377438 44331 377440
rect 44265 377435 44331 377438
rect 675753 377362 675819 377365
rect 676622 377362 676628 377364
rect 675753 377360 676628 377362
rect 675753 377304 675758 377360
rect 675814 377304 676628 377360
rect 675753 377302 676628 377304
rect 675753 377299 675819 377302
rect 676622 377300 676628 377302
rect 676692 377300 676698 377364
rect 35758 376549 35818 377060
rect 40401 376954 40467 376957
rect 43069 376954 43135 376957
rect 40401 376952 43135 376954
rect 40401 376896 40406 376952
rect 40462 376896 43074 376952
rect 43130 376896 43135 376952
rect 40401 376894 43135 376896
rect 40401 376891 40467 376894
rect 43069 376891 43135 376894
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 41462 376546 41522 376652
rect 41462 376486 41890 376546
rect 35801 376483 35867 376486
rect 35801 376138 35867 376141
rect 41830 376138 41890 376486
rect 672625 376274 672691 376277
rect 675385 376274 675451 376277
rect 672625 376272 675451 376274
rect 672625 376216 672630 376272
rect 672686 376216 675390 376272
rect 675446 376216 675451 376272
rect 672625 376214 675451 376216
rect 672625 376211 672691 376214
rect 675385 376211 675451 376214
rect 46381 376138 46447 376141
rect 35801 376136 46447 376138
rect 35801 376080 35806 376136
rect 35862 376080 46386 376136
rect 46442 376080 46447 376136
rect 35801 376078 46447 376080
rect 35801 376075 35867 376078
rect 46381 376075 46447 376078
rect 673729 375458 673795 375461
rect 675109 375458 675175 375461
rect 673729 375456 675175 375458
rect 673729 375400 673734 375456
rect 673790 375400 675114 375456
rect 675170 375400 675175 375456
rect 673729 375398 675175 375400
rect 673729 375395 673795 375398
rect 675109 375395 675175 375398
rect 35433 374642 35499 374645
rect 41822 374642 41828 374644
rect 35433 374640 41828 374642
rect 35433 374584 35438 374640
rect 35494 374584 41828 374640
rect 35433 374582 41828 374584
rect 35433 374579 35499 374582
rect 41822 374580 41828 374582
rect 41892 374580 41898 374644
rect 652201 373962 652267 373965
rect 649950 373960 652267 373962
rect 649950 373904 652206 373960
rect 652262 373904 652267 373960
rect 649950 373902 652267 373904
rect 649950 373892 650010 373902
rect 652201 373899 652267 373902
rect 675753 373690 675819 373693
rect 676070 373690 676076 373692
rect 675753 373688 676076 373690
rect 675753 373632 675758 373688
rect 675814 373632 676076 373688
rect 675753 373630 676076 373632
rect 675753 373627 675819 373630
rect 676070 373628 676076 373630
rect 676140 373628 676146 373692
rect 651465 373282 651531 373285
rect 649950 373280 651531 373282
rect 649950 373224 651470 373280
rect 651526 373224 651531 373280
rect 649950 373222 651531 373224
rect 649950 372710 650010 373222
rect 651465 373219 651531 373222
rect 675385 372468 675451 372469
rect 675334 372404 675340 372468
rect 675404 372466 675451 372468
rect 675404 372464 675496 372466
rect 675446 372408 675496 372464
rect 675404 372406 675496 372408
rect 675404 372404 675451 372406
rect 675385 372403 675451 372404
rect 652017 372194 652083 372197
rect 649950 372192 652083 372194
rect 649950 372136 652022 372192
rect 652078 372136 652083 372192
rect 649950 372134 652083 372136
rect 649950 371528 650010 372134
rect 652017 372131 652083 372134
rect 651465 370698 651531 370701
rect 649950 370696 651531 370698
rect 649950 370640 651470 370696
rect 651526 370640 651531 370696
rect 649950 370638 651531 370640
rect 649950 370346 650010 370638
rect 651465 370635 651531 370638
rect 655513 366346 655579 366349
rect 675334 366346 675340 366348
rect 655513 366344 675340 366346
rect 655513 366288 655518 366344
rect 655574 366288 675340 366344
rect 655513 366286 675340 366288
rect 655513 366283 655579 366286
rect 675334 366284 675340 366286
rect 675404 366284 675410 366348
rect 40902 364788 40908 364852
rect 40972 364850 40978 364852
rect 41781 364850 41847 364853
rect 40972 364848 41847 364850
rect 40972 364792 41786 364848
rect 41842 364792 41847 364848
rect 40972 364790 41847 364792
rect 40972 364788 40978 364790
rect 41781 364787 41847 364790
rect 40718 364108 40724 364172
rect 40788 364170 40794 364172
rect 41781 364170 41847 364173
rect 40788 364168 41847 364170
rect 40788 364112 41786 364168
rect 41842 364112 41847 364168
rect 40788 364110 41847 364112
rect 40788 364108 40794 364110
rect 41781 364107 41847 364110
rect 42057 363626 42123 363629
rect 43989 363626 44055 363629
rect 42057 363624 44055 363626
rect 42057 363568 42062 363624
rect 42118 363568 43994 363624
rect 44050 363568 44055 363624
rect 42057 363566 44055 363568
rect 42057 363563 42123 363566
rect 43989 363563 44055 363566
rect 42701 363082 42767 363085
rect 45645 363082 45711 363085
rect 42701 363080 45711 363082
rect 42701 363024 42706 363080
rect 42762 363024 45650 363080
rect 45706 363024 45711 363080
rect 42701 363022 45711 363024
rect 42701 363019 42767 363022
rect 45645 363019 45711 363022
rect 42425 362266 42491 362269
rect 51073 362266 51139 362269
rect 42425 362264 51139 362266
rect 42425 362208 42430 362264
rect 42486 362208 51078 362264
rect 51134 362208 51139 362264
rect 42425 362206 51139 362208
rect 42425 362203 42491 362206
rect 51073 362203 51139 362206
rect 62113 360906 62179 360909
rect 62113 360904 64706 360906
rect 62113 360848 62118 360904
rect 62174 360848 64706 360904
rect 62113 360846 64706 360848
rect 62113 360843 62179 360846
rect 64646 360328 64706 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 42149 359954 42215 359957
rect 43805 359954 43871 359957
rect 42149 359952 43871 359954
rect 42149 359896 42154 359952
rect 42210 359896 43810 359952
rect 43866 359896 43871 359952
rect 42149 359894 43871 359896
rect 42149 359891 42215 359894
rect 43805 359891 43871 359894
rect 62113 359818 62179 359821
rect 62113 359816 64706 359818
rect 62113 359760 62118 359816
rect 62174 359760 64706 359816
rect 62113 359758 64706 359760
rect 62113 359755 62179 359758
rect 64646 359146 64706 359758
rect 42425 359002 42491 359005
rect 44633 359002 44699 359005
rect 42425 359000 44699 359002
rect 42425 358944 42430 359000
rect 42486 358944 44638 359000
rect 44694 358944 44699 359000
rect 42425 358942 44699 358944
rect 42425 358939 42491 358942
rect 44633 358939 44699 358942
rect 41873 358732 41939 358733
rect 41822 358730 41828 358732
rect 41782 358670 41828 358730
rect 41892 358728 41939 358732
rect 41934 358672 41939 358728
rect 41822 358668 41828 358670
rect 41892 358668 41939 358672
rect 41873 358667 41939 358668
rect 663750 358670 676292 358730
rect 654777 358594 654843 358597
rect 663750 358594 663810 358670
rect 654777 358592 663810 358594
rect 654777 358536 654782 358592
rect 654838 358536 663810 358592
rect 654777 358534 663810 358536
rect 654777 358531 654843 358534
rect 674465 358322 674531 358325
rect 674465 358320 676292 358322
rect 674465 358264 674470 358320
rect 674526 358264 676292 358320
rect 674465 358262 676292 358264
rect 674465 358259 674531 358262
rect 62113 357778 62179 357781
rect 64646 357778 64706 357964
rect 675937 357914 676003 357917
rect 675937 357912 676292 357914
rect 675937 357856 675942 357912
rect 675998 357856 676292 357912
rect 675937 357854 676292 357856
rect 675937 357851 676003 357854
rect 62113 357776 64706 357778
rect 62113 357720 62118 357776
rect 62174 357720 64706 357776
rect 62113 357718 64706 357720
rect 62113 357715 62179 357718
rect 673177 357506 673243 357509
rect 673177 357504 676292 357506
rect 673177 357448 673182 357504
rect 673238 357448 676292 357504
rect 673177 357446 676292 357448
rect 673177 357443 673243 357446
rect 62481 357370 62547 357373
rect 62481 357368 64706 357370
rect 62481 357312 62486 357368
rect 62542 357312 64706 357368
rect 62481 357310 64706 357312
rect 62481 357307 62547 357310
rect 41454 356900 41460 356964
rect 41524 356962 41530 356964
rect 41781 356962 41847 356965
rect 41524 356960 41847 356962
rect 41524 356904 41786 356960
rect 41842 356904 41847 356960
rect 41524 356902 41847 356904
rect 41524 356900 41530 356902
rect 41781 356899 41847 356902
rect 64646 356782 64706 357310
rect 672349 357098 672415 357101
rect 672349 357096 676292 357098
rect 672349 357040 672354 357096
rect 672410 357040 676292 357096
rect 672349 357038 676292 357040
rect 672349 357035 672415 357038
rect 675937 356826 676003 356829
rect 669270 356824 676003 356826
rect 669270 356768 675942 356824
rect 675998 356768 676003 356824
rect 669270 356766 676003 356768
rect 652017 356690 652083 356693
rect 669270 356690 669330 356766
rect 675937 356763 676003 356766
rect 652017 356688 669330 356690
rect 652017 356632 652022 356688
rect 652078 356632 669330 356688
rect 652017 356630 669330 356632
rect 676170 356630 676292 356690
rect 652017 356627 652083 356630
rect 673913 356554 673979 356557
rect 676170 356554 676230 356630
rect 673913 356552 676230 356554
rect 673913 356496 673918 356552
rect 673974 356496 676230 356552
rect 673913 356494 676230 356496
rect 673913 356491 673979 356494
rect 672533 356282 672599 356285
rect 672533 356280 676292 356282
rect 672533 356224 672538 356280
rect 672594 356224 676292 356280
rect 672533 356222 676292 356224
rect 672533 356219 672599 356222
rect 42425 356010 42491 356013
rect 44633 356010 44699 356013
rect 42425 356008 44699 356010
rect 42425 355952 42430 356008
rect 42486 355952 44638 356008
rect 44694 355952 44699 356008
rect 42425 355950 44699 355952
rect 42425 355947 42491 355950
rect 44633 355947 44699 355950
rect 62113 356010 62179 356013
rect 62113 356008 64706 356010
rect 62113 355952 62118 356008
rect 62174 355952 64706 356008
rect 62113 355950 64706 355952
rect 62113 355947 62179 355950
rect 41873 355740 41939 355741
rect 41822 355738 41828 355740
rect 41782 355678 41828 355738
rect 41892 355736 41939 355740
rect 41934 355680 41939 355736
rect 41822 355676 41828 355678
rect 41892 355676 41939 355680
rect 41873 355675 41939 355676
rect 64646 355600 64706 355950
rect 673361 355874 673427 355877
rect 673361 355872 676292 355874
rect 673361 355816 673366 355872
rect 673422 355816 676292 355872
rect 673361 355814 676292 355816
rect 673361 355811 673427 355814
rect 673269 355466 673335 355469
rect 673269 355464 676292 355466
rect 673269 355408 673274 355464
rect 673330 355408 676292 355464
rect 673269 355406 676292 355408
rect 673269 355403 673335 355406
rect 672809 355058 672875 355061
rect 672809 355056 676292 355058
rect 672809 355000 672814 355056
rect 672870 355000 676292 355056
rect 672809 354998 676292 355000
rect 672809 354995 672875 354998
rect 43621 354786 43687 354789
rect 45829 354786 45895 354789
rect 43621 354784 45895 354786
rect 43621 354728 43626 354784
rect 43682 354728 45834 354784
rect 45890 354728 45895 354784
rect 43621 354726 45895 354728
rect 43621 354723 43687 354726
rect 45829 354723 45895 354726
rect 674649 354650 674715 354653
rect 674649 354648 676292 354650
rect 674649 354592 674654 354648
rect 674710 354592 676292 354648
rect 674649 354590 676292 354592
rect 674649 354587 674715 354590
rect 43294 354452 43300 354516
rect 43364 354514 43370 354516
rect 44449 354514 44515 354517
rect 43364 354512 44515 354514
rect 43364 354456 44454 354512
rect 44510 354456 44515 354512
rect 43364 354454 44515 354456
rect 43364 354452 43370 354454
rect 44449 354451 44515 354454
rect 63309 354514 63375 354517
rect 63309 354512 64706 354514
rect 63309 354456 63314 354512
rect 63370 354456 64706 354512
rect 63309 354454 64706 354456
rect 63309 354451 63375 354454
rect 64646 354418 64706 354454
rect 45645 354378 45711 354381
rect 47761 354378 47827 354381
rect 45645 354376 47827 354378
rect 45645 354320 45650 354376
rect 45706 354320 47766 354376
rect 47822 354320 47827 354376
rect 45645 354318 47827 354320
rect 45645 354315 45711 354318
rect 47761 354315 47827 354318
rect 43437 354242 43503 354245
rect 44725 354242 44791 354245
rect 43437 354240 44791 354242
rect 43437 354184 43442 354240
rect 43498 354184 44730 354240
rect 44786 354184 44791 354240
rect 43437 354182 44791 354184
rect 43437 354179 43503 354182
rect 44725 354179 44791 354182
rect 675518 354180 675524 354244
rect 675588 354242 675594 354244
rect 675588 354182 676292 354242
rect 675588 354180 675594 354182
rect 675886 353772 675892 353836
rect 675956 353834 675962 353836
rect 675956 353774 676292 353834
rect 675956 353772 675962 353774
rect 45461 353698 45527 353701
rect 51901 353698 51967 353701
rect 45461 353696 51967 353698
rect 45461 353640 45466 353696
rect 45522 353640 51906 353696
rect 51962 353640 51967 353696
rect 45461 353638 51967 353640
rect 45461 353635 45527 353638
rect 51901 353635 51967 353638
rect 45461 353426 45527 353429
rect 64321 353426 64387 353429
rect 45461 353424 64387 353426
rect 45461 353368 45466 353424
rect 45522 353368 64326 353424
rect 64382 353368 64387 353424
rect 45461 353366 64387 353368
rect 45461 353363 45527 353366
rect 64321 353363 64387 353366
rect 673085 353426 673151 353429
rect 673085 353424 676292 353426
rect 673085 353368 673090 353424
rect 673146 353368 676292 353424
rect 673085 353366 676292 353368
rect 673085 353363 673151 353366
rect 44265 353154 44331 353157
rect 45415 353154 45481 353157
rect 44265 353152 45481 353154
rect 44265 353096 44270 353152
rect 44326 353096 45420 353152
rect 45476 353096 45481 353152
rect 44265 353094 45481 353096
rect 44265 353091 44331 353094
rect 45415 353091 45481 353094
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 673729 352610 673795 352613
rect 673729 352608 676292 352610
rect 673729 352552 673734 352608
rect 673790 352552 676292 352608
rect 673729 352550 676292 352552
rect 673729 352547 673795 352550
rect 673913 352202 673979 352205
rect 673913 352200 676292 352202
rect 673913 352144 673918 352200
rect 673974 352144 676292 352200
rect 673913 352142 676292 352144
rect 673913 352139 673979 352142
rect 675886 351732 675892 351796
rect 675956 351794 675962 351796
rect 675956 351734 676292 351794
rect 675956 351732 675962 351734
rect 674281 351386 674347 351389
rect 674281 351384 676292 351386
rect 674281 351328 674286 351384
rect 674342 351328 676292 351384
rect 674281 351326 676292 351328
rect 674281 351323 674347 351326
rect 652385 351114 652451 351117
rect 674465 351114 674531 351117
rect 652385 351112 674531 351114
rect 652385 351056 652390 351112
rect 652446 351056 674470 351112
rect 674526 351056 674531 351112
rect 652385 351054 674531 351056
rect 652385 351051 652451 351054
rect 674465 351051 674531 351054
rect 676029 350978 676095 350981
rect 676029 350976 676292 350978
rect 676029 350920 676034 350976
rect 676090 350920 676292 350976
rect 676029 350918 676292 350920
rect 676029 350915 676095 350918
rect 674465 350570 674531 350573
rect 674465 350568 676292 350570
rect 674465 350512 674470 350568
rect 674526 350512 676292 350568
rect 674465 350510 676292 350512
rect 674465 350507 674531 350510
rect 672165 350162 672231 350165
rect 672165 350160 676292 350162
rect 672165 350104 672170 350160
rect 672226 350104 676292 350160
rect 672165 350102 676292 350104
rect 672165 350099 672231 350102
rect 672901 349754 672967 349757
rect 672901 349752 676292 349754
rect 672901 349696 672906 349752
rect 672962 349696 676292 349752
rect 672901 349694 676292 349696
rect 672901 349691 672967 349694
rect 673545 349346 673611 349349
rect 673545 349344 676292 349346
rect 673545 349288 673550 349344
rect 673606 349288 676292 349344
rect 673545 349286 676292 349288
rect 673545 349283 673611 349286
rect 671705 348938 671771 348941
rect 671705 348936 676292 348938
rect 671705 348880 671710 348936
rect 671766 348880 676292 348936
rect 671705 348878 676292 348880
rect 671705 348875 671771 348878
rect 672717 348530 672783 348533
rect 672717 348528 676292 348530
rect 672717 348472 672722 348528
rect 672778 348472 676292 348528
rect 672717 348470 676292 348472
rect 672717 348467 672783 348470
rect 675334 347652 675340 347716
rect 675404 347714 675410 347716
rect 683070 347714 683130 348092
rect 675404 347684 683130 347714
rect 675404 347654 683100 347684
rect 675404 347652 675410 347654
rect 669405 347306 669471 347309
rect 669405 347304 676292 347306
rect 669405 347248 669410 347304
rect 669466 347248 676292 347304
rect 669405 347246 676292 347248
rect 669405 347243 669471 347246
rect 676029 346626 676095 346629
rect 676438 346626 676444 346628
rect 676029 346624 676444 346626
rect 676029 346568 676034 346624
rect 676090 346568 676444 346624
rect 676029 346566 676444 346568
rect 676029 346563 676095 346566
rect 676438 346564 676444 346566
rect 676508 346564 676514 346628
rect 40217 345538 40283 345541
rect 43253 345538 43319 345541
rect 40217 345536 43319 345538
rect 40217 345480 40222 345536
rect 40278 345480 43258 345536
rect 43314 345480 43319 345536
rect 40217 345478 43319 345480
rect 40217 345475 40283 345478
rect 43253 345475 43319 345478
rect 35758 344317 35818 344556
rect 35758 344312 35867 344317
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35758 344254 35867 344256
rect 35801 344251 35867 344254
rect 35574 343909 35634 344148
rect 35574 343904 35683 343909
rect 35574 343848 35622 343904
rect 35678 343848 35683 343904
rect 35574 343846 35683 343848
rect 35617 343843 35683 343846
rect 32998 343501 33058 343740
rect 32998 343496 33107 343501
rect 32998 343440 33046 343496
rect 33102 343440 33107 343496
rect 32998 343438 33107 343440
rect 33041 343435 33107 343438
rect 44909 343362 44975 343365
rect 41492 343360 44975 343362
rect 41492 343304 44914 343360
rect 44970 343304 44975 343360
rect 41492 343302 44975 343304
rect 44909 343299 44975 343302
rect 44582 342954 44588 342956
rect 41492 342894 44588 342954
rect 44582 342892 44588 342894
rect 44652 342892 44658 342956
rect 35758 342277 35818 342516
rect 35758 342272 35867 342277
rect 35758 342216 35806 342272
rect 35862 342216 35867 342272
rect 35758 342214 35867 342216
rect 35801 342211 35867 342214
rect 39849 342274 39915 342277
rect 39849 342272 42810 342274
rect 39849 342216 39854 342272
rect 39910 342216 42810 342272
rect 39849 342214 42810 342216
rect 39849 342211 39915 342214
rect 42750 342138 42810 342214
rect 39622 341866 39682 342108
rect 42750 342078 55230 342138
rect 39849 341866 39915 341869
rect 39622 341864 39915 341866
rect 39622 341808 39854 341864
rect 39910 341808 39915 341864
rect 39622 341806 39915 341808
rect 39849 341803 39915 341806
rect 40033 341866 40099 341869
rect 40033 341864 50354 341866
rect 40033 341808 40038 341864
rect 40094 341808 50354 341864
rect 40033 341806 50354 341808
rect 40033 341803 40099 341806
rect 35758 341461 35818 341700
rect 35758 341456 35867 341461
rect 35758 341400 35806 341456
rect 35862 341400 35867 341456
rect 35758 341398 35867 341400
rect 35801 341395 35867 341398
rect 40217 341458 40283 341461
rect 45461 341458 45527 341461
rect 40217 341456 45527 341458
rect 40217 341400 40222 341456
rect 40278 341400 45466 341456
rect 45522 341400 45527 341456
rect 40217 341398 45527 341400
rect 50294 341458 50354 341806
rect 55170 341730 55230 342078
rect 62481 341730 62547 341733
rect 55170 341728 62547 341730
rect 55170 341672 62486 341728
rect 62542 341672 62547 341728
rect 55170 341670 62547 341672
rect 62481 341667 62547 341670
rect 63125 341458 63191 341461
rect 50294 341456 63191 341458
rect 50294 341400 63130 341456
rect 63186 341400 63191 341456
rect 50294 341398 63191 341400
rect 40217 341395 40283 341398
rect 45461 341395 45527 341398
rect 63125 341395 63191 341398
rect 39438 341053 39498 341292
rect 35801 341050 35867 341053
rect 35758 341048 35867 341050
rect 35758 340992 35806 341048
rect 35862 340992 35867 341048
rect 35758 340987 35867 340992
rect 39438 341048 39547 341053
rect 39438 340992 39486 341048
rect 39542 340992 39547 341048
rect 39438 340990 39547 340992
rect 39481 340987 39547 340990
rect 40217 341050 40283 341053
rect 45093 341050 45159 341053
rect 40217 341048 45159 341050
rect 40217 340992 40222 341048
rect 40278 340992 45098 341048
rect 45154 340992 45159 341048
rect 40217 340990 45159 340992
rect 40217 340987 40283 340990
rect 45093 340987 45159 340990
rect 35758 340884 35818 340987
rect 673085 340778 673151 340781
rect 675109 340778 675175 340781
rect 673085 340776 675175 340778
rect 673085 340720 673090 340776
rect 673146 340720 675114 340776
rect 675170 340720 675175 340776
rect 673085 340718 675175 340720
rect 673085 340715 673151 340718
rect 675109 340715 675175 340718
rect 40033 340642 40099 340645
rect 45277 340642 45343 340645
rect 40033 340640 45343 340642
rect 40033 340584 40038 340640
rect 40094 340584 45282 340640
rect 45338 340584 45343 340640
rect 40033 340582 45343 340584
rect 40033 340579 40099 340582
rect 45277 340579 45343 340582
rect 39622 340237 39682 340476
rect 39622 340232 39731 340237
rect 39622 340176 39670 340232
rect 39726 340176 39731 340232
rect 39622 340174 39731 340176
rect 39665 340171 39731 340174
rect 39849 340234 39915 340237
rect 42742 340234 42748 340236
rect 39849 340232 42748 340234
rect 39849 340176 39854 340232
rect 39910 340176 42748 340232
rect 39849 340174 42748 340176
rect 39849 340171 39915 340174
rect 42742 340172 42748 340174
rect 42812 340172 42818 340236
rect 675753 340234 675819 340237
rect 676254 340234 676260 340236
rect 675753 340232 676260 340234
rect 675753 340176 675758 340232
rect 675814 340176 676260 340232
rect 675753 340174 676260 340176
rect 675753 340171 675819 340174
rect 676254 340172 676260 340174
rect 676324 340172 676330 340236
rect 35574 339829 35634 340068
rect 35525 339824 35634 339829
rect 35801 339826 35867 339829
rect 35525 339768 35530 339824
rect 35586 339768 35634 339824
rect 35525 339766 35634 339768
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35525 339763 35591 339766
rect 35758 339763 35867 339768
rect 39665 339826 39731 339829
rect 44398 339826 44404 339828
rect 39665 339824 44404 339826
rect 39665 339768 39670 339824
rect 39726 339768 44404 339824
rect 39665 339766 44404 339768
rect 39665 339763 39731 339766
rect 44398 339764 44404 339766
rect 44468 339764 44474 339828
rect 35758 339660 35818 339763
rect 675477 339420 675543 339421
rect 675477 339416 675524 339420
rect 675588 339418 675594 339420
rect 675477 339360 675482 339416
rect 675477 339356 675524 339360
rect 675588 339358 675634 339418
rect 675588 339356 675594 339358
rect 675477 339355 675543 339356
rect 45645 339282 45711 339285
rect 41492 339280 45711 339282
rect 41492 339224 45650 339280
rect 45706 339224 45711 339280
rect 41492 339222 45711 339224
rect 45645 339219 45711 339222
rect 46933 338874 46999 338877
rect 41492 338872 46999 338874
rect 41492 338816 46938 338872
rect 46994 338816 46999 338872
rect 41492 338814 46999 338816
rect 46933 338811 46999 338814
rect 653397 338738 653463 338741
rect 674925 338738 674991 338741
rect 653397 338736 674991 338738
rect 653397 338680 653402 338736
rect 653458 338680 674930 338736
rect 674986 338680 674991 338736
rect 653397 338678 674991 338680
rect 653397 338675 653463 338678
rect 674925 338675 674991 338678
rect 41462 338194 41522 338436
rect 41638 338194 41644 338196
rect 41462 338134 41644 338194
rect 41638 338132 41644 338134
rect 41708 338132 41714 338196
rect 674281 338058 674347 338061
rect 675109 338058 675175 338061
rect 674281 338056 675175 338058
rect 41462 337922 41522 338028
rect 674281 338000 674286 338056
rect 674342 338000 675114 338056
rect 675170 338000 675175 338056
rect 674281 337998 675175 338000
rect 674281 337995 674347 337998
rect 675109 337995 675175 337998
rect 47117 337922 47183 337925
rect 41462 337920 47183 337922
rect 41462 337864 47122 337920
rect 47178 337864 47183 337920
rect 41462 337862 47183 337864
rect 47117 337859 47183 337862
rect 675753 337922 675819 337925
rect 676070 337922 676076 337924
rect 675753 337920 676076 337922
rect 675753 337864 675758 337920
rect 675814 337864 676076 337920
rect 675753 337862 676076 337864
rect 675753 337859 675819 337862
rect 676070 337860 676076 337862
rect 676140 337860 676146 337924
rect 45461 337650 45527 337653
rect 41492 337648 45527 337650
rect 41492 337592 45466 337648
rect 45522 337592 45527 337648
rect 41492 337590 45527 337592
rect 45461 337587 45527 337590
rect 39481 337378 39547 337381
rect 44766 337378 44772 337380
rect 39481 337376 44772 337378
rect 39481 337320 39486 337376
rect 39542 337320 44772 337376
rect 39481 337318 44772 337320
rect 39481 337315 39547 337318
rect 44766 337316 44772 337318
rect 44836 337316 44842 337380
rect 40542 336972 40602 337212
rect 40534 336908 40540 336972
rect 40604 336908 40610 336972
rect 42926 336834 42932 336836
rect 41492 336774 42932 336834
rect 42926 336772 42932 336774
rect 42996 336772 43002 336836
rect 38653 336562 38719 336565
rect 41454 336562 41460 336564
rect 38653 336560 41460 336562
rect 38653 336504 38658 336560
rect 38714 336504 41460 336560
rect 38653 336502 41460 336504
rect 38653 336499 38719 336502
rect 41454 336500 41460 336502
rect 41524 336500 41530 336564
rect 675753 336562 675819 336565
rect 676438 336562 676444 336564
rect 675753 336560 676444 336562
rect 675753 336504 675758 336560
rect 675814 336504 676444 336560
rect 675753 336502 676444 336504
rect 675753 336499 675819 336502
rect 676438 336500 676444 336502
rect 676508 336500 676514 336564
rect 35758 336157 35818 336396
rect 35758 336152 35867 336157
rect 35758 336096 35806 336152
rect 35862 336096 35867 336152
rect 35758 336094 35867 336096
rect 35801 336091 35867 336094
rect 40910 335748 40970 335988
rect 672165 335882 672231 335885
rect 674925 335882 674991 335885
rect 672165 335880 674991 335882
rect 672165 335824 672170 335880
rect 672226 335824 674930 335880
rect 674986 335824 674991 335880
rect 672165 335822 674991 335824
rect 672165 335819 672231 335822
rect 674925 335819 674991 335822
rect 40902 335684 40908 335748
rect 40972 335684 40978 335748
rect 672901 335610 672967 335613
rect 675109 335610 675175 335613
rect 672901 335608 675175 335610
rect 40726 335340 40786 335580
rect 672901 335552 672906 335608
rect 672962 335552 675114 335608
rect 675170 335552 675175 335608
rect 672901 335550 675175 335552
rect 672901 335547 672967 335550
rect 675109 335547 675175 335550
rect 40718 335276 40724 335340
rect 40788 335276 40794 335340
rect 41462 334930 41522 335172
rect 41462 334870 44282 334930
rect 35758 334525 35818 334764
rect 44222 334661 44282 334870
rect 43294 334596 43300 334660
rect 43364 334658 43370 334660
rect 43989 334658 44055 334661
rect 43364 334656 44055 334658
rect 43364 334600 43994 334656
rect 44050 334600 44055 334656
rect 43364 334598 44055 334600
rect 44222 334656 44331 334661
rect 44222 334600 44270 334656
rect 44326 334600 44331 334656
rect 44222 334598 44331 334600
rect 43364 334596 43370 334598
rect 43989 334595 44055 334598
rect 44265 334595 44331 334598
rect 35758 334520 35867 334525
rect 35758 334464 35806 334520
rect 35862 334464 35867 334520
rect 35758 334462 35867 334464
rect 35801 334459 35867 334462
rect 40217 334522 40283 334525
rect 43069 334522 43135 334525
rect 40217 334520 43135 334522
rect 40217 334464 40222 334520
rect 40278 334464 43074 334520
rect 43130 334464 43135 334520
rect 40217 334462 43135 334464
rect 40217 334459 40283 334462
rect 43069 334459 43135 334462
rect 41462 334114 41522 334356
rect 49141 334114 49207 334117
rect 41462 334112 49207 334114
rect 41462 334056 49146 334112
rect 49202 334056 49207 334112
rect 41462 334054 49207 334056
rect 49141 334051 49207 334054
rect 673729 333978 673795 333981
rect 675109 333978 675175 333981
rect 673729 333976 675175 333978
rect 41278 333570 41338 333948
rect 673729 333920 673734 333976
rect 673790 333920 675114 333976
rect 675170 333920 675175 333976
rect 673729 333918 675175 333920
rect 673729 333915 673795 333918
rect 675109 333915 675175 333918
rect 41278 333540 41492 333570
rect 41308 333510 41522 333540
rect 41462 333298 41522 333510
rect 41462 333238 51090 333298
rect 39757 332890 39823 332893
rect 42885 332890 42951 332893
rect 39757 332888 42951 332890
rect 39757 332832 39762 332888
rect 39818 332832 42890 332888
rect 42946 332832 42951 332888
rect 39757 332830 42951 332832
rect 39757 332827 39823 332830
rect 42885 332827 42951 332830
rect 51030 332618 51090 333238
rect 673545 332754 673611 332757
rect 675109 332754 675175 332757
rect 673545 332752 675175 332754
rect 673545 332696 673550 332752
rect 673606 332696 675114 332752
rect 675170 332696 675175 332752
rect 673545 332694 675175 332696
rect 673545 332691 673611 332694
rect 675109 332691 675175 332694
rect 63401 332618 63467 332621
rect 51030 332616 63467 332618
rect 51030 332560 63406 332616
rect 63462 332560 63467 332616
rect 51030 332558 63467 332560
rect 63401 332555 63467 332558
rect 37917 331258 37983 331261
rect 41822 331258 41828 331260
rect 37917 331256 41828 331258
rect 37917 331200 37922 331256
rect 37978 331200 41828 331256
rect 37917 331198 41828 331200
rect 37917 331195 37983 331198
rect 41822 331196 41828 331198
rect 41892 331196 41898 331260
rect 671705 331258 671771 331261
rect 675109 331258 675175 331261
rect 671705 331256 675175 331258
rect 671705 331200 671710 331256
rect 671766 331200 675114 331256
rect 675170 331200 675175 331256
rect 671705 331198 675175 331200
rect 671705 331195 671771 331198
rect 675109 331195 675175 331198
rect 652385 329762 652451 329765
rect 649950 329760 652451 329762
rect 649950 329704 652390 329760
rect 652446 329704 652451 329760
rect 649950 329702 652451 329704
rect 649950 329234 650010 329702
rect 652385 329699 652451 329702
rect 651373 328130 651439 328133
rect 649950 328128 651439 328130
rect 649950 328072 651378 328128
rect 651434 328072 651439 328128
rect 649950 328070 651439 328072
rect 649950 328052 650010 328070
rect 651373 328067 651439 328070
rect 675017 327994 675083 327997
rect 675385 327996 675451 327997
rect 675334 327994 675340 327996
rect 675017 327992 675340 327994
rect 675404 327994 675451 327996
rect 675404 327992 675496 327994
rect 675017 327936 675022 327992
rect 675078 327936 675340 327992
rect 675446 327936 675496 327992
rect 675017 327934 675340 327936
rect 675017 327931 675083 327934
rect 675334 327932 675340 327934
rect 675404 327934 675496 327936
rect 675404 327932 675451 327934
rect 675385 327931 675451 327932
rect 652017 326906 652083 326909
rect 650502 326904 652083 326906
rect 650502 326900 652022 326904
rect 649980 326848 652022 326900
rect 652078 326848 652083 326904
rect 649980 326846 652083 326848
rect 649980 326840 650562 326846
rect 652017 326843 652083 326846
rect 673913 326906 673979 326909
rect 675385 326906 675451 326909
rect 673913 326904 675451 326906
rect 673913 326848 673918 326904
rect 673974 326848 675390 326904
rect 675446 326848 675451 326904
rect 673913 326846 675451 326848
rect 673913 326843 673979 326846
rect 675385 326843 675451 326846
rect 649950 325682 650010 325710
rect 651373 325682 651439 325685
rect 649950 325680 651439 325682
rect 649950 325624 651378 325680
rect 651434 325624 651439 325680
rect 649950 325622 651439 325624
rect 651373 325619 651439 325622
rect 675201 325682 675267 325685
rect 676622 325682 676628 325684
rect 675201 325680 676628 325682
rect 675201 325624 675206 325680
rect 675262 325624 676628 325680
rect 675201 325622 676628 325624
rect 675201 325619 675267 325622
rect 676622 325620 676628 325622
rect 676692 325620 676698 325684
rect 672901 325002 672967 325005
rect 675017 325002 675083 325005
rect 672901 325000 675083 325002
rect 672901 324944 672906 325000
rect 672962 324944 675022 325000
rect 675078 324944 675083 325000
rect 672901 324942 675083 324944
rect 672901 324939 672967 324942
rect 675017 324939 675083 324942
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 42241 324322 42307 324325
rect 47117 324322 47183 324325
rect 42241 324320 47183 324322
rect 42241 324264 42246 324320
rect 42302 324264 47122 324320
rect 47178 324264 47183 324320
rect 42241 324262 47183 324264
rect 42241 324259 42307 324262
rect 47117 324259 47183 324262
rect 40902 321132 40908 321196
rect 40972 321194 40978 321196
rect 41781 321194 41847 321197
rect 40972 321192 41847 321194
rect 40972 321136 41786 321192
rect 41842 321136 41847 321192
rect 40972 321134 41847 321136
rect 40972 321132 40978 321134
rect 41781 321131 41847 321134
rect 42609 320650 42675 320653
rect 45277 320650 45343 320653
rect 42609 320648 45343 320650
rect 42609 320592 42614 320648
rect 42670 320592 45282 320648
rect 45338 320592 45343 320648
rect 42609 320590 45343 320592
rect 42609 320587 42675 320590
rect 45277 320587 45343 320590
rect 41781 319972 41847 319973
rect 41781 319968 41828 319972
rect 41892 319970 41898 319972
rect 42241 319970 42307 319973
rect 44265 319970 44331 319973
rect 41781 319912 41786 319968
rect 41781 319908 41828 319912
rect 41892 319910 41938 319970
rect 42241 319968 44331 319970
rect 42241 319912 42246 319968
rect 42302 319912 44270 319968
rect 44326 319912 44331 319968
rect 42241 319910 44331 319912
rect 41892 319908 41898 319910
rect 41781 319907 41847 319908
rect 42241 319907 42307 319910
rect 44265 319907 44331 319910
rect 42425 319426 42491 319429
rect 61561 319426 61627 319429
rect 42425 319424 61627 319426
rect 42425 319368 42430 319424
rect 42486 319368 61566 319424
rect 61622 319368 61627 319424
rect 42425 319366 61627 319368
rect 42425 319363 42491 319366
rect 61561 319363 61627 319366
rect 40718 317324 40724 317388
rect 40788 317386 40794 317388
rect 41781 317386 41847 317389
rect 40788 317384 41847 317386
rect 40788 317328 41786 317384
rect 41842 317328 41847 317384
rect 40788 317326 41847 317328
rect 40788 317324 40794 317326
rect 41781 317323 41847 317326
rect 62113 317386 62179 317389
rect 62113 317384 64706 317386
rect 62113 317328 62118 317384
rect 62174 317328 64706 317384
rect 62113 317326 64706 317328
rect 62113 317323 62179 317326
rect 64646 317106 64706 317326
rect 42425 316434 42491 316437
rect 42926 316434 42932 316436
rect 42425 316432 42932 316434
rect 42425 316376 42430 316432
rect 42486 316376 42932 316432
rect 42425 316374 42932 316376
rect 42425 316371 42491 316374
rect 42926 316372 42932 316374
rect 42996 316372 43002 316436
rect 40534 315964 40540 316028
rect 40604 316026 40610 316028
rect 41781 316026 41847 316029
rect 40604 316024 41847 316026
rect 40604 315968 41786 316024
rect 41842 315968 41847 316024
rect 40604 315966 41847 315968
rect 40604 315964 40610 315966
rect 41781 315963 41847 315966
rect 61561 316026 61627 316029
rect 61561 316024 64706 316026
rect 61561 315968 61566 316024
rect 61622 315968 64706 316024
rect 61561 315966 64706 315968
rect 61561 315963 61627 315966
rect 64646 315924 64706 315966
rect 62113 314802 62179 314805
rect 62113 314800 64706 314802
rect 62113 314744 62118 314800
rect 62174 314744 64706 314800
rect 62113 314742 64706 314744
rect 62113 314739 62179 314742
rect 62297 314122 62363 314125
rect 62297 314120 64706 314122
rect 62297 314064 62302 314120
rect 62358 314064 64706 314120
rect 62297 314062 64706 314064
rect 62297 314059 62363 314062
rect 41454 313652 41460 313716
rect 41524 313714 41530 313716
rect 41781 313714 41847 313717
rect 41524 313712 41847 313714
rect 41524 313656 41786 313712
rect 41842 313656 41847 313712
rect 41524 313654 41847 313656
rect 41524 313652 41530 313654
rect 41781 313651 41847 313654
rect 64646 313560 64706 314062
rect 676213 313986 676279 313989
rect 676213 313984 676322 313986
rect 676213 313928 676218 313984
rect 676274 313928 676322 313984
rect 676213 313923 676322 313928
rect 676262 313684 676322 313923
rect 653397 313306 653463 313309
rect 653397 313304 676292 313306
rect 653397 313248 653402 313304
rect 653458 313248 676292 313304
rect 653397 313246 676292 313248
rect 653397 313243 653463 313246
rect 42425 313170 42491 313173
rect 46933 313170 46999 313173
rect 42425 313168 46999 313170
rect 42425 313112 42430 313168
rect 42486 313112 46938 313168
rect 46994 313112 46999 313168
rect 42425 313110 46999 313112
rect 42425 313107 42491 313110
rect 46933 313107 46999 313110
rect 62481 313034 62547 313037
rect 62481 313032 64706 313034
rect 62481 312976 62486 313032
rect 62542 312976 64706 313032
rect 62481 312974 64706 312976
rect 62481 312971 62547 312974
rect 42425 312898 42491 312901
rect 45277 312898 45343 312901
rect 42425 312896 45343 312898
rect 42425 312840 42430 312896
rect 42486 312840 45282 312896
rect 45338 312840 45343 312896
rect 42425 312838 45343 312840
rect 42425 312835 42491 312838
rect 45277 312835 45343 312838
rect 42149 312626 42215 312629
rect 45645 312626 45711 312629
rect 42149 312624 45711 312626
rect 42149 312568 42154 312624
rect 42210 312568 45650 312624
rect 45706 312568 45711 312624
rect 42149 312566 45711 312568
rect 42149 312563 42215 312566
rect 45645 312563 45711 312566
rect 64646 312378 64706 312974
rect 674833 312898 674899 312901
rect 674833 312896 676292 312898
rect 674833 312840 674838 312896
rect 674894 312840 676292 312896
rect 674833 312838 676292 312840
rect 674833 312835 674899 312838
rect 672349 312490 672415 312493
rect 672349 312488 676292 312490
rect 672349 312432 672354 312488
rect 672410 312432 676292 312488
rect 672349 312430 676292 312432
rect 672349 312427 672415 312430
rect 675477 312082 675543 312085
rect 675477 312080 676292 312082
rect 675477 312024 675482 312080
rect 675538 312024 676292 312080
rect 675477 312022 676292 312024
rect 675477 312019 675543 312022
rect 658917 311946 658983 311949
rect 674833 311946 674899 311949
rect 658917 311944 674899 311946
rect 658917 311888 658922 311944
rect 658978 311888 674838 311944
rect 674894 311888 674899 311944
rect 658917 311886 674899 311888
rect 658917 311883 658983 311886
rect 674833 311883 674899 311886
rect 42149 311810 42215 311813
rect 45461 311810 45527 311813
rect 42149 311808 45527 311810
rect 42149 311752 42154 311808
rect 42210 311752 45466 311808
rect 45522 311752 45527 311808
rect 42149 311750 45527 311752
rect 42149 311747 42215 311750
rect 45461 311747 45527 311750
rect 63125 311810 63191 311813
rect 63125 311808 64706 311810
rect 63125 311752 63130 311808
rect 63186 311752 64706 311808
rect 63125 311750 64706 311752
rect 63125 311747 63191 311750
rect 64646 311196 64706 311750
rect 672533 311674 672599 311677
rect 672533 311672 676292 311674
rect 672533 311616 672538 311672
rect 672594 311616 676292 311672
rect 672533 311614 676292 311616
rect 672533 311611 672599 311614
rect 673913 311266 673979 311269
rect 673913 311264 676292 311266
rect 673913 311208 673918 311264
rect 673974 311208 676292 311264
rect 673913 311206 676292 311208
rect 673913 311203 673979 311206
rect 673269 310858 673335 310861
rect 673269 310856 676292 310858
rect 673269 310800 673274 310856
rect 673330 310800 676292 310856
rect 673269 310798 676292 310800
rect 673269 310795 673335 310798
rect 675477 310450 675543 310453
rect 675477 310448 676292 310450
rect 675477 310392 675482 310448
rect 675538 310392 676292 310448
rect 675477 310390 676292 310392
rect 675477 310387 675543 310390
rect 674649 310042 674715 310045
rect 674649 310040 676292 310042
rect 674649 309984 674654 310040
rect 674710 309984 676292 310040
rect 674649 309982 676292 309984
rect 674649 309979 674715 309982
rect 652293 309906 652359 309909
rect 652293 309904 663810 309906
rect 652293 309848 652298 309904
rect 652354 309848 663810 309904
rect 652293 309846 663810 309848
rect 652293 309843 652359 309846
rect 663750 309770 663810 309846
rect 675937 309770 676003 309773
rect 663750 309768 676003 309770
rect 663750 309712 675942 309768
rect 675998 309712 676003 309768
rect 663750 309710 676003 309712
rect 675937 309707 676003 309710
rect 676170 309574 676292 309634
rect 673361 309498 673427 309501
rect 676170 309498 676230 309574
rect 673361 309496 676230 309498
rect 673361 309440 673366 309496
rect 673422 309440 676230 309496
rect 673361 309438 676230 309440
rect 673361 309435 673427 309438
rect 675334 309164 675340 309228
rect 675404 309226 675410 309228
rect 675404 309166 676292 309226
rect 675404 309164 675410 309166
rect 675886 308756 675892 308820
rect 675956 308818 675962 308820
rect 675956 308758 676292 308818
rect 675956 308756 675962 308758
rect 675109 308410 675175 308413
rect 675109 308408 676292 308410
rect 675109 308352 675114 308408
rect 675170 308352 676292 308408
rect 675109 308350 676292 308352
rect 675109 308347 675175 308350
rect 674925 308002 674991 308005
rect 674925 308000 676292 308002
rect 674925 307944 674930 308000
rect 674986 307944 676292 308000
rect 674925 307942 676292 307944
rect 674925 307939 674991 307942
rect 676029 307594 676095 307597
rect 676029 307592 676292 307594
rect 676029 307536 676034 307592
rect 676090 307536 676292 307592
rect 676029 307534 676292 307536
rect 676029 307531 676095 307534
rect 676029 307186 676095 307189
rect 676029 307184 676292 307186
rect 676029 307128 676034 307184
rect 676090 307128 676292 307184
rect 676029 307126 676292 307128
rect 676029 307123 676095 307126
rect 678237 306778 678303 306781
rect 678237 306776 678316 306778
rect 678237 306720 678242 306776
rect 678298 306720 678316 306776
rect 678237 306718 678316 306720
rect 678237 306715 678303 306718
rect 678973 306370 679039 306373
rect 678973 306368 679052 306370
rect 678973 306312 678978 306368
rect 679034 306312 679052 306368
rect 678973 306310 679052 306312
rect 678973 306307 679039 306310
rect 673545 305962 673611 305965
rect 673545 305960 676292 305962
rect 673545 305904 673550 305960
rect 673606 305904 676292 305960
rect 673545 305902 676292 305904
rect 673545 305899 673611 305902
rect 672533 305554 672599 305557
rect 672533 305552 676292 305554
rect 672533 305496 672538 305552
rect 672594 305496 676292 305552
rect 672533 305494 676292 305496
rect 672533 305491 672599 305494
rect 675894 305086 676292 305146
rect 675894 304602 675954 305086
rect 676581 304738 676647 304741
rect 676581 304736 676660 304738
rect 676581 304680 676586 304736
rect 676642 304680 676660 304736
rect 676581 304678 676660 304680
rect 676581 304675 676647 304678
rect 676070 304602 676076 304604
rect 675894 304542 676076 304602
rect 676070 304540 676076 304542
rect 676140 304540 676146 304604
rect 673177 304330 673243 304333
rect 673177 304328 676292 304330
rect 673177 304272 673182 304328
rect 673238 304272 676292 304328
rect 673177 304270 676292 304272
rect 673177 304267 673243 304270
rect 674649 303922 674715 303925
rect 674649 303920 676292 303922
rect 674649 303864 674654 303920
rect 674710 303864 676292 303920
rect 674649 303862 676292 303864
rect 674649 303859 674715 303862
rect 676029 303514 676095 303517
rect 676029 303512 676292 303514
rect 676029 303456 676034 303512
rect 676090 303456 676292 303512
rect 676029 303454 676292 303456
rect 676029 303451 676095 303454
rect 651373 303378 651439 303381
rect 649950 303376 651439 303378
rect 649950 303320 651378 303376
rect 651434 303320 651439 303376
rect 649950 303318 651439 303320
rect 649950 302776 650010 303318
rect 651373 303315 651439 303318
rect 675886 302636 675892 302700
rect 675956 302698 675962 302700
rect 676262 302698 676322 303076
rect 675956 302668 676322 302698
rect 675956 302638 676292 302668
rect 675956 302636 675962 302638
rect 671521 302290 671587 302293
rect 671521 302288 676292 302290
rect 671521 302232 671526 302288
rect 671582 302232 676292 302288
rect 671521 302230 676292 302232
rect 671521 302227 671587 302230
rect 652293 302154 652359 302157
rect 649950 302152 652359 302154
rect 649950 302096 652298 302152
rect 652354 302096 652359 302152
rect 649950 302094 652359 302096
rect 41321 301610 41387 301613
rect 41278 301608 41387 301610
rect 41278 301552 41326 301608
rect 41382 301552 41387 301608
rect 649950 301594 650010 302094
rect 652293 302091 652359 302094
rect 669865 302018 669931 302021
rect 676029 302018 676095 302021
rect 669865 302016 676095 302018
rect 669865 301960 669870 302016
rect 669926 301960 676034 302016
rect 676090 301960 676095 302016
rect 669865 301958 676095 301960
rect 669865 301955 669931 301958
rect 676029 301955 676095 301958
rect 676581 301612 676647 301613
rect 676581 301608 676628 301612
rect 676692 301610 676698 301612
rect 41278 301547 41387 301552
rect 676581 301552 676586 301608
rect 676581 301548 676628 301552
rect 676692 301550 676738 301610
rect 676692 301548 676698 301550
rect 676581 301547 676647 301548
rect 41278 301308 41338 301547
rect 41137 300930 41203 300933
rect 41124 300928 41203 300930
rect 41124 300872 41142 300928
rect 41198 300872 41203 300928
rect 41124 300870 41203 300872
rect 41137 300867 41203 300870
rect 651465 300658 651531 300661
rect 649950 300656 651531 300658
rect 649950 300600 651470 300656
rect 651526 300600 651531 300656
rect 649950 300598 651531 300600
rect 45185 300522 45251 300525
rect 41492 300520 45251 300522
rect 41492 300464 45190 300520
rect 45246 300464 45251 300520
rect 41492 300462 45251 300464
rect 45185 300459 45251 300462
rect 649950 300412 650010 300598
rect 651465 300595 651531 300598
rect 44582 300114 44588 300116
rect 41492 300054 44588 300114
rect 44582 300052 44588 300054
rect 44652 300052 44658 300116
rect 44357 299706 44423 299709
rect 41492 299704 44423 299706
rect 41492 299648 44362 299704
rect 44418 299648 44423 299704
rect 41492 299646 44423 299648
rect 44357 299643 44423 299646
rect 42742 299298 42748 299300
rect 41492 299238 42748 299298
rect 42742 299236 42748 299238
rect 42812 299236 42818 299300
rect 44173 299026 44239 299029
rect 41784 299024 44239 299026
rect 41784 298968 44178 299024
rect 44234 298968 44239 299024
rect 41784 298966 44239 298968
rect 41784 298890 41844 298966
rect 44173 298963 44239 298966
rect 41492 298830 41844 298890
rect 42149 298754 42215 298757
rect 63125 298754 63191 298757
rect 42149 298752 63191 298754
rect 42149 298696 42154 298752
rect 42210 298696 63130 298752
rect 63186 298696 63191 298752
rect 42149 298694 63191 298696
rect 649950 298754 650010 299230
rect 651465 298754 651531 298757
rect 649950 298752 651531 298754
rect 649950 298696 651470 298752
rect 651526 298696 651531 298752
rect 649950 298694 651531 298696
rect 42149 298691 42215 298694
rect 63125 298691 63191 298694
rect 651465 298691 651531 298694
rect 44766 298482 44772 298484
rect 41492 298422 44772 298482
rect 44766 298420 44772 298422
rect 44836 298420 44842 298484
rect 44633 298074 44699 298077
rect 41492 298072 44699 298074
rect 41492 298016 44638 298072
rect 44694 298016 44699 298072
rect 41492 298014 44699 298016
rect 44633 298011 44699 298014
rect 44398 297666 44404 297668
rect 41492 297606 44404 297666
rect 44398 297604 44404 297606
rect 44468 297604 44474 297668
rect 649950 297530 650010 298048
rect 652385 297530 652451 297533
rect 649950 297528 652451 297530
rect 649950 297472 652390 297528
rect 652446 297472 652451 297528
rect 649950 297470 652451 297472
rect 652385 297467 652451 297470
rect 42333 297394 42399 297397
rect 62481 297394 62547 297397
rect 42333 297392 62547 297394
rect 42333 297336 42338 297392
rect 42394 297336 62486 297392
rect 62542 297336 62547 297392
rect 42333 297334 62547 297336
rect 42333 297331 42399 297334
rect 62481 297331 62547 297334
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 676857 297394 676923 297397
rect 675772 297392 676923 297394
rect 675772 297336 676862 297392
rect 676918 297336 676923 297392
rect 675772 297334 676923 297336
rect 675772 297332 675778 297334
rect 676857 297331 676923 297334
rect 41492 297198 41844 297258
rect 41784 297122 41844 297198
rect 43161 297122 43227 297125
rect 41784 297120 43227 297122
rect 41784 297064 43166 297120
rect 43222 297064 43227 297120
rect 41784 297062 43227 297064
rect 43161 297059 43227 297062
rect 42190 296850 42196 296852
rect 41492 296790 42196 296850
rect 42190 296788 42196 296790
rect 42260 296788 42266 296852
rect 649950 296850 650010 296866
rect 652201 296850 652267 296853
rect 649950 296848 652267 296850
rect 649950 296792 652206 296848
rect 652262 296792 652267 296848
rect 649950 296790 652267 296792
rect 652201 296787 652267 296790
rect 675518 296516 675524 296580
rect 675588 296578 675594 296580
rect 676029 296578 676095 296581
rect 675588 296576 676095 296578
rect 675588 296520 676034 296576
rect 676090 296520 676095 296576
rect 675588 296518 676095 296520
rect 675588 296516 675594 296518
rect 676029 296515 676095 296518
rect 41137 296442 41203 296445
rect 41124 296440 41203 296442
rect 41124 296384 41142 296440
rect 41198 296384 41203 296440
rect 41124 296382 41203 296384
rect 41137 296379 41203 296382
rect 42793 296034 42859 296037
rect 41492 296032 42859 296034
rect 41492 295976 42798 296032
rect 42854 295976 42859 296032
rect 41492 295974 42859 295976
rect 42793 295971 42859 295974
rect 62113 295762 62179 295765
rect 670969 295762 671035 295765
rect 675569 295762 675635 295765
rect 62113 295760 64706 295762
rect 62113 295704 62118 295760
rect 62174 295704 64706 295760
rect 62113 295702 64706 295704
rect 62113 295699 62179 295702
rect 64646 295684 64706 295702
rect 670969 295760 675635 295762
rect 670969 295704 670974 295760
rect 671030 295704 675574 295760
rect 675630 295704 675635 295760
rect 670969 295702 675635 295704
rect 670969 295699 671035 295702
rect 675569 295699 675635 295702
rect 42006 295626 42012 295628
rect 41492 295566 42012 295626
rect 42006 295564 42012 295566
rect 42076 295564 42082 295628
rect 649950 295354 650010 295684
rect 651649 295354 651715 295357
rect 649950 295352 651715 295354
rect 649950 295296 651654 295352
rect 651710 295296 651715 295352
rect 649950 295294 651715 295296
rect 651649 295291 651715 295294
rect 41321 295218 41387 295221
rect 41308 295216 41387 295218
rect 41308 295160 41326 295216
rect 41382 295160 41387 295216
rect 41308 295158 41387 295160
rect 41321 295155 41387 295158
rect 33777 294810 33843 294813
rect 33764 294808 33843 294810
rect 33764 294752 33782 294808
rect 33838 294752 33843 294808
rect 33764 294750 33843 294752
rect 33777 294747 33843 294750
rect 675753 294674 675819 294677
rect 676438 294674 676444 294676
rect 675753 294672 676444 294674
rect 675753 294616 675758 294672
rect 675814 294616 676444 294672
rect 675753 294614 676444 294616
rect 675753 294611 675819 294614
rect 676438 294612 676444 294614
rect 676508 294612 676514 294676
rect 41822 294402 41828 294404
rect 41492 294342 41828 294402
rect 41822 294340 41828 294342
rect 41892 294340 41898 294404
rect 62113 294130 62179 294133
rect 64646 294130 64706 294502
rect 649950 294266 650010 294502
rect 651465 294266 651531 294269
rect 649950 294264 651531 294266
rect 649950 294208 651470 294264
rect 651526 294208 651531 294264
rect 649950 294206 651531 294208
rect 651465 294203 651531 294206
rect 62113 294128 64706 294130
rect 62113 294072 62118 294128
rect 62174 294072 64706 294128
rect 62113 294070 64706 294072
rect 62113 294067 62179 294070
rect 32397 293994 32463 293997
rect 32397 293992 32476 293994
rect 32397 293936 32402 293992
rect 32458 293936 32476 293992
rect 32397 293934 32476 293936
rect 32397 293931 32463 293934
rect 660573 293858 660639 293861
rect 670969 293858 671035 293861
rect 660573 293856 671035 293858
rect 660573 293800 660578 293856
rect 660634 293800 670974 293856
rect 671030 293800 671035 293856
rect 660573 293798 671035 293800
rect 660573 293795 660639 293798
rect 670969 293795 671035 293798
rect 41321 293586 41387 293589
rect 41308 293584 41387 293586
rect 41308 293528 41326 293584
rect 41382 293528 41387 293584
rect 41308 293526 41387 293528
rect 41321 293523 41387 293526
rect 42977 293178 43043 293181
rect 41492 293176 43043 293178
rect 41492 293120 42982 293176
rect 43038 293120 43043 293176
rect 41492 293118 43043 293120
rect 42977 293115 43043 293118
rect 43345 292770 43411 292773
rect 41492 292768 43411 292770
rect 41492 292712 43350 292768
rect 43406 292712 43411 292768
rect 41492 292710 43411 292712
rect 43345 292707 43411 292710
rect 62297 292770 62363 292773
rect 64646 292770 64706 293320
rect 649950 293042 650010 293320
rect 651465 293042 651531 293045
rect 649950 293040 651531 293042
rect 649950 292984 651470 293040
rect 651526 292984 651531 293040
rect 649950 292982 651531 292984
rect 651465 292979 651531 292982
rect 62297 292768 64706 292770
rect 62297 292712 62302 292768
rect 62358 292712 64706 292768
rect 62297 292710 64706 292712
rect 62297 292707 62363 292710
rect 45001 292634 45067 292637
rect 45461 292634 45527 292637
rect 45001 292632 45527 292634
rect 40718 292528 40724 292592
rect 40788 292528 40794 292592
rect 45001 292576 45006 292632
rect 45062 292576 45466 292632
rect 45522 292576 45527 292632
rect 45001 292574 45527 292576
rect 45001 292571 45067 292574
rect 45461 292571 45527 292574
rect 40726 292332 40786 292528
rect 62113 292498 62179 292501
rect 62113 292496 64706 292498
rect 62113 292440 62118 292496
rect 62174 292440 64706 292496
rect 62113 292438 64706 292440
rect 62113 292435 62179 292438
rect 64646 292138 64706 292438
rect 675569 292228 675635 292229
rect 675518 292164 675524 292228
rect 675588 292226 675635 292228
rect 675588 292224 675680 292226
rect 675630 292168 675680 292224
rect 675588 292166 675680 292168
rect 675588 292164 675635 292166
rect 675569 292163 675635 292164
rect 41492 291894 41844 291954
rect 41784 291820 41844 291894
rect 41784 291758 41828 291820
rect 41822 291756 41828 291758
rect 41892 291756 41898 291820
rect 45185 291546 45251 291549
rect 41492 291544 45251 291546
rect 41492 291488 45190 291544
rect 45246 291488 45251 291544
rect 41492 291486 45251 291488
rect 649950 291546 650010 292138
rect 651649 291818 651715 291821
rect 673821 291818 673887 291821
rect 651649 291816 673887 291818
rect 651649 291760 651654 291816
rect 651710 291760 673826 291816
rect 673882 291760 673887 291816
rect 651649 291758 673887 291760
rect 651649 291755 651715 291758
rect 673821 291755 673887 291758
rect 652109 291546 652175 291549
rect 649950 291544 652175 291546
rect 649950 291488 652114 291544
rect 652170 291488 652175 291544
rect 649950 291486 652175 291488
rect 45185 291483 45251 291486
rect 652109 291483 652175 291486
rect 673545 291546 673611 291549
rect 675385 291546 675451 291549
rect 673545 291544 675451 291546
rect 673545 291488 673550 291544
rect 673606 291488 675390 291544
rect 675446 291488 675451 291544
rect 673545 291486 675451 291488
rect 673545 291483 673611 291486
rect 675385 291483 675451 291486
rect 50521 291138 50587 291141
rect 41492 291136 50587 291138
rect 41492 291080 50526 291136
rect 50582 291080 50587 291136
rect 41492 291078 50587 291080
rect 50521 291075 50587 291078
rect 62481 291002 62547 291005
rect 675753 291002 675819 291005
rect 676622 291002 676628 291004
rect 62481 291000 64154 291002
rect 62481 290944 62486 291000
rect 62542 290986 64154 291000
rect 675753 291000 676628 291002
rect 62542 290944 64676 290986
rect 62481 290942 64676 290944
rect 62481 290939 62547 290942
rect 64094 290926 64676 290942
rect 47577 290730 47643 290733
rect 41492 290728 47643 290730
rect 41492 290672 47582 290728
rect 47638 290672 47643 290728
rect 41492 290670 47643 290672
rect 47577 290667 47643 290670
rect 649950 290458 650010 290956
rect 675753 290944 675758 291000
rect 675814 290944 676628 291000
rect 675753 290942 676628 290944
rect 675753 290939 675819 290942
rect 676622 290940 676628 290942
rect 676692 290940 676698 291004
rect 651465 290458 651531 290461
rect 649950 290456 651531 290458
rect 649950 290400 651470 290456
rect 651526 290400 651531 290456
rect 649950 290398 651531 290400
rect 651465 290395 651531 290398
rect 39941 290322 40007 290325
rect 39941 290320 40020 290322
rect 39941 290264 39946 290320
rect 40002 290264 40020 290320
rect 39941 290262 40020 290264
rect 39941 290259 40007 290262
rect 41822 289988 41828 290052
rect 41892 290050 41898 290052
rect 42190 290050 42196 290052
rect 41892 289990 42196 290050
rect 41892 289988 41898 289990
rect 42190 289988 42196 289990
rect 42260 289988 42266 290052
rect 63125 289778 63191 289781
rect 63125 289776 64706 289778
rect 63125 289720 63130 289776
rect 63186 289720 64706 289776
rect 63125 289718 64706 289720
rect 63125 289715 63191 289718
rect 649950 289234 650010 289774
rect 651649 289234 651715 289237
rect 649950 289232 651715 289234
rect 649950 289176 651654 289232
rect 651710 289176 651715 289232
rect 649950 289174 651715 289176
rect 651649 289171 651715 289174
rect 651465 288690 651531 288693
rect 649950 288688 651531 288690
rect 649950 288632 651470 288688
rect 651526 288632 651531 288688
rect 649950 288630 651531 288632
rect 649950 288592 650010 288630
rect 651465 288627 651531 288630
rect 62205 288554 62271 288557
rect 64646 288554 64706 288592
rect 62205 288552 64706 288554
rect 62205 288496 62210 288552
rect 62266 288496 64706 288552
rect 62205 288494 64706 288496
rect 62205 288491 62271 288494
rect 673177 287874 673243 287877
rect 675109 287874 675175 287877
rect 673177 287872 675175 287874
rect 673177 287816 673182 287872
rect 673238 287816 675114 287872
rect 675170 287816 675175 287872
rect 673177 287814 675175 287816
rect 673177 287811 673243 287814
rect 675109 287811 675175 287814
rect 651649 287738 651715 287741
rect 651649 287736 663810 287738
rect 651649 287680 651654 287736
rect 651710 287680 663810 287736
rect 651649 287678 663810 287680
rect 651649 287675 651715 287678
rect 663750 287602 663810 287678
rect 673637 287602 673703 287605
rect 663750 287600 673703 287602
rect 663750 287544 673642 287600
rect 673698 287544 673703 287600
rect 663750 287542 673703 287544
rect 673637 287539 673703 287542
rect 651465 287466 651531 287469
rect 649766 287464 651531 287466
rect 62389 287194 62455 287197
rect 64646 287194 64706 287410
rect 649766 287408 651470 287464
rect 651526 287408 651531 287464
rect 649766 287406 651531 287408
rect 651465 287403 651531 287406
rect 62389 287192 64706 287194
rect 62389 287136 62394 287192
rect 62450 287136 64706 287192
rect 62389 287134 64706 287136
rect 62389 287131 62455 287134
rect 675753 287058 675819 287061
rect 676254 287058 676260 287060
rect 675753 287056 676260 287058
rect 675753 287000 675758 287056
rect 675814 287000 676260 287056
rect 675753 286998 676260 287000
rect 675753 286995 675819 286998
rect 676254 286996 676260 286998
rect 676324 286996 676330 287060
rect 62113 285970 62179 285973
rect 64646 285970 64706 286228
rect 62113 285968 64706 285970
rect 62113 285912 62118 285968
rect 62174 285912 64706 285968
rect 62113 285910 64706 285912
rect 649950 285970 650010 286228
rect 651465 285970 651531 285973
rect 649950 285968 651531 285970
rect 649950 285912 651470 285968
rect 651526 285912 651531 285968
rect 649950 285910 651531 285912
rect 62113 285907 62179 285910
rect 651465 285907 651531 285910
rect 672533 285562 672599 285565
rect 675109 285562 675175 285565
rect 672533 285560 675175 285562
rect 672533 285504 672538 285560
rect 672594 285504 675114 285560
rect 675170 285504 675175 285560
rect 672533 285502 675175 285504
rect 672533 285499 672599 285502
rect 675109 285499 675175 285502
rect 32397 284882 32463 284885
rect 41822 284882 41828 284884
rect 32397 284880 41828 284882
rect 32397 284824 32402 284880
rect 32458 284824 41828 284880
rect 32397 284822 41828 284824
rect 32397 284819 32463 284822
rect 41822 284820 41828 284822
rect 41892 284820 41898 284884
rect 63217 284610 63283 284613
rect 64646 284610 64706 285046
rect 649950 284746 650010 285046
rect 651465 284746 651531 284749
rect 649950 284744 651531 284746
rect 649950 284688 651470 284744
rect 651526 284688 651531 284744
rect 649950 284686 651531 284688
rect 651465 284683 651531 284686
rect 63217 284608 64706 284610
rect 63217 284552 63222 284608
rect 63278 284552 64706 284608
rect 63217 284550 64706 284552
rect 63217 284547 63283 284550
rect 62113 283250 62179 283253
rect 64646 283250 64706 283864
rect 649950 283386 650010 283864
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 651465 283386 651531 283389
rect 649950 283384 651531 283386
rect 649950 283328 651470 283384
rect 651526 283328 651531 283384
rect 649950 283326 651531 283328
rect 651465 283323 651531 283326
rect 62113 283248 64706 283250
rect 62113 283192 62118 283248
rect 62174 283192 64706 283248
rect 62113 283190 64706 283192
rect 62113 283187 62179 283190
rect 675753 282706 675819 282709
rect 676070 282706 676076 282708
rect 675753 282704 676076 282706
rect 62849 282162 62915 282165
rect 64646 282162 64706 282682
rect 62849 282160 64706 282162
rect 62849 282104 62854 282160
rect 62910 282104 64706 282160
rect 62849 282102 64706 282104
rect 649950 282162 650010 282682
rect 675753 282648 675758 282704
rect 675814 282648 676076 282704
rect 675753 282646 676076 282648
rect 675753 282643 675819 282646
rect 676070 282644 676076 282646
rect 676140 282644 676146 282708
rect 652017 282162 652083 282165
rect 649950 282160 652083 282162
rect 649950 282104 652022 282160
rect 652078 282104 652083 282160
rect 649950 282102 652083 282104
rect 62849 282099 62915 282102
rect 652017 282099 652083 282102
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 42425 281482 42491 281485
rect 45001 281482 45067 281485
rect 42425 281480 45067 281482
rect 42425 281424 42430 281480
rect 42486 281424 45006 281480
rect 45062 281424 45067 281480
rect 42425 281422 45067 281424
rect 42425 281419 42491 281422
rect 45001 281419 45067 281422
rect 62113 280938 62179 280941
rect 64646 280938 64706 281500
rect 62113 280936 64706 280938
rect 62113 280880 62118 280936
rect 62174 280880 64706 280936
rect 62113 280878 64706 280880
rect 649950 280938 650010 281500
rect 651465 280938 651531 280941
rect 649950 280936 651531 280938
rect 649950 280880 651470 280936
rect 651526 280880 651531 280936
rect 649950 280878 651531 280880
rect 62113 280875 62179 280878
rect 651465 280875 651531 280878
rect 63125 280394 63191 280397
rect 652385 280394 652451 280397
rect 63125 280392 64706 280394
rect 63125 280336 63130 280392
rect 63186 280336 64706 280392
rect 63125 280334 64706 280336
rect 63125 280331 63191 280334
rect 64646 280318 64706 280334
rect 649950 280392 652451 280394
rect 649950 280336 652390 280392
rect 652446 280336 652451 280392
rect 649950 280334 652451 280336
rect 649950 280318 650010 280334
rect 652385 280331 652451 280334
rect 652569 279442 652635 279445
rect 676857 279442 676923 279445
rect 652569 279440 676923 279442
rect 652569 279384 652574 279440
rect 652630 279384 676862 279440
rect 676918 279384 676923 279440
rect 652569 279382 676923 279384
rect 652569 279379 652635 279382
rect 676857 279379 676923 279382
rect 62062 278836 62068 278900
rect 62132 278898 62138 278900
rect 62941 278898 63007 278901
rect 62132 278896 63007 278898
rect 62132 278840 62946 278896
rect 63002 278840 63007 278896
rect 62132 278838 63007 278840
rect 62132 278836 62138 278838
rect 62941 278835 63007 278838
rect 671705 278626 671771 278629
rect 672901 278626 672967 278629
rect 671705 278624 672967 278626
rect 671705 278568 671710 278624
rect 671766 278568 672906 278624
rect 672962 278568 672967 278624
rect 671705 278566 672967 278568
rect 671705 278563 671771 278566
rect 672901 278563 672967 278566
rect 42057 278490 42123 278493
rect 45185 278490 45251 278493
rect 42057 278488 45251 278490
rect 42057 278432 42062 278488
rect 42118 278432 45190 278488
rect 45246 278432 45251 278488
rect 42057 278430 45251 278432
rect 42057 278427 42123 278430
rect 45185 278427 45251 278430
rect 59997 278354 60063 278357
rect 674833 278354 674899 278357
rect 59997 278352 674899 278354
rect 59997 278296 60002 278352
rect 60058 278296 674838 278352
rect 674894 278296 674899 278352
rect 59997 278294 674899 278296
rect 59997 278291 60063 278294
rect 674833 278291 674899 278294
rect 57237 278082 57303 278085
rect 675477 278082 675543 278085
rect 57237 278080 675543 278082
rect 57237 278024 57242 278080
rect 57298 278024 675482 278080
rect 675538 278024 675543 278080
rect 57237 278022 675543 278024
rect 57237 278019 57303 278022
rect 675477 278019 675543 278022
rect 42149 277946 42215 277949
rect 43437 277946 43503 277949
rect 42149 277944 43503 277946
rect 42149 277888 42154 277944
rect 42210 277888 43442 277944
rect 43498 277888 43503 277944
rect 42149 277886 43503 277888
rect 42149 277883 42215 277886
rect 43437 277883 43503 277886
rect 60181 277402 60247 277405
rect 675293 277402 675359 277405
rect 60181 277400 675359 277402
rect 60181 277344 60186 277400
rect 60242 277344 675298 277400
rect 675354 277344 675359 277400
rect 60181 277342 675359 277344
rect 60181 277339 60247 277342
rect 675293 277339 675359 277342
rect 40902 277068 40908 277132
rect 40972 277130 40978 277132
rect 41781 277130 41847 277133
rect 40972 277128 41847 277130
rect 40972 277072 41786 277128
rect 41842 277072 41847 277128
rect 40972 277070 41847 277072
rect 40972 277068 40978 277070
rect 41781 277067 41847 277070
rect 42609 275906 42675 275909
rect 57421 275906 57487 275909
rect 42609 275904 57487 275906
rect 42609 275848 42614 275904
rect 42670 275848 57426 275904
rect 57482 275848 57487 275904
rect 42609 275846 57487 275848
rect 42609 275843 42675 275846
rect 57421 275843 57487 275846
rect 40718 274212 40724 274276
rect 40788 274274 40794 274276
rect 41781 274274 41847 274277
rect 40788 274272 41847 274274
rect 40788 274216 41786 274272
rect 41842 274216 41847 274272
rect 40788 274214 41847 274216
rect 40788 274212 40794 274214
rect 41781 274211 41847 274214
rect 539317 274002 539383 274005
rect 545941 274002 546007 274005
rect 539317 274000 546007 274002
rect 539317 273944 539322 274000
rect 539378 273944 545946 274000
rect 546002 273944 546007 274000
rect 539317 273942 546007 273944
rect 539317 273939 539383 273942
rect 545941 273939 546007 273942
rect 674833 273866 674899 273869
rect 675334 273866 675340 273868
rect 674833 273864 675340 273866
rect 674833 273808 674838 273864
rect 674894 273808 675340 273864
rect 674833 273806 675340 273808
rect 674833 273803 674899 273806
rect 675334 273804 675340 273806
rect 675404 273804 675410 273868
rect 42333 273186 42399 273189
rect 43621 273186 43687 273189
rect 42333 273184 43687 273186
rect 42333 273128 42338 273184
rect 42394 273128 43626 273184
rect 43682 273128 43687 273184
rect 42333 273126 43687 273128
rect 42333 273123 42399 273126
rect 43621 273123 43687 273126
rect 41781 273052 41847 273053
rect 41781 273048 41828 273052
rect 41892 273050 41898 273052
rect 41781 272992 41786 273048
rect 41781 272988 41828 272992
rect 41892 272990 41938 273050
rect 41892 272988 41898 272990
rect 41781 272987 41847 272988
rect 536373 272914 536439 272917
rect 538121 272914 538187 272917
rect 536373 272912 538187 272914
rect 536373 272856 536378 272912
rect 536434 272856 538126 272912
rect 538182 272856 538187 272912
rect 536373 272854 538187 272856
rect 536373 272851 536439 272854
rect 538121 272851 538187 272854
rect 459369 272642 459435 272645
rect 466085 272642 466151 272645
rect 459369 272640 466151 272642
rect 459369 272584 459374 272640
rect 459430 272584 466090 272640
rect 466146 272584 466151 272640
rect 459369 272582 466151 272584
rect 459369 272579 459435 272582
rect 466085 272579 466151 272582
rect 537937 272642 538003 272645
rect 538673 272642 538739 272645
rect 537937 272640 538739 272642
rect 537937 272584 537942 272640
rect 537998 272584 538678 272640
rect 538734 272584 538739 272640
rect 537937 272582 538739 272584
rect 537937 272579 538003 272582
rect 538673 272579 538739 272582
rect 470685 272506 470751 272509
rect 466410 272504 470751 272506
rect 466410 272448 470690 272504
rect 470746 272448 470751 272504
rect 466410 272446 470751 272448
rect 41781 272372 41847 272373
rect 41781 272368 41828 272372
rect 41892 272370 41898 272372
rect 464705 272370 464771 272373
rect 466410 272370 466470 272446
rect 470685 272443 470751 272446
rect 41781 272312 41786 272368
rect 41781 272308 41828 272312
rect 41892 272310 41938 272370
rect 464705 272368 466470 272370
rect 464705 272312 464710 272368
rect 464766 272312 466470 272368
rect 464705 272310 466470 272312
rect 538213 272370 538279 272373
rect 547689 272370 547755 272373
rect 538213 272368 547755 272370
rect 538213 272312 538218 272368
rect 538274 272312 547694 272368
rect 547750 272312 547755 272368
rect 538213 272310 547755 272312
rect 41892 272308 41898 272310
rect 41781 272307 41847 272308
rect 464705 272307 464771 272310
rect 538213 272307 538279 272310
rect 547689 272307 547755 272310
rect 500861 272234 500927 272237
rect 504541 272234 504607 272237
rect 500861 272232 504607 272234
rect 500861 272176 500866 272232
rect 500922 272176 504546 272232
rect 504602 272176 504607 272232
rect 500861 272174 504607 272176
rect 500861 272171 500927 272174
rect 504541 272171 504607 272174
rect 547505 272098 547571 272101
rect 547873 272098 547939 272101
rect 547505 272096 547939 272098
rect 547505 272040 547510 272096
rect 547566 272040 547878 272096
rect 547934 272040 547939 272096
rect 547505 272038 547939 272040
rect 547505 272035 547571 272038
rect 547873 272035 547939 272038
rect 470593 271962 470659 271965
rect 478045 271962 478111 271965
rect 470593 271960 478111 271962
rect 470593 271904 470598 271960
rect 470654 271904 478050 271960
rect 478106 271904 478111 271960
rect 470593 271902 478111 271904
rect 470593 271899 470659 271902
rect 478045 271899 478111 271902
rect 479517 271962 479583 271965
rect 483013 271962 483079 271965
rect 479517 271960 483079 271962
rect 479517 271904 479522 271960
rect 479578 271904 483018 271960
rect 483074 271904 483079 271960
rect 479517 271902 483079 271904
rect 479517 271899 479583 271902
rect 483013 271899 483079 271902
rect 501597 271962 501663 271965
rect 504541 271962 504607 271965
rect 501597 271960 504607 271962
rect 501597 271904 501602 271960
rect 501658 271904 504546 271960
rect 504602 271904 504607 271960
rect 501597 271902 504607 271904
rect 501597 271899 501663 271902
rect 504541 271899 504607 271902
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 136633 270466 136699 270469
rect 137829 270466 137895 270469
rect 136633 270464 137895 270466
rect 136633 270408 136638 270464
rect 136694 270408 137834 270464
rect 137890 270408 137895 270464
rect 136633 270406 137895 270408
rect 136633 270403 136699 270406
rect 137829 270403 137895 270406
rect 530393 270194 530459 270197
rect 534073 270194 534139 270197
rect 530393 270192 534139 270194
rect 530393 270136 530398 270192
rect 530454 270136 534078 270192
rect 534134 270136 534139 270192
rect 530393 270134 534139 270136
rect 530393 270131 530459 270134
rect 534073 270131 534139 270134
rect 509233 269922 509299 269925
rect 516501 269922 516567 269925
rect 509233 269920 516567 269922
rect 509233 269864 509238 269920
rect 509294 269864 516506 269920
rect 516562 269864 516567 269920
rect 509233 269862 516567 269864
rect 509233 269859 509299 269862
rect 516501 269859 516567 269862
rect 537845 269922 537911 269925
rect 538305 269922 538371 269925
rect 537845 269920 538371 269922
rect 537845 269864 537850 269920
rect 537906 269864 538310 269920
rect 538366 269864 538371 269920
rect 537845 269862 538371 269864
rect 537845 269859 537911 269862
rect 538305 269859 538371 269862
rect 40534 269724 40540 269788
rect 40604 269786 40610 269788
rect 41781 269786 41847 269789
rect 40604 269784 41847 269786
rect 40604 269728 41786 269784
rect 41842 269728 41847 269784
rect 40604 269726 41847 269728
rect 40604 269724 40610 269726
rect 41781 269723 41847 269726
rect 43437 269786 43503 269789
rect 62389 269786 62455 269789
rect 43437 269784 62455 269786
rect 43437 269728 43442 269784
rect 43498 269728 62394 269784
rect 62450 269728 62455 269784
rect 43437 269726 62455 269728
rect 43437 269723 43503 269726
rect 62389 269723 62455 269726
rect 509141 269514 509207 269517
rect 509877 269514 509943 269517
rect 509141 269512 509943 269514
rect 509141 269456 509146 269512
rect 509202 269456 509882 269512
rect 509938 269456 509943 269512
rect 509141 269454 509943 269456
rect 509141 269451 509207 269454
rect 509877 269451 509943 269454
rect 676262 268562 676322 268668
rect 676857 268562 676923 268565
rect 663750 268502 676322 268562
rect 676814 268560 676923 268562
rect 676814 268504 676862 268560
rect 676918 268504 676923 268560
rect 658917 268154 658983 268157
rect 663750 268154 663810 268502
rect 676814 268499 676923 268504
rect 676814 268260 676874 268499
rect 658917 268152 663810 268154
rect 658917 268096 658922 268152
rect 658978 268096 663810 268152
rect 658917 268094 663810 268096
rect 673821 268154 673887 268157
rect 676213 268154 676279 268157
rect 673821 268152 676279 268154
rect 673821 268096 673826 268152
rect 673882 268096 676218 268152
rect 676274 268096 676279 268152
rect 673821 268094 676279 268096
rect 658917 268091 658983 268094
rect 673821 268091 673887 268094
rect 676213 268091 676279 268094
rect 676262 267749 676322 267852
rect 42149 267746 42215 267749
rect 60365 267746 60431 267749
rect 42149 267744 60431 267746
rect 42149 267688 42154 267744
rect 42210 267688 60370 267744
rect 60426 267688 60431 267744
rect 42149 267686 60431 267688
rect 42149 267683 42215 267686
rect 60365 267683 60431 267686
rect 676213 267744 676322 267749
rect 676213 267688 676218 267744
rect 676274 267688 676322 267744
rect 676213 267686 676322 267688
rect 676213 267683 676279 267686
rect 674373 267474 674439 267477
rect 674373 267472 676292 267474
rect 674373 267416 674378 267472
rect 674434 267416 676292 267472
rect 674373 267414 676292 267416
rect 674373 267411 674439 267414
rect 674281 267066 674347 267069
rect 674281 267064 676292 267066
rect 674281 267008 674286 267064
rect 674342 267008 676292 267064
rect 674281 267006 676292 267008
rect 674281 267003 674347 267006
rect 674097 266658 674163 266661
rect 674097 266656 676292 266658
rect 674097 266600 674102 266656
rect 674158 266600 676292 266656
rect 674097 266598 676292 266600
rect 674097 266595 674163 266598
rect 673177 266114 673243 266117
rect 676262 266114 676322 266220
rect 673177 266112 676322 266114
rect 673177 266056 673182 266112
rect 673238 266056 676322 266112
rect 673177 266054 676322 266056
rect 673177 266051 673243 266054
rect 674649 265842 674715 265845
rect 674649 265840 676292 265842
rect 674649 265784 674654 265840
rect 674710 265784 676292 265840
rect 674649 265782 676292 265784
rect 674649 265779 674715 265782
rect 672533 265298 672599 265301
rect 676262 265298 676322 265404
rect 672533 265296 676322 265298
rect 672533 265240 672538 265296
rect 672594 265240 676322 265296
rect 672533 265238 676322 265240
rect 672533 265235 672599 265238
rect 673361 265026 673427 265029
rect 673361 265024 676292 265026
rect 673361 264968 673366 265024
rect 673422 264968 676292 265024
rect 673361 264966 676292 264968
rect 673361 264963 673427 264966
rect 53097 264754 53163 264757
rect 675109 264754 675175 264757
rect 53097 264752 675175 264754
rect 53097 264696 53102 264752
rect 53158 264696 675114 264752
rect 675170 264696 675175 264752
rect 53097 264694 675175 264696
rect 53097 264691 53163 264694
rect 675109 264691 675175 264694
rect 673453 264482 673519 264485
rect 676262 264482 676322 264588
rect 673453 264480 676322 264482
rect 673453 264424 673458 264480
rect 673514 264424 676322 264480
rect 673453 264422 676322 264424
rect 673453 264419 673519 264422
rect 676446 264077 676506 264180
rect 676397 264072 676506 264077
rect 676397 264016 676402 264072
rect 676458 264016 676506 264072
rect 676397 264014 676506 264016
rect 676397 264011 676463 264014
rect 671705 263802 671771 263805
rect 671705 263800 673470 263802
rect 671705 263744 671710 263800
rect 671766 263744 673470 263800
rect 671705 263742 673470 263744
rect 671705 263739 671771 263742
rect 673410 263666 673470 263742
rect 676262 263666 676322 263772
rect 673410 263606 676322 263666
rect 673085 263394 673151 263397
rect 673085 263392 676292 263394
rect 673085 263336 673090 263392
rect 673146 263336 676292 263392
rect 673085 263334 676292 263336
rect 673085 263331 673151 263334
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 674649 262578 674715 262581
rect 674649 262576 676292 262578
rect 674649 262520 674654 262576
rect 674710 262520 676292 262576
rect 674649 262518 676292 262520
rect 674649 262515 674715 262518
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 670325 262170 670391 262173
rect 670325 262168 676292 262170
rect 670325 262112 670330 262168
rect 670386 262112 676292 262168
rect 670325 262110 676292 262112
rect 670325 262107 670391 262110
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 676814 261220 676874 261324
rect 676806 261156 676812 261220
rect 676876 261156 676882 261220
rect 674189 260946 674255 260949
rect 674189 260944 676292 260946
rect 674189 260888 674194 260944
rect 674250 260888 676292 260944
rect 674189 260886 676292 260888
rect 674189 260883 674255 260886
rect 674833 260538 674899 260541
rect 674833 260536 676292 260538
rect 674833 260480 674838 260536
rect 674894 260480 676292 260536
rect 674833 260478 676292 260480
rect 674833 260475 674899 260478
rect 674189 260130 674255 260133
rect 674189 260128 676292 260130
rect 674189 260072 674194 260128
rect 674250 260072 676292 260128
rect 674189 260070 676292 260072
rect 674189 260067 674255 260070
rect 554313 259994 554379 259997
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 671245 259586 671311 259589
rect 676262 259586 676322 259692
rect 671245 259584 676322 259586
rect 671245 259528 671250 259584
rect 671306 259528 676322 259584
rect 671245 259526 676322 259528
rect 671245 259523 671311 259526
rect 672901 259314 672967 259317
rect 672901 259312 676292 259314
rect 672901 259256 672906 259312
rect 672962 259256 676292 259312
rect 672901 259254 676292 259256
rect 672901 259251 672967 259254
rect 674373 258906 674439 258909
rect 674373 258904 676292 258906
rect 674373 258848 674378 258904
rect 674434 258848 676292 258904
rect 674373 258846 676292 258848
rect 674373 258843 674439 258846
rect 670141 258498 670207 258501
rect 670141 258496 676292 258498
rect 670141 258440 670146 258496
rect 670202 258440 676292 258496
rect 670141 258438 676292 258440
rect 670141 258435 670207 258438
rect 44817 258090 44883 258093
rect 675477 258092 675543 258093
rect 675477 258090 675524 258092
rect 41492 258088 44883 258090
rect 41492 258032 44822 258088
rect 44878 258032 44883 258088
rect 41492 258030 44883 258032
rect 675396 258088 675524 258090
rect 675588 258090 675594 258092
rect 675396 258032 675482 258088
rect 675588 258060 676292 258090
rect 675396 258030 675524 258032
rect 44817 258027 44883 258030
rect 675477 258028 675524 258030
rect 675588 258030 676322 258060
rect 675588 258028 675594 258030
rect 675477 258027 675543 258028
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 46381 257682 46447 257685
rect 41492 257680 46447 257682
rect 41492 257624 46386 257680
rect 46442 257624 46447 257680
rect 676262 257652 676322 258030
rect 41492 257622 46447 257624
rect 46381 257619 46447 257622
rect 670693 257274 670759 257277
rect 670693 257272 676292 257274
rect 35758 257141 35818 257244
rect 670693 257216 670698 257272
rect 670754 257216 676292 257272
rect 670693 257214 676292 257216
rect 670693 257211 670759 257214
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 40493 257138 40559 257141
rect 43345 257138 43411 257141
rect 40493 257136 43411 257138
rect 40493 257080 40498 257136
rect 40554 257080 43350 257136
rect 43406 257080 43411 257136
rect 40493 257078 43411 257080
rect 40493 257075 40559 257078
rect 43345 257075 43411 257078
rect 44357 256866 44423 256869
rect 41492 256864 44423 256866
rect 41492 256808 44362 256864
rect 44418 256808 44423 256864
rect 41492 256806 44423 256808
rect 44357 256803 44423 256806
rect 35574 256325 35634 256428
rect 35574 256320 35683 256325
rect 35574 256264 35622 256320
rect 35678 256264 35683 256320
rect 35574 256262 35683 256264
rect 35617 256259 35683 256262
rect 40217 256322 40283 256325
rect 42977 256322 43043 256325
rect 40217 256320 43043 256322
rect 40217 256264 40222 256320
rect 40278 256264 42982 256320
rect 43038 256264 43043 256320
rect 40217 256262 43043 256264
rect 40217 256259 40283 256262
rect 42977 256259 43043 256262
rect 671613 256322 671679 256325
rect 674833 256322 674899 256325
rect 671613 256320 674899 256322
rect 671613 256264 671618 256320
rect 671674 256264 674838 256320
rect 674894 256264 674899 256320
rect 671613 256262 674899 256264
rect 671613 256259 671679 256262
rect 674833 256259 674899 256262
rect 44173 256050 44239 256053
rect 41492 256048 44239 256050
rect 41492 255992 44178 256048
rect 44234 255992 44239 256048
rect 41492 255990 44239 255992
rect 44173 255987 44239 255990
rect 35801 255914 35867 255917
rect 35758 255912 35867 255914
rect 35758 255856 35806 255912
rect 35862 255856 35867 255912
rect 35758 255851 35867 255856
rect 35758 255612 35818 255851
rect 554497 255642 554563 255645
rect 552460 255640 554563 255642
rect 552460 255584 554502 255640
rect 554558 255584 554563 255640
rect 552460 255582 554563 255584
rect 554497 255579 554563 255582
rect 39573 255506 39639 255509
rect 43069 255506 43135 255509
rect 39573 255504 43135 255506
rect 39573 255448 39578 255504
rect 39634 255448 43074 255504
rect 43130 255448 43135 255504
rect 39573 255446 43135 255448
rect 39573 255443 39639 255446
rect 43069 255443 43135 255446
rect 44633 255234 44699 255237
rect 41492 255232 44699 255234
rect 41492 255176 44638 255232
rect 44694 255176 44699 255232
rect 41492 255174 44699 255176
rect 44633 255171 44699 255174
rect 674833 254962 674899 254965
rect 675845 254962 675911 254965
rect 674833 254960 675911 254962
rect 674833 254904 674838 254960
rect 674894 254904 675850 254960
rect 675906 254904 675911 254960
rect 674833 254902 675911 254904
rect 674833 254899 674899 254902
rect 675845 254899 675911 254902
rect 44265 254826 44331 254829
rect 41492 254824 44331 254826
rect 41492 254768 44270 254824
rect 44326 254768 44331 254824
rect 41492 254766 44331 254768
rect 44265 254763 44331 254766
rect 35758 254285 35818 254388
rect 35758 254280 35867 254285
rect 35758 254224 35806 254280
rect 35862 254224 35867 254280
rect 35758 254222 35867 254224
rect 35801 254219 35867 254222
rect 39849 254282 39915 254285
rect 42885 254282 42951 254285
rect 39849 254280 42951 254282
rect 39849 254224 39854 254280
rect 39910 254224 42890 254280
rect 42946 254224 42951 254280
rect 39849 254222 42951 254224
rect 39849 254219 39915 254222
rect 42885 254219 42951 254222
rect 44909 254010 44975 254013
rect 41492 254008 44975 254010
rect 41492 253952 44914 254008
rect 44970 253952 44975 254008
rect 41492 253950 44975 253952
rect 44909 253947 44975 253950
rect 35574 253469 35634 253572
rect 35574 253464 35683 253469
rect 554405 253466 554471 253469
rect 35574 253408 35622 253464
rect 35678 253408 35683 253464
rect 35574 253406 35683 253408
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 35617 253403 35683 253406
rect 554405 253403 554471 253406
rect 35758 253061 35818 253164
rect 35758 253056 35867 253061
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35758 252998 35867 253000
rect 35801 252995 35867 252998
rect 45553 252786 45619 252789
rect 41492 252784 45619 252786
rect 41492 252728 45558 252784
rect 45614 252728 45619 252784
rect 41492 252726 45619 252728
rect 45553 252723 45619 252726
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 47209 251970 47275 251973
rect 41492 251968 47275 251970
rect 41492 251912 47214 251968
rect 47270 251912 47275 251968
rect 41492 251910 47275 251912
rect 47209 251907 47275 251910
rect 44541 251562 44607 251565
rect 41492 251560 44607 251562
rect 41492 251504 44546 251560
rect 44602 251504 44607 251560
rect 41492 251502 44607 251504
rect 44541 251499 44607 251502
rect 554129 251290 554195 251293
rect 552460 251288 554195 251290
rect 552460 251232 554134 251288
rect 554190 251232 554195 251288
rect 552460 251230 554195 251232
rect 554129 251227 554195 251230
rect 46933 251154 46999 251157
rect 41492 251152 46999 251154
rect 41492 251096 46938 251152
rect 46994 251096 46999 251152
rect 41492 251094 46999 251096
rect 46933 251091 46999 251094
rect 673085 250746 673151 250749
rect 675477 250746 675543 250749
rect 673085 250744 675543 250746
rect 35758 250613 35818 250716
rect 673085 250688 673090 250744
rect 673146 250688 675482 250744
rect 675538 250688 675543 250744
rect 673085 250686 675543 250688
rect 673085 250683 673151 250686
rect 675477 250683 675543 250686
rect 35758 250608 35867 250613
rect 35758 250552 35806 250608
rect 35862 250552 35867 250608
rect 35758 250550 35867 250552
rect 35801 250547 35867 250550
rect 44725 250338 44791 250341
rect 41492 250336 44791 250338
rect 41492 250280 44730 250336
rect 44786 250280 44791 250336
rect 41492 250278 44791 250280
rect 44725 250275 44791 250278
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 669221 250202 669287 250205
rect 675293 250202 675359 250205
rect 669221 250200 675359 250202
rect 669221 250144 669226 250200
rect 669282 250144 675298 250200
rect 675354 250144 675359 250200
rect 669221 250142 675359 250144
rect 669221 250139 669287 250142
rect 675293 250139 675359 250142
rect 675477 250068 675543 250069
rect 675477 250066 675524 250068
rect 675432 250064 675524 250066
rect 675432 250008 675482 250064
rect 675432 250006 675524 250008
rect 675477 250004 675524 250006
rect 675588 250004 675594 250068
rect 675477 250003 675543 250004
rect 40542 249796 40602 249900
rect 40534 249732 40540 249796
rect 40604 249732 40610 249796
rect 673085 249658 673151 249661
rect 675334 249658 675340 249660
rect 673085 249656 675340 249658
rect 673085 249600 673090 249656
rect 673146 249600 675340 249656
rect 673085 249598 675340 249600
rect 673085 249595 673151 249598
rect 675334 249596 675340 249598
rect 675404 249596 675410 249660
rect 40726 249388 40786 249492
rect 40718 249324 40724 249388
rect 40788 249324 40794 249388
rect 45093 249114 45159 249117
rect 554037 249114 554103 249117
rect 41492 249112 45159 249114
rect 41492 249056 45098 249112
rect 45154 249056 45159 249112
rect 41492 249054 45159 249056
rect 552460 249112 554103 249114
rect 552460 249056 554042 249112
rect 554098 249056 554103 249112
rect 552460 249054 554103 249056
rect 45093 249051 45159 249054
rect 554037 249051 554103 249054
rect 45829 248706 45895 248709
rect 41492 248704 45895 248706
rect 41492 248648 45834 248704
rect 45890 248648 45895 248704
rect 41492 248646 45895 248648
rect 45829 248643 45895 248646
rect 46013 248298 46079 248301
rect 41492 248296 46079 248298
rect 41492 248240 46018 248296
rect 46074 248240 46079 248296
rect 41492 248238 46079 248240
rect 46013 248235 46079 248238
rect 35758 247757 35818 247860
rect 35758 247752 35867 247757
rect 35758 247696 35806 247752
rect 35862 247696 35867 247752
rect 35758 247694 35867 247696
rect 35801 247691 35867 247694
rect 664437 247754 664503 247757
rect 669221 247754 669287 247757
rect 664437 247752 669287 247754
rect 664437 247696 664442 247752
rect 664498 247696 669226 247752
rect 669282 247696 669287 247752
rect 664437 247694 669287 247696
rect 664437 247691 664503 247694
rect 669221 247691 669287 247694
rect 47761 247482 47827 247485
rect 41492 247480 47827 247482
rect 41492 247424 47766 247480
rect 47822 247424 47827 247480
rect 41492 247422 47827 247424
rect 47761 247419 47827 247422
rect 47393 247074 47459 247077
rect 41492 247072 47459 247074
rect 41492 247016 47398 247072
rect 47454 247016 47459 247072
rect 41492 247014 47459 247016
rect 47393 247011 47459 247014
rect 553853 246938 553919 246941
rect 552460 246936 553919 246938
rect 552460 246880 553858 246936
rect 553914 246880 553919 246936
rect 552460 246878 553919 246880
rect 553853 246875 553919 246878
rect 675753 246666 675819 246669
rect 676806 246666 676812 246668
rect 675753 246664 676812 246666
rect 675753 246608 675758 246664
rect 675814 246608 676812 246664
rect 675753 246606 676812 246608
rect 675753 246603 675819 246606
rect 676806 246604 676812 246606
rect 676876 246604 676882 246668
rect 41689 246530 41755 246533
rect 43437 246530 43503 246533
rect 41689 246528 43503 246530
rect 41689 246472 41694 246528
rect 41750 246472 43442 246528
rect 43498 246472 43503 246528
rect 41689 246470 43503 246472
rect 41689 246467 41755 246470
rect 43437 246467 43503 246470
rect 672165 246258 672231 246261
rect 673310 246258 673316 246260
rect 672165 246256 673316 246258
rect 672165 246200 672170 246256
rect 672226 246200 673316 246256
rect 672165 246198 673316 246200
rect 672165 246195 672231 246198
rect 673310 246196 673316 246198
rect 673380 246196 673386 246260
rect 673729 246258 673795 246261
rect 674598 246258 674604 246260
rect 673729 246256 674604 246258
rect 673729 246200 673734 246256
rect 673790 246200 674604 246256
rect 673729 246198 674604 246200
rect 673729 246195 673795 246198
rect 674598 246196 674604 246198
rect 674668 246196 674674 246260
rect 673821 245850 673887 245853
rect 675201 245850 675267 245853
rect 673821 245848 675267 245850
rect 673821 245792 673826 245848
rect 673882 245792 675206 245848
rect 675262 245792 675267 245848
rect 673821 245790 675267 245792
rect 673821 245787 673887 245790
rect 675201 245787 675267 245790
rect 39757 245714 39823 245717
rect 43253 245714 43319 245717
rect 39757 245712 43319 245714
rect 39757 245656 39762 245712
rect 39818 245656 43258 245712
rect 43314 245656 43319 245712
rect 39757 245654 43319 245656
rect 39757 245651 39823 245654
rect 43253 245651 43319 245654
rect 666553 245714 666619 245717
rect 667790 245714 667796 245716
rect 666553 245712 667796 245714
rect 666553 245656 666558 245712
rect 666614 245656 667796 245712
rect 666553 245654 667796 245656
rect 666553 245651 666619 245654
rect 667790 245652 667796 245654
rect 667860 245652 667866 245716
rect 671153 245578 671219 245581
rect 675201 245578 675267 245581
rect 671153 245576 675267 245578
rect 671153 245520 671158 245576
rect 671214 245520 675206 245576
rect 675262 245520 675267 245576
rect 671153 245518 675267 245520
rect 671153 245515 671219 245518
rect 675201 245515 675267 245518
rect 673085 245306 673151 245309
rect 675518 245306 675524 245308
rect 673085 245304 675524 245306
rect 673085 245248 673090 245304
rect 673146 245248 675524 245304
rect 673085 245246 675524 245248
rect 673085 245243 673151 245246
rect 675518 245244 675524 245246
rect 675588 245244 675594 245308
rect 553485 244762 553551 244765
rect 552460 244760 553551 244762
rect 552460 244704 553490 244760
rect 553546 244704 553551 244760
rect 552460 244702 553551 244704
rect 553485 244699 553551 244702
rect 674649 243538 674715 243541
rect 675385 243538 675451 243541
rect 674649 243536 675451 243538
rect 674649 243480 674654 243536
rect 674710 243480 675390 243536
rect 675446 243480 675451 243536
rect 674649 243478 675451 243480
rect 674649 243475 674715 243478
rect 675385 243475 675451 243478
rect 672901 242722 672967 242725
rect 675477 242722 675543 242725
rect 672901 242720 675543 242722
rect 672901 242664 672906 242720
rect 672962 242664 675482 242720
rect 675538 242664 675543 242720
rect 672901 242662 675543 242664
rect 672901 242659 672967 242662
rect 675477 242659 675543 242662
rect 553669 242586 553735 242589
rect 552460 242584 553735 242586
rect 552460 242528 553674 242584
rect 553730 242528 553735 242584
rect 552460 242526 553735 242528
rect 553669 242523 553735 242526
rect 674189 242178 674255 242181
rect 675385 242178 675451 242181
rect 674189 242176 675451 242178
rect 674189 242120 674194 242176
rect 674250 242120 675390 242176
rect 675446 242120 675451 242176
rect 674189 242118 675451 242120
rect 674189 242115 674255 242118
rect 675385 242115 675451 242118
rect 673545 241906 673611 241909
rect 676806 241906 676812 241908
rect 673545 241904 676812 241906
rect 673545 241848 673550 241904
rect 673606 241848 676812 241904
rect 673545 241846 676812 241848
rect 673545 241843 673611 241846
rect 676806 241844 676812 241846
rect 676876 241844 676882 241908
rect 673269 241634 673335 241637
rect 675017 241634 675083 241637
rect 673269 241632 675083 241634
rect 673269 241576 673274 241632
rect 673330 241576 675022 241632
rect 675078 241576 675083 241632
rect 673269 241574 675083 241576
rect 673269 241571 673335 241574
rect 675017 241571 675083 241574
rect 674465 241090 674531 241093
rect 675385 241090 675451 241093
rect 674465 241088 675451 241090
rect 674465 241032 674470 241088
rect 674526 241032 675390 241088
rect 675446 241032 675451 241088
rect 674465 241030 675451 241032
rect 674465 241027 674531 241030
rect 675385 241027 675451 241030
rect 554497 240410 554563 240413
rect 552460 240408 554563 240410
rect 552460 240352 554502 240408
rect 554558 240352 554563 240408
rect 552460 240350 554563 240352
rect 554497 240347 554563 240350
rect 672165 240274 672231 240277
rect 675385 240274 675451 240277
rect 672165 240272 675451 240274
rect 672165 240216 672170 240272
rect 672226 240216 675390 240272
rect 675446 240216 675451 240272
rect 672165 240214 675451 240216
rect 672165 240211 672231 240214
rect 675385 240211 675451 240214
rect 42057 240138 42123 240141
rect 44541 240138 44607 240141
rect 42057 240136 44607 240138
rect 42057 240080 42062 240136
rect 42118 240080 44546 240136
rect 44602 240080 44607 240136
rect 42057 240078 44607 240080
rect 42057 240075 42123 240078
rect 44541 240075 44607 240078
rect 671705 238642 671771 238645
rect 675385 238642 675451 238645
rect 671705 238640 675451 238642
rect 671705 238584 671710 238640
rect 671766 238584 675390 238640
rect 675446 238584 675451 238640
rect 671705 238582 675451 238584
rect 671705 238579 671771 238582
rect 675385 238579 675451 238582
rect 41965 238506 42031 238509
rect 47393 238506 47459 238509
rect 41965 238504 47459 238506
rect 41965 238448 41970 238504
rect 42026 238448 47398 238504
rect 47454 238448 47459 238504
rect 41965 238446 47459 238448
rect 41965 238443 42031 238446
rect 47393 238443 47459 238446
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 42006 238036 42012 238100
rect 42076 238098 42082 238100
rect 42333 238098 42399 238101
rect 42076 238096 42399 238098
rect 42076 238040 42338 238096
rect 42394 238040 42399 238096
rect 42076 238038 42399 238040
rect 42076 238036 42082 238038
rect 42333 238035 42399 238038
rect 674833 237282 674899 237285
rect 675477 237282 675543 237285
rect 674833 237280 675543 237282
rect 674833 237224 674838 237280
rect 674894 237224 675482 237280
rect 675538 237224 675543 237280
rect 674833 237222 675543 237224
rect 674833 237219 674899 237222
rect 675477 237219 675543 237222
rect 672947 236738 673013 236741
rect 674189 236738 674255 236741
rect 672947 236736 674255 236738
rect 672947 236680 672952 236736
rect 673008 236680 674194 236736
rect 674250 236680 674255 236736
rect 672947 236678 674255 236680
rect 672947 236675 673013 236678
rect 674189 236675 674255 236678
rect 40534 236540 40540 236604
rect 40604 236602 40610 236604
rect 41781 236602 41847 236605
rect 40604 236600 41847 236602
rect 40604 236544 41786 236600
rect 41842 236544 41847 236600
rect 40604 236542 41847 236544
rect 40604 236540 40610 236542
rect 41781 236539 41847 236542
rect 670325 236194 670391 236197
rect 675477 236194 675543 236197
rect 670325 236192 675543 236194
rect 670325 236136 670330 236192
rect 670386 236136 675482 236192
rect 675538 236136 675543 236192
rect 670325 236134 675543 236136
rect 670325 236131 670391 236134
rect 675477 236131 675543 236134
rect 553761 236058 553827 236061
rect 552460 236056 553827 236058
rect 552460 236000 553766 236056
rect 553822 236000 553827 236056
rect 552460 235998 553827 236000
rect 553761 235995 553827 235998
rect 675477 235516 675543 235517
rect 675477 235514 675524 235516
rect 675432 235512 675524 235514
rect 675432 235456 675482 235512
rect 675432 235454 675524 235456
rect 675477 235452 675524 235454
rect 675588 235452 675594 235516
rect 675477 235451 675543 235452
rect 40718 234636 40724 234700
rect 40788 234698 40794 234700
rect 41781 234698 41847 234701
rect 40788 234696 41847 234698
rect 40788 234640 41786 234696
rect 41842 234640 41847 234696
rect 40788 234638 41847 234640
rect 40788 234636 40794 234638
rect 41781 234635 41847 234638
rect 42333 233882 42399 233885
rect 554405 233882 554471 233885
rect 42333 233880 42442 233882
rect 42333 233824 42338 233880
rect 42394 233824 42442 233880
rect 42333 233819 42442 233824
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 670877 233882 670943 233885
rect 675845 233882 675911 233885
rect 670877 233880 675911 233882
rect 670877 233824 670882 233880
rect 670938 233824 675850 233880
rect 675906 233824 675911 233880
rect 670877 233822 675911 233824
rect 670877 233819 670943 233822
rect 675845 233819 675911 233822
rect 42382 233202 42442 233819
rect 46013 233202 46079 233205
rect 42382 233200 46079 233202
rect 42382 233144 46018 233200
rect 46074 233144 46079 233200
rect 42382 233142 46079 233144
rect 46013 233139 46079 233142
rect 674373 232658 674439 232661
rect 675845 232658 675911 232661
rect 674373 232656 675911 232658
rect 674373 232600 674378 232656
rect 674434 232600 675850 232656
rect 675906 232600 675911 232656
rect 674373 232598 675911 232600
rect 674373 232595 674439 232598
rect 675845 232595 675911 232598
rect 668761 232522 668827 232525
rect 673545 232522 673611 232525
rect 668761 232520 673611 232522
rect 668761 232464 668766 232520
rect 668822 232464 673550 232520
rect 673606 232464 673611 232520
rect 668761 232462 673611 232464
rect 668761 232459 668827 232462
rect 673545 232459 673611 232462
rect 674557 232386 674623 232389
rect 676029 232386 676095 232389
rect 674557 232384 676095 232386
rect 674557 232328 674562 232384
rect 674618 232328 676034 232384
rect 676090 232328 676095 232384
rect 674557 232326 676095 232328
rect 674557 232323 674623 232326
rect 676029 232323 676095 232326
rect 42425 232250 42491 232253
rect 47209 232250 47275 232253
rect 42425 232248 47275 232250
rect 42425 232192 42430 232248
rect 42486 232192 47214 232248
rect 47270 232192 47275 232248
rect 42425 232190 47275 232192
rect 42425 232187 42491 232190
rect 47209 232187 47275 232190
rect 670734 231916 670740 231980
rect 670804 231978 670810 231980
rect 671889 231978 671955 231981
rect 670804 231976 671955 231978
rect 670804 231920 671894 231976
rect 671950 231920 671955 231976
rect 670804 231918 671955 231920
rect 670804 231916 670810 231918
rect 671889 231915 671955 231918
rect 42425 231842 42491 231845
rect 45829 231842 45895 231845
rect 42425 231840 45895 231842
rect 42425 231784 42430 231840
rect 42486 231784 45834 231840
rect 45890 231784 45895 231840
rect 42425 231782 45895 231784
rect 42425 231779 42491 231782
rect 45829 231779 45895 231782
rect 42425 231570 42491 231573
rect 45001 231570 45067 231573
rect 42425 231568 45067 231570
rect 42425 231512 42430 231568
rect 42486 231512 45006 231568
rect 45062 231512 45067 231568
rect 42425 231510 45067 231512
rect 42425 231507 42491 231510
rect 45001 231507 45067 231510
rect 43989 231162 44055 231165
rect 669129 231162 669195 231165
rect 43989 231160 669195 231162
rect 43989 231104 43994 231160
rect 44050 231104 669134 231160
rect 669190 231104 669195 231160
rect 43989 231102 669195 231104
rect 43989 231099 44055 231102
rect 669129 231099 669195 231102
rect 42149 230482 42215 230485
rect 44633 230482 44699 230485
rect 42149 230480 44699 230482
rect 42149 230424 42154 230480
rect 42210 230424 44638 230480
rect 44694 230424 44699 230480
rect 42149 230422 44699 230424
rect 42149 230419 42215 230422
rect 44633 230419 44699 230422
rect 144637 230482 144703 230485
rect 151077 230482 151143 230485
rect 144637 230480 151143 230482
rect 144637 230424 144642 230480
rect 144698 230424 151082 230480
rect 151138 230424 151143 230480
rect 144637 230422 151143 230424
rect 144637 230419 144703 230422
rect 151077 230419 151143 230422
rect 664897 230346 664963 230349
rect 674669 230346 674735 230349
rect 664897 230344 674735 230346
rect 664897 230288 664902 230344
rect 664958 230288 674674 230344
rect 674730 230288 674735 230344
rect 664897 230286 674735 230288
rect 664897 230283 664963 230286
rect 674669 230283 674735 230286
rect 157609 230210 157675 230213
rect 162301 230210 162367 230213
rect 676489 230210 676555 230213
rect 157609 230208 162367 230210
rect 157609 230152 157614 230208
rect 157670 230152 162306 230208
rect 162362 230152 162367 230208
rect 157609 230150 162367 230152
rect 157609 230147 157675 230150
rect 162301 230147 162367 230150
rect 674974 230208 676555 230210
rect 674974 230152 676494 230208
rect 676550 230152 676555 230208
rect 674974 230150 676555 230152
rect 156781 230074 156847 230077
rect 157425 230074 157491 230077
rect 156781 230072 157491 230074
rect 156781 230016 156786 230072
rect 156842 230016 157430 230072
rect 157486 230016 157491 230072
rect 156781 230014 157491 230016
rect 156781 230011 156847 230014
rect 157425 230011 157491 230014
rect 674327 230074 674393 230077
rect 674974 230074 675034 230150
rect 676489 230147 676555 230150
rect 674327 230072 675034 230074
rect 674327 230016 674332 230072
rect 674388 230016 675034 230072
rect 674327 230014 675034 230016
rect 674327 230011 674393 230014
rect 185393 229938 185459 229941
rect 186037 229938 186103 229941
rect 185393 229936 186103 229938
rect 185393 229880 185398 229936
rect 185454 229880 186042 229936
rect 186098 229880 186103 229936
rect 185393 229878 186103 229880
rect 185393 229875 185459 229878
rect 186037 229875 186103 229878
rect 144453 229802 144519 229805
rect 148133 229802 148199 229805
rect 144453 229800 148199 229802
rect 144453 229744 144458 229800
rect 144514 229744 148138 229800
rect 148194 229744 148199 229800
rect 144453 229742 148199 229744
rect 144453 229739 144519 229742
rect 148133 229739 148199 229742
rect 156781 229802 156847 229805
rect 156781 229800 157442 229802
rect 156781 229744 156786 229800
rect 156842 229744 157442 229800
rect 156781 229742 157442 229744
rect 156781 229739 156847 229742
rect 157382 229666 157442 229742
rect 157977 229666 158043 229669
rect 157382 229664 158043 229666
rect 157382 229608 157982 229664
rect 158038 229608 158043 229664
rect 157382 229606 158043 229608
rect 157977 229603 158043 229606
rect 150341 229530 150407 229533
rect 150341 229528 154590 229530
rect 150341 229472 150346 229528
rect 150402 229472 154590 229528
rect 150341 229470 154590 229472
rect 150341 229467 150407 229470
rect 145833 229394 145899 229397
rect 147949 229394 148015 229397
rect 145833 229392 148015 229394
rect 145833 229336 145838 229392
rect 145894 229336 147954 229392
rect 148010 229336 148015 229392
rect 145833 229334 148015 229336
rect 154530 229394 154590 229470
rect 162485 229394 162551 229397
rect 154530 229392 162551 229394
rect 154530 229336 162490 229392
rect 162546 229336 162551 229392
rect 154530 229334 162551 229336
rect 145833 229331 145899 229334
rect 147949 229331 148015 229334
rect 162485 229331 162551 229334
rect 148133 229258 148199 229261
rect 150985 229258 151051 229261
rect 674465 229258 674531 229261
rect 148133 229256 151051 229258
rect 148133 229200 148138 229256
rect 148194 229200 150990 229256
rect 151046 229200 151051 229256
rect 148133 229198 151051 229200
rect 148133 229195 148199 229198
rect 150985 229195 151051 229198
rect 663750 229256 674531 229258
rect 663750 229200 674470 229256
rect 674526 229200 674531 229256
rect 663750 229198 674531 229200
rect 663750 229125 663810 229198
rect 674465 229195 674531 229198
rect 140037 229122 140103 229125
rect 143533 229122 143599 229125
rect 140037 229120 143599 229122
rect 140037 229064 140042 229120
rect 140098 229064 143538 229120
rect 143594 229064 143599 229120
rect 140037 229062 143599 229064
rect 140037 229059 140103 229062
rect 143533 229059 143599 229062
rect 663701 229120 663810 229125
rect 663701 229064 663706 229120
rect 663762 229064 663810 229120
rect 663701 229062 663810 229064
rect 663701 229059 663767 229062
rect 193029 228986 193095 228989
rect 195421 228986 195487 228989
rect 193029 228984 195487 228986
rect 193029 228928 193034 228984
rect 193090 228928 195426 228984
rect 195482 228928 195487 228984
rect 193029 228926 195487 228928
rect 193029 228923 193095 228926
rect 195421 228923 195487 228926
rect 159357 228850 159423 228853
rect 162485 228850 162551 228853
rect 159357 228848 162551 228850
rect 159357 228792 159362 228848
rect 159418 228792 162490 228848
rect 162546 228792 162551 228848
rect 159357 228790 162551 228792
rect 159357 228787 159423 228790
rect 162485 228787 162551 228790
rect 173157 228850 173223 228853
rect 176101 228850 176167 228853
rect 173157 228848 176167 228850
rect 173157 228792 173162 228848
rect 173218 228792 176106 228848
rect 176162 228792 176167 228848
rect 173157 228790 176167 228792
rect 173157 228787 173223 228790
rect 176101 228787 176167 228790
rect 662137 228578 662203 228581
rect 673453 228578 673519 228581
rect 675477 228580 675543 228581
rect 675477 228578 675524 228580
rect 662137 228576 673519 228578
rect 662137 228520 662142 228576
rect 662198 228520 673458 228576
rect 673514 228520 673519 228576
rect 662137 228518 673519 228520
rect 675432 228576 675524 228578
rect 675432 228520 675482 228576
rect 675432 228518 675524 228520
rect 662137 228515 662203 228518
rect 673453 228515 673519 228518
rect 675477 228516 675524 228518
rect 675588 228516 675594 228580
rect 675477 228515 675543 228516
rect 160001 228442 160067 228445
rect 166809 228442 166875 228445
rect 160001 228440 166875 228442
rect 160001 228384 160006 228440
rect 160062 228384 166814 228440
rect 166870 228384 166875 228440
rect 160001 228382 166875 228384
rect 160001 228379 160067 228382
rect 166809 228379 166875 228382
rect 146109 228034 146175 228037
rect 147121 228034 147187 228037
rect 146109 228032 147187 228034
rect 146109 227976 146114 228032
rect 146170 227976 147126 228032
rect 147182 227976 147187 228032
rect 146109 227974 147187 227976
rect 146109 227971 146175 227974
rect 147121 227971 147187 227974
rect 136633 227898 136699 227901
rect 141509 227898 141575 227901
rect 136633 227896 141575 227898
rect 136633 227840 136638 227896
rect 136694 227840 141514 227896
rect 141570 227840 141575 227896
rect 136633 227838 141575 227840
rect 136633 227835 136699 227838
rect 141509 227835 141575 227838
rect 175181 227626 175247 227629
rect 177205 227626 177271 227629
rect 175181 227624 177271 227626
rect 175181 227568 175186 227624
rect 175242 227568 177210 227624
rect 177266 227568 177271 227624
rect 175181 227566 177271 227568
rect 175181 227563 175247 227566
rect 177205 227563 177271 227566
rect 157333 227490 157399 227493
rect 166533 227490 166599 227493
rect 157333 227488 166599 227490
rect 157333 227432 157338 227488
rect 157394 227432 166538 227488
rect 166594 227432 166599 227488
rect 157333 227430 166599 227432
rect 157333 227427 157399 227430
rect 166533 227427 166599 227430
rect 170765 227490 170831 227493
rect 171685 227490 171751 227493
rect 170765 227488 171751 227490
rect 170765 227432 170770 227488
rect 170826 227432 171690 227488
rect 171746 227432 171751 227488
rect 170765 227430 171751 227432
rect 170765 227427 170831 227430
rect 171685 227427 171751 227430
rect 41965 227356 42031 227357
rect 41965 227352 42012 227356
rect 42076 227354 42082 227356
rect 175917 227354 175983 227357
rect 176745 227354 176811 227357
rect 41965 227296 41970 227352
rect 41965 227292 42012 227296
rect 42076 227294 42122 227354
rect 175917 227352 176811 227354
rect 175917 227296 175922 227352
rect 175978 227296 176750 227352
rect 176806 227296 176811 227352
rect 175917 227294 176811 227296
rect 42076 227292 42082 227294
rect 41965 227291 42031 227292
rect 175917 227291 175983 227294
rect 176745 227291 176811 227294
rect 169569 227218 169635 227221
rect 171087 227218 171153 227221
rect 169569 227216 171153 227218
rect 169569 227160 169574 227216
rect 169630 227160 171092 227216
rect 171148 227160 171153 227216
rect 169569 227158 171153 227160
rect 169569 227155 169635 227158
rect 171087 227155 171153 227158
rect 155585 227082 155651 227085
rect 157517 227082 157583 227085
rect 155585 227080 157583 227082
rect 155585 227024 155590 227080
rect 155646 227024 157522 227080
rect 157578 227024 157583 227080
rect 155585 227022 157583 227024
rect 155585 227019 155651 227022
rect 157517 227019 157583 227022
rect 672349 227082 672415 227085
rect 672574 227082 672580 227084
rect 672349 227080 672580 227082
rect 672349 227024 672354 227080
rect 672410 227024 672580 227080
rect 672349 227022 672580 227024
rect 672349 227019 672415 227022
rect 672574 227020 672580 227022
rect 672644 227020 672650 227084
rect 673269 227082 673335 227085
rect 676765 227082 676831 227085
rect 673269 227080 676831 227082
rect 673269 227024 673274 227080
rect 673330 227024 676770 227080
rect 676826 227024 676831 227080
rect 673269 227022 676831 227024
rect 673269 227019 673335 227022
rect 676765 227019 676831 227022
rect 652385 226946 652451 226949
rect 652385 226944 663810 226946
rect 652385 226888 652390 226944
rect 652446 226888 663810 226944
rect 652385 226886 663810 226888
rect 652385 226883 652451 226886
rect 221825 226810 221891 226813
rect 223113 226810 223179 226813
rect 221825 226808 223179 226810
rect 221825 226752 221830 226808
rect 221886 226752 223118 226808
rect 223174 226752 223179 226808
rect 221825 226750 223179 226752
rect 663750 226810 663810 226886
rect 673545 226810 673611 226813
rect 676949 226810 677015 226813
rect 663750 226750 673010 226810
rect 221825 226747 221891 226750
rect 223113 226747 223179 226750
rect 141601 226538 141667 226541
rect 142245 226538 142311 226541
rect 141601 226536 142311 226538
rect 141601 226480 141606 226536
rect 141662 226480 142250 226536
rect 142306 226480 142311 226536
rect 141601 226478 142311 226480
rect 672950 226538 673010 226750
rect 673545 226808 677015 226810
rect 673545 226752 673550 226808
rect 673606 226752 676954 226808
rect 677010 226752 677015 226808
rect 673545 226750 677015 226752
rect 673545 226747 673611 226750
rect 676949 226747 677015 226750
rect 674046 226538 674052 226540
rect 672950 226478 674052 226538
rect 141601 226475 141667 226478
rect 142245 226475 142311 226478
rect 674046 226476 674052 226478
rect 674116 226476 674122 226540
rect 658917 226402 658983 226405
rect 672717 226402 672783 226405
rect 658917 226400 672783 226402
rect 658917 226344 658922 226400
rect 658978 226344 672722 226400
rect 672778 226344 672783 226400
rect 658917 226342 672783 226344
rect 658917 226339 658983 226342
rect 672717 226339 672783 226342
rect 151445 226266 151511 226269
rect 157149 226266 157215 226269
rect 151445 226264 157215 226266
rect 151445 226208 151450 226264
rect 151506 226208 157154 226264
rect 157210 226208 157215 226264
rect 151445 226206 157215 226208
rect 151445 226203 151511 226206
rect 157149 226203 157215 226206
rect 672597 226130 672663 226133
rect 674833 226130 674899 226133
rect 672597 226128 674899 226130
rect 672597 226072 672602 226128
rect 672658 226072 674838 226128
rect 674894 226072 674899 226128
rect 672597 226070 674899 226072
rect 672597 226067 672663 226070
rect 674833 226067 674899 226070
rect 142613 225994 142679 225997
rect 149789 225994 149855 225997
rect 672487 225994 672553 225997
rect 142613 225992 149855 225994
rect 142613 225936 142618 225992
rect 142674 225936 149794 225992
rect 149850 225936 149855 225992
rect 142613 225934 149855 225936
rect 142613 225931 142679 225934
rect 149789 225931 149855 225934
rect 663750 225992 672553 225994
rect 663750 225936 672492 225992
rect 672548 225936 672553 225992
rect 663750 225934 672553 225936
rect 156597 225858 156663 225861
rect 158161 225858 158227 225861
rect 156597 225856 158227 225858
rect 156597 225800 156602 225856
rect 156658 225800 158166 225856
rect 158222 225800 158227 225856
rect 156597 225798 158227 225800
rect 156597 225795 156663 225798
rect 158161 225795 158227 225798
rect 42425 225722 42491 225725
rect 45553 225722 45619 225725
rect 42425 225720 45619 225722
rect 42425 225664 42430 225720
rect 42486 225664 45558 225720
rect 45614 225664 45619 225720
rect 42425 225662 45619 225664
rect 42425 225659 42491 225662
rect 45553 225659 45619 225662
rect 656157 225586 656223 225589
rect 663750 225586 663810 225934
rect 672487 225931 672553 225934
rect 672373 225722 672439 225725
rect 675477 225722 675543 225725
rect 672373 225720 675543 225722
rect 672373 225664 672378 225720
rect 672434 225664 675482 225720
rect 675538 225664 675543 225720
rect 672373 225662 675543 225664
rect 672373 225659 672439 225662
rect 675477 225659 675543 225662
rect 656157 225584 663810 225586
rect 656157 225528 656162 225584
rect 656218 225528 663810 225584
rect 656157 225526 663810 225528
rect 656157 225523 656223 225526
rect 148869 225450 148935 225453
rect 157149 225450 157215 225453
rect 148869 225448 157215 225450
rect 148869 225392 148874 225448
rect 148930 225392 157154 225448
rect 157210 225392 157215 225448
rect 148869 225390 157215 225392
rect 148869 225387 148935 225390
rect 157149 225387 157215 225390
rect 652753 225314 652819 225317
rect 672027 225314 672093 225317
rect 652753 225312 672093 225314
rect 652753 225256 652758 225312
rect 652814 225256 672032 225312
rect 672088 225256 672093 225312
rect 652753 225254 672093 225256
rect 652753 225251 652819 225254
rect 672027 225251 672093 225254
rect 672149 225178 672215 225181
rect 675845 225178 675911 225181
rect 672149 225176 675911 225178
rect 672149 225120 672154 225176
rect 672210 225120 675850 225176
rect 675906 225120 675911 225176
rect 672149 225118 675911 225120
rect 672149 225115 672215 225118
rect 675845 225115 675911 225118
rect 650637 225042 650703 225045
rect 671889 225042 671955 225045
rect 650637 225040 671955 225042
rect 650637 224984 650642 225040
rect 650698 224984 671894 225040
rect 671950 224984 671955 225040
rect 650637 224982 671955 224984
rect 650637 224979 650703 224982
rect 671889 224979 671955 224982
rect 42609 224906 42675 224909
rect 46933 224906 46999 224909
rect 42609 224904 46999 224906
rect 42609 224848 42614 224904
rect 42670 224848 46938 224904
rect 46994 224848 46999 224904
rect 42609 224846 46999 224848
rect 42609 224843 42675 224846
rect 46933 224843 46999 224846
rect 548057 224770 548123 224773
rect 549989 224770 550055 224773
rect 550449 224770 550515 224773
rect 548057 224768 550515 224770
rect 548057 224712 548062 224768
rect 548118 224712 549994 224768
rect 550050 224712 550454 224768
rect 550510 224712 550515 224768
rect 548057 224710 550515 224712
rect 548057 224707 548123 224710
rect 549989 224707 550055 224710
rect 550449 224707 550515 224710
rect 562133 224770 562199 224773
rect 563697 224770 563763 224773
rect 562133 224768 563763 224770
rect 562133 224712 562138 224768
rect 562194 224712 563702 224768
rect 563758 224712 563763 224768
rect 562133 224710 563763 224712
rect 562133 224707 562199 224710
rect 563697 224707 563763 224710
rect 671813 224770 671879 224773
rect 673453 224770 673519 224773
rect 671813 224768 673519 224770
rect 671813 224712 671818 224768
rect 671874 224712 673458 224768
rect 673514 224712 673519 224768
rect 671813 224710 673519 224712
rect 671813 224707 671879 224710
rect 673453 224707 673519 224710
rect 557993 224634 558059 224637
rect 557766 224632 558059 224634
rect 557766 224576 557998 224632
rect 558054 224576 558059 224632
rect 557766 224574 558059 224576
rect 41689 224498 41755 224501
rect 63125 224498 63191 224501
rect 41689 224496 63191 224498
rect 41689 224440 41694 224496
rect 41750 224440 63130 224496
rect 63186 224440 63191 224496
rect 41689 224438 63191 224440
rect 41689 224435 41755 224438
rect 63125 224435 63191 224438
rect 151629 224498 151695 224501
rect 152365 224498 152431 224501
rect 151629 224496 152431 224498
rect 151629 224440 151634 224496
rect 151690 224440 152370 224496
rect 152426 224440 152431 224496
rect 151629 224438 152431 224440
rect 151629 224435 151695 224438
rect 152365 224435 152431 224438
rect 542445 224498 542511 224501
rect 543181 224498 543247 224501
rect 542445 224496 543247 224498
rect 542445 224440 542450 224496
rect 542506 224440 543186 224496
rect 543242 224440 543247 224496
rect 542445 224438 543247 224440
rect 542445 224435 542511 224438
rect 543181 224435 543247 224438
rect 554865 224498 554931 224501
rect 556061 224498 556127 224501
rect 557766 224498 557826 224574
rect 557993 224571 558059 224574
rect 554865 224496 557826 224498
rect 554865 224440 554870 224496
rect 554926 224440 556066 224496
rect 556122 224440 557826 224496
rect 554865 224438 557826 224440
rect 554865 224435 554931 224438
rect 556061 224435 556127 224438
rect 62665 224226 62731 224229
rect 591481 224226 591547 224229
rect 667749 224226 667815 224229
rect 62665 224224 591547 224226
rect 62665 224168 62670 224224
rect 62726 224168 591486 224224
rect 591542 224168 591547 224224
rect 62665 224166 591547 224168
rect 62665 224163 62731 224166
rect 591481 224163 591547 224166
rect 663750 224224 667815 224226
rect 663750 224168 667754 224224
rect 667810 224168 667815 224224
rect 663750 224166 667815 224168
rect 136725 223954 136791 223957
rect 142245 223954 142311 223957
rect 136725 223952 142311 223954
rect 136725 223896 136730 223952
rect 136786 223896 142250 223952
rect 142306 223896 142311 223952
rect 136725 223894 142311 223896
rect 136725 223891 136791 223894
rect 142245 223891 142311 223894
rect 142429 223954 142495 223957
rect 151629 223954 151695 223957
rect 142429 223952 151695 223954
rect 142429 223896 142434 223952
rect 142490 223896 151634 223952
rect 151690 223896 151695 223952
rect 142429 223894 151695 223896
rect 142429 223891 142495 223894
rect 151629 223891 151695 223894
rect 654777 223954 654843 223957
rect 663750 223954 663810 224166
rect 667749 224163 667815 224166
rect 671475 224090 671541 224093
rect 672073 224090 672139 224093
rect 671475 224088 672139 224090
rect 671475 224032 671480 224088
rect 671536 224032 672078 224088
rect 672134 224032 672139 224088
rect 671475 224030 672139 224032
rect 671475 224027 671541 224030
rect 672073 224027 672139 224030
rect 654777 223952 663810 223954
rect 654777 223896 654782 223952
rect 654838 223896 663810 223952
rect 654777 223894 663810 223896
rect 654777 223891 654843 223894
rect 678237 223818 678303 223821
rect 678237 223816 678346 223818
rect 678237 223760 678242 223816
rect 678298 223760 678346 223816
rect 678237 223755 678346 223760
rect 657537 223682 657603 223685
rect 667749 223682 667815 223685
rect 657537 223680 667815 223682
rect 657537 223624 657542 223680
rect 657598 223624 667754 223680
rect 667810 223624 667815 223680
rect 657537 223622 667815 223624
rect 657537 223619 657603 223622
rect 667749 223619 667815 223622
rect 42149 223546 42215 223549
rect 58617 223546 58683 223549
rect 42149 223544 58683 223546
rect 42149 223488 42154 223544
rect 42210 223488 58622 223544
rect 58678 223488 58683 223544
rect 42149 223486 58683 223488
rect 42149 223483 42215 223486
rect 58617 223483 58683 223486
rect 62941 223546 63007 223549
rect 62941 223544 582390 223546
rect 62941 223488 62946 223544
rect 63002 223488 582390 223544
rect 678286 223516 678346 223755
rect 62941 223486 582390 223488
rect 62941 223483 63007 223486
rect 582330 223410 582390 223486
rect 591982 223410 591988 223412
rect 582330 223350 591988 223410
rect 591982 223348 591988 223350
rect 592052 223348 592058 223412
rect 669267 223410 669333 223413
rect 669446 223410 669452 223412
rect 669267 223408 669452 223410
rect 669267 223352 669272 223408
rect 669328 223352 669452 223408
rect 669267 223350 669452 223352
rect 669267 223347 669333 223350
rect 669446 223348 669452 223350
rect 669516 223348 669522 223412
rect 142153 223274 142219 223277
rect 149513 223274 149579 223277
rect 142153 223272 149579 223274
rect 142153 223216 142158 223272
rect 142214 223216 149518 223272
rect 149574 223216 149579 223272
rect 142153 223214 149579 223216
rect 142153 223211 142219 223214
rect 149513 223211 149579 223214
rect 665817 223138 665883 223141
rect 667749 223138 667815 223141
rect 665817 223136 667815 223138
rect 665817 223080 665822 223136
rect 665878 223080 667754 223136
rect 667810 223080 667815 223136
rect 665817 223078 667815 223080
rect 665817 223075 665883 223078
rect 667749 223075 667815 223078
rect 683389 223138 683455 223141
rect 683389 223136 683468 223138
rect 683389 223080 683394 223136
rect 683450 223080 683468 223136
rect 683389 223078 683468 223080
rect 683389 223075 683455 223078
rect 145925 223002 145991 223005
rect 147121 223002 147187 223005
rect 145925 223000 147187 223002
rect 145925 222944 145930 223000
rect 145986 222944 147126 223000
rect 147182 222944 147187 223000
rect 145925 222942 147187 222944
rect 145925 222939 145991 222942
rect 147121 222939 147187 222942
rect 649574 222940 649580 223004
rect 649644 223002 649650 223004
rect 651966 223002 651972 223004
rect 649644 222942 651972 223002
rect 649644 222940 649650 222942
rect 651966 222940 651972 222942
rect 652036 222940 652042 223004
rect 141969 222866 142035 222869
rect 142429 222866 142495 222869
rect 141969 222864 142495 222866
rect 141969 222808 141974 222864
rect 142030 222808 142434 222864
rect 142490 222808 142495 222864
rect 141969 222806 142495 222808
rect 141969 222803 142035 222806
rect 142429 222803 142495 222806
rect 653397 222866 653463 222869
rect 673269 222866 673335 222869
rect 653397 222864 673335 222866
rect 653397 222808 653402 222864
rect 653458 222808 673274 222864
rect 673330 222808 673335 222864
rect 653397 222806 673335 222808
rect 653397 222803 653463 222806
rect 673269 222803 673335 222806
rect 683205 222730 683271 222733
rect 683205 222728 683284 222730
rect 683205 222672 683210 222728
rect 683266 222672 683284 222728
rect 683205 222670 683284 222672
rect 683205 222667 683271 222670
rect 172237 222458 172303 222461
rect 175825 222458 175891 222461
rect 172237 222456 175891 222458
rect 172237 222400 172242 222456
rect 172298 222400 175830 222456
rect 175886 222400 175891 222456
rect 172237 222398 175891 222400
rect 172237 222395 172303 222398
rect 175825 222395 175891 222398
rect 674281 222458 674347 222461
rect 674281 222456 676230 222458
rect 674281 222400 674286 222456
rect 674342 222400 676230 222456
rect 674281 222398 676230 222400
rect 674281 222395 674347 222398
rect 118417 222322 118483 222325
rect 141969 222322 142035 222325
rect 118417 222320 142035 222322
rect 118417 222264 118422 222320
rect 118478 222264 141974 222320
rect 142030 222264 142035 222320
rect 118417 222262 142035 222264
rect 118417 222259 118483 222262
rect 141969 222259 142035 222262
rect 553301 222322 553367 222325
rect 557349 222322 557415 222325
rect 553301 222320 557415 222322
rect 553301 222264 553306 222320
rect 553362 222264 557354 222320
rect 557410 222264 557415 222320
rect 553301 222262 557415 222264
rect 676170 222322 676230 222398
rect 676170 222262 676292 222322
rect 553301 222259 553367 222262
rect 557349 222259 557415 222262
rect 157609 222050 157675 222053
rect 158345 222050 158411 222053
rect 157609 222048 158411 222050
rect 157609 221992 157614 222048
rect 157670 221992 158350 222048
rect 158406 221992 158411 222048
rect 157609 221990 158411 221992
rect 157609 221987 157675 221990
rect 158345 221987 158411 221990
rect 166809 222050 166875 222053
rect 166993 222050 167059 222053
rect 166809 222048 167059 222050
rect 166809 221992 166814 222048
rect 166870 221992 166998 222048
rect 167054 221992 167059 222048
rect 166809 221990 167059 221992
rect 166809 221987 166875 221990
rect 166993 221987 167059 221990
rect 559373 222050 559439 222053
rect 561489 222050 561555 222053
rect 559373 222048 561555 222050
rect 559373 221992 559378 222048
rect 559434 221992 561494 222048
rect 561550 221992 561555 222048
rect 559373 221990 561555 221992
rect 559373 221987 559439 221990
rect 561489 221987 561555 221990
rect 176561 221914 176627 221917
rect 177389 221914 177455 221917
rect 176561 221912 177455 221914
rect 176561 221856 176566 221912
rect 176622 221856 177394 221912
rect 177450 221856 177455 221912
rect 176561 221854 177455 221856
rect 176561 221851 176627 221854
rect 177389 221851 177455 221854
rect 556981 221914 557047 221917
rect 557533 221914 557599 221917
rect 556981 221912 557599 221914
rect 556981 221856 556986 221912
rect 557042 221856 557538 221912
rect 557594 221856 557599 221912
rect 556981 221854 557599 221856
rect 556981 221851 557047 221854
rect 557533 221851 557599 221854
rect 676029 221914 676095 221917
rect 676029 221912 676292 221914
rect 676029 221856 676034 221912
rect 676090 221856 676292 221912
rect 676029 221854 676292 221856
rect 676029 221851 676095 221854
rect 545757 221778 545823 221781
rect 549253 221778 549319 221781
rect 545757 221776 549319 221778
rect 545757 221720 545762 221776
rect 545818 221720 549258 221776
rect 549314 221720 549319 221776
rect 545757 221718 549319 221720
rect 545757 221715 545823 221718
rect 549253 221715 549319 221718
rect 563697 221778 563763 221781
rect 572621 221778 572687 221781
rect 563697 221776 572687 221778
rect 563697 221720 563702 221776
rect 563758 221720 572626 221776
rect 572682 221720 572687 221776
rect 563697 221718 572687 221720
rect 563697 221715 563763 221718
rect 572621 221715 572687 221718
rect 660757 221778 660823 221781
rect 674833 221778 674899 221781
rect 660757 221776 674899 221778
rect 660757 221720 660762 221776
rect 660818 221720 674838 221776
rect 674894 221720 674899 221776
rect 660757 221718 674899 221720
rect 660757 221715 660823 221718
rect 674833 221715 674899 221718
rect 157425 221642 157491 221645
rect 158161 221642 158227 221645
rect 157425 221640 158227 221642
rect 157425 221584 157430 221640
rect 157486 221584 158166 221640
rect 158222 221584 158227 221640
rect 157425 221582 158227 221584
rect 157425 221579 157491 221582
rect 158161 221579 158227 221582
rect 522573 221506 522639 221509
rect 618253 221506 618319 221509
rect 522573 221504 618319 221506
rect 522573 221448 522578 221504
rect 522634 221448 618258 221504
rect 618314 221448 618319 221504
rect 522573 221446 618319 221448
rect 522573 221443 522639 221446
rect 618253 221443 618319 221446
rect 651465 221506 651531 221509
rect 666829 221506 666895 221509
rect 651465 221504 666895 221506
rect 651465 221448 651470 221504
rect 651526 221448 666834 221504
rect 666890 221448 666895 221504
rect 651465 221446 666895 221448
rect 651465 221443 651531 221446
rect 666829 221443 666895 221446
rect 675017 221506 675083 221509
rect 675017 221504 676292 221506
rect 675017 221448 675022 221504
rect 675078 221448 676292 221504
rect 675017 221446 676292 221448
rect 675017 221443 675083 221446
rect 171409 221370 171475 221373
rect 171961 221370 172027 221373
rect 171409 221368 172027 221370
rect 171409 221312 171414 221368
rect 171470 221312 171966 221368
rect 172022 221312 172027 221368
rect 171409 221310 172027 221312
rect 171409 221307 171475 221310
rect 171961 221307 172027 221310
rect 161013 221234 161079 221237
rect 162301 221234 162367 221237
rect 161013 221232 162367 221234
rect 161013 221176 161018 221232
rect 161074 221176 162306 221232
rect 162362 221176 162367 221232
rect 161013 221174 162367 221176
rect 161013 221171 161079 221174
rect 162301 221171 162367 221174
rect 515765 221234 515831 221237
rect 600865 221234 600931 221237
rect 515765 221232 600931 221234
rect 515765 221176 515770 221232
rect 515826 221176 600870 221232
rect 600926 221176 600931 221232
rect 515765 221174 600931 221176
rect 515765 221171 515831 221174
rect 600865 221171 600931 221174
rect 673269 221098 673335 221101
rect 673269 221096 676292 221098
rect 673269 221040 673274 221096
rect 673330 221040 676292 221096
rect 673269 221038 676292 221040
rect 673269 221035 673335 221038
rect 142107 220962 142173 220965
rect 148501 220962 148567 220965
rect 142107 220960 148567 220962
rect 142107 220904 142112 220960
rect 142168 220904 148506 220960
rect 148562 220904 148567 220960
rect 142107 220902 148567 220904
rect 142107 220899 142173 220902
rect 148501 220899 148567 220902
rect 160645 220962 160711 220965
rect 164509 220962 164575 220965
rect 160645 220960 164575 220962
rect 160645 220904 160650 220960
rect 160706 220904 164514 220960
rect 164570 220904 164575 220960
rect 160645 220902 164575 220904
rect 160645 220899 160711 220902
rect 164509 220899 164575 220902
rect 180793 220962 180859 220965
rect 185025 220962 185091 220965
rect 180793 220960 185091 220962
rect 180793 220904 180798 220960
rect 180854 220904 185030 220960
rect 185086 220904 185091 220960
rect 180793 220902 185091 220904
rect 180793 220899 180859 220902
rect 185025 220899 185091 220902
rect 513557 220962 513623 220965
rect 599485 220962 599551 220965
rect 513557 220960 599551 220962
rect 513557 220904 513562 220960
rect 513618 220904 599490 220960
rect 599546 220904 599551 220960
rect 513557 220902 599551 220904
rect 513557 220899 513623 220902
rect 599485 220899 599551 220902
rect 185853 220826 185919 220829
rect 190407 220826 190473 220829
rect 185853 220824 190473 220826
rect 185853 220768 185858 220824
rect 185914 220768 190412 220824
rect 190468 220768 190473 220824
rect 185853 220766 190473 220768
rect 185853 220763 185919 220766
rect 190407 220763 190473 220766
rect 176561 220690 176627 220693
rect 181069 220690 181135 220693
rect 176561 220688 181135 220690
rect 176561 220632 176566 220688
rect 176622 220632 181074 220688
rect 181130 220632 181135 220688
rect 176561 220630 181135 220632
rect 176561 220627 176627 220630
rect 181069 220627 181135 220630
rect 673085 220690 673151 220693
rect 673085 220688 676292 220690
rect 673085 220632 673090 220688
rect 673146 220632 676292 220688
rect 673085 220630 676292 220632
rect 673085 220627 673151 220630
rect 150709 220554 150775 220557
rect 151905 220554 151971 220557
rect 150709 220552 151971 220554
rect 150709 220496 150714 220552
rect 150770 220496 151910 220552
rect 151966 220496 151971 220552
rect 150709 220494 151971 220496
rect 150709 220491 150775 220494
rect 151905 220491 151971 220494
rect 561765 220554 561831 220557
rect 563145 220554 563211 220557
rect 561765 220552 563211 220554
rect 561765 220496 561770 220552
rect 561826 220496 563150 220552
rect 563206 220496 563211 220552
rect 561765 220494 563211 220496
rect 561765 220491 561831 220494
rect 563145 220491 563211 220494
rect 565629 220554 565695 220557
rect 569953 220554 570019 220557
rect 565629 220552 570019 220554
rect 565629 220496 565634 220552
rect 565690 220496 569958 220552
rect 570014 220496 570019 220552
rect 565629 220494 570019 220496
rect 565629 220491 565695 220494
rect 569953 220491 570019 220494
rect 654133 220418 654199 220421
rect 667013 220418 667079 220421
rect 654133 220416 667079 220418
rect 654133 220360 654138 220416
rect 654194 220360 667018 220416
rect 667074 220360 667079 220416
rect 654133 220358 667079 220360
rect 654133 220355 654199 220358
rect 667013 220355 667079 220358
rect 486969 220282 487035 220285
rect 611629 220282 611695 220285
rect 486969 220280 611695 220282
rect 486969 220224 486974 220280
rect 487030 220224 611634 220280
rect 611690 220224 611695 220280
rect 486969 220222 611695 220224
rect 486969 220219 487035 220222
rect 611629 220219 611695 220222
rect 672441 220282 672507 220285
rect 672441 220280 676292 220282
rect 672441 220224 672446 220280
rect 672502 220224 676292 220280
rect 672441 220222 676292 220224
rect 672441 220219 672507 220222
rect 152181 220146 152247 220149
rect 154389 220146 154455 220149
rect 152181 220144 154455 220146
rect 152181 220088 152186 220144
rect 152242 220088 154394 220144
rect 154450 220088 154455 220144
rect 152181 220086 154455 220088
rect 152181 220083 152247 220086
rect 154389 220083 154455 220086
rect 190269 220010 190335 220013
rect 190637 220010 190703 220013
rect 190269 220008 190703 220010
rect 190269 219952 190274 220008
rect 190330 219952 190642 220008
rect 190698 219952 190703 220008
rect 190269 219950 190703 219952
rect 190269 219947 190335 219950
rect 190637 219947 190703 219950
rect 515121 220010 515187 220013
rect 617149 220010 617215 220013
rect 515121 220008 617215 220010
rect 515121 219952 515126 220008
rect 515182 219952 617154 220008
rect 617210 219952 617215 220008
rect 515121 219950 617215 219952
rect 515121 219947 515187 219950
rect 617149 219947 617215 219950
rect 151813 219874 151879 219877
rect 156321 219874 156387 219877
rect 151813 219872 156387 219874
rect 151813 219816 151818 219872
rect 151874 219816 156326 219872
rect 156382 219816 156387 219872
rect 151813 219814 156387 219816
rect 151813 219811 151879 219814
rect 156321 219811 156387 219814
rect 645853 219874 645919 219877
rect 675477 219874 675543 219877
rect 645853 219872 675543 219874
rect 645853 219816 645858 219872
rect 645914 219816 675482 219872
rect 675538 219816 675543 219872
rect 645853 219814 675543 219816
rect 645853 219811 645919 219814
rect 675477 219811 675543 219814
rect 676024 219812 676030 219876
rect 676094 219874 676100 219876
rect 676094 219814 676292 219874
rect 676094 219812 676100 219814
rect 492949 219738 493015 219741
rect 493685 219738 493751 219741
rect 612733 219738 612799 219741
rect 492949 219736 612799 219738
rect 492949 219680 492954 219736
rect 493010 219680 493690 219736
rect 493746 219680 612738 219736
rect 612794 219680 612799 219736
rect 492949 219678 612799 219680
rect 492949 219675 493015 219678
rect 493685 219675 493751 219678
rect 612733 219675 612799 219678
rect 520181 219466 520247 219469
rect 618437 219466 618503 219469
rect 520181 219464 618503 219466
rect 520181 219408 520186 219464
rect 520242 219408 618442 219464
rect 618498 219408 618503 219464
rect 520181 219406 618503 219408
rect 520181 219403 520247 219406
rect 618437 219403 618503 219406
rect 666829 219466 666895 219469
rect 666829 219464 676292 219466
rect 666829 219408 666834 219464
rect 666890 219408 676292 219464
rect 666829 219406 676292 219408
rect 666829 219403 666895 219406
rect 572529 219194 572595 219197
rect 574737 219194 574803 219197
rect 572529 219192 574803 219194
rect 572529 219136 572534 219192
rect 572590 219136 574742 219192
rect 574798 219136 574803 219192
rect 572529 219134 574803 219136
rect 572529 219131 572595 219134
rect 574737 219131 574803 219134
rect 563007 219058 563073 219061
rect 675109 219058 675175 219061
rect 563007 219056 568498 219058
rect 563007 219000 563012 219056
rect 563068 219000 568498 219056
rect 563007 218998 568498 219000
rect 563007 218995 563073 218998
rect 568438 218922 568498 218998
rect 675109 219056 676292 219058
rect 675109 219000 675114 219056
rect 675170 219000 676292 219056
rect 675109 218998 676292 219000
rect 675109 218995 675175 218998
rect 572529 218922 572595 218925
rect 568438 218920 572595 218922
rect 568438 218864 572534 218920
rect 572590 218864 572595 218920
rect 568438 218862 572595 218864
rect 572529 218859 572595 218862
rect 656801 218922 656867 218925
rect 669446 218922 669452 218924
rect 656801 218920 669452 218922
rect 656801 218864 656806 218920
rect 656862 218864 669452 218920
rect 656801 218862 669452 218864
rect 656801 218859 656867 218862
rect 669446 218860 669452 218862
rect 669516 218860 669522 218924
rect 547413 218786 547479 218789
rect 548609 218786 548675 218789
rect 547413 218784 548675 218786
rect 547413 218728 547418 218784
rect 547474 218728 548614 218784
rect 548670 218728 548675 218784
rect 547413 218726 548675 218728
rect 547413 218723 547479 218726
rect 548609 218723 548675 218726
rect 567653 218786 567719 218789
rect 568297 218786 568363 218789
rect 567653 218784 568363 218786
rect 567653 218728 567658 218784
rect 567714 218728 568302 218784
rect 568358 218728 568363 218784
rect 567653 218726 568363 218728
rect 567653 218723 567719 218726
rect 568297 218723 568363 218726
rect 560293 218650 560359 218653
rect 561673 218650 561739 218653
rect 560293 218648 561739 218650
rect 560293 218592 560298 218648
rect 560354 218592 561678 218648
rect 561734 218592 561739 218648
rect 560293 218590 561739 218592
rect 560293 218587 560359 218590
rect 561673 218587 561739 218590
rect 648429 218650 648495 218653
rect 675477 218650 675543 218653
rect 648429 218648 675543 218650
rect 648429 218592 648434 218648
rect 648490 218592 675482 218648
rect 675538 218592 675543 218648
rect 648429 218590 675543 218592
rect 648429 218587 648495 218590
rect 675477 218587 675543 218590
rect 675702 218588 675708 218652
rect 675772 218650 675778 218652
rect 675772 218590 676292 218650
rect 675772 218588 675778 218590
rect 142429 218514 142495 218517
rect 146569 218514 146635 218517
rect 142429 218512 146635 218514
rect 142429 218456 142434 218512
rect 142490 218456 146574 218512
rect 146630 218456 146635 218512
rect 142429 218454 146635 218456
rect 142429 218451 142495 218454
rect 146569 218451 146635 218454
rect 132493 218378 132559 218381
rect 136725 218378 136791 218381
rect 132493 218376 136791 218378
rect 132493 218320 132498 218376
rect 132554 218320 136730 218376
rect 136786 218320 136791 218376
rect 132493 218318 136791 218320
rect 132493 218315 132559 218318
rect 136725 218315 136791 218318
rect 494697 218378 494763 218381
rect 630673 218378 630739 218381
rect 494697 218376 630739 218378
rect 494697 218320 494702 218376
rect 494758 218320 630678 218376
rect 630734 218320 630739 218376
rect 494697 218318 630739 218320
rect 494697 218315 494763 218318
rect 630673 218315 630739 218318
rect 669630 218180 669636 218244
rect 669700 218242 669706 218244
rect 670601 218242 670667 218245
rect 669700 218240 670667 218242
rect 669700 218184 670606 218240
rect 670662 218184 670667 218240
rect 669700 218182 670667 218184
rect 669700 218180 669706 218182
rect 670601 218179 670667 218182
rect 674925 218242 674991 218245
rect 674925 218240 676292 218242
rect 674925 218184 674930 218240
rect 674986 218184 676292 218240
rect 674925 218182 676292 218184
rect 674925 218179 674991 218182
rect 487797 218106 487863 218109
rect 623957 218106 624023 218109
rect 487797 218104 624023 218106
rect 487797 218048 487802 218104
rect 487858 218048 623962 218104
rect 624018 218048 624023 218104
rect 487797 218046 624023 218048
rect 487797 218043 487863 218046
rect 623957 218043 624023 218046
rect 35525 217970 35591 217973
rect 56041 217970 56107 217973
rect 35525 217968 56107 217970
rect 35525 217912 35530 217968
rect 35586 217912 56046 217968
rect 56102 217912 56107 217968
rect 35525 217910 56107 217912
rect 35525 217907 35591 217910
rect 56041 217907 56107 217910
rect 667013 217970 667079 217973
rect 670366 217970 670372 217972
rect 667013 217968 670372 217970
rect 667013 217912 667018 217968
rect 667074 217912 670372 217968
rect 667013 217910 670372 217912
rect 667013 217907 667079 217910
rect 670366 217908 670372 217910
rect 670436 217908 670442 217972
rect 672625 217970 672691 217973
rect 675661 217970 675727 217973
rect 672625 217968 675727 217970
rect 672625 217912 672630 217968
rect 672686 217912 675666 217968
rect 675722 217912 675727 217968
rect 672625 217910 675727 217912
rect 672625 217907 672691 217910
rect 675661 217907 675727 217910
rect 675886 217908 675892 217972
rect 675956 217970 675962 217972
rect 675956 217910 676230 217970
rect 675956 217908 675962 217910
rect 564801 217834 564867 217837
rect 571885 217834 571951 217837
rect 564801 217832 571951 217834
rect 564801 217776 564806 217832
rect 564862 217776 571890 217832
rect 571946 217776 571951 217832
rect 564801 217774 571951 217776
rect 564801 217771 564867 217774
rect 571885 217771 571951 217774
rect 572069 217834 572135 217837
rect 574369 217834 574435 217837
rect 572069 217832 574435 217834
rect 572069 217776 572074 217832
rect 572130 217776 574374 217832
rect 574430 217776 574435 217832
rect 572069 217774 574435 217776
rect 676170 217834 676230 217910
rect 676170 217774 676292 217834
rect 572069 217771 572135 217774
rect 574369 217771 574435 217774
rect 510981 217564 511047 217565
rect 519997 217564 520063 217565
rect 510981 217562 511028 217564
rect 510936 217560 511028 217562
rect 510936 217504 510986 217560
rect 510936 217502 511028 217504
rect 510981 217500 511028 217502
rect 511092 217500 511098 217564
rect 519997 217562 520044 217564
rect 519952 217560 520044 217562
rect 519952 217504 520002 217560
rect 519952 217502 520044 217504
rect 519997 217500 520044 217502
rect 520108 217500 520114 217564
rect 531497 217562 531563 217565
rect 532509 217564 532575 217565
rect 532509 217562 532556 217564
rect 531497 217560 532556 217562
rect 531497 217504 531502 217560
rect 531558 217504 532514 217560
rect 531497 217502 532556 217504
rect 510981 217499 511047 217500
rect 519997 217499 520063 217500
rect 531497 217499 531563 217502
rect 532509 217500 532556 217502
rect 532620 217500 532626 217564
rect 560753 217562 560819 217565
rect 560937 217562 561003 217565
rect 563145 217562 563211 217565
rect 560753 217560 563211 217562
rect 560753 217504 560758 217560
rect 560814 217504 560942 217560
rect 560998 217504 563150 217560
rect 563206 217504 563211 217560
rect 560753 217502 563211 217504
rect 532509 217499 532575 217500
rect 560753 217499 560819 217502
rect 560937 217499 561003 217502
rect 563145 217499 563211 217502
rect 572529 217562 572595 217565
rect 574185 217562 574251 217565
rect 572529 217560 574251 217562
rect 572529 217504 572534 217560
rect 572590 217504 574190 217560
rect 574246 217504 574251 217560
rect 572529 217502 574251 217504
rect 572529 217499 572595 217502
rect 574185 217499 574251 217502
rect 653765 217562 653831 217565
rect 672073 217562 672139 217565
rect 653765 217560 672139 217562
rect 653765 217504 653770 217560
rect 653826 217504 672078 217560
rect 672134 217504 672139 217560
rect 653765 217502 672139 217504
rect 653765 217499 653831 217502
rect 672073 217499 672139 217502
rect 673085 217426 673151 217429
rect 673085 217424 676292 217426
rect 673085 217368 673090 217424
rect 673146 217368 676292 217424
rect 673085 217366 676292 217368
rect 673085 217363 673151 217366
rect 500953 217290 501019 217293
rect 595161 217290 595227 217293
rect 500953 217288 595227 217290
rect 500953 217232 500958 217288
rect 501014 217232 595166 217288
rect 595222 217232 595227 217288
rect 500953 217230 595227 217232
rect 500953 217227 501019 217230
rect 595161 217227 595227 217230
rect 651097 217290 651163 217293
rect 651097 217288 663810 217290
rect 651097 217232 651102 217288
rect 651158 217232 663810 217288
rect 651097 217230 663810 217232
rect 651097 217227 651163 217230
rect 488809 217154 488875 217157
rect 495157 217154 495223 217157
rect 488809 217152 491034 217154
rect 488809 217096 488814 217152
rect 488870 217096 491034 217152
rect 488809 217094 491034 217096
rect 488809 217091 488875 217094
rect 490974 216746 491034 217094
rect 495157 217152 500234 217154
rect 495157 217096 495162 217152
rect 495218 217096 500234 217152
rect 495157 217094 500234 217096
rect 495157 217091 495223 217094
rect 500174 217018 500234 217094
rect 595713 217018 595779 217021
rect 500174 217016 595779 217018
rect 500174 216960 595718 217016
rect 595774 216960 595779 217016
rect 500174 216958 595779 216960
rect 595713 216955 595779 216958
rect 663750 216882 663810 217230
rect 670366 217092 670372 217156
rect 670436 217154 670442 217156
rect 670436 217094 676230 217154
rect 670436 217092 670442 217094
rect 676170 217018 676230 217094
rect 676170 216958 676292 217018
rect 673453 216882 673519 216885
rect 663750 216880 673519 216882
rect 663750 216824 673458 216880
rect 673514 216824 673519 216880
rect 663750 216822 673519 216824
rect 673453 216819 673519 216822
rect 575473 216746 575539 216749
rect 490974 216744 575539 216746
rect 490974 216688 575478 216744
rect 575534 216688 575539 216744
rect 490974 216686 575539 216688
rect 575473 216683 575539 216686
rect 669405 216612 669471 216613
rect 669405 216610 669452 216612
rect 669360 216608 669452 216610
rect 669360 216552 669410 216608
rect 669360 216550 669452 216552
rect 669405 216548 669452 216550
rect 669516 216548 669522 216612
rect 673453 216610 673519 216613
rect 673453 216608 676292 216610
rect 673453 216552 673458 216608
rect 673514 216552 676292 216608
rect 673453 216550 676292 216552
rect 669405 216547 669471 216548
rect 673453 216547 673519 216550
rect 39941 216474 40007 216477
rect 43069 216474 43135 216477
rect 39941 216472 43135 216474
rect 39941 216416 39946 216472
rect 40002 216416 43074 216472
rect 43130 216416 43135 216472
rect 39941 216414 43135 216416
rect 39941 216411 40007 216414
rect 43069 216411 43135 216414
rect 670509 216474 670575 216477
rect 673085 216474 673151 216477
rect 670509 216472 673151 216474
rect 670509 216416 670514 216472
rect 670570 216416 673090 216472
rect 673146 216416 673151 216472
rect 670509 216414 673151 216416
rect 670509 216411 670575 216414
rect 673085 216411 673151 216414
rect 39573 216202 39639 216205
rect 42885 216202 42951 216205
rect 672073 216202 672139 216205
rect 39573 216200 42951 216202
rect 39573 216144 39578 216200
rect 39634 216144 42890 216200
rect 42946 216144 42951 216200
rect 39573 216142 42951 216144
rect 39573 216139 39639 216142
rect 42885 216139 42951 216142
rect 663750 216200 672139 216202
rect 663750 216144 672078 216200
rect 672134 216144 672139 216200
rect 663750 216142 672139 216144
rect 520038 215868 520044 215932
rect 520108 215930 520114 215932
rect 617793 215930 617859 215933
rect 520108 215928 617859 215930
rect 520108 215872 617798 215928
rect 617854 215872 617859 215928
rect 520108 215870 617859 215872
rect 520108 215868 520114 215870
rect 617793 215867 617859 215870
rect 511022 215596 511028 215660
rect 511092 215658 511098 215660
rect 599025 215658 599091 215661
rect 511092 215656 599091 215658
rect 511092 215600 599030 215656
rect 599086 215600 599091 215656
rect 511092 215598 599091 215600
rect 511092 215596 511098 215598
rect 599025 215595 599091 215598
rect 532550 215324 532556 215388
rect 532620 215386 532626 215388
rect 621105 215386 621171 215389
rect 532620 215384 621171 215386
rect 532620 215328 621110 215384
rect 621166 215328 621171 215384
rect 532620 215326 621171 215328
rect 532620 215324 532626 215326
rect 621105 215323 621171 215326
rect 659561 215386 659627 215389
rect 663750 215386 663810 216142
rect 672073 216139 672139 216142
rect 673085 216202 673151 216205
rect 673085 216200 676292 216202
rect 673085 216144 673090 216200
rect 673146 216144 676292 216200
rect 673085 216142 676292 216144
rect 673085 216139 673151 216142
rect 666645 215930 666711 215933
rect 666645 215928 676230 215930
rect 666645 215872 666650 215928
rect 666706 215872 676230 215928
rect 666645 215870 676230 215872
rect 666645 215867 666711 215870
rect 676170 215794 676230 215870
rect 676170 215734 676292 215794
rect 664621 215658 664687 215661
rect 669589 215658 669655 215661
rect 664621 215656 669655 215658
rect 664621 215600 664626 215656
rect 664682 215600 669594 215656
rect 669650 215600 669655 215656
rect 664621 215598 669655 215600
rect 664621 215595 664687 215598
rect 669589 215595 669655 215598
rect 672073 215658 672139 215661
rect 675661 215658 675727 215661
rect 672073 215656 675727 215658
rect 672073 215600 672078 215656
rect 672134 215600 675666 215656
rect 675722 215600 675727 215656
rect 672073 215598 675727 215600
rect 672073 215595 672139 215598
rect 675661 215595 675727 215598
rect 675886 215460 675892 215524
rect 675956 215522 675962 215524
rect 675956 215462 676230 215522
rect 675956 215460 675962 215462
rect 673453 215386 673519 215389
rect 659561 215384 663810 215386
rect 659561 215328 659566 215384
rect 659622 215328 663810 215384
rect 659561 215326 663810 215328
rect 669638 215384 673519 215386
rect 669638 215328 673458 215384
rect 673514 215328 673519 215384
rect 669638 215326 673519 215328
rect 676170 215386 676230 215462
rect 676170 215326 676292 215386
rect 659561 215323 659627 215326
rect 53281 215114 53347 215117
rect 41462 215112 53347 215114
rect 41462 215056 53286 215112
rect 53342 215056 53347 215112
rect 41462 215054 53347 215056
rect 41462 214948 41522 215054
rect 53281 215051 53347 215054
rect 669405 215114 669471 215117
rect 669638 215114 669698 215326
rect 673453 215323 673519 215326
rect 669405 215112 669698 215114
rect 669405 215056 669410 215112
rect 669466 215056 669698 215112
rect 669405 215054 669698 215056
rect 669405 215051 669471 215054
rect 674465 214978 674531 214981
rect 674465 214976 676292 214978
rect 674465 214920 674470 214976
rect 674526 214920 676292 214976
rect 674465 214918 676292 214920
rect 674465 214915 674531 214918
rect 675661 214706 675727 214709
rect 663750 214704 675727 214706
rect 663750 214648 675666 214704
rect 675722 214648 675727 214704
rect 663750 214646 675727 214648
rect 660389 214570 660455 214573
rect 663750 214570 663810 214646
rect 675661 214643 675727 214646
rect 660389 214568 663810 214570
rect 35758 214301 35818 214540
rect 660389 214512 660394 214568
rect 660450 214512 663810 214568
rect 660389 214510 663810 214512
rect 676029 214570 676095 214573
rect 676029 214568 676292 214570
rect 676029 214512 676034 214568
rect 676090 214512 676292 214568
rect 676029 214510 676292 214512
rect 660389 214507 660455 214510
rect 676029 214507 676095 214510
rect 673913 214434 673979 214437
rect 675845 214434 675911 214437
rect 673913 214432 675911 214434
rect 35525 214298 35591 214301
rect 35525 214296 35634 214298
rect 35525 214240 35530 214296
rect 35586 214240 35634 214296
rect 35525 214235 35634 214240
rect 35758 214296 35867 214301
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214238 35867 214240
rect 35801 214235 35867 214238
rect 35574 214132 35634 214235
rect 575982 214026 576042 214404
rect 673913 214376 673918 214432
rect 673974 214376 675850 214432
rect 675906 214376 675911 214432
rect 673913 214374 675911 214376
rect 673913 214371 673979 214374
rect 675845 214371 675911 214374
rect 672073 214162 672139 214165
rect 672073 214160 676292 214162
rect 672073 214104 672078 214160
rect 672134 214104 676292 214160
rect 672073 214102 676292 214104
rect 672073 214099 672139 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 674649 213754 674715 213757
rect 674649 213752 676292 213754
rect 35574 213485 35634 213724
rect 674649 213696 674654 213752
rect 674710 213696 676292 213752
rect 674649 213694 676292 213696
rect 674649 213691 674715 213694
rect 672717 213618 672783 213621
rect 663750 213616 672783 213618
rect 663750 213560 672722 213616
rect 672778 213560 672783 213616
rect 663750 213558 672783 213560
rect 35574 213480 35683 213485
rect 35574 213424 35622 213480
rect 35678 213424 35683 213480
rect 35574 213422 35683 213424
rect 35617 213419 35683 213422
rect 661493 213482 661559 213485
rect 663750 213482 663810 213558
rect 672717 213555 672783 213558
rect 661493 213480 663810 213482
rect 661493 213424 661498 213480
rect 661554 213424 663810 213480
rect 661493 213422 663810 213424
rect 661493 213419 661559 213422
rect 672809 213346 672875 213349
rect 672809 213344 676292 213346
rect 672809 213288 672814 213344
rect 672870 213288 676292 213344
rect 672809 213286 676292 213288
rect 672809 213283 672875 213286
rect 658733 213210 658799 213213
rect 672533 213210 672599 213213
rect 658733 213208 672599 213210
rect 658733 213152 658738 213208
rect 658794 213152 672538 213208
rect 672594 213152 672599 213208
rect 658733 213150 672599 213152
rect 658733 213147 658799 213150
rect 672533 213147 672599 213150
rect 35801 213074 35867 213077
rect 35758 213072 35867 213074
rect 35758 213016 35806 213072
rect 35862 213016 35867 213072
rect 35758 213011 35867 213016
rect 35758 212908 35818 213011
rect 675293 212530 675359 212533
rect 675886 212530 675892 212532
rect 675293 212528 675892 212530
rect 675293 212472 675298 212528
rect 675354 212472 675892 212528
rect 675293 212470 675892 212472
rect 675293 212467 675359 212470
rect 675886 212468 675892 212470
rect 675956 212530 675962 212532
rect 683070 212530 683130 212908
rect 675956 212500 683130 212530
rect 675956 212470 683100 212500
rect 675956 212468 675962 212470
rect 44265 212122 44331 212125
rect 41492 212120 44331 212122
rect 41492 212064 44270 212120
rect 44326 212064 44331 212120
rect 41492 212062 44331 212064
rect 44265 212059 44331 212062
rect 575982 211714 576042 212228
rect 672625 212122 672691 212125
rect 672625 212120 676292 212122
rect 672625 212064 672630 212120
rect 672686 212064 676292 212120
rect 672625 212062 676292 212064
rect 672625 212059 672691 212062
rect 578509 211714 578575 211717
rect 575982 211712 578575 211714
rect 575982 211656 578514 211712
rect 578570 211656 578575 211712
rect 575982 211654 578575 211656
rect 578509 211651 578575 211654
rect 676029 211442 676095 211445
rect 676622 211442 676628 211444
rect 676029 211440 676628 211442
rect 676029 211384 676034 211440
rect 676090 211384 676628 211440
rect 676029 211382 676628 211384
rect 676029 211379 676095 211382
rect 676622 211380 676628 211382
rect 676692 211380 676698 211444
rect 44817 211306 44883 211309
rect 41492 211304 44883 211306
rect 41492 211248 44822 211304
rect 44878 211248 44883 211304
rect 41492 211246 44883 211248
rect 44817 211243 44883 211246
rect 35758 210221 35818 210460
rect 35758 210216 35867 210221
rect 35758 210160 35806 210216
rect 35862 210160 35867 210216
rect 35758 210158 35867 210160
rect 35801 210155 35867 210158
rect 41822 210082 41828 210084
rect 41492 210022 41828 210082
rect 41822 210020 41828 210022
rect 41892 210020 41898 210084
rect 575982 209810 576042 210052
rect 579521 209810 579587 209813
rect 575982 209808 579587 209810
rect 575982 209752 579526 209808
rect 579582 209752 579587 209808
rect 575982 209750 579587 209752
rect 579521 209747 579587 209750
rect 35574 209405 35634 209644
rect 35574 209400 35683 209405
rect 35574 209344 35622 209400
rect 35678 209344 35683 209400
rect 35574 209342 35683 209344
rect 35617 209339 35683 209342
rect 35758 208997 35818 209236
rect 35758 208992 35867 208997
rect 35758 208936 35806 208992
rect 35862 208936 35867 208992
rect 35758 208934 35867 208936
rect 35801 208931 35867 208934
rect 40401 208994 40467 208997
rect 42885 208994 42951 208997
rect 40401 208992 42951 208994
rect 40401 208936 40406 208992
rect 40462 208936 42890 208992
rect 42946 208936 42951 208992
rect 40401 208934 42951 208936
rect 40401 208931 40467 208934
rect 42885 208931 42951 208934
rect 35758 208589 35818 208828
rect 35758 208584 35867 208589
rect 35758 208528 35806 208584
rect 35862 208528 35867 208584
rect 35758 208526 35867 208528
rect 35801 208523 35867 208526
rect 44449 208450 44515 208453
rect 41492 208448 44515 208450
rect 41492 208392 44454 208448
rect 44510 208392 44515 208448
rect 41492 208390 44515 208392
rect 44449 208387 44515 208390
rect 40033 208178 40099 208181
rect 41638 208178 41644 208180
rect 40033 208176 41644 208178
rect 40033 208120 40038 208176
rect 40094 208120 41644 208176
rect 40033 208118 41644 208120
rect 40033 208115 40099 208118
rect 41638 208116 41644 208118
rect 41708 208116 41714 208180
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 41462 207770 41522 208012
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 44173 207770 44239 207773
rect 41462 207768 44239 207770
rect 41462 207712 44178 207768
rect 44234 207712 44239 207768
rect 41462 207710 44239 207712
rect 44173 207707 44239 207710
rect 35801 207362 35867 207365
rect 40542 207364 40602 207604
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 35758 207360 35867 207362
rect 35758 207304 35806 207360
rect 35862 207304 35867 207360
rect 35758 207299 35867 207304
rect 40534 207300 40540 207364
rect 40604 207300 40610 207364
rect 35758 207196 35818 207299
rect 40585 206954 40651 206957
rect 42701 206954 42767 206957
rect 40585 206952 42767 206954
rect 40585 206896 40590 206952
rect 40646 206896 42706 206952
rect 42762 206896 42767 206952
rect 40585 206894 42767 206896
rect 40585 206891 40651 206894
rect 42701 206891 42767 206894
rect 674598 206892 674604 206956
rect 674668 206954 674674 206956
rect 675109 206954 675175 206957
rect 674668 206952 675175 206954
rect 674668 206896 675114 206952
rect 675170 206896 675175 206952
rect 674668 206894 675175 206896
rect 674668 206892 674674 206894
rect 675109 206891 675175 206894
rect 40726 206548 40786 206788
rect 40718 206484 40724 206548
rect 40788 206484 40794 206548
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 40910 206140 40970 206380
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 40902 206076 40908 206140
rect 40972 206076 40978 206140
rect 44633 206002 44699 206005
rect 41492 206000 44699 206002
rect 41492 205944 44638 206000
rect 44694 205944 44699 206000
rect 41492 205942 44699 205944
rect 44633 205939 44699 205942
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 669262 205668 669268 205732
rect 669332 205730 669338 205732
rect 669630 205730 669636 205732
rect 669332 205670 669636 205730
rect 669332 205668 669338 205670
rect 669630 205668 669636 205670
rect 669700 205668 669706 205732
rect 35758 205325 35818 205564
rect 669262 205396 669268 205460
rect 669332 205458 669338 205460
rect 669630 205458 669636 205460
rect 669332 205398 669636 205458
rect 669332 205396 669338 205398
rect 669630 205396 669636 205398
rect 669700 205396 669706 205460
rect 35758 205320 35867 205325
rect 35758 205264 35806 205320
rect 35862 205264 35867 205320
rect 35758 205262 35867 205264
rect 35801 205259 35867 205262
rect 44817 205186 44883 205189
rect 41492 205184 44883 205186
rect 41492 205128 44822 205184
rect 44878 205128 44883 205184
rect 41492 205126 44883 205128
rect 44817 205123 44883 205126
rect 674741 205050 674807 205053
rect 675385 205050 675451 205053
rect 674741 205048 675451 205050
rect 674741 204992 674746 205048
rect 674802 204992 675390 205048
rect 675446 204992 675451 205048
rect 674741 204990 675451 204992
rect 674741 204987 674807 204990
rect 675385 204987 675451 204990
rect 41454 204852 41460 204916
rect 41524 204914 41530 204916
rect 46197 204914 46263 204917
rect 41524 204912 46263 204914
rect 41524 204856 46202 204912
rect 46258 204856 46263 204912
rect 41524 204854 46263 204856
rect 41524 204852 41530 204854
rect 46197 204851 46263 204854
rect 589457 204778 589523 204781
rect 589457 204776 592572 204778
rect 35758 204509 35818 204748
rect 589457 204720 589462 204776
rect 589518 204720 592572 204776
rect 589457 204718 592572 204720
rect 589457 204715 589523 204718
rect 35758 204504 35867 204509
rect 35758 204448 35806 204504
rect 35862 204448 35867 204504
rect 35758 204446 35867 204448
rect 35801 204443 35867 204446
rect 41505 204506 41571 204509
rect 43713 204506 43779 204509
rect 41505 204504 43779 204506
rect 41505 204448 41510 204504
rect 41566 204448 43718 204504
rect 43774 204448 43779 204504
rect 41505 204446 43779 204448
rect 41505 204443 41571 204446
rect 43713 204443 43779 204446
rect 41462 204100 41522 204340
rect 674925 204234 674991 204237
rect 675385 204234 675451 204237
rect 674925 204232 675451 204234
rect 674925 204176 674930 204232
rect 674986 204176 675390 204232
rect 675446 204176 675451 204232
rect 674925 204174 675451 204176
rect 674925 204171 674991 204174
rect 675385 204171 675451 204174
rect 41454 204036 41460 204100
rect 41524 204036 41530 204100
rect 41689 204098 41755 204101
rect 43437 204098 43503 204101
rect 669129 204098 669195 204101
rect 41689 204096 43503 204098
rect 41689 204040 41694 204096
rect 41750 204040 43442 204096
rect 43498 204040 43503 204096
rect 41689 204038 43503 204040
rect 41689 204035 41755 204038
rect 43437 204035 43503 204038
rect 666694 204096 669195 204098
rect 666694 204040 669134 204096
rect 669190 204040 669195 204096
rect 666694 204038 669195 204040
rect 666694 204030 666754 204038
rect 669129 204035 669195 204038
rect 666356 203970 666754 204030
rect 35758 203693 35818 203932
rect 35758 203688 35867 203693
rect 35758 203632 35806 203688
rect 35862 203632 35867 203688
rect 35758 203630 35867 203632
rect 35801 203627 35867 203630
rect 39941 203690 40007 203693
rect 43253 203690 43319 203693
rect 39941 203688 43319 203690
rect 39941 203632 39946 203688
rect 40002 203632 43258 203688
rect 43314 203632 43319 203688
rect 39941 203630 43319 203632
rect 39941 203627 40007 203630
rect 43253 203627 43319 203630
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 578325 203219 578391 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 669405 202874 669471 202877
rect 674925 202874 674991 202877
rect 669405 202872 674991 202874
rect 669405 202816 669410 202872
rect 669466 202816 674930 202872
rect 674986 202816 674991 202872
rect 669405 202814 674991 202816
rect 669405 202811 669471 202814
rect 674925 202811 674991 202814
rect 675753 202738 675819 202741
rect 676438 202738 676444 202740
rect 675753 202736 676444 202738
rect 675753 202680 675758 202736
rect 675814 202680 676444 202736
rect 675753 202678 676444 202680
rect 675753 202675 675819 202678
rect 676438 202676 676444 202678
rect 676508 202676 676514 202740
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 672993 201378 673059 201381
rect 675477 201378 675543 201381
rect 672993 201376 675543 201378
rect 575982 200834 576042 201348
rect 672993 201320 672998 201376
rect 673054 201320 675482 201376
rect 675538 201320 675543 201376
rect 672993 201318 675543 201320
rect 672993 201315 673059 201318
rect 675477 201315 675543 201318
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 672574 200772 672580 200836
rect 672644 200834 672650 200836
rect 672993 200834 673059 200837
rect 672644 200832 673059 200834
rect 672644 200776 672998 200832
rect 673054 200776 673059 200832
rect 672644 200774 673059 200776
rect 672644 200772 672650 200774
rect 672993 200771 673059 200774
rect 675753 200018 675819 200021
rect 676622 200018 676628 200020
rect 675753 200016 676628 200018
rect 675753 199960 675758 200016
rect 675814 199960 676628 200016
rect 675753 199958 676628 199960
rect 675753 199955 675819 199958
rect 676622 199956 676628 199958
rect 676692 199956 676698 200020
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 672073 199746 672139 199749
rect 674925 199746 674991 199749
rect 672073 199744 674991 199746
rect 672073 199688 672078 199744
rect 672134 199688 674930 199744
rect 674986 199688 674991 199744
rect 672073 199686 674991 199688
rect 672073 199683 672139 199686
rect 674925 199683 674991 199686
rect 668393 199202 668459 199205
rect 666694 199200 668459 199202
rect 575982 198930 576042 199172
rect 666694 199144 668398 199200
rect 668454 199144 668459 199200
rect 666694 199142 668459 199144
rect 666694 199134 666754 199142
rect 668393 199139 668459 199142
rect 666356 199074 666754 199134
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 37917 198794 37983 198797
rect 42006 198794 42012 198796
rect 37917 198792 42012 198794
rect 37917 198736 37922 198792
rect 37978 198736 42012 198792
rect 37917 198734 42012 198736
rect 37917 198731 37983 198734
rect 42006 198732 42012 198734
rect 42076 198732 42082 198796
rect 669129 198794 669195 198797
rect 670734 198794 670740 198796
rect 669129 198792 670740 198794
rect 669129 198736 669134 198792
rect 669190 198736 670740 198792
rect 669129 198734 670740 198736
rect 669129 198731 669195 198734
rect 670734 198732 670740 198734
rect 670804 198732 670810 198796
rect 666645 198522 666711 198525
rect 675109 198522 675175 198525
rect 666645 198520 675175 198522
rect 666645 198464 666650 198520
rect 666706 198464 675114 198520
rect 675170 198464 675175 198520
rect 666645 198462 675175 198464
rect 666645 198459 666711 198462
rect 675109 198459 675175 198462
rect 590377 198250 590443 198253
rect 670509 198250 670575 198253
rect 675477 198250 675543 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 670509 198248 675543 198250
rect 670509 198192 670514 198248
rect 670570 198192 675482 198248
rect 675538 198192 675543 198248
rect 670509 198190 675543 198192
rect 590377 198187 590443 198190
rect 670509 198187 670575 198190
rect 675477 198187 675543 198190
rect 673269 197978 673335 197981
rect 676806 197978 676812 197980
rect 673269 197976 676812 197978
rect 673269 197920 673274 197976
rect 673330 197920 676812 197976
rect 673269 197918 676812 197920
rect 673269 197915 673335 197918
rect 676806 197916 676812 197918
rect 676876 197916 676882 197980
rect 42425 197298 42491 197301
rect 44449 197298 44515 197301
rect 42425 197296 44515 197298
rect 42425 197240 42430 197296
rect 42486 197240 44454 197296
rect 44510 197240 44515 197296
rect 42425 197238 44515 197240
rect 42425 197235 42491 197238
rect 44449 197235 44515 197238
rect 674465 197162 674531 197165
rect 675385 197162 675451 197165
rect 674465 197160 675451 197162
rect 674465 197104 674470 197160
rect 674526 197104 675390 197160
rect 675446 197104 675451 197160
rect 674465 197102 675451 197104
rect 674465 197099 674531 197102
rect 675385 197099 675451 197102
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 578509 196419 578575 196422
rect 669262 196012 669268 196076
rect 669332 196074 669338 196076
rect 669630 196074 669636 196076
rect 669332 196014 669636 196074
rect 669332 196012 669338 196014
rect 669630 196012 669636 196014
rect 669700 196012 669706 196076
rect 41965 195668 42031 195669
rect 41965 195664 42012 195668
rect 42076 195666 42082 195668
rect 41965 195608 41970 195664
rect 41965 195604 42012 195608
rect 42076 195606 42122 195666
rect 42076 195604 42082 195606
rect 41965 195603 42031 195604
rect 41781 195260 41847 195261
rect 41781 195256 41828 195260
rect 41892 195258 41898 195260
rect 41781 195200 41786 195256
rect 41781 195196 41828 195200
rect 41892 195198 41938 195258
rect 41892 195196 41898 195198
rect 41781 195195 41847 195196
rect 40902 194924 40908 194988
rect 40972 194986 40978 194988
rect 42241 194986 42307 194989
rect 579521 194986 579587 194989
rect 40972 194984 42307 194986
rect 40972 194928 42246 194984
rect 42302 194928 42307 194984
rect 40972 194926 42307 194928
rect 40972 194924 40978 194926
rect 42241 194923 42307 194926
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 675753 194578 675819 194581
rect 676254 194578 676260 194580
rect 675753 194576 676260 194578
rect 675753 194520 675758 194576
rect 675814 194520 676260 194576
rect 675753 194518 676260 194520
rect 675753 194515 675819 194518
rect 676254 194516 676260 194518
rect 676324 194516 676330 194580
rect 668117 194306 668183 194309
rect 666694 194304 668183 194306
rect 666694 194248 668122 194304
rect 668178 194248 668183 194304
rect 666694 194246 668183 194248
rect 666694 194238 666754 194246
rect 668117 194243 668183 194246
rect 666356 194178 666754 194238
rect 40718 193428 40724 193492
rect 40788 193490 40794 193492
rect 41781 193490 41847 193493
rect 40788 193488 41847 193490
rect 40788 193432 41786 193488
rect 41842 193432 41847 193488
rect 40788 193430 41847 193432
rect 40788 193428 40794 193430
rect 41781 193427 41847 193430
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 675753 193218 675819 193221
rect 676070 193218 676076 193220
rect 675753 193216 676076 193218
rect 675753 193160 675758 193216
rect 675814 193160 676076 193216
rect 675753 193158 676076 193160
rect 675753 193155 675819 193158
rect 676070 193156 676076 193158
rect 676140 193156 676146 193220
rect 675661 192810 675727 192813
rect 675886 192810 675892 192812
rect 675661 192808 675892 192810
rect 675661 192752 675666 192808
rect 675722 192752 675892 192808
rect 675661 192750 675892 192752
rect 675661 192747 675727 192750
rect 675886 192748 675892 192750
rect 675956 192748 675962 192812
rect 575982 192266 576042 192644
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 589457 191722 589523 191725
rect 668393 191722 668459 191725
rect 669446 191722 669452 191724
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 668393 191720 669452 191722
rect 668393 191664 668398 191720
rect 668454 191664 669452 191720
rect 668393 191662 669452 191664
rect 589457 191659 589523 191662
rect 668393 191659 668459 191662
rect 669446 191660 669452 191662
rect 669516 191660 669522 191724
rect 42057 191586 42123 191589
rect 44817 191586 44883 191589
rect 42057 191584 44883 191586
rect 42057 191528 42062 191584
rect 42118 191528 44822 191584
rect 44878 191528 44883 191584
rect 42057 191526 44883 191528
rect 42057 191523 42123 191526
rect 44817 191523 44883 191526
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 43713 190498 43779 190501
rect 42425 190496 43779 190498
rect 42425 190440 42430 190496
rect 42486 190440 43718 190496
rect 43774 190440 43779 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 42425 190438 43779 190440
rect 42425 190435 42491 190438
rect 43713 190435 43779 190438
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 668945 189410 669011 189413
rect 666694 189408 669011 189410
rect 666694 189352 668950 189408
rect 669006 189352 669011 189408
rect 666694 189350 669011 189352
rect 666694 189342 666754 189350
rect 668945 189347 669011 189350
rect 666356 189282 666754 189342
rect 675334 189076 675340 189140
rect 675404 189138 675410 189140
rect 676029 189138 676095 189141
rect 675404 189136 676095 189138
rect 675404 189080 676034 189136
rect 676090 189080 676095 189136
rect 675404 189078 676095 189080
rect 675404 189076 675410 189078
rect 676029 189075 676095 189078
rect 667013 188866 667079 188869
rect 675109 188866 675175 188869
rect 667013 188864 675175 188866
rect 667013 188808 667018 188864
rect 667074 188808 675114 188864
rect 675170 188808 675175 188864
rect 667013 188806 675175 188808
rect 667013 188803 667079 188806
rect 675109 188803 675175 188806
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42241 187642 42307 187645
rect 44633 187642 44699 187645
rect 42241 187640 44699 187642
rect 42241 187584 42246 187640
rect 42302 187584 44638 187640
rect 44694 187584 44699 187640
rect 42241 187582 44699 187584
rect 42241 187579 42307 187582
rect 44633 187579 44699 187582
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 40534 186356 40540 186420
rect 40604 186418 40610 186420
rect 41781 186418 41847 186421
rect 40604 186416 41847 186418
rect 40604 186360 41786 186416
rect 41842 186360 41847 186416
rect 40604 186358 41847 186360
rect 40604 186356 40610 186358
rect 41781 186355 41847 186358
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 41454 185948 41460 186012
rect 41524 186010 41530 186012
rect 41781 186010 41847 186013
rect 41524 186008 41847 186010
rect 41524 185952 41786 186008
rect 41842 185952 41847 186008
rect 41524 185950 41847 185952
rect 41524 185948 41530 185950
rect 41781 185947 41847 185950
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 667933 184514 667999 184517
rect 666694 184512 667999 184514
rect 666694 184456 667938 184512
rect 667994 184456 667999 184512
rect 666694 184454 667999 184456
rect 666694 184446 666754 184454
rect 667933 184451 667999 184454
rect 666356 184386 666754 184446
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 42425 183562 42491 183565
rect 43897 183562 43963 183565
rect 42425 183560 43963 183562
rect 42425 183504 42430 183560
rect 42486 183504 43902 183560
rect 43958 183504 43963 183560
rect 42425 183502 43963 183504
rect 42425 183499 42491 183502
rect 43897 183499 43963 183502
rect 589457 183562 589523 183565
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 589457 183499 589523 183502
rect 42241 183290 42307 183293
rect 44173 183290 44239 183293
rect 42241 183288 44239 183290
rect 42241 183232 42246 183288
rect 42302 183232 44178 183288
rect 44234 183232 44239 183288
rect 42241 183230 44239 183232
rect 42241 183227 42307 183230
rect 44173 183227 44239 183230
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 673085 181524 673151 181525
rect 673085 181522 673132 181524
rect 673040 181520 673132 181522
rect 673040 181464 673090 181520
rect 673040 181462 673132 181464
rect 673085 181460 673132 181462
rect 673196 181460 673202 181524
rect 673085 181459 673151 181460
rect 667565 181386 667631 181389
rect 667565 181384 669330 181386
rect 667565 181328 667570 181384
rect 667626 181328 669330 181384
rect 667565 181326 669330 181328
rect 667565 181323 667631 181326
rect 669270 181250 669330 181326
rect 676213 181250 676279 181253
rect 669270 181248 676279 181250
rect 669270 181192 676218 181248
rect 676274 181192 676279 181248
rect 669270 181190 676279 181192
rect 676213 181187 676279 181190
rect 42057 180842 42123 180845
rect 51717 180842 51783 180845
rect 42057 180840 51783 180842
rect 42057 180784 42062 180840
rect 42118 180784 51722 180840
rect 51778 180784 51783 180840
rect 42057 180782 51783 180784
rect 42057 180779 42123 180782
rect 51717 180779 51783 180782
rect 589641 180298 589707 180301
rect 667381 180298 667447 180301
rect 675845 180298 675911 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 667381 180296 675911 180298
rect 667381 180240 667386 180296
rect 667442 180240 675850 180296
rect 675906 180240 675911 180296
rect 667381 180238 675911 180240
rect 589641 180235 589707 180238
rect 667381 180235 667447 180238
rect 675845 180235 675911 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 668158 179618 668164 179620
rect 666694 179558 668164 179618
rect 666694 179550 666754 179558
rect 668158 179556 668164 179558
rect 668228 179556 668234 179620
rect 666356 179490 666754 179550
rect 676213 178938 676279 178941
rect 676213 178936 676322 178938
rect 676213 178880 676218 178936
rect 676274 178880 676322 178936
rect 676213 178875 676322 178880
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 676262 178500 676322 178875
rect 673310 178060 673316 178124
rect 673380 178122 673386 178124
rect 673380 178062 676292 178122
rect 673380 178060 673386 178062
rect 668209 177986 668275 177989
rect 666694 177984 668275 177986
rect 666694 177928 668214 177984
rect 668270 177928 668275 177984
rect 666694 177926 668275 177928
rect 666694 177918 666754 177926
rect 668209 177923 668275 177926
rect 670785 177986 670851 177989
rect 671337 177986 671403 177989
rect 670785 177984 671403 177986
rect 670785 177928 670790 177984
rect 670846 177928 671342 177984
rect 671398 177928 671403 177984
rect 670785 177926 671403 177928
rect 670785 177923 670851 177926
rect 671337 177923 671403 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 675845 177714 675911 177717
rect 675845 177712 676292 177714
rect 675845 177656 675850 177712
rect 675906 177656 676292 177712
rect 675845 177654 676292 177656
rect 675845 177651 675911 177654
rect 673913 177306 673979 177309
rect 673913 177304 676292 177306
rect 673913 177248 673918 177304
rect 673974 177248 676292 177304
rect 673913 177246 676292 177248
rect 673913 177243 673979 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 673361 176898 673427 176901
rect 673361 176896 676292 176898
rect 673361 176840 673366 176896
rect 673422 176840 676292 176896
rect 673361 176838 676292 176840
rect 673361 176835 673427 176838
rect 676806 176608 676812 176672
rect 676876 176608 676882 176672
rect 676814 176460 676874 176608
rect 674741 176082 674807 176085
rect 674741 176080 676292 176082
rect 674741 176024 674746 176080
rect 674802 176024 676292 176080
rect 674741 176022 676292 176024
rect 674741 176019 674807 176022
rect 672441 175674 672507 175677
rect 672441 175672 676292 175674
rect 672441 175616 672446 175672
rect 672502 175616 676292 175672
rect 672441 175614 676292 175616
rect 672441 175611 672507 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 674557 175266 674623 175269
rect 674557 175264 676292 175266
rect 575982 175130 576042 175236
rect 674557 175208 674562 175264
rect 674618 175208 676292 175264
rect 674557 175206 676292 175208
rect 674557 175203 674623 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 666829 174994 666895 174997
rect 666829 174992 669330 174994
rect 666829 174936 666834 174992
rect 666890 174936 669330 174992
rect 666829 174934 669330 174936
rect 666829 174931 666895 174934
rect 669270 174858 669330 174934
rect 669270 174798 676292 174858
rect 668025 174722 668091 174725
rect 666694 174720 668091 174722
rect 666694 174664 668030 174720
rect 668086 174664 668091 174720
rect 666694 174662 668091 174664
rect 666694 174654 666754 174662
rect 668025 174659 668091 174662
rect 666356 174594 666754 174654
rect 673913 174450 673979 174453
rect 673913 174448 676292 174450
rect 673913 174392 673918 174448
rect 673974 174392 676292 174448
rect 673913 174390 676292 174392
rect 673913 174387 673979 174390
rect 674833 174042 674899 174045
rect 674833 174040 676292 174042
rect 674833 173984 674838 174040
rect 674894 173984 676292 174040
rect 674833 173982 676292 173984
rect 674833 173979 674899 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 680997 173634 681063 173637
rect 680997 173632 681076 173634
rect 680997 173576 681002 173632
rect 681058 173576 681076 173632
rect 680997 173574 681076 173576
rect 680997 173571 681063 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 676029 173226 676095 173229
rect 676029 173224 676292 173226
rect 676029 173168 676034 173224
rect 676090 173168 676292 173224
rect 676029 173166 676292 173168
rect 676029 173163 676095 173166
rect 666356 172962 666938 173022
rect 666878 172954 666938 172962
rect 674097 172954 674163 172957
rect 666878 172952 674163 172954
rect 666878 172896 674102 172952
rect 674158 172896 674163 172952
rect 666878 172894 674163 172896
rect 674097 172891 674163 172894
rect 675886 172756 675892 172820
rect 675956 172818 675962 172820
rect 675956 172758 676292 172818
rect 675956 172756 675962 172758
rect 669497 172410 669563 172413
rect 669497 172408 676292 172410
rect 669497 172352 669502 172408
rect 669558 172352 676292 172408
rect 669497 172350 676292 172352
rect 669497 172347 669563 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 671981 172002 672047 172005
rect 671981 172000 676292 172002
rect 671981 171944 671986 172000
rect 672042 171944 676292 172000
rect 671981 171942 676292 171944
rect 671981 171939 672047 171942
rect 682377 171594 682443 171597
rect 682364 171592 682443 171594
rect 682364 171536 682382 171592
rect 682438 171536 682443 171592
rect 682364 171534 682443 171536
rect 682377 171531 682443 171534
rect 670417 171186 670483 171189
rect 670417 171184 676292 171186
rect 670417 171128 670422 171184
rect 670478 171128 676292 171184
rect 670417 171126 676292 171128
rect 670417 171123 670483 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 673729 170778 673795 170781
rect 673729 170776 676292 170778
rect 673729 170720 673734 170776
rect 673790 170720 676292 170776
rect 673729 170718 676292 170720
rect 673729 170715 673795 170718
rect 589641 170506 589707 170509
rect 589641 170504 592572 170506
rect 589641 170448 589646 170504
rect 589702 170448 592572 170504
rect 589641 170446 592572 170448
rect 589641 170443 589707 170446
rect 670601 170370 670667 170373
rect 670601 170368 676292 170370
rect 670601 170312 670606 170368
rect 670662 170312 676292 170368
rect 670601 170310 676292 170312
rect 670601 170307 670667 170310
rect 676581 169962 676647 169965
rect 676581 169960 676660 169962
rect 676581 169904 676586 169960
rect 676642 169904 676660 169960
rect 676581 169902 676660 169904
rect 676581 169899 676647 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 667933 169690 667999 169693
rect 666694 169688 667999 169690
rect 666694 169632 667938 169688
rect 667994 169632 667999 169688
rect 666694 169630 667999 169632
rect 667933 169627 667999 169630
rect 676170 169494 676292 169554
rect 675886 169356 675892 169420
rect 675956 169418 675962 169420
rect 676170 169418 676230 169494
rect 675956 169358 676230 169418
rect 675956 169356 675962 169358
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 672993 169146 673059 169149
rect 672993 169144 676292 169146
rect 672993 169088 672998 169144
rect 673054 169088 676292 169144
rect 672993 169086 676292 169088
rect 672993 169083 673059 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 673085 168738 673151 168741
rect 673085 168736 676292 168738
rect 673085 168680 673090 168736
rect 673146 168680 676292 168736
rect 673085 168678 676292 168680
rect 673085 168675 673151 168678
rect 672349 168330 672415 168333
rect 672349 168328 676292 168330
rect 672349 168272 672354 168328
rect 672410 168272 676292 168328
rect 672349 168270 676292 168272
rect 672349 168267 672415 168270
rect 666356 168066 666754 168126
rect 666694 168058 666754 168066
rect 672165 168058 672231 168061
rect 666694 168056 672231 168058
rect 666694 168000 672170 168056
rect 672226 168000 672231 168056
rect 666694 167998 672231 168000
rect 672165 167995 672231 167998
rect 683113 167922 683179 167925
rect 683100 167920 683179 167922
rect 683100 167864 683118 167920
rect 683174 167864 683179 167920
rect 683100 167862 683179 167864
rect 683113 167859 683179 167862
rect 675334 167452 675340 167516
rect 675404 167514 675410 167516
rect 675661 167514 675727 167517
rect 675404 167512 676292 167514
rect 675404 167456 675666 167512
rect 675722 167456 676292 167512
rect 675404 167454 676292 167456
rect 675404 167452 675410 167454
rect 675661 167451 675727 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 578233 166970 578299 166973
rect 575798 166968 578299 166970
rect 575798 166912 578238 166968
rect 578294 166912 578299 166968
rect 575798 166910 578299 166912
rect 575798 166532 575858 166910
rect 578233 166907 578299 166910
rect 672349 166970 672415 166973
rect 676170 166970 676230 167046
rect 672349 166968 676230 166970
rect 672349 166912 672354 166968
rect 672410 166912 676230 166968
rect 672349 166910 676230 166912
rect 672349 166907 672415 166910
rect 676581 166428 676647 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676581 166363 676647 166364
rect 589457 165610 589523 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 589457 165547 589523 165550
rect 667933 164930 667999 164933
rect 666694 164928 667999 164930
rect 666694 164872 667938 164928
rect 667994 164872 667999 164928
rect 666694 164870 667999 164872
rect 666694 164862 666754 164870
rect 667933 164867 667999 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668761 163298 668827 163301
rect 666694 163296 668827 163298
rect 666694 163240 668766 163296
rect 668822 163240 668827 163296
rect 666694 163238 668827 163240
rect 666694 163230 666754 163238
rect 668761 163235 668827 163238
rect 666356 163170 666754 163230
rect 579337 162754 579403 162757
rect 575798 162752 579403 162754
rect 575798 162696 579342 162752
rect 579398 162696 579403 162752
rect 575798 162694 579403 162696
rect 575798 162180 575858 162694
rect 579337 162691 579403 162694
rect 676070 162692 676076 162756
rect 676140 162754 676146 162756
rect 680997 162754 681063 162757
rect 676140 162752 681063 162754
rect 676140 162696 681002 162752
rect 681058 162696 681063 162752
rect 676140 162694 681063 162696
rect 676140 162692 676146 162694
rect 680997 162691 681063 162694
rect 668761 162482 668827 162485
rect 673453 162482 673519 162485
rect 668761 162480 673519 162482
rect 668761 162424 668766 162480
rect 668822 162424 673458 162480
rect 673514 162424 673519 162480
rect 668761 162422 673519 162424
rect 668761 162419 668827 162422
rect 673453 162419 673519 162422
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 675201 162074 675267 162077
rect 675845 162074 675911 162077
rect 683113 162074 683179 162077
rect 675201 162072 675911 162074
rect 675201 162016 675206 162072
rect 675262 162016 675850 162072
rect 675906 162016 675911 162072
rect 675201 162014 675911 162016
rect 675201 162011 675267 162014
rect 675845 162011 675911 162014
rect 678930 162072 683179 162074
rect 678930 162016 683118 162072
rect 683174 162016 683179 162072
rect 678930 162014 683179 162016
rect 674097 161802 674163 161805
rect 678930 161802 678990 162014
rect 683113 162011 683179 162014
rect 674097 161800 678990 161802
rect 674097 161744 674102 161800
rect 674158 161744 678990 161800
rect 674097 161742 678990 161744
rect 674097 161739 674163 161742
rect 673126 161468 673132 161532
rect 673196 161530 673202 161532
rect 675477 161530 675543 161533
rect 673196 161528 675543 161530
rect 673196 161472 675482 161528
rect 675538 161472 675543 161528
rect 673196 161470 675543 161472
rect 673196 161468 673202 161470
rect 675477 161467 675543 161470
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 668209 160034 668275 160037
rect 666694 160032 668275 160034
rect 575982 159898 576042 160004
rect 666694 159976 668214 160032
rect 668270 159976 668275 160032
rect 666694 159974 668275 159976
rect 666694 159966 666754 159974
rect 668209 159971 668275 159974
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 673729 158810 673795 158813
rect 667982 158808 673795 158810
rect 667982 158752 673734 158808
rect 673790 158752 673795 158808
rect 667982 158750 673795 158752
rect 578417 158402 578483 158405
rect 667982 158402 668042 158750
rect 673729 158747 673795 158750
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666878 158342 668042 158402
rect 666878 158334 666938 158342
rect 666356 158274 666938 158334
rect 589273 157450 589339 157453
rect 589273 157448 592572 157450
rect 589273 157392 589278 157448
rect 589334 157392 592572 157448
rect 589273 157390 592572 157392
rect 589273 157387 589339 157390
rect 675753 157042 675819 157045
rect 676438 157042 676444 157044
rect 675753 157040 676444 157042
rect 675753 156984 675758 157040
rect 675814 156984 676444 157040
rect 675753 156982 676444 156984
rect 675753 156979 675819 156982
rect 676438 156980 676444 156982
rect 676508 156980 676514 157044
rect 673545 156498 673611 156501
rect 675293 156498 675359 156501
rect 673545 156496 675359 156498
rect 673545 156440 673550 156496
rect 673606 156440 675298 156496
rect 675354 156440 675359 156496
rect 673545 156438 675359 156440
rect 673545 156435 673611 156438
rect 675293 156435 675359 156438
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 670417 155954 670483 155957
rect 675109 155954 675175 155957
rect 670417 155952 675175 155954
rect 670417 155896 670422 155952
rect 670478 155896 675114 155952
rect 675170 155896 675175 155952
rect 670417 155894 675175 155896
rect 670417 155891 670483 155894
rect 675109 155891 675175 155894
rect 589457 155818 589523 155821
rect 675753 155818 675819 155821
rect 676254 155818 676260 155820
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 675753 155816 676260 155818
rect 675753 155760 675758 155816
rect 675814 155760 676260 155816
rect 675753 155758 676260 155760
rect 589457 155755 589523 155758
rect 675753 155755 675819 155758
rect 676254 155756 676260 155758
rect 676324 155756 676330 155820
rect 668209 155138 668275 155141
rect 666694 155136 668275 155138
rect 666694 155080 668214 155136
rect 668270 155080 668275 155136
rect 666694 155078 668275 155080
rect 666694 155070 666754 155078
rect 668209 155075 668275 155078
rect 666356 155010 666754 155070
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 154050 578391 154053
rect 575798 154048 578391 154050
rect 575798 153992 578330 154048
rect 578386 153992 578391 154048
rect 575798 153990 578391 153992
rect 575798 153476 575858 153990
rect 578325 153987 578391 153990
rect 666356 153378 666938 153438
rect 666878 153370 666938 153378
rect 666878 153310 673470 153370
rect 673410 153234 673470 153310
rect 674281 153234 674347 153237
rect 673410 153232 674347 153234
rect 673410 153176 674286 153232
rect 674342 153176 674347 153232
rect 673410 153174 674347 153176
rect 674281 153171 674347 153174
rect 673085 152690 673151 152693
rect 675109 152690 675175 152693
rect 673085 152688 675175 152690
rect 673085 152632 673090 152688
rect 673146 152632 675114 152688
rect 675170 152632 675175 152688
rect 673085 152630 675175 152632
rect 673085 152627 673151 152630
rect 675109 152627 675175 152630
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 675753 151466 675819 151469
rect 676622 151466 676628 151468
rect 675753 151464 676628 151466
rect 675753 151408 675758 151464
rect 675814 151408 676628 151464
rect 675753 151406 676628 151408
rect 675753 151403 675819 151406
rect 676622 151404 676628 151406
rect 676692 151404 676698 151468
rect 673177 151330 673243 151333
rect 675109 151330 675175 151333
rect 673177 151328 675175 151330
rect 673177 151272 673182 151328
rect 673238 151272 675114 151328
rect 675170 151272 675175 151328
rect 673177 151270 675175 151272
rect 673177 151267 673243 151270
rect 675109 151267 675175 151270
rect 590009 150922 590075 150925
rect 590009 150920 592572 150922
rect 590009 150864 590014 150920
rect 590070 150864 592572 150920
rect 590009 150862 592572 150864
rect 590009 150859 590075 150862
rect 669589 150378 669655 150381
rect 674925 150378 674991 150381
rect 669589 150376 674991 150378
rect 669589 150320 669594 150376
rect 669650 150320 674930 150376
rect 674986 150320 674991 150376
rect 669589 150318 674991 150320
rect 669589 150315 669655 150318
rect 674925 150315 674991 150318
rect 666356 150114 666754 150174
rect 666694 150106 666754 150114
rect 671705 150106 671771 150109
rect 666694 150104 671771 150106
rect 666694 150048 671710 150104
rect 671766 150048 671771 150104
rect 666694 150046 671771 150048
rect 671705 150043 671771 150046
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 668761 148610 668827 148613
rect 666694 148608 668827 148610
rect 666694 148552 668766 148608
rect 668822 148552 668827 148608
rect 666694 148550 668827 148552
rect 666694 148542 666754 148550
rect 668761 148547 668827 148550
rect 666356 148482 666754 148542
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 588537 147658 588603 147661
rect 670601 147658 670667 147661
rect 675109 147658 675175 147661
rect 675385 147660 675451 147661
rect 588537 147656 592572 147658
rect 588537 147600 588542 147656
rect 588598 147600 592572 147656
rect 588537 147598 592572 147600
rect 670601 147656 675175 147658
rect 670601 147600 670606 147656
rect 670662 147600 675114 147656
rect 675170 147600 675175 147656
rect 670601 147598 675175 147600
rect 588537 147595 588603 147598
rect 670601 147595 670667 147598
rect 675109 147595 675175 147598
rect 675334 147596 675340 147660
rect 675404 147658 675451 147660
rect 675404 147656 675496 147658
rect 675446 147600 675496 147656
rect 675404 147598 675496 147600
rect 675404 147596 675451 147598
rect 675385 147595 675451 147596
rect 579521 147522 579587 147525
rect 575798 147520 579587 147522
rect 575798 147464 579526 147520
rect 579582 147464 579587 147520
rect 575798 147462 579587 147464
rect 575798 146948 575858 147462
rect 579521 147459 579587 147462
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 668761 145346 668827 145349
rect 666694 145344 668827 145346
rect 666694 145288 668766 145344
rect 668822 145288 668827 145344
rect 666694 145286 668827 145288
rect 666694 145278 666754 145286
rect 668761 145283 668827 145286
rect 666356 145218 666754 145278
rect 671981 144938 672047 144941
rect 675109 144938 675175 144941
rect 671981 144936 675175 144938
rect 671981 144880 671986 144936
rect 672042 144880 675114 144936
rect 675170 144880 675175 144936
rect 671981 144878 675175 144880
rect 671981 144875 672047 144878
rect 675109 144875 675175 144878
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 669129 143714 669195 143717
rect 666694 143712 669195 143714
rect 666694 143656 669134 143712
rect 669190 143656 669195 143712
rect 666694 143654 669195 143656
rect 666694 143646 666754 143654
rect 669129 143651 669195 143654
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589825 142762 589891 142765
rect 589825 142760 592572 142762
rect 589825 142704 589830 142760
rect 589886 142704 592572 142760
rect 589825 142702 592572 142704
rect 589825 142699 589891 142702
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 669262 140450 669268 140452
rect 666694 140390 669268 140450
rect 666694 140382 666754 140390
rect 669262 140388 669268 140390
rect 669332 140388 669338 140452
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 668577 138818 668643 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 668643 138818
rect 666694 138760 668582 138816
rect 668638 138760 668643 138816
rect 666694 138758 668643 138760
rect 666694 138750 666754 138758
rect 668577 138755 668643 138758
rect 666356 138690 666754 138750
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 668393 135554 668459 135557
rect 666694 135552 668459 135554
rect 666694 135496 668398 135552
rect 668454 135496 668459 135552
rect 666694 135494 668459 135496
rect 666694 135486 666754 135494
rect 668393 135491 668459 135494
rect 666356 135426 666754 135486
rect 668761 135146 668827 135149
rect 672165 135146 672231 135149
rect 668761 135144 672231 135146
rect 668761 135088 668766 135144
rect 668822 135088 672170 135144
rect 672226 135088 672231 135144
rect 668761 135086 672231 135088
rect 668761 135083 668827 135086
rect 672165 135083 672231 135086
rect 590377 134602 590443 134605
rect 590377 134600 592572 134602
rect 590377 134544 590382 134600
rect 590438 134544 592572 134600
rect 590377 134542 592572 134544
rect 590377 134539 590443 134542
rect 667790 134540 667796 134604
rect 667860 134602 667866 134604
rect 675845 134602 675911 134605
rect 667860 134600 675911 134602
rect 667860 134544 675850 134600
rect 675906 134544 675911 134600
rect 667860 134542 675911 134544
rect 667860 134540 667866 134542
rect 675845 134539 675911 134542
rect 579521 134466 579587 134469
rect 575798 134464 579587 134466
rect 575798 134408 579526 134464
rect 579582 134408 579587 134464
rect 575798 134406 579587 134408
rect 575798 133892 575858 134406
rect 579521 134403 579587 134406
rect 666356 133794 666754 133854
rect 666694 133786 666754 133794
rect 667933 133786 667999 133789
rect 666694 133784 667999 133786
rect 666694 133728 667938 133784
rect 667994 133728 667999 133784
rect 666694 133726 667999 133728
rect 667933 133723 667999 133726
rect 667749 133106 667815 133109
rect 676262 133106 676322 133348
rect 676489 133106 676555 133109
rect 667749 133104 676322 133106
rect 667749 133048 667754 133104
rect 667810 133048 676322 133104
rect 667749 133046 676322 133048
rect 676446 133104 676555 133106
rect 676446 133048 676494 133104
rect 676550 133048 676555 133104
rect 667749 133043 667815 133046
rect 676446 133043 676555 133048
rect 589457 132970 589523 132973
rect 589457 132968 592572 132970
rect 589457 132912 589462 132968
rect 589518 132912 592572 132968
rect 676446 132940 676506 133043
rect 589457 132910 592572 132912
rect 589457 132907 589523 132910
rect 667197 132562 667263 132565
rect 667197 132560 676292 132562
rect 667197 132504 667202 132560
rect 667258 132504 676292 132560
rect 667197 132502 676292 132504
rect 667197 132499 667263 132502
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 673361 132154 673427 132157
rect 673361 132152 676292 132154
rect 673361 132096 673366 132152
rect 673422 132096 676292 132152
rect 673361 132094 676292 132096
rect 673361 132091 673427 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 589457 131338 589523 131341
rect 674649 131338 674715 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 589457 131278 592572 131280
rect 674649 131336 676292 131338
rect 674649 131280 674654 131336
rect 674710 131280 676292 131336
rect 674649 131278 676292 131280
rect 589457 131275 589523 131278
rect 674649 131275 674715 131278
rect 669957 130930 670023 130933
rect 669957 130928 676292 130930
rect 669957 130872 669962 130928
rect 670018 130872 676292 130928
rect 669957 130870 676292 130872
rect 669957 130867 670023 130870
rect 668485 130658 668551 130661
rect 666694 130656 668551 130658
rect 666694 130600 668490 130656
rect 668546 130600 668551 130656
rect 666694 130598 668551 130600
rect 666694 130590 666754 130598
rect 668485 130595 668551 130598
rect 666356 130530 666754 130590
rect 674465 130522 674531 130525
rect 674465 130520 676292 130522
rect 674465 130464 674470 130520
rect 674526 130464 676292 130520
rect 674465 130462 676292 130464
rect 674465 130459 674531 130462
rect 676213 130250 676279 130253
rect 676213 130248 676322 130250
rect 676213 130192 676218 130248
rect 676274 130192 676322 130248
rect 676213 130187 676322 130192
rect 676262 130084 676322 130187
rect 578877 129706 578943 129709
rect 575798 129704 578943 129706
rect 575798 129648 578882 129704
rect 578938 129648 578943 129704
rect 575798 129646 578943 129648
rect 575798 129540 575858 129646
rect 578877 129643 578943 129646
rect 588537 129706 588603 129709
rect 673913 129706 673979 129709
rect 588537 129704 592572 129706
rect 588537 129648 588542 129704
rect 588598 129648 592572 129704
rect 588537 129646 592572 129648
rect 673913 129704 676292 129706
rect 673913 129648 673918 129704
rect 673974 129648 676292 129704
rect 673913 129646 676292 129648
rect 588537 129643 588603 129646
rect 673913 129643 673979 129646
rect 671521 129298 671587 129301
rect 671521 129296 676292 129298
rect 671521 129240 671526 129296
rect 671582 129240 676292 129296
rect 671521 129238 676292 129240
rect 671521 129235 671587 129238
rect 668025 129026 668091 129029
rect 666694 129024 668091 129026
rect 666694 128968 668030 129024
rect 668086 128968 668091 129024
rect 666694 128966 668091 128968
rect 666694 128958 666754 128966
rect 668025 128963 668091 128966
rect 666356 128898 666754 128958
rect 675017 128890 675083 128893
rect 675017 128888 676292 128890
rect 675017 128832 675022 128888
rect 675078 128832 676292 128888
rect 675017 128830 676292 128832
rect 675017 128827 675083 128830
rect 674373 128482 674439 128485
rect 674373 128480 676292 128482
rect 674373 128424 674378 128480
rect 674434 128424 676292 128480
rect 674373 128422 676292 128424
rect 674373 128419 674439 128422
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 579521 127938 579587 127941
rect 575798 127936 579587 127938
rect 575798 127880 579526 127936
rect 579582 127880 579587 127936
rect 575798 127878 579587 127880
rect 575798 127364 575858 127878
rect 579521 127875 579587 127878
rect 676446 127805 676506 128044
rect 668577 127802 668643 127805
rect 676213 127802 676279 127805
rect 668577 127800 676279 127802
rect 668577 127744 668582 127800
rect 668638 127744 676218 127800
rect 676274 127744 676279 127800
rect 668577 127742 676279 127744
rect 668577 127739 668643 127742
rect 676213 127739 676279 127742
rect 676397 127800 676506 127805
rect 676397 127744 676402 127800
rect 676458 127744 676506 127800
rect 676397 127742 676506 127744
rect 676397 127739 676463 127742
rect 676814 127396 676874 127636
rect 676806 127332 676812 127396
rect 676876 127332 676882 127396
rect 676070 126924 676076 126988
rect 676140 126986 676146 126988
rect 676262 126986 676322 127228
rect 676140 126926 676322 126986
rect 676140 126924 676146 126926
rect 673361 126578 673427 126581
rect 676262 126578 676322 126820
rect 673361 126576 676322 126578
rect 673361 126520 673366 126576
rect 673422 126520 676322 126576
rect 673361 126518 676322 126520
rect 673361 126515 673427 126518
rect 589917 126442 589983 126445
rect 589917 126440 592572 126442
rect 589917 126384 589922 126440
rect 589978 126384 592572 126440
rect 589917 126382 592572 126384
rect 589917 126379 589983 126382
rect 679574 126173 679634 126412
rect 679574 126168 679683 126173
rect 679574 126112 679622 126168
rect 679678 126112 679683 126168
rect 679574 126110 679683 126112
rect 679617 126107 679683 126110
rect 668945 125762 669011 125765
rect 676262 125764 676322 126004
rect 666694 125760 669011 125762
rect 666694 125704 668950 125760
rect 669006 125704 669011 125760
rect 666694 125702 669011 125704
rect 666694 125694 666754 125702
rect 668945 125699 669011 125702
rect 676254 125700 676260 125764
rect 676324 125700 676330 125764
rect 666356 125634 666754 125694
rect 682334 125357 682394 125596
rect 578325 125354 578391 125357
rect 575798 125352 578391 125354
rect 575798 125296 578330 125352
rect 578386 125296 578391 125352
rect 575798 125294 578391 125296
rect 682334 125352 682443 125357
rect 682334 125296 682382 125352
rect 682438 125296 682443 125352
rect 682334 125294 682443 125296
rect 575798 125188 575858 125294
rect 578325 125291 578391 125294
rect 682377 125291 682443 125294
rect 673177 124946 673243 124949
rect 676262 124946 676322 125188
rect 673177 124944 676322 124946
rect 673177 124888 673182 124944
rect 673238 124888 676322 124944
rect 673177 124886 676322 124888
rect 673177 124883 673243 124886
rect 589457 124810 589523 124813
rect 589457 124808 592572 124810
rect 589457 124752 589462 124808
rect 589518 124752 592572 124808
rect 589457 124750 592572 124752
rect 589457 124747 589523 124750
rect 673913 124538 673979 124541
rect 676262 124538 676322 124780
rect 673913 124536 676322 124538
rect 673913 124480 673918 124536
rect 673974 124480 676322 124536
rect 673913 124478 676322 124480
rect 673913 124475 673979 124478
rect 672809 124130 672875 124133
rect 666694 124128 672875 124130
rect 666694 124072 672814 124128
rect 672870 124072 672875 124128
rect 666694 124070 672875 124072
rect 666694 124062 666754 124070
rect 672809 124067 672875 124070
rect 674649 124130 674715 124133
rect 676630 124132 676690 124372
rect 676438 124130 676444 124132
rect 674649 124128 676444 124130
rect 674649 124072 674654 124128
rect 674710 124072 676444 124128
rect 674649 124070 676444 124072
rect 674649 124067 674715 124070
rect 676438 124068 676444 124070
rect 676508 124068 676514 124132
rect 676622 124068 676628 124132
rect 676692 124068 676698 124132
rect 666356 124002 666754 124062
rect 674833 123722 674899 123725
rect 676262 123722 676322 123964
rect 674833 123720 676322 123722
rect 674833 123664 674838 123720
rect 674894 123664 676322 123720
rect 674833 123662 676322 123664
rect 674833 123659 674899 123662
rect 676438 123660 676444 123724
rect 676508 123660 676514 123724
rect 578417 123586 578483 123589
rect 575798 123584 578483 123586
rect 575798 123528 578422 123584
rect 578478 123528 578483 123584
rect 676446 123556 676506 123660
rect 575798 123526 578483 123528
rect 575798 123012 575858 123526
rect 578417 123523 578483 123526
rect 672073 123314 672139 123317
rect 672073 123312 676322 123314
rect 672073 123256 672078 123312
rect 672134 123256 676322 123312
rect 672073 123254 676322 123256
rect 672073 123251 672139 123254
rect 589457 123178 589523 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 676262 123148 676322 123254
rect 589457 123118 592572 123120
rect 589457 123115 589523 123118
rect 673085 123042 673151 123045
rect 674833 123042 674899 123045
rect 673085 123040 674899 123042
rect 673085 122984 673090 123040
rect 673146 122984 674838 123040
rect 674894 122984 674899 123040
rect 673085 122982 674899 122984
rect 673085 122979 673151 122982
rect 674833 122979 674899 122982
rect 676254 122844 676260 122908
rect 676324 122906 676330 122908
rect 676806 122906 676812 122908
rect 676324 122846 676812 122906
rect 676324 122844 676330 122846
rect 676806 122844 676812 122846
rect 676876 122844 676882 122908
rect 670601 122498 670667 122501
rect 676262 122498 676322 122740
rect 670601 122496 676322 122498
rect 670601 122440 670606 122496
rect 670662 122440 676322 122496
rect 670601 122438 676322 122440
rect 670601 122435 670667 122438
rect 675334 122028 675340 122092
rect 675404 122090 675410 122092
rect 676262 122090 676322 122332
rect 675404 122030 676322 122090
rect 675404 122028 675410 122030
rect 676262 121682 676322 121924
rect 676032 121622 676322 121682
rect 590009 121546 590075 121549
rect 590009 121544 592572 121546
rect 590009 121488 590014 121544
rect 590070 121488 592572 121544
rect 590009 121486 592572 121488
rect 590009 121483 590075 121486
rect 578877 121410 578943 121413
rect 575798 121408 578943 121410
rect 575798 121352 578882 121408
rect 578938 121352 578943 121408
rect 575798 121350 578943 121352
rect 575798 120836 575858 121350
rect 578877 121347 578943 121350
rect 672625 120866 672691 120869
rect 666694 120864 672691 120866
rect 666694 120808 672630 120864
rect 672686 120808 672691 120864
rect 666694 120806 672691 120808
rect 666694 120798 666754 120806
rect 672625 120803 672691 120806
rect 666356 120738 666754 120798
rect 672901 120730 672967 120733
rect 676032 120730 676092 121622
rect 672901 120728 676092 120730
rect 672901 120672 672906 120728
rect 672962 120672 676092 120728
rect 672901 120670 676092 120672
rect 672901 120667 672967 120670
rect 589641 119914 589707 119917
rect 589641 119912 592572 119914
rect 589641 119856 589646 119912
rect 589702 119856 592572 119912
rect 589641 119854 592572 119856
rect 589641 119851 589707 119854
rect 668761 119234 668827 119237
rect 666694 119232 668827 119234
rect 666694 119176 668766 119232
rect 668822 119176 668827 119232
rect 666694 119174 668827 119176
rect 666694 119166 666754 119174
rect 668761 119171 668827 119174
rect 666356 119106 666754 119166
rect 668945 118826 669011 118829
rect 672073 118826 672139 118829
rect 668945 118824 672139 118826
rect 668945 118768 668950 118824
rect 669006 118768 672078 118824
rect 672134 118768 672139 118824
rect 668945 118766 672139 118768
rect 668945 118763 669011 118766
rect 672073 118763 672139 118766
rect 575982 118418 576042 118660
rect 578509 118418 578575 118421
rect 575982 118416 578575 118418
rect 575982 118360 578514 118416
rect 578570 118360 578575 118416
rect 575982 118358 578575 118360
rect 578509 118355 578575 118358
rect 590101 118282 590167 118285
rect 590101 118280 592572 118282
rect 590101 118224 590106 118280
rect 590162 118224 592572 118280
rect 590101 118222 592572 118224
rect 590101 118219 590167 118222
rect 666356 117474 666938 117534
rect 666878 117466 666938 117474
rect 674097 117466 674163 117469
rect 666878 117464 674163 117466
rect 666878 117408 674102 117464
rect 674158 117408 674163 117464
rect 666878 117406 674163 117408
rect 674097 117403 674163 117406
rect 675702 117268 675708 117332
rect 675772 117330 675778 117332
rect 682377 117330 682443 117333
rect 675772 117328 682443 117330
rect 675772 117272 682382 117328
rect 682438 117272 682443 117328
rect 675772 117270 682443 117272
rect 675772 117268 675778 117270
rect 682377 117267 682443 117270
rect 675201 117058 675267 117061
rect 675845 117058 675911 117061
rect 675201 117056 675911 117058
rect 675201 117000 675206 117056
rect 675262 117000 675850 117056
rect 675906 117000 675911 117056
rect 675201 116998 675911 117000
rect 675201 116995 675267 116998
rect 675845 116995 675911 116998
rect 579521 116922 579587 116925
rect 575798 116920 579587 116922
rect 575798 116864 579526 116920
rect 579582 116864 579587 116920
rect 575798 116862 579587 116864
rect 575798 116484 575858 116862
rect 579521 116859 579587 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 672349 115834 672415 115837
rect 666694 115832 672415 115834
rect 666694 115776 672354 115832
rect 672410 115776 672415 115832
rect 666694 115774 672415 115776
rect 672349 115771 672415 115774
rect 674046 115772 674052 115836
rect 674116 115834 674122 115836
rect 675477 115834 675543 115837
rect 674116 115832 675543 115834
rect 674116 115776 675482 115832
rect 675538 115776 675543 115832
rect 674116 115774 675543 115776
rect 674116 115772 674122 115774
rect 675477 115771 675543 115774
rect 590285 115018 590351 115021
rect 590285 115016 592572 115018
rect 590285 114960 590290 115016
rect 590346 114960 592572 115016
rect 590285 114958 592572 114960
rect 590285 114955 590351 114958
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 668945 114338 669011 114341
rect 666694 114336 669011 114338
rect 666694 114280 668950 114336
rect 669006 114280 669011 114336
rect 666694 114278 669011 114280
rect 666694 114270 666754 114278
rect 668945 114275 669011 114278
rect 666356 114210 666754 114270
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 668761 112706 668827 112709
rect 666694 112704 668827 112706
rect 666694 112648 668766 112704
rect 668822 112648 668827 112704
rect 666694 112646 668827 112648
rect 666694 112638 666754 112646
rect 668761 112643 668827 112646
rect 666356 112578 666754 112638
rect 579521 112570 579587 112573
rect 575798 112568 579587 112570
rect 575798 112512 579526 112568
rect 579582 112512 579587 112568
rect 575798 112510 579587 112512
rect 575798 112132 575858 112510
rect 579521 112507 579587 112510
rect 675753 112434 675819 112437
rect 676254 112434 676260 112436
rect 675753 112432 676260 112434
rect 675753 112376 675758 112432
rect 675814 112376 676260 112432
rect 675753 112374 676260 112376
rect 675753 112371 675819 112374
rect 676254 112372 676260 112374
rect 676324 112372 676330 112436
rect 589457 111754 589523 111757
rect 675753 111754 675819 111757
rect 676438 111754 676444 111756
rect 589457 111752 592572 111754
rect 589457 111696 589462 111752
rect 589518 111696 592572 111752
rect 589457 111694 592572 111696
rect 675753 111752 676444 111754
rect 675753 111696 675758 111752
rect 675814 111696 676444 111752
rect 675753 111694 676444 111696
rect 589457 111691 589523 111694
rect 675753 111691 675819 111694
rect 676438 111692 676444 111694
rect 676508 111692 676514 111756
rect 675753 111348 675819 111349
rect 675702 111284 675708 111348
rect 675772 111346 675819 111348
rect 675772 111344 675864 111346
rect 675814 111288 675864 111344
rect 675772 111286 675864 111288
rect 675772 111284 675819 111286
rect 675753 111283 675819 111284
rect 672901 111074 672967 111077
rect 666694 111072 672967 111074
rect 666694 111016 672906 111072
rect 672962 111016 672967 111072
rect 666694 111014 672967 111016
rect 666694 111006 666754 111014
rect 672901 111011 672967 111014
rect 666356 110946 666754 111006
rect 675753 110394 675819 110397
rect 676622 110394 676628 110396
rect 675753 110392 676628 110394
rect 675753 110336 675758 110392
rect 675814 110336 676628 110392
rect 675753 110334 676628 110336
rect 675753 110331 675819 110334
rect 676622 110332 676628 110334
rect 676692 110332 676698 110396
rect 579337 110122 579403 110125
rect 575798 110120 579403 110122
rect 575798 110064 579342 110120
rect 579398 110064 579403 110120
rect 575798 110062 579403 110064
rect 575798 109956 575858 110062
rect 579337 110059 579403 110062
rect 589273 110122 589339 110125
rect 589273 110120 592572 110122
rect 589273 110064 589278 110120
rect 589334 110064 592572 110120
rect 589273 110062 592572 110064
rect 589273 110059 589339 110062
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675753 108218 675819 108221
rect 676070 108218 676076 108220
rect 675753 108216 676076 108218
rect 675753 108160 675758 108216
rect 675814 108160 676076 108216
rect 675753 108158 676076 108160
rect 675753 108155 675819 108158
rect 676070 108156 676076 108158
rect 676140 108156 676146 108220
rect 667933 107810 667999 107813
rect 666694 107808 667999 107810
rect 666694 107752 667938 107808
rect 667994 107752 667999 107808
rect 666694 107750 667999 107752
rect 666694 107742 666754 107750
rect 667933 107747 667999 107750
rect 666356 107682 666754 107742
rect 673913 106994 673979 106997
rect 675385 106994 675451 106997
rect 673913 106992 675451 106994
rect 673913 106936 673918 106992
rect 673974 106936 675390 106992
rect 675446 106936 675451 106992
rect 673913 106934 675451 106936
rect 673913 106931 673979 106934
rect 675385 106931 675451 106934
rect 589825 106858 589891 106861
rect 589825 106856 592572 106858
rect 589825 106800 589830 106856
rect 589886 106800 592572 106856
rect 589825 106798 592572 106800
rect 589825 106795 589891 106798
rect 668393 106178 668459 106181
rect 666694 106176 668459 106178
rect 666694 106120 668398 106176
rect 668454 106120 668459 106176
rect 666694 106118 668459 106120
rect 666694 106110 666754 106118
rect 668393 106115 668459 106118
rect 672993 106178 673059 106181
rect 675109 106178 675175 106181
rect 672993 106176 675175 106178
rect 672993 106120 672998 106176
rect 673054 106120 675114 106176
rect 675170 106120 675175 106176
rect 672993 106118 675175 106120
rect 672993 106115 673059 106118
rect 675109 106115 675175 106118
rect 666356 106050 666754 106110
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 673177 104682 673243 104685
rect 675109 104682 675175 104685
rect 673177 104680 675175 104682
rect 673177 104624 673182 104680
rect 673238 104624 675114 104680
rect 675170 104624 675175 104680
rect 673177 104622 675175 104624
rect 673177 104619 673243 104622
rect 675109 104619 675175 104622
rect 668761 104546 668827 104549
rect 666694 104544 668827 104546
rect 666694 104488 668766 104544
rect 668822 104488 668827 104544
rect 666694 104486 668827 104488
rect 666694 104478 666754 104486
rect 668761 104483 668827 104486
rect 666356 104418 666754 104478
rect 588721 103594 588787 103597
rect 588721 103592 592572 103594
rect 588721 103536 588726 103592
rect 588782 103536 592572 103592
rect 588721 103534 592572 103536
rect 588721 103531 588787 103534
rect 575982 103322 576042 103428
rect 579521 103322 579587 103325
rect 575982 103320 579587 103322
rect 575982 103264 579526 103320
rect 579582 103264 579587 103320
rect 575982 103262 579587 103264
rect 579521 103259 579587 103262
rect 668577 102914 668643 102917
rect 666694 102912 668643 102914
rect 666694 102856 668582 102912
rect 668638 102856 668643 102912
rect 666694 102854 668643 102856
rect 666694 102846 666754 102854
rect 668577 102851 668643 102854
rect 666356 102786 666754 102846
rect 589457 101962 589523 101965
rect 675385 101964 675451 101965
rect 675334 101962 675340 101964
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 673410 101902 675340 101962
rect 675404 101962 675451 101964
rect 675404 101960 675496 101962
rect 675446 101904 675496 101960
rect 589457 101899 589523 101902
rect 673410 101826 673470 101902
rect 675334 101900 675340 101902
rect 675404 101902 675496 101904
rect 675404 101900 675451 101902
rect 675385 101899 675451 101900
rect 596130 101766 673470 101826
rect 579521 101690 579587 101693
rect 575798 101688 579587 101690
rect 575798 101632 579526 101688
rect 579582 101632 579587 101688
rect 575798 101630 579587 101632
rect 575798 101252 575858 101630
rect 579521 101627 579587 101630
rect 591481 101690 591547 101693
rect 596130 101690 596190 101766
rect 591481 101688 596190 101690
rect 591481 101632 591486 101688
rect 591542 101632 596190 101688
rect 591481 101630 596190 101632
rect 591481 101627 591547 101630
rect 673361 101010 673427 101013
rect 675109 101010 675175 101013
rect 673361 101008 675175 101010
rect 673361 100952 673366 101008
rect 673422 100952 675114 101008
rect 675170 100952 675175 101008
rect 673361 100950 675175 100952
rect 673361 100947 673427 100950
rect 675109 100947 675175 100950
rect 578601 99242 578667 99245
rect 575798 99240 578667 99242
rect 575798 99184 578606 99240
rect 578662 99184 578667 99240
rect 575798 99182 578667 99184
rect 575798 99076 575858 99182
rect 578601 99179 578667 99182
rect 578325 97474 578391 97477
rect 575798 97472 578391 97474
rect 575798 97416 578330 97472
rect 578386 97416 578391 97472
rect 575798 97414 578391 97416
rect 575798 96900 575858 97414
rect 578325 97411 578391 97414
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 641989 96522 642055 96525
rect 647182 96522 647188 96524
rect 641989 96520 647188 96522
rect 641989 96464 641994 96520
rect 642050 96464 647188 96520
rect 641989 96462 647188 96464
rect 641989 96459 642055 96462
rect 647182 96460 647188 96462
rect 647252 96460 647258 96524
rect 633934 95372 633940 95436
rect 634004 95434 634010 95436
rect 635733 95434 635799 95437
rect 634004 95432 635799 95434
rect 634004 95376 635738 95432
rect 635794 95376 635799 95432
rect 634004 95374 635799 95376
rect 634004 95372 634010 95374
rect 635733 95371 635799 95374
rect 579521 95026 579587 95029
rect 575798 95024 579587 95026
rect 575798 94968 579526 95024
rect 579582 94968 579587 95024
rect 575798 94966 579587 94968
rect 575798 94724 575858 94966
rect 579521 94963 579587 94966
rect 647141 95026 647207 95029
rect 647141 95024 647434 95026
rect 647141 94968 647146 95024
rect 647202 94968 647434 95024
rect 647141 94966 647434 94968
rect 647141 94963 647207 94966
rect 626441 94482 626507 94485
rect 626441 94480 628268 94482
rect 626441 94424 626446 94480
rect 626502 94424 628268 94480
rect 647374 94452 647434 94966
rect 626441 94422 628268 94424
rect 626441 94419 626507 94422
rect 655237 94210 655303 94213
rect 655237 94208 656788 94210
rect 655237 94152 655242 94208
rect 655298 94152 656788 94208
rect 655237 94150 656788 94152
rect 655237 94147 655303 94150
rect 625613 93666 625679 93669
rect 625613 93664 628268 93666
rect 625613 93608 625618 93664
rect 625674 93608 628268 93664
rect 625613 93606 628268 93608
rect 625613 93603 625679 93606
rect 655421 93394 655487 93397
rect 665173 93394 665239 93397
rect 655421 93392 656788 93394
rect 655421 93336 655426 93392
rect 655482 93336 656788 93392
rect 655421 93334 656788 93336
rect 663596 93392 665239 93394
rect 663596 93336 665178 93392
rect 665234 93336 665239 93392
rect 663596 93334 665239 93336
rect 655421 93331 655487 93334
rect 665173 93331 665239 93334
rect 578509 93122 578575 93125
rect 575798 93120 578575 93122
rect 575798 93064 578514 93120
rect 578570 93064 578575 93120
rect 575798 93062 578575 93064
rect 575798 92548 575858 93062
rect 578509 93059 578575 93062
rect 650310 93060 650316 93124
rect 650380 93122 650386 93124
rect 650380 93062 656818 93122
rect 650380 93060 650386 93062
rect 626441 92850 626507 92853
rect 626441 92848 628268 92850
rect 626441 92792 626446 92848
rect 626502 92792 628268 92848
rect 626441 92790 628268 92792
rect 626441 92787 626507 92790
rect 656758 92548 656818 93062
rect 663701 92850 663767 92853
rect 663382 92848 663767 92850
rect 663382 92792 663706 92848
rect 663762 92792 663767 92848
rect 663382 92790 663767 92792
rect 663382 92548 663442 92790
rect 663701 92787 663767 92790
rect 647509 92442 647575 92445
rect 647509 92440 647618 92442
rect 647509 92384 647514 92440
rect 647570 92384 647618 92440
rect 647509 92379 647618 92384
rect 625797 92034 625863 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 647558 92004 647618 92379
rect 625797 91974 628268 91976
rect 625797 91971 625863 91974
rect 665357 91762 665423 91765
rect 663596 91760 665423 91762
rect 663596 91704 665362 91760
rect 665418 91704 665423 91760
rect 663596 91702 665423 91704
rect 665357 91699 665423 91702
rect 654317 91490 654383 91493
rect 654317 91488 656788 91490
rect 654317 91432 654322 91488
rect 654378 91432 656788 91488
rect 654317 91430 656788 91432
rect 654317 91427 654383 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 579061 90946 579127 90949
rect 575798 90944 579127 90946
rect 575798 90888 579066 90944
rect 579122 90888 579127 90944
rect 575798 90886 579127 90888
rect 575798 90372 575858 90886
rect 579061 90883 579127 90886
rect 655421 90674 655487 90677
rect 665541 90674 665607 90677
rect 655421 90672 656788 90674
rect 655421 90616 655426 90672
rect 655482 90616 656788 90672
rect 655421 90614 656788 90616
rect 663596 90672 665607 90674
rect 663596 90616 665546 90672
rect 665602 90616 665607 90672
rect 663596 90614 665607 90616
rect 655421 90611 655487 90614
rect 665541 90611 665607 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 655789 89858 655855 89861
rect 664161 89858 664227 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664227 89858
rect 663596 89800 664166 89856
rect 664222 89800 664227 89856
rect 663596 89798 664227 89800
rect 655789 89795 655855 89798
rect 664161 89795 664227 89798
rect 625245 89586 625311 89589
rect 648245 89586 648311 89589
rect 625245 89584 628268 89586
rect 625245 89528 625250 89584
rect 625306 89528 628268 89584
rect 625245 89526 628268 89528
rect 648140 89584 648311 89586
rect 648140 89528 648250 89584
rect 648306 89528 648311 89584
rect 648140 89526 648311 89528
rect 625245 89523 625311 89526
rect 648245 89523 648311 89526
rect 664345 89042 664411 89045
rect 663596 89040 664411 89042
rect 663596 88984 664350 89040
rect 664406 88984 664411 89040
rect 663596 88982 664411 88984
rect 664345 88979 664411 88982
rect 624969 88770 625035 88773
rect 624969 88768 628268 88770
rect 624969 88712 624974 88768
rect 625030 88712 628268 88768
rect 624969 88710 628268 88712
rect 624969 88707 625035 88710
rect 575982 88090 576042 88196
rect 579521 88090 579587 88093
rect 575982 88088 579587 88090
rect 575982 88032 579526 88088
rect 579582 88032 579587 88088
rect 575982 88030 579587 88032
rect 579521 88027 579587 88030
rect 625153 87954 625219 87957
rect 625153 87952 628268 87954
rect 625153 87896 625158 87952
rect 625214 87896 628268 87952
rect 625153 87894 628268 87896
rect 625153 87891 625219 87894
rect 625337 87138 625403 87141
rect 649993 87138 650059 87141
rect 625337 87136 628268 87138
rect 625337 87080 625342 87136
rect 625398 87080 628268 87136
rect 625337 87078 628268 87080
rect 648140 87136 650059 87138
rect 648140 87080 649998 87136
rect 650054 87080 650059 87136
rect 648140 87078 650059 87080
rect 625337 87075 625403 87078
rect 649993 87075 650059 87078
rect 579337 86458 579403 86461
rect 575798 86456 579403 86458
rect 575798 86400 579342 86456
rect 579398 86400 579403 86456
rect 575798 86398 579403 86400
rect 575798 86020 575858 86398
rect 579337 86395 579403 86398
rect 625153 86322 625219 86325
rect 625153 86320 628268 86322
rect 625153 86264 625158 86320
rect 625214 86264 628268 86320
rect 625153 86262 628268 86264
rect 625153 86259 625219 86262
rect 625153 85506 625219 85509
rect 625153 85504 628268 85506
rect 625153 85448 625158 85504
rect 625214 85448 628268 85504
rect 625153 85446 628268 85448
rect 625153 85443 625219 85446
rect 625337 84690 625403 84693
rect 650545 84690 650611 84693
rect 625337 84688 628268 84690
rect 625337 84632 625342 84688
rect 625398 84632 628268 84688
rect 625337 84630 628268 84632
rect 648140 84688 650611 84690
rect 648140 84632 650550 84688
rect 650606 84632 650611 84688
rect 648140 84630 650611 84632
rect 625337 84627 625403 84630
rect 650545 84627 650611 84630
rect 579153 84010 579219 84013
rect 575798 84008 579219 84010
rect 575798 83952 579158 84008
rect 579214 83952 579219 84008
rect 575798 83950 579219 83952
rect 575798 83844 575858 83950
rect 579153 83947 579219 83950
rect 625153 83874 625219 83877
rect 625153 83872 628268 83874
rect 625153 83816 625158 83872
rect 625214 83816 628268 83872
rect 625153 83814 628268 83816
rect 625153 83811 625219 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 579061 82242 579127 82245
rect 650361 82242 650427 82245
rect 575798 82240 579127 82242
rect 575798 82184 579066 82240
rect 579122 82184 579127 82240
rect 648140 82240 650427 82242
rect 575798 82182 579127 82184
rect 575798 81668 575858 82182
rect 579061 82179 579127 82182
rect 628790 81698 628850 82212
rect 648140 82184 650366 82240
rect 650422 82184 650427 82240
rect 648140 82182 650427 82184
rect 650361 82179 650427 82182
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 578877 80066 578943 80069
rect 575798 80064 578943 80066
rect 575798 80008 578882 80064
rect 578938 80008 578943 80064
rect 575798 80006 578943 80008
rect 575798 79492 575858 80006
rect 578877 80003 578943 80006
rect 633893 78572 633959 78573
rect 633893 78570 633940 78572
rect 633848 78568 633940 78570
rect 633848 78512 633898 78568
rect 633848 78510 633940 78512
rect 633893 78508 633940 78510
rect 634004 78508 634010 78572
rect 633893 78507 633959 78508
rect 637062 78162 637068 78164
rect 625110 78102 637068 78162
rect 579521 77890 579587 77893
rect 575798 77888 579587 77890
rect 575798 77832 579526 77888
rect 579582 77832 579587 77888
rect 575798 77830 579587 77832
rect 575798 77316 575858 77830
rect 579521 77827 579587 77830
rect 581637 77890 581703 77893
rect 625110 77890 625170 78102
rect 637062 78100 637068 78102
rect 637132 78162 637138 78164
rect 639597 78162 639663 78165
rect 637132 78160 639663 78162
rect 637132 78104 639602 78160
rect 639658 78104 639663 78160
rect 637132 78102 639663 78104
rect 637132 78100 637138 78102
rect 639597 78099 639663 78102
rect 581637 77888 625170 77890
rect 581637 77832 581642 77888
rect 581698 77832 625170 77888
rect 581637 77830 625170 77832
rect 581637 77827 581703 77830
rect 624417 77346 624483 77349
rect 633893 77346 633959 77349
rect 624417 77344 633959 77346
rect 624417 77288 624422 77344
rect 624478 77288 633898 77344
rect 633954 77288 633959 77344
rect 624417 77286 633959 77288
rect 624417 77283 624483 77286
rect 633893 77283 633959 77286
rect 578233 75578 578299 75581
rect 575798 75576 578299 75578
rect 575798 75520 578238 75576
rect 578294 75520 578299 75576
rect 575798 75518 578299 75520
rect 575798 75140 575858 75518
rect 578233 75515 578299 75518
rect 646129 74218 646195 74221
rect 646086 74216 646195 74218
rect 646086 74160 646134 74216
rect 646190 74160 646195 74216
rect 646086 74155 646195 74160
rect 646086 73848 646146 74155
rect 579061 73130 579127 73133
rect 575798 73128 579127 73130
rect 575798 73072 579066 73128
rect 579122 73072 579127 73128
rect 575798 73070 579127 73072
rect 575798 72964 575858 73070
rect 579061 73067 579127 73070
rect 646313 71770 646379 71773
rect 646270 71768 646379 71770
rect 646270 71712 646318 71768
rect 646374 71712 646379 71768
rect 646270 71707 646379 71712
rect 646270 71400 646330 71707
rect 579061 71226 579127 71229
rect 575798 71224 579127 71226
rect 575798 71168 579066 71224
rect 579122 71168 579127 71224
rect 575798 71166 579127 71168
rect 575798 70788 575858 71166
rect 579061 71163 579127 71166
rect 646638 68914 646698 68952
rect 647233 68914 647299 68917
rect 646638 68912 647299 68914
rect 646638 68856 647238 68912
rect 647294 68856 647299 68912
rect 646638 68854 647299 68856
rect 647233 68851 647299 68854
rect 646497 67146 646563 67149
rect 646454 67144 646563 67146
rect 646454 67088 646502 67144
rect 646558 67088 646563 67144
rect 646454 67083 646563 67088
rect 646454 66504 646514 67083
rect 646129 64426 646195 64429
rect 646086 64424 646195 64426
rect 646086 64368 646134 64424
rect 646190 64368 646195 64424
rect 646086 64363 646195 64368
rect 646086 64056 646146 64363
rect 648613 62114 648679 62117
rect 646638 62112 648679 62114
rect 646638 62056 648618 62112
rect 648674 62056 648679 62112
rect 646638 62054 648679 62056
rect 646638 61608 646698 62054
rect 648613 62051 648679 62054
rect 647233 59258 647299 59261
rect 646638 59256 647299 59258
rect 646638 59200 647238 59256
rect 647294 59200 647299 59256
rect 646638 59198 647299 59200
rect 646638 59160 646698 59198
rect 647233 59195 647299 59198
rect 648797 57354 648863 57357
rect 646638 57352 648863 57354
rect 646638 57296 648802 57352
rect 648858 57296 648863 57352
rect 646638 57294 648863 57296
rect 646638 56712 646698 57294
rect 648797 57291 648863 57294
rect 460790 54980 460796 55044
rect 460860 55042 460866 55044
rect 576117 55042 576183 55045
rect 460860 55040 576183 55042
rect 460860 54984 576122 55040
rect 576178 54984 576183 55040
rect 460860 54982 576183 54984
rect 460860 54980 460866 54982
rect 576117 54979 576183 54982
rect 462630 54708 462636 54772
rect 462700 54770 462706 54772
rect 580257 54770 580323 54773
rect 462700 54768 580323 54770
rect 462700 54712 580262 54768
rect 580318 54712 580323 54768
rect 462700 54710 580323 54712
rect 462700 54708 462706 54710
rect 580257 54707 580323 54710
rect 578877 54498 578943 54501
rect 466410 54496 578943 54498
rect 466410 54440 578882 54496
rect 578938 54440 578943 54496
rect 466410 54438 578943 54440
rect 466410 54226 466470 54438
rect 578877 54435 578943 54438
rect 577497 54226 577563 54229
rect 459878 54166 466470 54226
rect 476070 54224 577563 54226
rect 476070 54168 577502 54224
rect 577558 54168 577563 54224
rect 476070 54166 577563 54168
rect 459878 53685 459938 54166
rect 460790 53892 460796 53956
rect 460860 53892 460866 53956
rect 476070 53954 476130 54166
rect 577497 54163 577563 54166
rect 461718 53894 476130 53954
rect 460798 53685 460858 53892
rect 461718 53685 461778 53894
rect 459829 53680 459938 53685
rect 459829 53624 459834 53680
rect 459890 53624 459938 53680
rect 459829 53622 459938 53624
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 462589 53684 462655 53685
rect 462589 53682 462636 53684
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462544 53680 462636 53682
rect 462544 53624 462594 53680
rect 462544 53622 462636 53624
rect 459829 53619 459895 53622
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53620 462636 53622
rect 462700 53620 462706 53684
rect 462589 53619 462655 53620
rect 471789 53546 471855 53549
rect 473537 53546 473603 53549
rect 471789 53544 473603 53546
rect 471789 53488 471794 53544
rect 471850 53488 473542 53544
rect 473598 53488 473603 53544
rect 471789 53486 473603 53488
rect 471789 53483 471855 53486
rect 473537 53483 473603 53486
rect 464153 53410 464219 53413
rect 464705 53410 464771 53413
rect 464153 53408 464771 53410
rect 464153 53352 464158 53408
rect 464214 53352 464710 53408
rect 464766 53352 464771 53408
rect 464153 53350 464771 53352
rect 464153 53347 464219 53350
rect 464705 53347 464771 53350
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 661585 48512 661651 48515
rect 661480 48510 661651 48512
rect 661480 48454 661590 48510
rect 661646 48454 661651 48510
rect 661480 48452 661651 48454
rect 661585 48449 661651 48452
rect 529606 48044 529612 48108
rect 529676 48106 529682 48108
rect 553669 48106 553735 48109
rect 529676 48104 553735 48106
rect 529676 48048 553674 48104
rect 553730 48048 553735 48104
rect 529676 48046 553735 48048
rect 529676 48044 529682 48046
rect 553669 48043 553735 48046
rect 515438 47772 515444 47836
rect 515508 47834 515514 47836
rect 522941 47834 523007 47837
rect 515508 47832 523007 47834
rect 515508 47776 522946 47832
rect 523002 47776 523007 47832
rect 515508 47774 523007 47776
rect 515508 47772 515514 47774
rect 522941 47771 523007 47774
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465073 47018 465139 47021
rect 458173 47016 465139 47018
rect 458173 46960 458178 47016
rect 458234 46960 465078 47016
rect 465134 46960 465139 47016
rect 458173 46958 465139 46960
rect 458173 46955 458239 46958
rect 465073 46955 465139 46958
rect 458357 46746 458423 46749
rect 465257 46746 465323 46749
rect 458357 46744 465323 46746
rect 458357 46688 458362 46744
rect 458418 46688 465262 46744
rect 465318 46688 465323 46744
rect 458357 46686 465323 46688
rect 458357 46683 458423 46686
rect 465257 46683 465323 46686
rect 461025 44436 461091 44437
rect 460974 44434 460980 44436
rect 460934 44374 460980 44434
rect 461044 44432 461091 44436
rect 461086 44376 461091 44432
rect 460974 44372 460980 44374
rect 461044 44372 461091 44376
rect 462262 44372 462268 44436
rect 462332 44434 462338 44436
rect 462865 44434 462931 44437
rect 463785 44436 463851 44437
rect 463734 44434 463740 44436
rect 462332 44432 462931 44434
rect 462332 44376 462870 44432
rect 462926 44376 462931 44432
rect 462332 44374 462931 44376
rect 463694 44374 463740 44434
rect 463804 44432 463851 44436
rect 463846 44376 463851 44432
rect 462332 44372 462338 44374
rect 461025 44371 461091 44372
rect 462865 44371 462931 44374
rect 463734 44372 463740 44374
rect 463804 44372 463851 44376
rect 463785 44371 463851 44372
rect 130377 44298 130443 44301
rect 132401 44298 132467 44301
rect 142613 44298 142679 44301
rect 130377 44296 132467 44298
rect 130377 44240 130382 44296
rect 130438 44240 132406 44296
rect 132462 44240 132467 44296
rect 130377 44238 132467 44240
rect 130377 44235 130443 44238
rect 132401 44235 132467 44238
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 255865 44162 255931 44165
rect 460105 44162 460171 44165
rect 464337 44162 464403 44165
rect 255865 44160 460171 44162
rect 255865 44104 255870 44160
rect 255926 44104 460110 44160
rect 460166 44104 460171 44160
rect 255865 44102 460171 44104
rect 255865 44099 255931 44102
rect 460105 44099 460171 44102
rect 460890 44160 464403 44162
rect 460890 44104 464342 44160
rect 464398 44104 464403 44160
rect 460890 44102 464403 44104
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 361757 43890 361823 43893
rect 440233 43890 440299 43893
rect 361757 43888 440299 43890
rect 361757 43832 361762 43888
rect 361818 43832 440238 43888
rect 440294 43832 440299 43888
rect 361757 43830 440299 43832
rect 361757 43827 361823 43830
rect 440233 43827 440299 43830
rect 441061 43890 441127 43893
rect 460890 43890 460950 44102
rect 464337 44099 464403 44102
rect 441061 43888 460950 43890
rect 441061 43832 441066 43888
rect 441122 43832 460950 43888
rect 441061 43830 460950 43832
rect 441061 43827 441127 43830
rect 460841 43482 460907 43485
rect 471053 43482 471119 43485
rect 460841 43480 471119 43482
rect 460841 43424 460846 43480
rect 460902 43424 471058 43480
rect 471114 43424 471119 43480
rect 460841 43422 471119 43424
rect 460841 43419 460907 43422
rect 471053 43419 471119 43422
rect 462681 43210 462747 43213
rect 465809 43210 465875 43213
rect 462681 43208 465875 43210
rect 462681 43152 462686 43208
rect 462742 43152 465814 43208
rect 465870 43152 465875 43208
rect 462681 43150 465875 43152
rect 462681 43147 462747 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463969 42938 464035 42941
rect 461761 42936 464035 42938
rect 461761 42880 461766 42936
rect 461822 42880 463974 42936
rect 464030 42880 464035 42936
rect 461761 42878 464035 42880
rect 461761 42875 461827 42878
rect 463969 42875 464035 42878
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 415577 42394 415643 42397
rect 415577 42392 422310 42394
rect 415577 42336 415582 42392
rect 415638 42336 422310 42392
rect 415577 42334 422310 42336
rect 415577 42331 415643 42334
rect 422250 42258 422310 42334
rect 446213 42258 446279 42261
rect 461945 42258 462011 42261
rect 422250 42198 427830 42258
rect 419206 42060 419212 42124
rect 419276 42122 419282 42124
rect 419276 42062 420194 42122
rect 419276 42060 419282 42062
rect 420134 41986 420194 42062
rect 420134 41926 424978 41986
rect 365069 41852 365135 41853
rect 416681 41852 416747 41853
rect 365069 41848 365116 41852
rect 365180 41850 365186 41852
rect 416630 41850 416636 41852
rect 365069 41792 365074 41848
rect 365069 41788 365116 41792
rect 365180 41790 365226 41850
rect 416590 41790 416636 41850
rect 416700 41848 416747 41852
rect 416742 41792 416747 41848
rect 365180 41788 365186 41790
rect 416630 41788 416636 41790
rect 416700 41788 416747 41792
rect 365069 41787 365135 41788
rect 416681 41787 416747 41788
rect 419901 41852 419967 41853
rect 419901 41848 419948 41852
rect 420012 41850 420018 41852
rect 424918 41850 424978 41926
rect 425094 41850 425100 41852
rect 419901 41792 419906 41848
rect 419901 41788 419948 41792
rect 420012 41790 420058 41850
rect 424918 41790 425100 41850
rect 420012 41788 420018 41790
rect 425094 41788 425100 41790
rect 425164 41788 425170 41852
rect 419901 41787 419967 41788
rect 427770 41578 427830 42198
rect 446213 42256 462011 42258
rect 446213 42200 446218 42256
rect 446274 42200 461950 42256
rect 462006 42200 462011 42256
rect 446213 42198 462011 42200
rect 446213 42195 446279 42198
rect 461945 42195 462011 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 529565 42124 529631 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529612 42124
rect 529520 42120 529612 42122
rect 529520 42064 529570 42120
rect 529520 42062 529612 42064
rect 529565 42060 529612 42062
rect 529676 42060 529682 42124
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42060
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 451958 41850 451964 41852
rect 441908 41790 451964 41850
rect 441908 41788 441914 41790
rect 451958 41788 451964 41790
rect 452028 41788 452034 41852
rect 446213 41578 446279 41581
rect 427770 41576 446279 41578
rect 427770 41520 446218 41576
rect 446274 41520 446279 41576
rect 427770 41518 446279 41520
rect 446213 41515 446279 41518
rect 141693 40356 141759 40357
rect 141693 40352 141740 40356
rect 141804 40354 141810 40356
rect 141693 40296 141698 40352
rect 141693 40292 141740 40296
rect 141804 40294 141850 40354
rect 141804 40292 141810 40294
rect 141693 40291 141759 40292
<< via3 >>
rect 233004 997384 233068 997388
rect 233004 997328 233018 997384
rect 233018 997328 233068 997384
rect 233004 997324 233068 997328
rect 285444 997384 285508 997388
rect 285444 997328 285458 997384
rect 285458 997328 285508 997384
rect 285444 997324 285508 997328
rect 387564 997384 387628 997388
rect 387564 997328 387578 997384
rect 387578 997328 387628 997384
rect 387564 997324 387628 997328
rect 233004 990932 233068 990996
rect 387564 990932 387628 990996
rect 285444 987940 285508 988004
rect 675892 892196 675956 892260
rect 675892 887708 675956 887772
rect 675708 885804 675772 885868
rect 675524 880636 675588 880700
rect 676260 880364 676324 880428
rect 675340 878460 675404 878524
rect 675156 877160 675220 877164
rect 675156 877104 675206 877160
rect 675206 877104 675220 877160
rect 675156 877100 675220 877104
rect 675340 874108 675404 874172
rect 676260 873020 676324 873084
rect 676444 872748 676508 872812
rect 675156 870436 675220 870500
rect 675708 865676 675772 865740
rect 676076 865404 676140 865468
rect 675892 864996 675956 865060
rect 41828 813180 41892 813244
rect 41828 809976 41892 809980
rect 41828 809920 41842 809976
rect 41842 809920 41892 809976
rect 41828 809916 41892 809920
rect 41828 807876 41892 807940
rect 40540 805564 40604 805628
rect 40724 805156 40788 805220
rect 40908 804748 40972 804812
rect 41828 804748 41892 804812
rect 41828 802436 41892 802500
rect 42196 801000 42260 801004
rect 42196 800944 42210 801000
rect 42210 800944 42260 801000
rect 42196 800940 42260 800944
rect 41092 800668 41156 800732
rect 40356 800532 40420 800596
rect 41092 796180 41156 796244
rect 40908 794820 40972 794884
rect 42196 794472 42260 794476
rect 42196 794416 42210 794472
rect 42210 794416 42260 794472
rect 42196 794412 42260 794416
rect 40356 793052 40420 793116
rect 40724 790604 40788 790668
rect 40540 789380 40604 789444
rect 41644 789108 41708 789172
rect 41828 788700 41892 788764
rect 41460 788156 41524 788220
rect 676076 788020 676140 788084
rect 674420 786660 674484 786724
rect 675340 786720 675404 786724
rect 675340 786664 675390 786720
rect 675390 786664 675404 786720
rect 675340 786660 675404 786664
rect 41644 769796 41708 769860
rect 41460 768980 41524 769044
rect 40540 766532 40604 766596
rect 40724 765308 40788 765372
rect 40908 764900 40972 764964
rect 41828 757692 41892 757756
rect 40908 754836 40972 754900
rect 42012 754836 42076 754900
rect 40724 754156 40788 754220
rect 42012 750408 42076 750412
rect 42012 750352 42062 750408
rect 42062 750352 42076 750408
rect 42012 750348 42076 750352
rect 40540 746676 40604 746740
rect 41828 745724 41892 745788
rect 41644 745452 41708 745516
rect 41460 745044 41524 745108
rect 674236 743276 674300 743340
rect 674604 738108 674668 738172
rect 675340 730824 675404 730828
rect 675340 730768 675354 730824
rect 675354 730768 675404 730824
rect 675340 730764 675404 730768
rect 676812 729812 676876 729876
rect 676076 726548 676140 726612
rect 674420 726276 674484 726340
rect 41828 725868 41892 725932
rect 41828 725656 41892 725660
rect 41828 725600 41842 725656
rect 41842 725600 41892 725656
rect 41828 725596 41892 725600
rect 674052 721848 674116 721852
rect 674052 721792 674066 721848
rect 674066 721792 674116 721848
rect 674052 721788 674116 721792
rect 40724 721708 40788 721772
rect 675156 721712 675220 721716
rect 675156 721656 675170 721712
rect 675170 721656 675220 721712
rect 675156 721652 675220 721656
rect 674052 719672 674116 719676
rect 674052 719616 674066 719672
rect 674066 719616 674116 719672
rect 674052 719612 674116 719616
rect 40540 718524 40604 718588
rect 41828 716892 41892 716956
rect 42196 714368 42260 714372
rect 42196 714312 42246 714368
rect 42246 714312 42260 714368
rect 42196 714308 42260 714312
rect 40356 714172 40420 714236
rect 40356 709820 40420 709884
rect 40724 707100 40788 707164
rect 42196 706284 42260 706348
rect 40540 704244 40604 704308
rect 41828 701796 41892 701860
rect 41460 701524 41524 701588
rect 41828 700496 41892 700500
rect 41828 700440 41878 700496
rect 41878 700440 41892 700496
rect 41828 700436 41892 700440
rect 675524 696824 675588 696828
rect 675524 696768 675538 696824
rect 675538 696768 675588 696824
rect 675524 696764 675588 696768
rect 674420 694588 674484 694652
rect 675524 683980 675588 684044
rect 675340 683768 675404 683772
rect 675340 683712 675354 683768
rect 675354 683712 675404 683768
rect 675340 683708 675404 683712
rect 42012 683572 42076 683636
rect 674236 682620 674300 682684
rect 42196 681396 42260 681460
rect 40540 678928 40604 678992
rect 41828 678268 41892 678332
rect 676076 676364 676140 676428
rect 41828 672692 41892 672756
rect 42196 672616 42260 672620
rect 42196 672560 42246 672616
rect 42246 672560 42260 672616
rect 42196 672556 42260 672560
rect 42196 668476 42260 668540
rect 676812 665756 676876 665820
rect 40724 665076 40788 665140
rect 40540 663988 40604 664052
rect 674604 662356 674668 662420
rect 41644 658548 41708 658612
rect 41828 658336 41892 658340
rect 41828 658280 41842 658336
rect 41842 658280 41892 658336
rect 41828 658276 41892 658280
rect 41460 657188 41524 657252
rect 674236 652836 674300 652900
rect 675524 645492 675588 645556
rect 675524 643648 675588 643652
rect 675524 643592 675574 643648
rect 675574 643592 675588 643648
rect 675524 643588 675588 643592
rect 41460 640596 41524 640660
rect 676076 637468 676140 637532
rect 40540 635292 40604 635356
rect 40724 634884 40788 634948
rect 675156 631348 675220 631412
rect 676076 631348 676140 631412
rect 41644 629852 41708 629916
rect 41828 629172 41892 629236
rect 40724 621964 40788 622028
rect 40540 620740 40604 620804
rect 674420 618972 674484 619036
rect 676812 617068 676876 617132
rect 673868 616116 673932 616180
rect 41460 615708 41524 615772
rect 41828 615436 41892 615500
rect 41828 613456 41892 613460
rect 41828 613400 41878 613456
rect 41878 613400 41892 613456
rect 41828 613396 41892 613400
rect 40540 612308 40604 612372
rect 674420 602924 674484 602988
rect 40540 601972 40604 602036
rect 43116 598436 43180 598500
rect 42012 597212 42076 597276
rect 43116 597000 43180 597004
rect 43116 596944 43130 597000
rect 43130 596944 43180 597000
rect 43116 596940 43180 596944
rect 674972 595308 675036 595372
rect 41828 593948 41892 594012
rect 675156 593132 675220 593196
rect 40724 592486 40788 592550
rect 41828 592316 41892 592380
rect 42196 592044 42260 592108
rect 676076 591636 676140 591700
rect 674236 591228 674300 591292
rect 674972 590472 675036 590476
rect 674972 590416 674986 590472
rect 674986 590416 675036 590472
rect 674972 590412 675036 590416
rect 676076 586196 676140 586260
rect 62068 585652 62132 585716
rect 41828 585108 41892 585172
rect 40356 584564 40420 584628
rect 40356 580212 40420 580276
rect 40908 577764 40972 577828
rect 676812 576812 676876 576876
rect 40724 575860 40788 575924
rect 40540 575452 40604 575516
rect 42012 575452 42076 575516
rect 42012 573880 42076 573884
rect 42012 573824 42026 573880
rect 42026 573824 42076 573880
rect 42012 573820 42076 573824
rect 41460 573276 41524 573340
rect 41644 571508 41708 571572
rect 41828 570208 41892 570212
rect 41828 570152 41842 570208
rect 41842 570152 41892 570208
rect 41828 570148 41892 570152
rect 675340 561912 675404 561916
rect 675340 561856 675390 561912
rect 675390 561856 675404 561912
rect 675340 561852 675404 561856
rect 41276 559268 41340 559332
rect 41276 557488 41340 557552
rect 676260 557500 676324 557564
rect 41828 553964 41892 554028
rect 676812 553828 676876 553892
rect 41828 552740 41892 552804
rect 676996 548252 677060 548316
rect 676260 547572 676324 547636
rect 674420 547028 674484 547092
rect 676076 546756 676140 546820
rect 675340 545668 675404 545732
rect 40724 545532 40788 545596
rect 40540 545320 40604 545324
rect 40540 545264 40554 545320
rect 40554 545264 40604 545320
rect 40540 545260 40604 545264
rect 44772 543628 44836 543692
rect 41828 542268 41892 542332
rect 40724 535196 40788 535260
rect 40540 533292 40604 533356
rect 41644 532612 41708 532676
rect 41460 530028 41524 530092
rect 41828 528668 41892 528732
rect 676996 503644 677060 503708
rect 676812 500924 676876 500988
rect 44772 489908 44836 489972
rect 676030 488820 676094 488884
rect 675892 487868 675956 487932
rect 673868 455228 673932 455292
rect 41782 423540 41846 423604
rect 42012 421908 42076 421972
rect 40908 418508 40972 418572
rect 40540 418236 40604 418300
rect 40724 417964 40788 418028
rect 42012 417964 42076 418028
rect 41460 417692 41524 417756
rect 41828 417692 41892 417756
rect 42012 415244 42076 415308
rect 41828 414564 41892 414628
rect 40908 406948 40972 407012
rect 40540 406676 40604 406740
rect 40724 404500 40788 404564
rect 677180 401236 677244 401300
rect 676812 400420 676876 400484
rect 41460 400012 41524 400076
rect 41828 399392 41892 399396
rect 41828 399336 41842 399392
rect 41842 399336 41892 399392
rect 41828 399332 41892 399336
rect 42012 398848 42076 398852
rect 42012 398792 42026 398848
rect 42026 398792 42076 398848
rect 42012 398788 42076 398792
rect 676076 398788 676140 398852
rect 676260 396748 676324 396812
rect 676444 396340 676508 396404
rect 676628 395116 676692 395180
rect 675892 392804 675956 392868
rect 675708 387636 675772 387700
rect 676260 384916 676324 384980
rect 676444 382196 676508 382260
rect 41460 381788 41524 381852
rect 41644 379340 41708 379404
rect 40724 378932 40788 378996
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 40908 377708 40972 377772
rect 676628 377300 676692 377364
rect 41828 374580 41892 374644
rect 676076 373628 676140 373692
rect 675340 372464 675404 372468
rect 675340 372408 675390 372464
rect 675390 372408 675404 372464
rect 675340 372404 675404 372408
rect 675340 366284 675404 366348
rect 40908 364788 40972 364852
rect 40724 364108 40788 364172
rect 40540 360028 40604 360092
rect 41828 358728 41892 358732
rect 41828 358672 41878 358728
rect 41878 358672 41892 358728
rect 41828 358668 41892 358672
rect 41460 356900 41524 356964
rect 41828 355736 41892 355740
rect 41828 355680 41878 355736
rect 41878 355680 41892 355736
rect 41828 355676 41892 355680
rect 43300 354452 43364 354516
rect 675524 354180 675588 354244
rect 675892 353772 675956 353836
rect 675708 352956 675772 353020
rect 675892 351732 675956 351796
rect 675340 347652 675404 347716
rect 676444 346564 676508 346628
rect 44588 342892 44652 342956
rect 42748 340172 42812 340236
rect 676260 340172 676324 340236
rect 44404 339764 44468 339828
rect 675524 339416 675588 339420
rect 675524 339360 675538 339416
rect 675538 339360 675588 339416
rect 675524 339356 675588 339360
rect 41644 338132 41708 338196
rect 676076 337860 676140 337924
rect 44772 337316 44836 337380
rect 40540 336908 40604 336972
rect 42932 336772 42996 336836
rect 41460 336500 41524 336564
rect 676444 336500 676508 336564
rect 40908 335684 40972 335748
rect 40724 335276 40788 335340
rect 43300 334596 43364 334660
rect 41828 331196 41892 331260
rect 675340 327992 675404 327996
rect 675340 327936 675390 327992
rect 675390 327936 675404 327992
rect 675340 327932 675404 327936
rect 676628 325620 676692 325684
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 40908 321132 40972 321196
rect 41828 319968 41892 319972
rect 41828 319912 41842 319968
rect 41842 319912 41892 319968
rect 41828 319908 41892 319912
rect 40724 317324 40788 317388
rect 42932 316372 42996 316436
rect 40540 315964 40604 316028
rect 41460 313652 41524 313716
rect 675340 309164 675404 309228
rect 675892 308756 675956 308820
rect 676076 304540 676140 304604
rect 675892 302636 675956 302700
rect 676628 301608 676692 301612
rect 676628 301552 676642 301608
rect 676642 301552 676692 301608
rect 676628 301548 676692 301552
rect 44588 300052 44652 300116
rect 42748 299236 42812 299300
rect 44772 298420 44836 298484
rect 44404 297604 44468 297668
rect 675708 297332 675772 297396
rect 42196 296788 42260 296852
rect 675524 296516 675588 296580
rect 42012 295564 42076 295628
rect 676444 294612 676508 294676
rect 41828 294340 41892 294404
rect 40724 292528 40788 292592
rect 675524 292224 675588 292228
rect 675524 292168 675574 292224
rect 675574 292168 675588 292224
rect 675524 292164 675588 292168
rect 41828 291756 41892 291820
rect 676628 290940 676692 291004
rect 41828 289988 41892 290052
rect 42196 289988 42260 290052
rect 676260 286996 676324 287060
rect 41828 284820 41892 284884
rect 676076 283596 676140 283660
rect 676076 282644 676140 282708
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 62068 278836 62132 278900
rect 40908 277068 40972 277132
rect 40724 274212 40788 274276
rect 675340 273804 675404 273868
rect 41828 273048 41892 273052
rect 41828 272992 41842 273048
rect 41842 272992 41892 273048
rect 41828 272988 41892 272992
rect 41828 272368 41892 272372
rect 41828 272312 41842 272368
rect 41842 272312 41892 272368
rect 41828 272308 41892 272312
rect 41460 270404 41524 270468
rect 40540 269724 40604 269788
rect 676996 261564 677060 261628
rect 676812 261156 676876 261220
rect 675524 258088 675588 258092
rect 675524 258032 675538 258088
rect 675538 258032 675588 258088
rect 675524 258028 675588 258032
rect 676996 250276 677060 250340
rect 675524 250064 675588 250068
rect 675524 250008 675538 250064
rect 675538 250008 675588 250064
rect 675524 250004 675588 250008
rect 40540 249732 40604 249796
rect 675340 249596 675404 249660
rect 40724 249324 40788 249388
rect 676812 246604 676876 246668
rect 673316 246196 673380 246260
rect 674604 246196 674668 246260
rect 667796 245652 667860 245716
rect 675524 245244 675588 245308
rect 676812 241844 676876 241908
rect 42012 238036 42076 238100
rect 40540 236540 40604 236604
rect 675524 235512 675588 235516
rect 675524 235456 675538 235512
rect 675538 235456 675588 235512
rect 675524 235452 675588 235456
rect 40724 234636 40788 234700
rect 670740 231916 670804 231980
rect 675524 228576 675588 228580
rect 675524 228520 675538 228576
rect 675538 228520 675588 228576
rect 675524 228516 675588 228520
rect 42012 227352 42076 227356
rect 42012 227296 42026 227352
rect 42026 227296 42076 227352
rect 42012 227292 42076 227296
rect 672580 227020 672644 227084
rect 674052 226476 674116 226540
rect 591988 223348 592052 223412
rect 669452 223348 669516 223412
rect 649580 222940 649644 223004
rect 651972 222940 652036 223004
rect 676030 219812 676094 219876
rect 669452 218860 669516 218924
rect 675708 218588 675772 218652
rect 669636 218180 669700 218244
rect 670372 217908 670436 217972
rect 675892 217908 675956 217972
rect 511028 217560 511092 217564
rect 511028 217504 511042 217560
rect 511042 217504 511092 217560
rect 511028 217500 511092 217504
rect 520044 217560 520108 217564
rect 520044 217504 520058 217560
rect 520058 217504 520108 217560
rect 520044 217500 520108 217504
rect 532556 217560 532620 217564
rect 532556 217504 532570 217560
rect 532570 217504 532620 217560
rect 532556 217500 532620 217504
rect 670372 217092 670436 217156
rect 669452 216608 669516 216612
rect 669452 216552 669466 216608
rect 669466 216552 669516 216608
rect 669452 216548 669516 216552
rect 520044 215868 520108 215932
rect 511028 215596 511092 215660
rect 532556 215324 532620 215388
rect 675892 215460 675956 215524
rect 675892 212468 675956 212532
rect 676628 211380 676692 211444
rect 41828 210020 41892 210084
rect 41644 208116 41708 208180
rect 40540 207300 40604 207364
rect 674604 206892 674668 206956
rect 40724 206484 40788 206548
rect 40908 206076 40972 206140
rect 669268 205668 669332 205732
rect 669636 205668 669700 205732
rect 669268 205396 669332 205460
rect 669636 205396 669700 205460
rect 41460 204852 41524 204916
rect 41460 204036 41524 204100
rect 676444 202676 676508 202740
rect 672580 200772 672644 200836
rect 676628 199956 676692 200020
rect 42012 198732 42076 198796
rect 670740 198732 670804 198796
rect 676812 197916 676876 197980
rect 669268 196012 669332 196076
rect 669636 196012 669700 196076
rect 42012 195664 42076 195668
rect 42012 195608 42026 195664
rect 42026 195608 42076 195664
rect 42012 195604 42076 195608
rect 41828 195256 41892 195260
rect 41828 195200 41842 195256
rect 41842 195200 41892 195256
rect 41828 195196 41892 195200
rect 40908 194924 40972 194988
rect 676260 194516 676324 194580
rect 40724 193428 40788 193492
rect 676076 193156 676140 193220
rect 675892 192748 675956 192812
rect 669452 191660 669516 191724
rect 675340 189076 675404 189140
rect 40540 186356 40604 186420
rect 41460 185948 41524 186012
rect 673132 181520 673196 181524
rect 673132 181464 673146 181520
rect 673146 181464 673196 181520
rect 673132 181460 673196 181464
rect 668164 179556 668228 179620
rect 673316 178060 673380 178124
rect 676812 176608 676876 176672
rect 675892 172756 675956 172820
rect 675892 169356 675956 169420
rect 675340 167452 675404 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 676076 162692 676140 162756
rect 673132 161468 673196 161532
rect 676444 156980 676508 157044
rect 676260 155756 676324 155820
rect 676628 151404 676692 151468
rect 676076 148412 676140 148476
rect 675340 147656 675404 147660
rect 675340 147600 675390 147656
rect 675390 147600 675404 147656
rect 675340 147596 675404 147600
rect 669268 140388 669332 140452
rect 667796 134540 667860 134604
rect 676812 127332 676876 127396
rect 676076 126924 676140 126988
rect 676260 125700 676324 125764
rect 676444 124068 676508 124132
rect 676628 124068 676692 124132
rect 676444 123660 676508 123724
rect 676260 122844 676324 122908
rect 676812 122844 676876 122908
rect 675340 122028 675404 122092
rect 675708 117268 675772 117332
rect 674052 115772 674116 115836
rect 676260 112372 676324 112436
rect 676444 111692 676508 111756
rect 675708 111344 675772 111348
rect 675708 111288 675758 111344
rect 675758 111288 675772 111344
rect 675708 111284 675772 111288
rect 676628 110332 676692 110396
rect 676076 108156 676140 108220
rect 675340 101960 675404 101964
rect 675340 101904 675390 101960
rect 675390 101904 675404 101960
rect 675340 101900 675404 101904
rect 637252 96868 637316 96932
rect 647188 96460 647252 96524
rect 633940 95372 634004 95436
rect 650316 93060 650380 93124
rect 633940 78568 634004 78572
rect 633940 78512 633954 78568
rect 633954 78512 634004 78568
rect 633940 78508 634004 78512
rect 637068 78100 637132 78164
rect 460796 54980 460860 55044
rect 462636 54708 462700 54772
rect 460796 53892 460860 53956
rect 462636 53680 462700 53684
rect 462636 53624 462650 53680
rect 462650 53624 462700 53680
rect 462636 53620 462700 53624
rect 518756 48860 518820 48924
rect 529612 48044 529676 48108
rect 515444 47772 515508 47836
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 522068 47228 522132 47292
rect 460980 44432 461044 44436
rect 460980 44376 461030 44432
rect 461030 44376 461044 44432
rect 460980 44372 461044 44376
rect 462268 44372 462332 44436
rect 463740 44432 463804 44436
rect 463740 44376 463790 44432
rect 463790 44376 463804 44432
rect 463740 44372 463804 44376
rect 141740 43964 141804 44028
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 419212 42060 419276 42124
rect 365116 41848 365180 41852
rect 365116 41792 365130 41848
rect 365130 41792 365180 41848
rect 365116 41788 365180 41792
rect 416636 41848 416700 41852
rect 416636 41792 416686 41848
rect 416686 41792 416700 41848
rect 416636 41788 416700 41792
rect 419948 41848 420012 41852
rect 419948 41792 419962 41848
rect 419962 41792 420012 41848
rect 419948 41788 420012 41792
rect 425100 41788 425164 41852
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529612 42120 529676 42124
rect 529612 42064 529626 42120
rect 529626 42064 529676 42120
rect 529612 42060 529676 42064
rect 441844 41788 441908 41852
rect 451964 41788 452028 41852
rect 141740 40352 141804 40356
rect 141740 40296 141754 40352
rect 141754 40296 141804 40352
rect 141740 40292 141804 40296
<< metal4 >>
rect 233003 997388 233069 997389
rect 233003 997324 233004 997388
rect 233068 997324 233069 997388
rect 233003 997323 233069 997324
rect 285443 997388 285509 997389
rect 285443 997324 285444 997388
rect 285508 997324 285509 997388
rect 285443 997323 285509 997324
rect 387563 997388 387629 997389
rect 387563 997324 387564 997388
rect 387628 997324 387629 997388
rect 387563 997323 387629 997324
rect 233006 990997 233066 997323
rect 233003 990996 233069 990997
rect 233003 990932 233004 990996
rect 233068 990932 233069 990996
rect 233003 990931 233069 990932
rect 285446 988005 285506 997323
rect 387566 990997 387626 997323
rect 387563 990996 387629 990997
rect 387563 990932 387564 990996
rect 387628 990932 387629 990996
rect 387563 990931 387629 990932
rect 285443 988004 285509 988005
rect 285443 987940 285444 988004
rect 285508 987940 285509 988004
rect 285443 987939 285509 987940
rect 675891 892260 675957 892261
rect 675891 892196 675892 892260
rect 675956 892196 675957 892260
rect 675891 892195 675957 892196
rect 675894 891510 675954 892195
rect 675710 891450 675954 891510
rect 675710 887090 675770 891450
rect 675891 887772 675957 887773
rect 675891 887708 675892 887772
rect 675956 887770 675957 887772
rect 675956 887710 676322 887770
rect 675956 887708 675957 887710
rect 675891 887707 675957 887708
rect 675710 887030 675954 887090
rect 675707 885868 675773 885869
rect 675707 885804 675708 885868
rect 675772 885804 675773 885868
rect 675707 885803 675773 885804
rect 675523 880700 675589 880701
rect 675523 880636 675524 880700
rect 675588 880636 675589 880700
rect 675523 880635 675589 880636
rect 675339 878524 675405 878525
rect 675339 878460 675340 878524
rect 675404 878460 675405 878524
rect 675339 878459 675405 878460
rect 675155 877164 675221 877165
rect 675155 877100 675156 877164
rect 675220 877100 675221 877164
rect 675155 877099 675221 877100
rect 675158 870501 675218 877099
rect 675342 874173 675402 878459
rect 675339 874172 675405 874173
rect 675339 874108 675340 874172
rect 675404 874108 675405 874172
rect 675339 874107 675405 874108
rect 675526 872190 675586 880635
rect 675710 876890 675770 885803
rect 675894 881850 675954 887030
rect 676262 881850 676322 887710
rect 675894 881790 676138 881850
rect 676262 881790 676506 881850
rect 675710 876830 675954 876890
rect 675526 872130 675770 872190
rect 675155 870500 675221 870501
rect 675155 870436 675156 870500
rect 675220 870436 675221 870500
rect 675155 870435 675221 870436
rect 675710 865741 675770 872130
rect 675707 865740 675773 865741
rect 675707 865676 675708 865740
rect 675772 865676 675773 865740
rect 675707 865675 675773 865676
rect 675894 865061 675954 876830
rect 676078 865469 676138 881790
rect 676259 880428 676325 880429
rect 676259 880364 676260 880428
rect 676324 880364 676325 880428
rect 676259 880363 676325 880364
rect 676262 873085 676322 880363
rect 676259 873084 676325 873085
rect 676259 873020 676260 873084
rect 676324 873020 676325 873084
rect 676259 873019 676325 873020
rect 676446 872813 676506 881790
rect 676443 872812 676509 872813
rect 676443 872748 676444 872812
rect 676508 872748 676509 872812
rect 676443 872747 676509 872748
rect 676075 865468 676141 865469
rect 676075 865404 676076 865468
rect 676140 865404 676141 865468
rect 676075 865403 676141 865404
rect 675891 865060 675957 865061
rect 675891 864996 675892 865060
rect 675956 864996 675957 865060
rect 675891 864995 675957 864996
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40539 805628 40605 805629
rect 40539 805564 40540 805628
rect 40604 805564 40605 805628
rect 40539 805563 40605 805564
rect 40355 800596 40421 800597
rect 40355 800532 40356 800596
rect 40420 800532 40421 800596
rect 40355 800531 40421 800532
rect 40358 793117 40418 800531
rect 40355 793116 40421 793117
rect 40355 793052 40356 793116
rect 40420 793052 40421 793116
rect 40355 793051 40421 793052
rect 40542 789445 40602 805563
rect 40723 805220 40789 805221
rect 40723 805156 40724 805220
rect 40788 805156 40789 805220
rect 40723 805155 40789 805156
rect 40726 790669 40786 805155
rect 40907 804812 40973 804813
rect 40907 804748 40908 804812
rect 40972 804748 40973 804812
rect 40907 804747 40973 804748
rect 40910 794885 40970 804747
rect 41091 800732 41157 800733
rect 41091 800668 41092 800732
rect 41156 800668 41157 800732
rect 41091 800667 41157 800668
rect 41094 796245 41154 800667
rect 41091 796244 41157 796245
rect 41091 796180 41092 796244
rect 41156 796180 41157 796244
rect 41091 796179 41157 796180
rect 40907 794884 40973 794885
rect 40907 794820 40908 794884
rect 40972 794820 40973 794884
rect 40907 794819 40973 794820
rect 40723 790668 40789 790669
rect 40723 790604 40724 790668
rect 40788 790604 40789 790668
rect 40723 790603 40789 790604
rect 40539 789444 40605 789445
rect 40539 789380 40540 789444
rect 40604 789380 40605 789444
rect 40539 789379 40605 789380
rect 41462 788221 41522 812910
rect 41827 809980 41893 809981
rect 41827 809916 41828 809980
rect 41892 809916 41893 809980
rect 41827 809915 41893 809916
rect 41830 808710 41890 809915
rect 41646 808650 41890 808710
rect 41646 789173 41706 808650
rect 41827 807940 41893 807941
rect 41827 807876 41828 807940
rect 41892 807876 41893 807940
rect 41827 807875 41893 807876
rect 41830 804813 41890 807875
rect 41827 804812 41893 804813
rect 41827 804748 41828 804812
rect 41892 804748 41893 804812
rect 41827 804747 41893 804748
rect 41827 802500 41893 802501
rect 41827 802436 41828 802500
rect 41892 802436 41893 802500
rect 41827 802435 41893 802436
rect 41643 789172 41709 789173
rect 41643 789108 41644 789172
rect 41708 789108 41709 789172
rect 41643 789107 41709 789108
rect 41830 788765 41890 802435
rect 42195 801004 42261 801005
rect 42195 800940 42196 801004
rect 42260 800940 42261 801004
rect 42195 800939 42261 800940
rect 42198 794477 42258 800939
rect 42195 794476 42261 794477
rect 42195 794412 42196 794476
rect 42260 794412 42261 794476
rect 42195 794411 42261 794412
rect 41827 788764 41893 788765
rect 41827 788700 41828 788764
rect 41892 788700 41893 788764
rect 41827 788699 41893 788700
rect 41459 788220 41525 788221
rect 41459 788156 41460 788220
rect 41524 788156 41525 788220
rect 41459 788155 41525 788156
rect 676075 788084 676141 788085
rect 676075 788020 676076 788084
rect 676140 788020 676141 788084
rect 676075 788019 676141 788020
rect 674419 786724 674485 786725
rect 674419 786660 674420 786724
rect 674484 786660 674485 786724
rect 674419 786659 674485 786660
rect 675339 786724 675405 786725
rect 675339 786660 675340 786724
rect 675404 786660 675405 786724
rect 675339 786659 675405 786660
rect 41643 769860 41709 769861
rect 41643 769796 41644 769860
rect 41708 769796 41709 769860
rect 41643 769795 41709 769796
rect 41459 769044 41525 769045
rect 41459 768980 41460 769044
rect 41524 768980 41525 769044
rect 41459 768979 41525 768980
rect 40539 766596 40605 766597
rect 40539 766532 40540 766596
rect 40604 766532 40605 766596
rect 40539 766531 40605 766532
rect 40542 746741 40602 766531
rect 40723 765372 40789 765373
rect 40723 765308 40724 765372
rect 40788 765308 40789 765372
rect 40723 765307 40789 765308
rect 40726 754221 40786 765307
rect 40907 764964 40973 764965
rect 40907 764900 40908 764964
rect 40972 764900 40973 764964
rect 40907 764899 40973 764900
rect 40910 754901 40970 764899
rect 40907 754900 40973 754901
rect 40907 754836 40908 754900
rect 40972 754836 40973 754900
rect 40907 754835 40973 754836
rect 40723 754220 40789 754221
rect 40723 754156 40724 754220
rect 40788 754156 40789 754220
rect 40723 754155 40789 754156
rect 40539 746740 40605 746741
rect 40539 746676 40540 746740
rect 40604 746676 40605 746740
rect 40539 746675 40605 746676
rect 41462 745109 41522 768979
rect 41646 745517 41706 769795
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41830 745789 41890 757691
rect 42011 754900 42077 754901
rect 42011 754836 42012 754900
rect 42076 754836 42077 754900
rect 42011 754835 42077 754836
rect 42014 750413 42074 754835
rect 42011 750412 42077 750413
rect 42011 750348 42012 750412
rect 42076 750348 42077 750412
rect 42011 750347 42077 750348
rect 41827 745788 41893 745789
rect 41827 745724 41828 745788
rect 41892 745724 41893 745788
rect 41827 745723 41893 745724
rect 41643 745516 41709 745517
rect 41643 745452 41644 745516
rect 41708 745452 41709 745516
rect 41643 745451 41709 745452
rect 41459 745108 41525 745109
rect 41459 745044 41460 745108
rect 41524 745044 41525 745108
rect 41459 745043 41525 745044
rect 674235 743340 674301 743341
rect 674235 743276 674236 743340
rect 674300 743276 674301 743340
rect 674235 743275 674301 743276
rect 41827 725932 41893 725933
rect 41827 725930 41828 725932
rect 41646 725870 41828 725930
rect 41646 724530 41706 725870
rect 41827 725868 41828 725870
rect 41892 725868 41893 725932
rect 41827 725867 41893 725868
rect 41827 725660 41893 725661
rect 41827 725596 41828 725660
rect 41892 725596 41893 725660
rect 41827 725595 41893 725596
rect 41462 724470 41706 724530
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40355 714236 40421 714237
rect 40355 714172 40356 714236
rect 40420 714172 40421 714236
rect 40355 714171 40421 714172
rect 40358 709885 40418 714171
rect 40355 709884 40421 709885
rect 40355 709820 40356 709884
rect 40420 709820 40421 709884
rect 40355 709819 40421 709820
rect 40542 704309 40602 718523
rect 40726 707165 40786 721707
rect 40723 707164 40789 707165
rect 40723 707100 40724 707164
rect 40788 707100 40789 707164
rect 40723 707099 40789 707100
rect 40539 704308 40605 704309
rect 40539 704244 40540 704308
rect 40604 704244 40605 704308
rect 40539 704243 40605 704244
rect 41462 701589 41522 724470
rect 41830 717630 41890 725595
rect 674051 721852 674117 721853
rect 674051 721788 674052 721852
rect 674116 721788 674117 721852
rect 674051 721787 674117 721788
rect 674054 719677 674114 721787
rect 674051 719676 674117 719677
rect 674051 719612 674052 719676
rect 674116 719612 674117 719676
rect 674051 719611 674117 719612
rect 41646 717570 41890 717630
rect 41459 701588 41525 701589
rect 41459 701524 41460 701588
rect 41524 701524 41525 701588
rect 41646 701586 41706 717570
rect 41827 716956 41893 716957
rect 41827 716892 41828 716956
rect 41892 716892 41893 716956
rect 41827 716891 41893 716892
rect 41830 701861 41890 716891
rect 42195 714372 42261 714373
rect 42195 714308 42196 714372
rect 42260 714308 42261 714372
rect 42195 714307 42261 714308
rect 42198 706349 42258 714307
rect 42195 706348 42261 706349
rect 42195 706284 42196 706348
rect 42260 706284 42261 706348
rect 42195 706283 42261 706284
rect 41827 701860 41893 701861
rect 41827 701796 41828 701860
rect 41892 701796 41893 701860
rect 41827 701795 41893 701796
rect 41646 701526 41890 701586
rect 41459 701523 41525 701524
rect 41830 700501 41890 701526
rect 41827 700500 41893 700501
rect 41827 700436 41828 700500
rect 41892 700436 41893 700500
rect 41827 700435 41893 700436
rect 42011 683636 42077 683637
rect 42011 683572 42012 683636
rect 42076 683572 42077 683636
rect 42011 683571 42077 683572
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40542 664053 40602 678927
rect 41827 678332 41893 678333
rect 41827 678330 41828 678332
rect 40726 678270 41828 678330
rect 40726 665141 40786 678270
rect 41827 678268 41828 678270
rect 41892 678268 41893 678332
rect 41827 678267 41893 678268
rect 42014 674930 42074 683571
rect 674238 682685 674298 743275
rect 674422 726341 674482 786659
rect 674603 738172 674669 738173
rect 674603 738108 674604 738172
rect 674668 738108 674669 738172
rect 674603 738107 674669 738108
rect 674419 726340 674485 726341
rect 674419 726276 674420 726340
rect 674484 726276 674485 726340
rect 674419 726275 674485 726276
rect 674419 694652 674485 694653
rect 674419 694588 674420 694652
rect 674484 694588 674485 694652
rect 674419 694587 674485 694588
rect 674235 682684 674301 682685
rect 674235 682620 674236 682684
rect 674300 682620 674301 682684
rect 674235 682619 674301 682620
rect 42195 681460 42261 681461
rect 42195 681396 42196 681460
rect 42260 681396 42261 681460
rect 42195 681395 42261 681396
rect 41462 674870 42074 674930
rect 40723 665140 40789 665141
rect 40723 665076 40724 665140
rect 40788 665076 40789 665140
rect 40723 665075 40789 665076
rect 40539 664052 40605 664053
rect 40539 663988 40540 664052
rect 40604 663988 40605 664052
rect 40539 663987 40605 663988
rect 41462 657253 41522 674870
rect 42198 674250 42258 681395
rect 41646 674190 42258 674250
rect 41646 658613 41706 674190
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 672691
rect 42195 672620 42261 672621
rect 42195 672556 42196 672620
rect 42260 672556 42261 672620
rect 42195 672555 42261 672556
rect 42198 668541 42258 672555
rect 42195 668540 42261 668541
rect 42195 668476 42196 668540
rect 42260 668476 42261 668540
rect 42195 668475 42261 668476
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 41459 657252 41525 657253
rect 41459 657188 41460 657252
rect 41524 657188 41525 657252
rect 41459 657187 41525 657188
rect 674235 652900 674301 652901
rect 674235 652836 674236 652900
rect 674300 652836 674301 652900
rect 674235 652835 674301 652836
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40539 635356 40605 635357
rect 40539 635292 40540 635356
rect 40604 635292 40605 635356
rect 40539 635291 40605 635292
rect 40542 620805 40602 635291
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40726 622029 40786 634883
rect 40723 622028 40789 622029
rect 40723 621964 40724 622028
rect 40788 621964 40789 622028
rect 40723 621963 40789 621964
rect 40539 620804 40605 620805
rect 40539 620740 40540 620804
rect 40604 620740 40605 620804
rect 40539 620739 40605 620740
rect 41462 615773 41522 640595
rect 41643 629916 41709 629917
rect 41643 629852 41644 629916
rect 41708 629852 41709 629916
rect 41643 629851 41709 629852
rect 41459 615772 41525 615773
rect 41459 615708 41460 615772
rect 41524 615708 41525 615772
rect 41459 615707 41525 615708
rect 41646 615090 41706 629851
rect 41827 629236 41893 629237
rect 41827 629172 41828 629236
rect 41892 629172 41893 629236
rect 41827 629171 41893 629172
rect 41830 615501 41890 629171
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 41827 615500 41893 615501
rect 41827 615436 41828 615500
rect 41892 615436 41893 615500
rect 41827 615435 41893 615436
rect 41646 615030 41890 615090
rect 41830 613461 41890 615030
rect 41827 613460 41893 613461
rect 41827 613396 41828 613460
rect 41892 613396 41893 613460
rect 41827 613395 41893 613396
rect 40539 612372 40605 612373
rect 40539 612308 40540 612372
rect 40604 612308 40605 612372
rect 40539 612307 40605 612308
rect 40542 602037 40602 612307
rect 40539 602036 40605 602037
rect 40539 601972 40540 602036
rect 40604 601972 40605 602036
rect 40539 601971 40605 601972
rect 43115 598500 43181 598501
rect 43115 598436 43116 598500
rect 43180 598436 43181 598500
rect 43115 598435 43181 598436
rect 42011 597276 42077 597277
rect 42011 597212 42012 597276
rect 42076 597212 42077 597276
rect 42011 597211 42077 597212
rect 41827 594012 41893 594013
rect 41827 594010 41828 594012
rect 40542 593950 41828 594010
rect 40355 584628 40421 584629
rect 40355 584564 40356 584628
rect 40420 584564 40421 584628
rect 40355 584563 40421 584564
rect 40358 580277 40418 584563
rect 40355 580276 40421 580277
rect 40355 580212 40356 580276
rect 40420 580212 40421 580276
rect 40355 580211 40421 580212
rect 40542 575517 40602 593950
rect 41827 593948 41828 593950
rect 41892 593948 41893 594012
rect 41827 593947 41893 593948
rect 40723 592550 40789 592551
rect 40723 592486 40724 592550
rect 40788 592486 40789 592550
rect 40723 592485 40789 592486
rect 40726 575925 40786 592485
rect 41827 592380 41893 592381
rect 41827 592316 41828 592380
rect 41892 592316 41893 592380
rect 41827 592315 41893 592316
rect 41830 592050 41890 592315
rect 41462 591990 41890 592050
rect 41462 591970 41522 591990
rect 40910 591910 41522 591970
rect 40910 577829 40970 591910
rect 42014 587890 42074 597211
rect 43118 597005 43178 598435
rect 43115 597004 43181 597005
rect 43115 596940 43116 597004
rect 43180 596940 43181 597004
rect 43115 596939 43181 596940
rect 42195 592108 42261 592109
rect 42195 592044 42196 592108
rect 42260 592044 42261 592108
rect 42195 592043 42261 592044
rect 41462 587830 42074 587890
rect 40907 577828 40973 577829
rect 40907 577764 40908 577828
rect 40972 577764 40973 577828
rect 40907 577763 40973 577764
rect 40723 575924 40789 575925
rect 40723 575860 40724 575924
rect 40788 575860 40789 575924
rect 40723 575859 40789 575860
rect 40539 575516 40605 575517
rect 40539 575452 40540 575516
rect 40604 575452 40605 575516
rect 40539 575451 40605 575452
rect 41462 573341 41522 587830
rect 42198 587210 42258 592043
rect 41646 587150 42258 587210
rect 41459 573340 41525 573341
rect 41459 573276 41460 573340
rect 41524 573276 41525 573340
rect 41459 573275 41525 573276
rect 41646 571573 41706 587150
rect 62067 585716 62133 585717
rect 62067 585652 62068 585716
rect 62132 585652 62133 585716
rect 62067 585651 62133 585652
rect 41827 585172 41893 585173
rect 41827 585108 41828 585172
rect 41892 585108 41893 585172
rect 41827 585107 41893 585108
rect 41643 571572 41709 571573
rect 41643 571508 41644 571572
rect 41708 571508 41709 571572
rect 41643 571507 41709 571508
rect 41830 570213 41890 585107
rect 42011 575516 42077 575517
rect 42011 575452 42012 575516
rect 42076 575452 42077 575516
rect 42011 575451 42077 575452
rect 42014 573885 42074 575451
rect 42011 573884 42077 573885
rect 42011 573820 42012 573884
rect 42076 573820 42077 573884
rect 42011 573819 42077 573820
rect 41827 570212 41893 570213
rect 41827 570148 41828 570212
rect 41892 570148 41893 570212
rect 41827 570147 41893 570148
rect 41275 559332 41341 559333
rect 41275 559268 41276 559332
rect 41340 559268 41341 559332
rect 41275 559267 41341 559268
rect 41278 557553 41338 559267
rect 41275 557552 41341 557553
rect 41275 557488 41276 557552
rect 41340 557488 41341 557552
rect 41275 557487 41341 557488
rect 41827 554028 41893 554029
rect 41827 553964 41828 554028
rect 41892 553964 41893 554028
rect 41827 553963 41893 553964
rect 41830 553410 41890 553963
rect 41462 553350 41890 553410
rect 40723 545596 40789 545597
rect 40723 545532 40724 545596
rect 40788 545532 40789 545596
rect 40723 545531 40789 545532
rect 40539 545324 40605 545325
rect 40539 545260 40540 545324
rect 40604 545260 40605 545324
rect 40539 545259 40605 545260
rect 40542 533357 40602 545259
rect 40726 535261 40786 545531
rect 40723 535260 40789 535261
rect 40723 535196 40724 535260
rect 40788 535196 40789 535260
rect 40723 535195 40789 535196
rect 40539 533356 40605 533357
rect 40539 533292 40540 533356
rect 40604 533292 40605 533356
rect 40539 533291 40605 533292
rect 41462 530093 41522 553350
rect 41827 552804 41893 552805
rect 41827 552740 41828 552804
rect 41892 552740 41893 552804
rect 41827 552739 41893 552740
rect 41830 543750 41890 552739
rect 41646 543690 41890 543750
rect 44771 543692 44837 543693
rect 41646 532677 41706 543690
rect 44771 543628 44772 543692
rect 44836 543628 44837 543692
rect 44771 543627 44837 543628
rect 41827 542332 41893 542333
rect 41827 542268 41828 542332
rect 41892 542268 41893 542332
rect 41827 542267 41893 542268
rect 41643 532676 41709 532677
rect 41643 532612 41644 532676
rect 41708 532612 41709 532676
rect 41643 532611 41709 532612
rect 41459 530092 41525 530093
rect 41459 530028 41460 530092
rect 41524 530028 41525 530092
rect 41459 530027 41525 530028
rect 41830 528733 41890 542267
rect 41827 528732 41893 528733
rect 41827 528668 41828 528732
rect 41892 528668 41893 528732
rect 41827 528667 41893 528668
rect 44774 489973 44834 543627
rect 44771 489972 44837 489973
rect 44771 489908 44772 489972
rect 44836 489908 44837 489972
rect 44771 489907 44837 489908
rect 41781 423604 41847 423605
rect 41781 423540 41782 423604
rect 41846 423602 41847 423604
rect 41846 423540 41890 423602
rect 41781 423539 41890 423540
rect 40907 418572 40973 418573
rect 40907 418508 40908 418572
rect 40972 418508 40973 418572
rect 40907 418507 40973 418508
rect 40539 418300 40605 418301
rect 40539 418236 40540 418300
rect 40604 418236 40605 418300
rect 40539 418235 40605 418236
rect 40542 406741 40602 418235
rect 40723 418028 40789 418029
rect 40723 417964 40724 418028
rect 40788 417964 40789 418028
rect 40723 417963 40789 417964
rect 40539 406740 40605 406741
rect 40539 406676 40540 406740
rect 40604 406676 40605 406740
rect 40539 406675 40605 406676
rect 40726 404565 40786 417963
rect 40910 407013 40970 418507
rect 41830 417757 41890 423539
rect 42011 421972 42077 421973
rect 42011 421908 42012 421972
rect 42076 421908 42077 421972
rect 42011 421907 42077 421908
rect 42014 418029 42074 421907
rect 42011 418028 42077 418029
rect 42011 417964 42012 418028
rect 42076 417964 42077 418028
rect 42011 417963 42077 417964
rect 41459 417756 41525 417757
rect 41459 417692 41460 417756
rect 41524 417692 41525 417756
rect 41459 417691 41525 417692
rect 41827 417756 41893 417757
rect 41827 417692 41828 417756
rect 41892 417692 41893 417756
rect 41827 417691 41893 417692
rect 40907 407012 40973 407013
rect 40907 406948 40908 407012
rect 40972 406948 40973 407012
rect 40907 406947 40973 406948
rect 40723 404564 40789 404565
rect 40723 404500 40724 404564
rect 40788 404500 40789 404564
rect 40723 404499 40789 404500
rect 41462 400077 41522 417691
rect 42011 415308 42077 415309
rect 42011 415244 42012 415308
rect 42076 415244 42077 415308
rect 42011 415243 42077 415244
rect 41827 414628 41893 414629
rect 41827 414564 41828 414628
rect 41892 414564 41893 414628
rect 41827 414563 41893 414564
rect 41459 400076 41525 400077
rect 41459 400012 41460 400076
rect 41524 400012 41525 400076
rect 41459 400011 41525 400012
rect 41830 399397 41890 414563
rect 41827 399396 41893 399397
rect 41827 399332 41828 399396
rect 41892 399332 41893 399396
rect 41827 399331 41893 399332
rect 42014 398853 42074 415243
rect 42011 398852 42077 398853
rect 42011 398788 42012 398852
rect 42076 398788 42077 398852
rect 42011 398787 42077 398788
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40723 378996 40789 378997
rect 40723 378932 40724 378996
rect 40788 378932 40789 378996
rect 40723 378931 40789 378932
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40542 360093 40602 378523
rect 40726 364173 40786 378931
rect 40907 377772 40973 377773
rect 40907 377708 40908 377772
rect 40972 377708 40973 377772
rect 40907 377707 40973 377708
rect 40910 364853 40970 377707
rect 40907 364852 40973 364853
rect 40907 364788 40908 364852
rect 40972 364788 40973 364852
rect 40907 364787 40973 364788
rect 40723 364172 40789 364173
rect 40723 364108 40724 364172
rect 40788 364108 40789 364172
rect 40723 364107 40789 364108
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 356965 41522 381787
rect 41643 379404 41709 379405
rect 41643 379340 41644 379404
rect 41708 379340 41709 379404
rect 41643 379339 41709 379340
rect 41646 358050 41706 379339
rect 41827 374644 41893 374645
rect 41827 374580 41828 374644
rect 41892 374580 41893 374644
rect 41827 374579 41893 374580
rect 41830 358733 41890 374579
rect 41827 358732 41893 358733
rect 41827 358668 41828 358732
rect 41892 358668 41893 358732
rect 41827 358667 41893 358668
rect 41646 357990 41890 358050
rect 41459 356964 41525 356965
rect 41459 356900 41460 356964
rect 41524 356900 41525 356964
rect 41459 356899 41525 356900
rect 41830 355741 41890 357990
rect 41827 355740 41893 355741
rect 41827 355676 41828 355740
rect 41892 355676 41893 355740
rect 41827 355675 41893 355676
rect 43299 354516 43365 354517
rect 43299 354452 43300 354516
rect 43364 354452 43365 354516
rect 43299 354451 43365 354452
rect 42747 340236 42813 340237
rect 42747 340172 42748 340236
rect 42812 340172 42813 340236
rect 42747 340171 42813 340172
rect 41643 338196 41709 338197
rect 41643 338132 41644 338196
rect 41708 338132 41709 338196
rect 41643 338131 41709 338132
rect 40539 336972 40605 336973
rect 40539 336908 40540 336972
rect 40604 336908 40605 336972
rect 40539 336907 40605 336908
rect 40542 316029 40602 336907
rect 41459 336564 41525 336565
rect 41459 336500 41460 336564
rect 41524 336500 41525 336564
rect 41459 336499 41525 336500
rect 40907 335748 40973 335749
rect 40907 335684 40908 335748
rect 40972 335684 40973 335748
rect 40907 335683 40973 335684
rect 40723 335340 40789 335341
rect 40723 335276 40724 335340
rect 40788 335276 40789 335340
rect 40723 335275 40789 335276
rect 40726 317389 40786 335275
rect 40910 321197 40970 335683
rect 40907 321196 40973 321197
rect 40907 321132 40908 321196
rect 40972 321132 40973 321196
rect 40907 321131 40973 321132
rect 40723 317388 40789 317389
rect 40723 317324 40724 317388
rect 40788 317324 40789 317388
rect 40723 317323 40789 317324
rect 40539 316028 40605 316029
rect 40539 315964 40540 316028
rect 40604 315964 40605 316028
rect 40539 315963 40605 315964
rect 41462 313717 41522 336499
rect 41646 319970 41706 338131
rect 41827 331260 41893 331261
rect 41827 331196 41828 331260
rect 41892 331196 41893 331260
rect 41827 331195 41893 331196
rect 41830 324869 41890 331195
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41827 319972 41893 319973
rect 41827 319970 41828 319972
rect 41646 319910 41828 319970
rect 41827 319908 41828 319910
rect 41892 319908 41893 319972
rect 41827 319907 41893 319908
rect 41459 313716 41525 313717
rect 41459 313652 41460 313716
rect 41524 313652 41525 313716
rect 41459 313651 41525 313652
rect 42750 299301 42810 340171
rect 42931 336836 42997 336837
rect 42931 336772 42932 336836
rect 42996 336772 42997 336836
rect 42931 336771 42997 336772
rect 42934 316437 42994 336771
rect 43302 334661 43362 354451
rect 44587 342956 44653 342957
rect 44587 342892 44588 342956
rect 44652 342892 44653 342956
rect 44587 342891 44653 342892
rect 44403 339828 44469 339829
rect 44403 339764 44404 339828
rect 44468 339764 44469 339828
rect 44403 339763 44469 339764
rect 43299 334660 43365 334661
rect 43299 334596 43300 334660
rect 43364 334596 43365 334660
rect 43299 334595 43365 334596
rect 42931 316436 42997 316437
rect 42931 316372 42932 316436
rect 42996 316372 42997 316436
rect 42931 316371 42997 316372
rect 42747 299300 42813 299301
rect 42747 299236 42748 299300
rect 42812 299236 42813 299300
rect 42747 299235 42813 299236
rect 44406 297669 44466 339763
rect 44590 300117 44650 342891
rect 44771 337380 44837 337381
rect 44771 337316 44772 337380
rect 44836 337316 44837 337380
rect 44771 337315 44837 337316
rect 44587 300116 44653 300117
rect 44587 300052 44588 300116
rect 44652 300052 44653 300116
rect 44587 300051 44653 300052
rect 44774 298485 44834 337315
rect 44771 298484 44837 298485
rect 44771 298420 44772 298484
rect 44836 298420 44837 298484
rect 44771 298419 44837 298420
rect 44403 297668 44469 297669
rect 44403 297604 44404 297668
rect 44468 297604 44469 297668
rect 44403 297603 44469 297604
rect 42195 296852 42261 296853
rect 42195 296788 42196 296852
rect 42260 296788 42261 296852
rect 42195 296787 42261 296788
rect 42011 295628 42077 295629
rect 42011 295564 42012 295628
rect 42076 295564 42077 295628
rect 42011 295563 42077 295564
rect 41827 294404 41893 294405
rect 41827 294340 41828 294404
rect 41892 294340 41893 294404
rect 41827 294339 41893 294340
rect 41830 292770 41890 294339
rect 40542 292710 41890 292770
rect 40542 269789 40602 292710
rect 40723 292592 40789 292593
rect 40723 292528 40724 292592
rect 40788 292528 40789 292592
rect 40723 292527 40789 292528
rect 40726 274277 40786 292527
rect 41827 291820 41893 291821
rect 41827 291818 41828 291820
rect 40910 291758 41828 291818
rect 40910 277133 40970 291758
rect 41827 291756 41828 291758
rect 41892 291756 41893 291820
rect 41827 291755 41893 291756
rect 41827 290052 41893 290053
rect 41827 290050 41828 290052
rect 41370 289990 41828 290050
rect 41370 289830 41430 289990
rect 41827 289988 41828 289990
rect 41892 289988 41893 290052
rect 41827 289987 41893 289988
rect 42014 289830 42074 295563
rect 42198 290053 42258 296787
rect 42195 290052 42261 290053
rect 42195 289988 42196 290052
rect 42260 289988 42261 290052
rect 42195 289987 42261 289988
rect 41370 289770 41522 289830
rect 40907 277132 40973 277133
rect 40907 277068 40908 277132
rect 40972 277068 40973 277132
rect 40907 277067 40973 277068
rect 40723 274276 40789 274277
rect 40723 274212 40724 274276
rect 40788 274212 40789 274276
rect 40723 274211 40789 274212
rect 41462 270469 41522 289770
rect 41646 289770 42074 289830
rect 41646 272370 41706 289770
rect 41827 284884 41893 284885
rect 41827 284820 41828 284884
rect 41892 284820 41893 284884
rect 41827 284819 41893 284820
rect 41830 273053 41890 284819
rect 62070 278901 62130 585651
rect 673870 455293 673930 616115
rect 674238 591293 674298 652835
rect 674422 619037 674482 694587
rect 674606 662421 674666 738107
rect 675342 730829 675402 786659
rect 675339 730828 675405 730829
rect 675339 730764 675340 730828
rect 675404 730764 675405 730828
rect 675339 730763 675405 730764
rect 676078 726613 676138 788019
rect 676811 729876 676877 729877
rect 676811 729812 676812 729876
rect 676876 729812 676877 729876
rect 676811 729811 676877 729812
rect 676075 726612 676141 726613
rect 676075 726548 676076 726612
rect 676140 726548 676141 726612
rect 676075 726547 676141 726548
rect 675155 721716 675221 721717
rect 675155 721652 675156 721716
rect 675220 721652 675221 721716
rect 675155 721651 675221 721652
rect 675158 717630 675218 721651
rect 675158 717570 675402 717630
rect 675342 683773 675402 717570
rect 675523 696828 675589 696829
rect 675523 696764 675524 696828
rect 675588 696764 675589 696828
rect 675523 696763 675589 696764
rect 675526 684045 675586 696763
rect 675523 684044 675589 684045
rect 675523 683980 675524 684044
rect 675588 683980 675589 684044
rect 675523 683979 675589 683980
rect 675339 683772 675405 683773
rect 675339 683708 675340 683772
rect 675404 683708 675405 683772
rect 675339 683707 675405 683708
rect 676075 676428 676141 676429
rect 676075 676364 676076 676428
rect 676140 676364 676141 676428
rect 676075 676363 676141 676364
rect 674603 662420 674669 662421
rect 674603 662356 674604 662420
rect 674668 662356 674669 662420
rect 674603 662355 674669 662356
rect 675523 645556 675589 645557
rect 675523 645492 675524 645556
rect 675588 645492 675589 645556
rect 675523 645491 675589 645492
rect 675526 643653 675586 645491
rect 675523 643652 675589 643653
rect 675523 643588 675524 643652
rect 675588 643588 675589 643652
rect 675523 643587 675589 643588
rect 676078 637533 676138 676363
rect 676814 665821 676874 729811
rect 676811 665820 676877 665821
rect 676811 665756 676812 665820
rect 676876 665756 676877 665820
rect 676811 665755 676877 665756
rect 676075 637532 676141 637533
rect 676075 637468 676076 637532
rect 676140 637468 676141 637532
rect 676075 637467 676141 637468
rect 675155 631412 675221 631413
rect 675155 631348 675156 631412
rect 675220 631348 675221 631412
rect 675155 631347 675221 631348
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 674419 619036 674485 619037
rect 674419 618972 674420 619036
rect 674484 618972 674485 619036
rect 674419 618971 674485 618972
rect 674419 602988 674485 602989
rect 674419 602924 674420 602988
rect 674484 602924 674485 602988
rect 674419 602923 674485 602924
rect 674235 591292 674301 591293
rect 674235 591228 674236 591292
rect 674300 591228 674301 591292
rect 674235 591227 674301 591228
rect 674422 547093 674482 602923
rect 674971 595372 675037 595373
rect 674971 595308 674972 595372
rect 675036 595308 675037 595372
rect 674971 595307 675037 595308
rect 674974 590477 675034 595307
rect 675158 593197 675218 631347
rect 675155 593196 675221 593197
rect 675155 593132 675156 593196
rect 675220 593132 675221 593196
rect 675155 593131 675221 593132
rect 676078 591701 676138 631347
rect 676811 617132 676877 617133
rect 676811 617068 676812 617132
rect 676876 617068 676877 617132
rect 676811 617067 676877 617068
rect 676075 591700 676141 591701
rect 676075 591636 676076 591700
rect 676140 591636 676141 591700
rect 676075 591635 676141 591636
rect 674971 590476 675037 590477
rect 674971 590412 674972 590476
rect 675036 590412 675037 590476
rect 674971 590411 675037 590412
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675339 561916 675405 561917
rect 675339 561852 675340 561916
rect 675404 561852 675405 561916
rect 675339 561851 675405 561852
rect 674419 547092 674485 547093
rect 674419 547028 674420 547092
rect 674484 547028 674485 547092
rect 674419 547027 674485 547028
rect 675342 545733 675402 561851
rect 676078 546821 676138 586195
rect 676814 576877 676874 617067
rect 676811 576876 676877 576877
rect 676811 576812 676812 576876
rect 676876 576812 676877 576876
rect 676811 576811 676877 576812
rect 676259 557564 676325 557565
rect 676259 557500 676260 557564
rect 676324 557500 676325 557564
rect 676259 557499 676325 557500
rect 676262 547637 676322 557499
rect 676811 553892 676877 553893
rect 676811 553828 676812 553892
rect 676876 553828 676877 553892
rect 676811 553827 676877 553828
rect 676259 547636 676325 547637
rect 676259 547572 676260 547636
rect 676324 547572 676325 547636
rect 676259 547571 676325 547572
rect 676075 546820 676141 546821
rect 676075 546756 676076 546820
rect 676140 546756 676141 546820
rect 676075 546755 676141 546756
rect 675339 545732 675405 545733
rect 675339 545668 675340 545732
rect 675404 545668 675405 545732
rect 675339 545667 675405 545668
rect 676814 500989 676874 553827
rect 676995 548316 677061 548317
rect 676995 548252 676996 548316
rect 677060 548252 677061 548316
rect 676995 548251 677061 548252
rect 676998 503709 677058 548251
rect 676995 503708 677061 503709
rect 676995 503644 676996 503708
rect 677060 503644 677061 503708
rect 676995 503643 677061 503644
rect 676811 500988 676877 500989
rect 676811 500924 676812 500988
rect 676876 500924 676877 500988
rect 676811 500923 676877 500924
rect 676029 488884 676095 488885
rect 676029 488820 676030 488884
rect 676094 488820 676095 488884
rect 676029 488819 676095 488820
rect 676032 488610 676092 488819
rect 676032 488550 677242 488610
rect 675891 487932 675957 487933
rect 675891 487868 675892 487932
rect 675956 487930 675957 487932
rect 675956 487870 676322 487930
rect 675956 487868 675957 487870
rect 675891 487867 675957 487868
rect 676262 483030 676322 487870
rect 676262 482970 676874 483030
rect 673867 455292 673933 455293
rect 673867 455228 673868 455292
rect 673932 455228 673933 455292
rect 673867 455227 673933 455228
rect 676814 400485 676874 482970
rect 677182 401301 677242 488550
rect 677179 401300 677245 401301
rect 677179 401236 677180 401300
rect 677244 401236 677245 401300
rect 677179 401235 677245 401236
rect 676811 400484 676877 400485
rect 676811 400420 676812 400484
rect 676876 400420 676877 400484
rect 676811 400419 676877 400420
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 392868 675957 392869
rect 675891 392804 675892 392868
rect 675956 392804 675957 392868
rect 675891 392803 675957 392804
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 675894 374010 675954 392803
rect 675342 373950 675954 374010
rect 675342 372469 675402 373950
rect 676078 373693 676138 398787
rect 676259 396812 676325 396813
rect 676259 396748 676260 396812
rect 676324 396748 676325 396812
rect 676259 396747 676325 396748
rect 676262 384981 676322 396747
rect 676443 396404 676509 396405
rect 676443 396340 676444 396404
rect 676508 396340 676509 396404
rect 676443 396339 676509 396340
rect 676259 384980 676325 384981
rect 676259 384916 676260 384980
rect 676324 384916 676325 384980
rect 676259 384915 676325 384916
rect 676446 382261 676506 396339
rect 676627 395180 676693 395181
rect 676627 395116 676628 395180
rect 676692 395116 676693 395180
rect 676627 395115 676693 395116
rect 676443 382260 676509 382261
rect 676443 382196 676444 382260
rect 676508 382196 676509 382260
rect 676443 382195 676509 382196
rect 676630 377365 676690 395115
rect 676627 377364 676693 377365
rect 676627 377300 676628 377364
rect 676692 377300 676693 377364
rect 676627 377299 676693 377300
rect 676075 373692 676141 373693
rect 676075 373628 676076 373692
rect 676140 373628 676141 373692
rect 676075 373627 676141 373628
rect 675339 372468 675405 372469
rect 675339 372404 675340 372468
rect 675404 372404 675405 372468
rect 675339 372403 675405 372404
rect 675342 366349 675402 372403
rect 675339 366348 675405 366349
rect 675339 366284 675340 366348
rect 675404 366284 675405 366348
rect 675339 366283 675405 366284
rect 675523 354244 675589 354245
rect 675523 354180 675524 354244
rect 675588 354180 675589 354244
rect 675523 354179 675589 354180
rect 675339 347716 675405 347717
rect 675339 347652 675340 347716
rect 675404 347652 675405 347716
rect 675339 347651 675405 347652
rect 675342 327997 675402 347651
rect 675526 339421 675586 354179
rect 675891 353836 675957 353837
rect 675891 353772 675892 353836
rect 675956 353772 675957 353836
rect 675891 353771 675957 353772
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 349210 675770 352955
rect 675894 352610 675954 353771
rect 675894 352550 676690 352610
rect 675891 351796 675957 351797
rect 675891 351732 675892 351796
rect 675956 351732 675957 351796
rect 675891 351731 675957 351732
rect 675894 349890 675954 351731
rect 675894 349830 676322 349890
rect 675710 349150 676138 349210
rect 675523 339420 675589 339421
rect 675523 339356 675524 339420
rect 675588 339356 675589 339420
rect 675523 339355 675589 339356
rect 676078 337925 676138 349150
rect 676262 340237 676322 349830
rect 676443 346628 676509 346629
rect 676443 346564 676444 346628
rect 676508 346564 676509 346628
rect 676443 346563 676509 346564
rect 676259 340236 676325 340237
rect 676259 340172 676260 340236
rect 676324 340172 676325 340236
rect 676259 340171 676325 340172
rect 676075 337924 676141 337925
rect 676075 337860 676076 337924
rect 676140 337860 676141 337924
rect 676075 337859 676141 337860
rect 676446 336565 676506 346563
rect 676443 336564 676509 336565
rect 676443 336500 676444 336564
rect 676508 336500 676509 336564
rect 676443 336499 676509 336500
rect 675339 327996 675405 327997
rect 675339 327932 675340 327996
rect 675404 327932 675405 327996
rect 675339 327931 675405 327932
rect 676630 325685 676690 352550
rect 676627 325684 676693 325685
rect 676627 325620 676628 325684
rect 676692 325620 676693 325684
rect 676627 325619 676693 325620
rect 675342 309710 675770 309770
rect 675342 309229 675402 309710
rect 675339 309228 675405 309229
rect 675339 309164 675340 309228
rect 675404 309164 675405 309228
rect 675339 309163 675405 309164
rect 675710 309090 675770 309710
rect 675710 309030 676506 309090
rect 675891 308820 675957 308821
rect 675891 308756 675892 308820
rect 675956 308756 675957 308820
rect 675891 308755 675957 308756
rect 675894 303650 675954 308755
rect 676075 304604 676141 304605
rect 676075 304540 676076 304604
rect 676140 304540 676141 304604
rect 676075 304539 676141 304540
rect 676078 304330 676138 304539
rect 676078 304270 676322 304330
rect 675894 303590 676138 303650
rect 675891 302700 675957 302701
rect 675891 302636 675892 302700
rect 675956 302636 675957 302700
rect 675891 302635 675957 302636
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 675523 296580 675589 296581
rect 675523 296516 675524 296580
rect 675588 296516 675589 296580
rect 675523 296515 675589 296516
rect 675526 292229 675586 296515
rect 675523 292228 675589 292229
rect 675523 292164 675524 292228
rect 675588 292164 675589 292228
rect 675523 292163 675589 292164
rect 675710 281621 675770 297331
rect 675894 282930 675954 302635
rect 676078 283661 676138 303590
rect 676262 287061 676322 304270
rect 676446 294677 676506 309030
rect 676627 301612 676693 301613
rect 676627 301548 676628 301612
rect 676692 301548 676693 301612
rect 676627 301547 676693 301548
rect 676443 294676 676509 294677
rect 676443 294612 676444 294676
rect 676508 294612 676509 294676
rect 676443 294611 676509 294612
rect 676630 291005 676690 301547
rect 676627 291004 676693 291005
rect 676627 290940 676628 291004
rect 676692 290940 676693 291004
rect 676627 290939 676693 290940
rect 676259 287060 676325 287061
rect 676259 286996 676260 287060
rect 676324 286996 676325 287060
rect 676259 286995 676325 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675894 282870 676138 282930
rect 676078 282709 676138 282870
rect 676075 282708 676141 282709
rect 676075 282644 676076 282708
rect 676140 282644 676141 282708
rect 676075 282643 676141 282644
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 62067 278900 62133 278901
rect 62067 278836 62068 278900
rect 62132 278836 62133 278900
rect 62067 278835 62133 278836
rect 675339 273868 675405 273869
rect 675339 273804 675340 273868
rect 675404 273804 675405 273868
rect 675339 273803 675405 273804
rect 41827 273052 41893 273053
rect 41827 272988 41828 273052
rect 41892 272988 41893 273052
rect 41827 272987 41893 272988
rect 41827 272372 41893 272373
rect 41827 272370 41828 272372
rect 41646 272310 41828 272370
rect 41827 272308 41828 272310
rect 41892 272308 41893 272372
rect 41827 272307 41893 272308
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 40539 269788 40605 269789
rect 40539 269724 40540 269788
rect 40604 269724 40605 269788
rect 40539 269723 40605 269724
rect 40539 249796 40605 249797
rect 40539 249732 40540 249796
rect 40604 249732 40605 249796
rect 40539 249731 40605 249732
rect 40542 236605 40602 249731
rect 675342 249661 675402 273803
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 261220 676877 261221
rect 676811 261156 676812 261220
rect 676876 261156 676877 261220
rect 676811 261155 676877 261156
rect 675523 258092 675589 258093
rect 675523 258028 675524 258092
rect 675588 258028 675589 258092
rect 675523 258027 675589 258028
rect 675526 250069 675586 258027
rect 675523 250068 675589 250069
rect 675523 250004 675524 250068
rect 675588 250004 675589 250068
rect 675523 250003 675589 250004
rect 675339 249660 675405 249661
rect 675339 249596 675340 249660
rect 675404 249596 675405 249660
rect 675339 249595 675405 249596
rect 40723 249388 40789 249389
rect 40723 249324 40724 249388
rect 40788 249324 40789 249388
rect 40723 249323 40789 249324
rect 40539 236604 40605 236605
rect 40539 236540 40540 236604
rect 40604 236540 40605 236604
rect 40539 236539 40605 236540
rect 40726 234701 40786 249323
rect 676814 246669 676874 261155
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 676811 246668 676877 246669
rect 676811 246604 676812 246668
rect 676876 246604 676877 246668
rect 676811 246603 676877 246604
rect 673315 246260 673381 246261
rect 673315 246196 673316 246260
rect 673380 246196 673381 246260
rect 673315 246195 673381 246196
rect 674603 246260 674669 246261
rect 674603 246196 674604 246260
rect 674668 246196 674669 246260
rect 674603 246195 674669 246196
rect 667795 245716 667861 245717
rect 667795 245652 667796 245716
rect 667860 245652 667861 245716
rect 667795 245651 667861 245652
rect 42011 238100 42077 238101
rect 42011 238036 42012 238100
rect 42076 238036 42077 238100
rect 42011 238035 42077 238036
rect 40723 234700 40789 234701
rect 40723 234636 40724 234700
rect 40788 234636 40789 234700
rect 40723 234635 40789 234636
rect 42014 227357 42074 238035
rect 42011 227356 42077 227357
rect 42011 227292 42012 227356
rect 42076 227292 42077 227356
rect 42011 227291 42077 227292
rect 649579 223004 649645 223005
rect 649579 222940 649580 223004
rect 649644 222940 649645 223004
rect 649579 222939 649645 222940
rect 651971 223004 652037 223005
rect 651971 222940 651972 223004
rect 652036 222940 652037 223004
rect 651971 222939 652037 222940
rect 649582 222818 649642 222939
rect 651974 222818 652034 222939
rect 511027 217564 511093 217565
rect 511027 217500 511028 217564
rect 511092 217500 511093 217564
rect 511027 217499 511093 217500
rect 520043 217564 520109 217565
rect 520043 217500 520044 217564
rect 520108 217500 520109 217564
rect 520043 217499 520109 217500
rect 532555 217564 532621 217565
rect 532555 217500 532556 217564
rect 532620 217500 532621 217564
rect 532555 217499 532621 217500
rect 511030 215661 511090 217499
rect 520046 215933 520106 217499
rect 520043 215932 520109 215933
rect 520043 215868 520044 215932
rect 520108 215868 520109 215932
rect 520043 215867 520109 215868
rect 511027 215660 511093 215661
rect 511027 215596 511028 215660
rect 511092 215596 511093 215660
rect 511027 215595 511093 215596
rect 532558 215389 532618 217499
rect 532555 215388 532621 215389
rect 532555 215324 532556 215388
rect 532620 215324 532621 215388
rect 532555 215323 532621 215324
rect 41827 210084 41893 210085
rect 41827 210020 41828 210084
rect 41892 210020 41893 210084
rect 41827 210019 41893 210020
rect 41643 208180 41709 208181
rect 41643 208116 41644 208180
rect 41708 208116 41709 208180
rect 41643 208115 41709 208116
rect 40539 207364 40605 207365
rect 40539 207300 40540 207364
rect 40604 207300 40605 207364
rect 40539 207299 40605 207300
rect 40542 186421 40602 207299
rect 40723 206548 40789 206549
rect 40723 206484 40724 206548
rect 40788 206484 40789 206548
rect 40723 206483 40789 206484
rect 40726 193493 40786 206483
rect 40907 206140 40973 206141
rect 40907 206076 40908 206140
rect 40972 206076 40973 206140
rect 40907 206075 40973 206076
rect 40910 194989 40970 206075
rect 41459 204916 41525 204917
rect 41459 204852 41460 204916
rect 41524 204852 41525 204916
rect 41459 204851 41525 204852
rect 41462 204101 41522 204851
rect 41459 204100 41525 204101
rect 41459 204036 41460 204100
rect 41524 204036 41525 204100
rect 41459 204035 41525 204036
rect 41646 195990 41706 208115
rect 41462 195930 41706 195990
rect 40907 194988 40973 194989
rect 40907 194924 40908 194988
rect 40972 194924 40973 194988
rect 40907 194923 40973 194924
rect 40723 193492 40789 193493
rect 40723 193428 40724 193492
rect 40788 193428 40789 193492
rect 40723 193427 40789 193428
rect 40539 186420 40605 186421
rect 40539 186356 40540 186420
rect 40604 186356 40605 186420
rect 40539 186355 40605 186356
rect 41462 186013 41522 195930
rect 41830 195261 41890 210019
rect 42011 198796 42077 198797
rect 42011 198732 42012 198796
rect 42076 198732 42077 198796
rect 42011 198731 42077 198732
rect 42014 195669 42074 198731
rect 42011 195668 42077 195669
rect 42011 195604 42012 195668
rect 42076 195604 42077 195668
rect 42011 195603 42077 195604
rect 41827 195260 41893 195261
rect 41827 195196 41828 195260
rect 41892 195196 41893 195260
rect 41827 195195 41893 195196
rect 41459 186012 41525 186013
rect 41459 185948 41460 186012
rect 41524 185948 41525 186012
rect 41459 185947 41525 185948
rect 667798 134605 667858 245651
rect 670739 231980 670805 231981
rect 670739 231916 670740 231980
rect 670804 231916 670805 231980
rect 670739 231915 670805 231916
rect 669451 223412 669517 223413
rect 669451 223348 669452 223412
rect 669516 223348 669517 223412
rect 669451 223347 669517 223348
rect 668166 179621 668226 222582
rect 669454 218925 669514 223347
rect 669451 218924 669517 218925
rect 669451 218860 669452 218924
rect 669516 218860 669517 218924
rect 669451 218859 669517 218860
rect 669635 218244 669701 218245
rect 669635 218180 669636 218244
rect 669700 218180 669701 218244
rect 669635 218179 669701 218180
rect 669451 216612 669517 216613
rect 669451 216548 669452 216612
rect 669516 216548 669517 216612
rect 669451 216547 669517 216548
rect 669267 205732 669333 205733
rect 669267 205668 669268 205732
rect 669332 205668 669333 205732
rect 669267 205667 669333 205668
rect 669270 205461 669330 205667
rect 669267 205460 669333 205461
rect 669267 205396 669268 205460
rect 669332 205396 669333 205460
rect 669267 205395 669333 205396
rect 669267 196076 669333 196077
rect 669267 196012 669268 196076
rect 669332 196012 669333 196076
rect 669267 196011 669333 196012
rect 669270 186330 669330 196011
rect 669454 191725 669514 216547
rect 669638 205733 669698 218179
rect 670371 217972 670437 217973
rect 670371 217908 670372 217972
rect 670436 217908 670437 217972
rect 670371 217907 670437 217908
rect 670374 217157 670434 217907
rect 670371 217156 670437 217157
rect 670371 217092 670372 217156
rect 670436 217092 670437 217156
rect 670371 217091 670437 217092
rect 669635 205732 669701 205733
rect 669635 205668 669636 205732
rect 669700 205668 669701 205732
rect 669635 205667 669701 205668
rect 669635 205460 669701 205461
rect 669635 205396 669636 205460
rect 669700 205396 669701 205460
rect 669635 205395 669701 205396
rect 669638 196077 669698 205395
rect 670742 198797 670802 231915
rect 672579 227084 672645 227085
rect 672579 227020 672580 227084
rect 672644 227020 672645 227084
rect 672579 227019 672645 227020
rect 672582 200837 672642 227019
rect 672579 200836 672645 200837
rect 672579 200772 672580 200836
rect 672644 200772 672645 200836
rect 672579 200771 672645 200772
rect 670739 198796 670805 198797
rect 670739 198732 670740 198796
rect 670804 198732 670805 198796
rect 670739 198731 670805 198732
rect 669635 196076 669701 196077
rect 669635 196012 669636 196076
rect 669700 196012 669701 196076
rect 669635 196011 669701 196012
rect 669451 191724 669517 191725
rect 669451 191660 669452 191724
rect 669516 191660 669517 191724
rect 669451 191659 669517 191660
rect 669270 186270 669514 186330
rect 668163 179620 668229 179621
rect 668163 179556 668164 179620
rect 668228 179556 668229 179620
rect 668163 179555 668229 179556
rect 669454 157350 669514 186270
rect 673131 181524 673197 181525
rect 673131 181460 673132 181524
rect 673196 181460 673197 181524
rect 673131 181459 673197 181460
rect 673134 161533 673194 181459
rect 673318 178125 673378 246195
rect 674051 226540 674117 226541
rect 674051 226476 674052 226540
rect 674116 226476 674117 226540
rect 674051 226475 674117 226476
rect 673315 178124 673381 178125
rect 673315 178060 673316 178124
rect 673380 178060 673381 178124
rect 673315 178059 673381 178060
rect 673131 161532 673197 161533
rect 673131 161468 673132 161532
rect 673196 161468 673197 161532
rect 673131 161467 673197 161468
rect 669270 157290 669514 157350
rect 669270 140453 669330 157290
rect 669267 140452 669333 140453
rect 669267 140388 669268 140452
rect 669332 140388 669333 140452
rect 669267 140387 669333 140388
rect 667795 134604 667861 134605
rect 667795 134540 667796 134604
rect 667860 134540 667861 134604
rect 667795 134539 667861 134540
rect 674054 115837 674114 226475
rect 674606 206957 674666 246195
rect 675523 245308 675589 245309
rect 675523 245244 675524 245308
rect 675588 245244 675589 245308
rect 675523 245243 675589 245244
rect 675526 235517 675586 245243
rect 676811 241908 676877 241909
rect 676811 241844 676812 241908
rect 676876 241844 676877 241908
rect 676811 241843 676877 241844
rect 675523 235516 675589 235517
rect 675523 235452 675524 235516
rect 675588 235452 675589 235516
rect 675523 235451 675589 235452
rect 675523 228580 675589 228581
rect 675523 228516 675524 228580
rect 675588 228516 675589 228580
rect 675523 228515 675589 228516
rect 675526 215310 675586 228515
rect 676814 220010 676874 241843
rect 676078 219950 676874 220010
rect 676078 219877 676138 219950
rect 676029 219876 676138 219877
rect 676029 219812 676030 219876
rect 676094 219814 676138 219876
rect 676094 219812 676095 219814
rect 676029 219811 676095 219812
rect 675707 218652 675773 218653
rect 675707 218588 675708 218652
rect 675772 218588 675773 218652
rect 675707 218587 675773 218588
rect 675342 215250 675586 215310
rect 675710 215310 675770 218587
rect 675891 217972 675957 217973
rect 675891 217908 675892 217972
rect 675956 217970 675957 217972
rect 675956 217910 676322 217970
rect 675956 217908 675957 217910
rect 675891 217907 675957 217908
rect 676262 217290 676322 217910
rect 676262 217230 676506 217290
rect 675894 215870 676322 215930
rect 675894 215525 675954 215870
rect 675891 215524 675957 215525
rect 675891 215460 675892 215524
rect 675956 215460 675957 215524
rect 675891 215459 675957 215460
rect 675710 215250 676138 215310
rect 674603 206956 674669 206957
rect 674603 206892 674604 206956
rect 674668 206892 674669 206956
rect 674603 206891 674669 206892
rect 675342 189141 675402 215250
rect 675891 212532 675957 212533
rect 675891 212468 675892 212532
rect 675956 212468 675957 212532
rect 675891 212467 675957 212468
rect 675894 192813 675954 212467
rect 676078 193221 676138 215250
rect 676262 194581 676322 215870
rect 676446 202741 676506 217230
rect 676627 211444 676693 211445
rect 676627 211380 676628 211444
rect 676692 211380 676693 211444
rect 676627 211379 676693 211380
rect 676443 202740 676509 202741
rect 676443 202676 676444 202740
rect 676508 202676 676509 202740
rect 676443 202675 676509 202676
rect 676630 200021 676690 211379
rect 676627 200020 676693 200021
rect 676627 199956 676628 200020
rect 676692 199956 676693 200020
rect 676627 199955 676693 199956
rect 676811 197980 676877 197981
rect 676811 197916 676812 197980
rect 676876 197916 676877 197980
rect 676811 197915 676877 197916
rect 676259 194580 676325 194581
rect 676259 194516 676260 194580
rect 676324 194516 676325 194580
rect 676259 194515 676325 194516
rect 676075 193220 676141 193221
rect 676075 193156 676076 193220
rect 676140 193156 676141 193220
rect 676075 193155 676141 193156
rect 675891 192812 675957 192813
rect 675891 192748 675892 192812
rect 675956 192748 675957 192812
rect 675891 192747 675957 192748
rect 675339 189140 675405 189141
rect 675339 189076 675340 189140
rect 675404 189076 675405 189140
rect 675339 189075 675405 189076
rect 676814 176673 676874 197915
rect 676811 176672 676877 176673
rect 676811 176608 676812 176672
rect 676876 176608 676877 176672
rect 676811 176607 676877 176608
rect 675891 172820 675957 172821
rect 675891 172756 675892 172820
rect 675956 172756 675957 172820
rect 675891 172755 675957 172756
rect 675894 172410 675954 172755
rect 675894 172350 676506 172410
rect 675891 169420 675957 169421
rect 675891 169356 675892 169420
rect 675956 169356 675957 169420
rect 675891 169355 675957 169356
rect 675894 169010 675954 169355
rect 675894 168950 676322 169010
rect 675339 167516 675405 167517
rect 675339 167452 675340 167516
rect 675404 167452 675405 167516
rect 675339 167451 675405 167452
rect 675342 147661 675402 167451
rect 676075 162756 676141 162757
rect 676075 162692 676076 162756
rect 676140 162692 676141 162756
rect 676075 162691 676141 162692
rect 676078 148477 676138 162691
rect 676262 155821 676322 168950
rect 676446 157045 676506 172350
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 157044 676509 157045
rect 676443 156980 676444 157044
rect 676508 156980 676509 157044
rect 676443 156979 676509 156980
rect 676259 155820 676325 155821
rect 676259 155756 676260 155820
rect 676324 155756 676325 155820
rect 676259 155755 676325 155756
rect 676630 151469 676690 166363
rect 676627 151468 676693 151469
rect 676627 151404 676628 151468
rect 676692 151404 676693 151468
rect 676627 151403 676693 151404
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675339 147660 675405 147661
rect 675339 147596 675340 147660
rect 675404 147596 675405 147660
rect 675339 147595 675405 147596
rect 676811 127396 676877 127397
rect 676811 127332 676812 127396
rect 676876 127332 676877 127396
rect 676811 127331 676877 127332
rect 676075 126988 676141 126989
rect 676075 126924 676076 126988
rect 676140 126924 676141 126988
rect 676075 126923 676141 126924
rect 675339 122092 675405 122093
rect 675339 122028 675340 122092
rect 675404 122028 675405 122092
rect 675339 122027 675405 122028
rect 674051 115836 674117 115837
rect 674051 115772 674052 115836
rect 674116 115772 674117 115836
rect 674051 115771 674117 115772
rect 675342 101965 675402 122027
rect 675707 117332 675773 117333
rect 675707 117268 675708 117332
rect 675772 117268 675773 117332
rect 675707 117267 675773 117268
rect 675710 111349 675770 117267
rect 675707 111348 675773 111349
rect 675707 111284 675708 111348
rect 675772 111284 675773 111348
rect 675707 111283 675773 111284
rect 676078 108221 676138 126923
rect 676259 125764 676325 125765
rect 676259 125700 676260 125764
rect 676324 125700 676325 125764
rect 676259 125699 676325 125700
rect 676262 123450 676322 125699
rect 676443 124132 676509 124133
rect 676443 124068 676444 124132
rect 676508 124068 676509 124132
rect 676443 124067 676509 124068
rect 676627 124132 676693 124133
rect 676627 124068 676628 124132
rect 676692 124068 676693 124132
rect 676627 124067 676693 124068
rect 676446 123725 676506 124067
rect 676443 123724 676509 123725
rect 676443 123660 676444 123724
rect 676508 123660 676509 123724
rect 676443 123659 676509 123660
rect 676262 123390 676506 123450
rect 676259 122908 676325 122909
rect 676259 122844 676260 122908
rect 676324 122844 676325 122908
rect 676259 122843 676325 122844
rect 676262 112437 676322 122843
rect 676259 112436 676325 112437
rect 676259 112372 676260 112436
rect 676324 112372 676325 112436
rect 676259 112371 676325 112372
rect 676446 111757 676506 123390
rect 676443 111756 676509 111757
rect 676443 111692 676444 111756
rect 676508 111692 676509 111756
rect 676443 111691 676509 111692
rect 676630 110397 676690 124067
rect 676814 122909 676874 127331
rect 676811 122908 676877 122909
rect 676811 122844 676812 122908
rect 676876 122844 676877 122908
rect 676811 122843 676877 122844
rect 676627 110396 676693 110397
rect 676627 110332 676628 110396
rect 676692 110332 676693 110396
rect 676627 110331 676693 110332
rect 676075 108220 676141 108221
rect 676075 108156 676076 108220
rect 676140 108156 676141 108220
rect 676075 108155 676141 108156
rect 675339 101964 675405 101965
rect 675339 101900 675340 101964
rect 675404 101900 675405 101964
rect 675339 101899 675405 101900
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 633939 95436 634005 95437
rect 633939 95372 633940 95436
rect 634004 95372 634005 95436
rect 633939 95371 634005 95372
rect 633942 78573 634002 95371
rect 637254 84210 637314 96867
rect 647187 96524 647253 96525
rect 647187 96460 647188 96524
rect 647252 96460 647253 96524
rect 647187 96459 647253 96460
rect 647190 94298 647250 96459
rect 650318 93125 650378 93382
rect 650315 93124 650381 93125
rect 650315 93060 650316 93124
rect 650380 93060 650381 93124
rect 650315 93059 650381 93060
rect 637070 84150 637314 84210
rect 633939 78572 634005 78573
rect 633939 78508 633940 78572
rect 634004 78508 634005 78572
rect 633939 78507 634005 78508
rect 637070 78165 637130 84150
rect 637067 78164 637133 78165
rect 637067 78100 637068 78164
rect 637132 78100 637133 78164
rect 637067 78099 637133 78100
rect 460795 55044 460861 55045
rect 460795 54980 460796 55044
rect 460860 54980 460861 55044
rect 460795 54979 460861 54980
rect 460798 53957 460858 54979
rect 462635 54772 462701 54773
rect 462635 54708 462636 54772
rect 462700 54708 462701 54772
rect 462635 54707 462701 54708
rect 460795 53956 460861 53957
rect 460795 53892 460796 53956
rect 460860 53892 460861 53956
rect 460795 53891 460861 53892
rect 462638 53685 462698 54707
rect 462635 53684 462701 53685
rect 462635 53620 462636 53684
rect 462700 53620 462701 53684
rect 462635 53619 462701 53620
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47836 515509 47837
rect 515443 47772 515444 47836
rect 515508 47772 515509 47836
rect 515443 47771 515509 47772
rect 460979 44436 461045 44437
rect 460979 44372 460980 44436
rect 461044 44372 461045 44436
rect 460979 44371 461045 44372
rect 462267 44436 462333 44437
rect 462267 44372 462268 44436
rect 462332 44372 462333 44436
rect 462267 44371 462333 44372
rect 463739 44436 463805 44437
rect 463739 44372 463740 44436
rect 463804 44372 463805 44436
rect 463739 44371 463805 44372
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40357 141802 43963
rect 419211 42124 419277 42125
rect 419211 42060 419212 42124
rect 419276 42060 419277 42124
rect 419211 42059 419277 42060
rect 419214 41938 419274 42059
rect 416635 41852 416701 41853
rect 416635 41788 416636 41852
rect 416700 41788 416701 41852
rect 416635 41787 416701 41788
rect 416638 40578 416698 41787
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 451963 41852 452029 41853
rect 451963 41788 451964 41852
rect 452028 41788 452029 41852
rect 451963 41787 452029 41788
rect 451966 41258 452026 41787
rect 458958 41170 459018 41702
rect 458958 41110 460342 41170
rect 460982 40578 461042 44371
rect 462270 41258 462330 44371
rect 463742 41938 463802 44371
rect 515446 42125 515506 47771
rect 518758 42805 518818 48859
rect 529611 48108 529677 48109
rect 529611 48044 529612 48108
rect 529676 48044 529677 48108
rect 529611 48043 529677 48044
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 47771
rect 529614 42125 529674 48043
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529611 42124 529677 42125
rect 529611 42060 529612 42124
rect 529676 42060 529677 42124
rect 529611 42059 529677 42060
rect 141739 40356 141805 40357
rect 141739 40292 141740 40356
rect 141804 40292 141805 40356
rect 141739 40291 141805 40292
<< via4 >>
rect 591902 223412 592138 223498
rect 591902 223348 591988 223412
rect 591988 223348 592052 223412
rect 592052 223348 592138 223412
rect 591902 223262 592138 223348
rect 649494 222582 649730 222818
rect 651886 222582 652122 222818
rect 668078 222582 668314 222818
rect 647102 94062 647338 94298
rect 650230 93382 650466 93618
rect 365030 41852 365266 41938
rect 365030 41788 365116 41852
rect 365116 41788 365180 41852
rect 365180 41788 365266 41852
rect 365030 41702 365266 41788
rect 419126 41702 419362 41938
rect 419862 41852 420098 41938
rect 419862 41788 419948 41852
rect 419948 41788 420012 41852
rect 420012 41788 420098 41852
rect 419862 41702 420098 41788
rect 425014 41852 425250 41938
rect 425014 41788 425100 41852
rect 425100 41788 425164 41852
rect 425164 41788 425250 41852
rect 425014 41702 425250 41788
rect 441390 41702 441626 41938
rect 458870 41702 459106 41938
rect 451878 41022 452114 41258
rect 460342 41022 460578 41258
rect 463654 41702 463890 41938
rect 462182 41022 462418 41258
rect 416550 40342 416786 40578
rect 460894 40342 461130 40578
<< metal5 >>
rect 78610 1018624 90778 1030789
rect 130010 1018624 142178 1030789
rect 181410 1018624 193578 1030789
rect 231810 1018624 243978 1030789
rect 284410 1018624 296578 1030789
rect 334810 1018624 346978 1030789
rect 386210 1018624 398378 1030789
rect 475210 1018624 487378 1030789
rect 526610 1018624 538778 1030789
rect 577010 1018624 589178 1030789
rect 628410 1018624 640578 1030789
rect 6811 956610 18976 968778
rect 698624 953022 710789 965190
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 591860 223498 592180 223540
rect 591860 223262 591902 223498
rect 592138 223262 592180 223498
rect 591860 222860 592180 223262
rect 591860 222818 649772 222860
rect 591860 222582 649494 222818
rect 649730 222582 649772 222818
rect 591860 222540 649772 222582
rect 651844 222818 668356 222860
rect 651844 222582 651886 222818
rect 652122 222582 668078 222818
rect 668314 222582 668356 222818
rect 651844 222540 668356 222582
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 647060 94298 647748 94340
rect 647060 94062 647102 94298
rect 647338 94062 647748 94298
rect 647060 94020 647748 94062
rect 647428 93660 647748 94020
rect 647428 93618 650508 93660
rect 647428 93382 650230 93618
rect 650466 93382 650508 93618
rect 647428 93340 650508 93382
rect 6167 70054 19620 80934
rect 364988 41938 419404 41980
rect 364988 41702 365030 41938
rect 365266 41702 419126 41938
rect 419362 41702 419404 41938
rect 364988 41660 419404 41702
rect 419820 41938 424556 41980
rect 419820 41702 419862 41938
rect 420098 41702 424556 41938
rect 419820 41660 424556 41702
rect 424972 41938 441668 41980
rect 424972 41702 425014 41938
rect 425250 41702 441390 41938
rect 441626 41702 441668 41938
rect 424972 41660 441668 41702
rect 442084 41660 450684 41980
rect 424236 41300 424556 41660
rect 442084 41300 442404 41660
rect 424236 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41938 459148 41980
rect 451100 41702 458870 41938
rect 459106 41702 459148 41938
rect 451100 41660 459148 41702
rect 459564 41938 463932 41980
rect 459564 41702 463654 41938
rect 463890 41702 463932 41938
rect 459564 41660 463932 41702
rect 451100 41300 451420 41660
rect 459564 41300 459884 41660
rect 450364 40980 451420 41300
rect 451836 41258 459884 41300
rect 451836 41022 451878 41258
rect 452114 41022 459884 41258
rect 451836 40980 459884 41022
rect 460300 41258 462460 41300
rect 460300 41022 460342 41258
rect 460578 41022 462182 41258
rect 462418 41022 462460 41258
rect 460300 40980 462460 41022
rect 416508 40578 461172 40620
rect 416508 40342 416550 40578
rect 416786 40342 460894 40578
rect 461130 40342 461172 40578
rect 416508 40300 461172 40342
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravan_logo  caravan_logo
timestamp 0
transform 1 0 255300 0 1 6032
box 0 0 1 1
use caravan_motto  caravan_motto
timestamp 0
transform 1 0 -54560 0 1 -52
box 0 0 1 1
use copyright_block_a  copyright_block_a
timestamp 0
transform 1 0 149582 0 1 16298
box 0 0 1 1
use open_source  open_source
timestamp 0
transform 1 0 206074 0 1 2336
box 0 0 1 1
use xres_buf  rstb_level
timestamp 1666265755
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 96272 0 1 6890
box 0 0 1 1
use caravel_clocking  clock_ctrl
timestamp 1666265755
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1666265755
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1666265755
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1666265755
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1666265755
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use digital_pll  pll
timestamp 1666265755
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por
timestamp 1666265755
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use user_id_programming  user_id_value
timestamp 1666265755
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1666265755
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666265755
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1666265755
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666265755
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666265755
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1666265755
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1666265755
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use spare_logic_block  spare_logic\[2\]
timestamp 1666265755
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666265755
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666265755
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1666265755
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use mgmt_protect  mgmt_buffers
timestamp 1666265755
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1666265755
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1666265755
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1666265755
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666265755
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1666265755
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666265755
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1666265755
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1666265755
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666265755
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666265755
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666265755
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1666265755
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1666265755
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1666265755
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666265755
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666265755
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666265755
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1666265755
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1666265755
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1666265755
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1666265755
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1666265755
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666265755
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666265755
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666265755
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666265755
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666265755
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666265755
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1666265755
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1666265755
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1666265755
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1666265755
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1666265755
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1666265755
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666265755
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666265755
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666265755
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666265755
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666265755
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1666265755
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1666265755
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1666265755
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1666265755
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666265755
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666265755
transform -1 0 710203 0 1 884800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1666265755
transform -1 0 709467 0 1 897800
box -38 0 6018 2224
use caravan_power_routing  caravan_power_routing
timestamp 1666265755
transform 1 0 0 0 1 0
box 6022 30806 711814 997678
use user_analog_project_wrapper  mprj
timestamp 1666265755
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use chip_io_alt  padframe
timestamp 1666265755
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use gpio_signal_buffering_alt  sigbuf
timestamp 1666265755
transform 1 0 0 0 1 0
box 40023 41960 677583 728321
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698624 953022 710789 965190 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030789 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526610 1018624 538778 1030789 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475210 1018624 487378 1030789 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386210 1018624 398378 1030789 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284410 1018624 296578 1030789 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 231810 1018624 243978 1030789 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181410 1018624 193578 1030789 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 130010 1018624 142178 1030789 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78610 1018624 90778 1030789 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6811 956610 18976 968778 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
