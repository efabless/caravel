magic
tech sky130A
timestamp 1637698689
<< fillblock >>
rect 183980 5102 199901 7384
use font_44  font_44_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763661
transform 1 0 184889 0 1 5633
box 0 0 540 1260
use font_22  font_22_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598785768
transform 1 0 184172 0 1 5938
box 0 540 540 1260
use font_72  font_72_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777237
transform 1 0 185611 0 1 5635
box 0 0 540 900
use font_69  font_69_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776260
transform 1 0 186331 0 1 5631
box 0 0 360 1260
use font_76  font_76_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777472
transform 1 0 186868 0 1 5640
box 0 0 540 900
use font_69  font_69_1
timestamp 1598776260
transform 1 0 187580 0 1 5644
box 0 0 360 1260
use font_67  font_67_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776042
transform 1 0 188833 0 1 5635
box 0 -360 540 900
use font_6E  font_6E_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776997
transform 1 0 188118 0 1 5635
box 0 0 540 900
use font_54  font_54_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768910
transform 1 0 190053 0 1 5644
box 0 0 540 1260
use font_68  font_68_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776130
transform 1 0 190781 0 1 5652
box 0 0 540 1260
use font_65  font_65_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775915
transform 1 0 191497 0 1 5652
box 0 0 540 900
use font_4F  font_4F_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598767855
transform 1 0 192784 0 1 5648
box 0 0 540 1260
use font_70  font_70_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777090
transform 1 0 193504 0 1 5652
box 0 -360 540 900
use font_65  font_65_1
timestamp 1598775915
transform 1 0 194228 0 1 5657
box 0 0 540 900
use font_6E  font_6E_1
timestamp 1598776997
transform 1 0 194952 0 1 5661
box 0 0 540 900
use font_52  font_52_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768719
transform 1 0 196295 0 1 5661
box 0 0 540 1260
use font_6F  font_6F_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777049
transform 1 0 197019 0 1 5661
box 0 0 540 900
use font_61  font_61_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775307
transform 1 0 197747 0 1 5665
box 0 0 540 900
use font_64  font_64_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775833
transform 1 0 198463 0 1 5665
box 0 0 540 1260
use font_22  font_22_1
timestamp 1598785768
transform 1 0 199183 0 1 5961
box 0 540 540 1260
<< end >>
