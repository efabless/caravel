magic
tech sky130A
magscale 1 2
timestamp 1638662846
<< nwell >>
rect -38 10053 18898 10619
rect -38 8965 18898 9531
rect -38 7877 18898 8443
rect -38 6789 18898 7355
rect -38 5701 18898 6267
rect -38 4613 18898 5179
rect -38 3525 18898 4091
rect -38 2437 18898 3003
rect -38 1349 18898 1915
rect -38 261 18898 827
<< pwell >>
rect 29 -17 63 17
rect 305 -17 339 17
rect 1043 -10 1075 12
rect 1317 -17 1351 17
rect 2513 -17 2547 17
rect 3709 -17 3743 17
rect 4905 -17 4939 17
rect 5272 -11 5296 11
rect 5917 -17 5951 17
rect 6100 -17 6134 17
rect 6377 -17 6411 17
rect 7112 -11 7136 11
rect 7297 -17 7331 17
rect 8493 -17 8527 17
rect 9044 -11 9068 11
rect 9412 -17 9446 17
rect 9504 -11 9528 11
rect 9689 -17 9723 17
rect 10885 -17 10919 17
rect 12356 -17 12390 17
rect 12449 -17 12483 17
rect 13460 -17 13494 17
rect 13554 -17 13588 17
rect 13829 -17 13863 17
rect 14473 -17 14507 17
rect 15761 -17 15795 17
rect 15852 -17 15886 17
rect 16497 -17 16531 17
rect 16591 -10 16623 12
rect 16865 -17 16899 17
rect 17509 -17 17543 17
rect 17876 -11 17900 11
rect 18061 -17 18095 17
rect 18797 -17 18831 17
<< obsli1 >>
rect 0 -17 18860 10897
<< obsm1 >>
rect 0 -48 18860 10928
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
<< obsm2 >>
rect 296 11144 1342 11257
rect 1510 11144 4194 11257
rect 4362 11144 7046 11257
rect 7214 11144 9898 11257
rect 10066 11144 12750 11257
rect 12918 11144 15602 11257
rect 15770 11144 18454 11257
rect 18622 11144 18842 11257
rect 296 0 18842 11144
rect 4660 -48 4968 0
rect 7760 -48 8068 0
rect 10860 -48 11168 0
rect 13960 -48 14268 0
rect 17060 -48 17368 0
<< metal3 >>
rect 19200 11160 20000 11280
rect 19200 9664 20000 9784
rect 19200 8168 20000 8288
rect 19200 6672 20000 6792
rect 19200 5176 20000 5296
rect 19200 3680 20000 3800
rect 19200 2184 20000 2304
rect 19200 688 20000 808
<< obsm3 >>
rect 2497 11080 19120 11253
rect 2497 9864 19200 11080
rect 2497 9584 19120 9864
rect 2497 8368 19200 9584
rect 2497 8088 19120 8368
rect 2497 6872 19200 8088
rect 2497 6592 19120 6872
rect 2497 5376 19200 6592
rect 2497 5096 19120 5376
rect 2497 3880 19200 5096
rect 2497 3600 19120 3880
rect 2497 2384 19200 3600
rect 2497 2104 19120 2384
rect 2497 888 19200 2104
rect 2497 608 19120 888
rect 2497 0 19200 608
rect 4654 -33 4974 0
rect 7754 -33 8074 0
rect 10854 -33 11174 0
rect 13954 -33 14274 0
rect 17054 -33 17374 0
<< metal4 >>
rect 3104 -48 3424 10928
rect 4654 -48 4974 10928
rect 6204 -48 6524 10928
rect 7754 -48 8074 10928
rect 9304 -48 9624 10928
rect 10854 -48 11174 10928
rect 12404 -48 12724 10928
rect 13954 -48 14274 10928
rect 15504 -48 15824 10928
rect 17054 -48 17374 10928
<< metal5 >>
rect 0 9882 18860 10202
rect 0 8192 18860 8512
rect 0 6502 18860 6822
rect 0 4812 18860 5132
rect 0 3122 18860 3442
<< labels >>
rlabel metal5 s 0 4812 18860 5132 6 VGND
port 1 nsew ground input
rlabel metal5 s 0 8192 18860 8512 6 VGND
port 1 nsew ground input
rlabel metal4 s 4654 -48 4974 10928 6 VGND
port 1 nsew ground input
rlabel metal4 s 7754 -48 8074 10928 6 VGND
port 1 nsew ground input
rlabel metal4 s 10854 -48 11174 10928 6 VGND
port 1 nsew ground input
rlabel metal4 s 13954 -48 14274 10928 6 VGND
port 1 nsew ground input
rlabel metal4 s 17054 -48 17374 10928 6 VGND
port 1 nsew ground input
rlabel metal5 s 0 3122 18860 3442 6 VPWR
port 2 nsew power input
rlabel metal5 s 0 6502 18860 6822 6 VPWR
port 2 nsew power input
rlabel metal5 s 0 9882 18860 10202 6 VPWR
port 2 nsew power input
rlabel metal4 s 3104 -48 3424 10928 6 VPWR
port 2 nsew power input
rlabel metal4 s 6204 -48 6524 10928 6 VPWR
port 2 nsew power input
rlabel metal4 s 9304 -48 9624 10928 6 VPWR
port 2 nsew power input
rlabel metal4 s 12404 -48 12724 10928 6 VPWR
port 2 nsew power input
rlabel metal4 s 15504 -48 15824 10928 6 VPWR
port 2 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 3 nsew signal output
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 4 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 5 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 6 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 7 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 8 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 9 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 10 nsew signal output
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 11 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 12 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 13 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 14 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 15 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 16 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 17 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 20000 12000
string LEFview TRUE
string GDS_FILE ../gds/caravel_clocking.gds
string GDS_END 1197054
string GDS_START 422960
<< end >>

