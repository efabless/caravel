VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_power_routing
  CLASS BLOCK ;
  FOREIGN caravel_power_routing ;
  ORIGIN 0.000 -69.495 ;
  SIZE 3588.000 BY 5118.505 ;
  PIN vccd_core
    PORT
      LAYER met3 ;
        RECT 197.280 390.755 229.220 413.720 ;
        RECT 197.280 341.280 229.220 364.500 ;
      LAYER via3 ;
        RECT 209.885 391.210 228.205 413.530 ;
        RECT 209.765 341.690 228.085 364.010 ;
      LAYER met4 ;
        RECT 220.930 1152.330 315.800 1167.330 ;
        RECT 448.500 1152.330 450.780 1170.320 ;
        RECT 468.500 1152.330 470.780 1170.320 ;
        RECT 548.500 1152.330 550.780 1170.320 ;
        RECT 568.500 1152.330 570.780 1170.320 ;
        RECT 665.300 1152.330 667.580 1167.320 ;
        RECT 740.550 1152.330 742.830 1167.320 ;
        RECT 815.800 1152.330 818.080 1167.320 ;
        RECT 891.050 1152.330 893.330 1167.320 ;
        RECT 966.300 1152.330 968.580 1167.320 ;
        RECT 1041.550 1152.330 1043.830 1167.320 ;
        RECT 1116.800 1152.330 1119.080 1167.320 ;
        RECT 1192.050 1152.330 1194.330 1167.320 ;
        RECT 1267.300 1152.330 1269.580 1167.320 ;
        RECT 1342.550 1152.330 1344.830 1167.320 ;
        RECT 1417.800 1152.330 1420.080 1167.320 ;
        RECT 1493.050 1152.330 1495.330 1167.320 ;
        RECT 1568.300 1152.330 1570.580 1167.320 ;
        RECT 1643.550 1152.330 1645.830 1167.320 ;
        RECT 1718.800 1152.330 1721.080 1167.320 ;
        RECT 1794.050 1152.330 1796.330 1167.320 ;
        RECT 1869.300 1152.330 1871.580 1167.320 ;
        RECT 1944.550 1152.330 1946.830 1167.320 ;
        RECT 2019.800 1152.330 2022.080 1167.320 ;
        RECT 2095.050 1152.330 2097.330 1167.320 ;
        RECT 2170.300 1152.330 2172.580 1167.320 ;
        RECT 2245.550 1152.330 2247.830 1167.320 ;
        RECT 2320.800 1152.330 2323.080 1167.320 ;
        RECT 2396.050 1152.330 2398.330 1167.320 ;
        RECT 2471.300 1152.330 2473.580 1167.320 ;
        RECT 2546.550 1152.330 2548.830 1167.320 ;
        RECT 2621.800 1152.330 2624.080 1167.320 ;
        RECT 2696.800 1152.330 2699.080 1167.320 ;
        RECT 2898.600 1152.330 2900.880 1170.320 ;
        RECT 2918.600 1152.330 2920.880 1170.320 ;
        RECT 220.990 1046.990 233.990 1152.330 ;
        RECT 2921.840 1047.520 2984.810 1062.520 ;
        RECT 3135.220 1047.640 3140.540 1062.300 ;
        RECT 3212.020 1047.640 3217.340 1062.300 ;
        RECT 3288.820 1047.640 3294.140 1062.300 ;
        RECT 220.990 1043.790 257.600 1046.990 ;
        RECT 220.990 996.990 233.990 1043.790 ;
        RECT 2983.210 1038.460 2984.810 1047.520 ;
        RECT 3136.810 1038.420 3138.410 1047.640 ;
        RECT 3213.610 1038.420 3215.210 1047.640 ;
        RECT 3290.410 1038.420 3292.010 1047.640 ;
        RECT 2922.480 997.300 2935.870 999.040 ;
        RECT 220.990 993.790 257.600 996.990 ;
        RECT 2922.480 995.700 2964.880 997.300 ;
        RECT 2922.480 994.620 2935.870 995.700 ;
        RECT 220.990 946.990 233.990 993.790 ;
        RECT 220.990 943.790 257.600 946.990 ;
        RECT 220.990 896.990 233.990 943.790 ;
        RECT 2922.480 919.100 2935.870 920.840 ;
        RECT 2922.480 917.500 2964.880 919.100 ;
        RECT 2922.480 916.420 2935.870 917.500 ;
        RECT 220.990 893.790 257.600 896.990 ;
        RECT 220.990 883.710 233.990 893.790 ;
        RECT 209.320 865.630 233.990 883.710 ;
        RECT 208.840 843.790 257.600 846.990 ;
        RECT 2922.480 840.900 2935.870 842.640 ;
        RECT 2922.480 839.300 2964.880 840.900 ;
        RECT 2922.480 838.220 2935.870 839.300 ;
        RECT 208.840 793.790 257.600 796.990 ;
        RECT 2922.480 762.700 2935.870 764.440 ;
        RECT 2922.480 761.100 2964.880 762.700 ;
        RECT 2922.480 760.020 2935.870 761.100 ;
        RECT 208.840 743.790 257.600 746.990 ;
        RECT 208.840 693.790 257.600 696.990 ;
        RECT 2922.480 684.500 2935.870 686.240 ;
        RECT 2922.480 682.900 2964.880 684.500 ;
        RECT 2922.480 681.820 2935.870 682.900 ;
        RECT 208.840 643.790 257.600 646.990 ;
        RECT 2922.480 600.300 2935.870 602.040 ;
        RECT 2959.660 600.300 2965.060 606.530 ;
        RECT 2922.480 598.700 2965.060 600.300 ;
        RECT 2922.480 597.620 2935.870 598.700 ;
        RECT 208.840 593.790 257.600 596.990 ;
        RECT 208.840 543.790 257.600 546.990 ;
        RECT 2922.480 528.100 2935.870 529.840 ;
        RECT 2922.480 526.500 2964.880 528.100 ;
        RECT 2922.480 525.420 2935.870 526.500 ;
        RECT 208.840 493.790 257.600 496.990 ;
        RECT 208.840 443.790 257.600 446.990 ;
        RECT 209.320 396.990 228.890 413.970 ;
        RECT 3161.770 404.620 3163.370 410.310 ;
        RECT 3201.770 405.080 3203.370 410.000 ;
        RECT 208.840 393.790 257.600 396.990 ;
        RECT 209.320 390.770 228.890 393.790 ;
        RECT 3160.360 390.990 3165.050 404.620 ;
        RECT 3200.490 390.670 3204.610 405.080 ;
        RECT 3149.340 370.520 3150.940 386.870 ;
        RECT 3164.840 370.520 3166.440 386.870 ;
        RECT 3180.340 370.520 3181.940 386.870 ;
        RECT 3195.840 370.520 3197.440 386.870 ;
        RECT 3211.340 370.520 3212.940 386.870 ;
        RECT 209.290 346.990 228.860 364.450 ;
        RECT 208.840 343.790 257.600 346.990 ;
        RECT 209.290 341.250 228.860 343.790 ;
        RECT 3149.340 302.550 3150.940 318.900 ;
        RECT 3164.840 302.550 3166.440 318.900 ;
        RECT 3180.340 302.550 3181.940 318.900 ;
        RECT 3195.840 302.550 3197.440 318.900 ;
        RECT 3211.340 302.550 3212.940 318.900 ;
        RECT 208.840 293.790 257.600 296.990 ;
        RECT 209.370 241.110 292.680 260.610 ;
        RECT 716.620 249.680 723.690 253.440 ;
        RECT 719.300 248.190 720.200 249.680 ;
        RECT 3306.350 234.955 3347.130 236.600 ;
      LAYER via4 ;
        RECT 282.770 1153.675 314.350 1166.055 ;
        RECT 448.900 1165.630 450.080 1166.810 ;
        RECT 448.900 1164.030 450.080 1165.210 ;
        RECT 448.900 1162.430 450.080 1163.610 ;
        RECT 448.900 1160.830 450.080 1162.010 ;
        RECT 448.900 1159.230 450.080 1160.410 ;
        RECT 448.900 1157.630 450.080 1158.810 ;
        RECT 448.900 1156.030 450.080 1157.210 ;
        RECT 448.900 1154.430 450.080 1155.610 ;
        RECT 448.900 1152.830 450.080 1154.010 ;
        RECT 468.900 1165.630 470.080 1166.810 ;
        RECT 468.900 1164.030 470.080 1165.210 ;
        RECT 468.900 1162.430 470.080 1163.610 ;
        RECT 468.900 1160.830 470.080 1162.010 ;
        RECT 468.900 1159.230 470.080 1160.410 ;
        RECT 468.900 1157.630 470.080 1158.810 ;
        RECT 468.900 1156.030 470.080 1157.210 ;
        RECT 468.900 1154.430 470.080 1155.610 ;
        RECT 468.900 1152.830 470.080 1154.010 ;
        RECT 548.900 1165.630 550.080 1166.810 ;
        RECT 548.900 1164.030 550.080 1165.210 ;
        RECT 548.900 1162.430 550.080 1163.610 ;
        RECT 548.900 1160.830 550.080 1162.010 ;
        RECT 548.900 1159.230 550.080 1160.410 ;
        RECT 548.900 1157.630 550.080 1158.810 ;
        RECT 548.900 1156.030 550.080 1157.210 ;
        RECT 548.900 1154.430 550.080 1155.610 ;
        RECT 548.900 1152.830 550.080 1154.010 ;
        RECT 568.900 1165.630 570.080 1166.810 ;
        RECT 568.900 1164.030 570.080 1165.210 ;
        RECT 568.900 1162.430 570.080 1163.610 ;
        RECT 568.900 1160.830 570.080 1162.010 ;
        RECT 568.900 1159.230 570.080 1160.410 ;
        RECT 568.900 1157.630 570.080 1158.810 ;
        RECT 568.900 1156.030 570.080 1157.210 ;
        RECT 568.900 1154.430 570.080 1155.610 ;
        RECT 568.900 1152.830 570.080 1154.010 ;
        RECT 665.700 1165.630 666.880 1166.810 ;
        RECT 665.700 1164.030 666.880 1165.210 ;
        RECT 665.700 1162.430 666.880 1163.610 ;
        RECT 665.700 1160.830 666.880 1162.010 ;
        RECT 665.700 1159.230 666.880 1160.410 ;
        RECT 665.700 1157.630 666.880 1158.810 ;
        RECT 665.700 1156.030 666.880 1157.210 ;
        RECT 665.700 1154.430 666.880 1155.610 ;
        RECT 665.700 1152.830 666.880 1154.010 ;
        RECT 740.950 1165.630 742.130 1166.810 ;
        RECT 740.950 1164.030 742.130 1165.210 ;
        RECT 740.950 1162.430 742.130 1163.610 ;
        RECT 740.950 1160.830 742.130 1162.010 ;
        RECT 740.950 1159.230 742.130 1160.410 ;
        RECT 740.950 1157.630 742.130 1158.810 ;
        RECT 740.950 1156.030 742.130 1157.210 ;
        RECT 740.950 1154.430 742.130 1155.610 ;
        RECT 740.950 1152.830 742.130 1154.010 ;
        RECT 816.200 1165.630 817.380 1166.810 ;
        RECT 816.200 1164.030 817.380 1165.210 ;
        RECT 816.200 1162.430 817.380 1163.610 ;
        RECT 816.200 1160.830 817.380 1162.010 ;
        RECT 816.200 1159.230 817.380 1160.410 ;
        RECT 816.200 1157.630 817.380 1158.810 ;
        RECT 816.200 1156.030 817.380 1157.210 ;
        RECT 816.200 1154.430 817.380 1155.610 ;
        RECT 816.200 1152.830 817.380 1154.010 ;
        RECT 891.450 1165.630 892.630 1166.810 ;
        RECT 891.450 1164.030 892.630 1165.210 ;
        RECT 891.450 1162.430 892.630 1163.610 ;
        RECT 891.450 1160.830 892.630 1162.010 ;
        RECT 891.450 1159.230 892.630 1160.410 ;
        RECT 891.450 1157.630 892.630 1158.810 ;
        RECT 891.450 1156.030 892.630 1157.210 ;
        RECT 891.450 1154.430 892.630 1155.610 ;
        RECT 891.450 1152.830 892.630 1154.010 ;
        RECT 966.700 1165.630 967.880 1166.810 ;
        RECT 966.700 1164.030 967.880 1165.210 ;
        RECT 966.700 1162.430 967.880 1163.610 ;
        RECT 966.700 1160.830 967.880 1162.010 ;
        RECT 966.700 1159.230 967.880 1160.410 ;
        RECT 966.700 1157.630 967.880 1158.810 ;
        RECT 966.700 1156.030 967.880 1157.210 ;
        RECT 966.700 1154.430 967.880 1155.610 ;
        RECT 966.700 1152.830 967.880 1154.010 ;
        RECT 1041.950 1165.630 1043.130 1166.810 ;
        RECT 1041.950 1164.030 1043.130 1165.210 ;
        RECT 1041.950 1162.430 1043.130 1163.610 ;
        RECT 1041.950 1160.830 1043.130 1162.010 ;
        RECT 1041.950 1159.230 1043.130 1160.410 ;
        RECT 1041.950 1157.630 1043.130 1158.810 ;
        RECT 1041.950 1156.030 1043.130 1157.210 ;
        RECT 1041.950 1154.430 1043.130 1155.610 ;
        RECT 1041.950 1152.830 1043.130 1154.010 ;
        RECT 1117.200 1165.630 1118.380 1166.810 ;
        RECT 1117.200 1164.030 1118.380 1165.210 ;
        RECT 1117.200 1162.430 1118.380 1163.610 ;
        RECT 1117.200 1160.830 1118.380 1162.010 ;
        RECT 1117.200 1159.230 1118.380 1160.410 ;
        RECT 1117.200 1157.630 1118.380 1158.810 ;
        RECT 1117.200 1156.030 1118.380 1157.210 ;
        RECT 1117.200 1154.430 1118.380 1155.610 ;
        RECT 1117.200 1152.830 1118.380 1154.010 ;
        RECT 1192.450 1165.630 1193.630 1166.810 ;
        RECT 1192.450 1164.030 1193.630 1165.210 ;
        RECT 1192.450 1162.430 1193.630 1163.610 ;
        RECT 1192.450 1160.830 1193.630 1162.010 ;
        RECT 1192.450 1159.230 1193.630 1160.410 ;
        RECT 1192.450 1157.630 1193.630 1158.810 ;
        RECT 1192.450 1156.030 1193.630 1157.210 ;
        RECT 1192.450 1154.430 1193.630 1155.610 ;
        RECT 1192.450 1152.830 1193.630 1154.010 ;
        RECT 1267.700 1165.630 1268.880 1166.810 ;
        RECT 1267.700 1164.030 1268.880 1165.210 ;
        RECT 1267.700 1162.430 1268.880 1163.610 ;
        RECT 1267.700 1160.830 1268.880 1162.010 ;
        RECT 1267.700 1159.230 1268.880 1160.410 ;
        RECT 1267.700 1157.630 1268.880 1158.810 ;
        RECT 1267.700 1156.030 1268.880 1157.210 ;
        RECT 1267.700 1154.430 1268.880 1155.610 ;
        RECT 1267.700 1152.830 1268.880 1154.010 ;
        RECT 1342.950 1165.630 1344.130 1166.810 ;
        RECT 1342.950 1164.030 1344.130 1165.210 ;
        RECT 1342.950 1162.430 1344.130 1163.610 ;
        RECT 1342.950 1160.830 1344.130 1162.010 ;
        RECT 1342.950 1159.230 1344.130 1160.410 ;
        RECT 1342.950 1157.630 1344.130 1158.810 ;
        RECT 1342.950 1156.030 1344.130 1157.210 ;
        RECT 1342.950 1154.430 1344.130 1155.610 ;
        RECT 1342.950 1152.830 1344.130 1154.010 ;
        RECT 1418.200 1165.630 1419.380 1166.810 ;
        RECT 1418.200 1164.030 1419.380 1165.210 ;
        RECT 1418.200 1162.430 1419.380 1163.610 ;
        RECT 1418.200 1160.830 1419.380 1162.010 ;
        RECT 1418.200 1159.230 1419.380 1160.410 ;
        RECT 1418.200 1157.630 1419.380 1158.810 ;
        RECT 1418.200 1156.030 1419.380 1157.210 ;
        RECT 1418.200 1154.430 1419.380 1155.610 ;
        RECT 1418.200 1152.830 1419.380 1154.010 ;
        RECT 1493.450 1165.630 1494.630 1166.810 ;
        RECT 1493.450 1164.030 1494.630 1165.210 ;
        RECT 1493.450 1162.430 1494.630 1163.610 ;
        RECT 1493.450 1160.830 1494.630 1162.010 ;
        RECT 1493.450 1159.230 1494.630 1160.410 ;
        RECT 1493.450 1157.630 1494.630 1158.810 ;
        RECT 1493.450 1156.030 1494.630 1157.210 ;
        RECT 1493.450 1154.430 1494.630 1155.610 ;
        RECT 1493.450 1152.830 1494.630 1154.010 ;
        RECT 1568.700 1165.630 1569.880 1166.810 ;
        RECT 1568.700 1164.030 1569.880 1165.210 ;
        RECT 1568.700 1162.430 1569.880 1163.610 ;
        RECT 1568.700 1160.830 1569.880 1162.010 ;
        RECT 1568.700 1159.230 1569.880 1160.410 ;
        RECT 1568.700 1157.630 1569.880 1158.810 ;
        RECT 1568.700 1156.030 1569.880 1157.210 ;
        RECT 1568.700 1154.430 1569.880 1155.610 ;
        RECT 1568.700 1152.830 1569.880 1154.010 ;
        RECT 1643.950 1165.630 1645.130 1166.810 ;
        RECT 1643.950 1164.030 1645.130 1165.210 ;
        RECT 1643.950 1162.430 1645.130 1163.610 ;
        RECT 1643.950 1160.830 1645.130 1162.010 ;
        RECT 1643.950 1159.230 1645.130 1160.410 ;
        RECT 1643.950 1157.630 1645.130 1158.810 ;
        RECT 1643.950 1156.030 1645.130 1157.210 ;
        RECT 1643.950 1154.430 1645.130 1155.610 ;
        RECT 1643.950 1152.830 1645.130 1154.010 ;
        RECT 1719.200 1165.630 1720.380 1166.810 ;
        RECT 1719.200 1164.030 1720.380 1165.210 ;
        RECT 1719.200 1162.430 1720.380 1163.610 ;
        RECT 1719.200 1160.830 1720.380 1162.010 ;
        RECT 1719.200 1159.230 1720.380 1160.410 ;
        RECT 1719.200 1157.630 1720.380 1158.810 ;
        RECT 1719.200 1156.030 1720.380 1157.210 ;
        RECT 1719.200 1154.430 1720.380 1155.610 ;
        RECT 1719.200 1152.830 1720.380 1154.010 ;
        RECT 1794.450 1165.630 1795.630 1166.810 ;
        RECT 1794.450 1164.030 1795.630 1165.210 ;
        RECT 1794.450 1162.430 1795.630 1163.610 ;
        RECT 1794.450 1160.830 1795.630 1162.010 ;
        RECT 1794.450 1159.230 1795.630 1160.410 ;
        RECT 1794.450 1157.630 1795.630 1158.810 ;
        RECT 1794.450 1156.030 1795.630 1157.210 ;
        RECT 1794.450 1154.430 1795.630 1155.610 ;
        RECT 1794.450 1152.830 1795.630 1154.010 ;
        RECT 1869.700 1165.630 1870.880 1166.810 ;
        RECT 1869.700 1164.030 1870.880 1165.210 ;
        RECT 1869.700 1162.430 1870.880 1163.610 ;
        RECT 1869.700 1160.830 1870.880 1162.010 ;
        RECT 1869.700 1159.230 1870.880 1160.410 ;
        RECT 1869.700 1157.630 1870.880 1158.810 ;
        RECT 1869.700 1156.030 1870.880 1157.210 ;
        RECT 1869.700 1154.430 1870.880 1155.610 ;
        RECT 1869.700 1152.830 1870.880 1154.010 ;
        RECT 1944.950 1165.630 1946.130 1166.810 ;
        RECT 1944.950 1164.030 1946.130 1165.210 ;
        RECT 1944.950 1162.430 1946.130 1163.610 ;
        RECT 1944.950 1160.830 1946.130 1162.010 ;
        RECT 1944.950 1159.230 1946.130 1160.410 ;
        RECT 1944.950 1157.630 1946.130 1158.810 ;
        RECT 1944.950 1156.030 1946.130 1157.210 ;
        RECT 1944.950 1154.430 1946.130 1155.610 ;
        RECT 1944.950 1152.830 1946.130 1154.010 ;
        RECT 2020.200 1165.630 2021.380 1166.810 ;
        RECT 2020.200 1164.030 2021.380 1165.210 ;
        RECT 2020.200 1162.430 2021.380 1163.610 ;
        RECT 2020.200 1160.830 2021.380 1162.010 ;
        RECT 2020.200 1159.230 2021.380 1160.410 ;
        RECT 2020.200 1157.630 2021.380 1158.810 ;
        RECT 2020.200 1156.030 2021.380 1157.210 ;
        RECT 2020.200 1154.430 2021.380 1155.610 ;
        RECT 2020.200 1152.830 2021.380 1154.010 ;
        RECT 2095.450 1165.630 2096.630 1166.810 ;
        RECT 2095.450 1164.030 2096.630 1165.210 ;
        RECT 2095.450 1162.430 2096.630 1163.610 ;
        RECT 2095.450 1160.830 2096.630 1162.010 ;
        RECT 2095.450 1159.230 2096.630 1160.410 ;
        RECT 2095.450 1157.630 2096.630 1158.810 ;
        RECT 2095.450 1156.030 2096.630 1157.210 ;
        RECT 2095.450 1154.430 2096.630 1155.610 ;
        RECT 2095.450 1152.830 2096.630 1154.010 ;
        RECT 2170.700 1165.630 2171.880 1166.810 ;
        RECT 2170.700 1164.030 2171.880 1165.210 ;
        RECT 2170.700 1162.430 2171.880 1163.610 ;
        RECT 2170.700 1160.830 2171.880 1162.010 ;
        RECT 2170.700 1159.230 2171.880 1160.410 ;
        RECT 2170.700 1157.630 2171.880 1158.810 ;
        RECT 2170.700 1156.030 2171.880 1157.210 ;
        RECT 2170.700 1154.430 2171.880 1155.610 ;
        RECT 2170.700 1152.830 2171.880 1154.010 ;
        RECT 2245.950 1165.630 2247.130 1166.810 ;
        RECT 2245.950 1164.030 2247.130 1165.210 ;
        RECT 2245.950 1162.430 2247.130 1163.610 ;
        RECT 2245.950 1160.830 2247.130 1162.010 ;
        RECT 2245.950 1159.230 2247.130 1160.410 ;
        RECT 2245.950 1157.630 2247.130 1158.810 ;
        RECT 2245.950 1156.030 2247.130 1157.210 ;
        RECT 2245.950 1154.430 2247.130 1155.610 ;
        RECT 2245.950 1152.830 2247.130 1154.010 ;
        RECT 2321.200 1165.630 2322.380 1166.810 ;
        RECT 2321.200 1164.030 2322.380 1165.210 ;
        RECT 2321.200 1162.430 2322.380 1163.610 ;
        RECT 2321.200 1160.830 2322.380 1162.010 ;
        RECT 2321.200 1159.230 2322.380 1160.410 ;
        RECT 2321.200 1157.630 2322.380 1158.810 ;
        RECT 2321.200 1156.030 2322.380 1157.210 ;
        RECT 2321.200 1154.430 2322.380 1155.610 ;
        RECT 2321.200 1152.830 2322.380 1154.010 ;
        RECT 2396.450 1165.630 2397.630 1166.810 ;
        RECT 2396.450 1164.030 2397.630 1165.210 ;
        RECT 2396.450 1162.430 2397.630 1163.610 ;
        RECT 2396.450 1160.830 2397.630 1162.010 ;
        RECT 2396.450 1159.230 2397.630 1160.410 ;
        RECT 2396.450 1157.630 2397.630 1158.810 ;
        RECT 2396.450 1156.030 2397.630 1157.210 ;
        RECT 2396.450 1154.430 2397.630 1155.610 ;
        RECT 2396.450 1152.830 2397.630 1154.010 ;
        RECT 2471.700 1165.630 2472.880 1166.810 ;
        RECT 2471.700 1164.030 2472.880 1165.210 ;
        RECT 2471.700 1162.430 2472.880 1163.610 ;
        RECT 2471.700 1160.830 2472.880 1162.010 ;
        RECT 2471.700 1159.230 2472.880 1160.410 ;
        RECT 2471.700 1157.630 2472.880 1158.810 ;
        RECT 2471.700 1156.030 2472.880 1157.210 ;
        RECT 2471.700 1154.430 2472.880 1155.610 ;
        RECT 2471.700 1152.830 2472.880 1154.010 ;
        RECT 2546.950 1165.630 2548.130 1166.810 ;
        RECT 2546.950 1164.030 2548.130 1165.210 ;
        RECT 2546.950 1162.430 2548.130 1163.610 ;
        RECT 2546.950 1160.830 2548.130 1162.010 ;
        RECT 2546.950 1159.230 2548.130 1160.410 ;
        RECT 2546.950 1157.630 2548.130 1158.810 ;
        RECT 2546.950 1156.030 2548.130 1157.210 ;
        RECT 2546.950 1154.430 2548.130 1155.610 ;
        RECT 2546.950 1152.830 2548.130 1154.010 ;
        RECT 2622.200 1165.630 2623.380 1166.810 ;
        RECT 2622.200 1164.030 2623.380 1165.210 ;
        RECT 2622.200 1162.430 2623.380 1163.610 ;
        RECT 2622.200 1160.830 2623.380 1162.010 ;
        RECT 2622.200 1159.230 2623.380 1160.410 ;
        RECT 2622.200 1157.630 2623.380 1158.810 ;
        RECT 2622.200 1156.030 2623.380 1157.210 ;
        RECT 2622.200 1154.430 2623.380 1155.610 ;
        RECT 2622.200 1152.830 2623.380 1154.010 ;
        RECT 2697.200 1165.630 2698.380 1166.810 ;
        RECT 2697.200 1164.030 2698.380 1165.210 ;
        RECT 2697.200 1162.430 2698.380 1163.610 ;
        RECT 2697.200 1160.830 2698.380 1162.010 ;
        RECT 2697.200 1159.230 2698.380 1160.410 ;
        RECT 2697.200 1157.630 2698.380 1158.810 ;
        RECT 2697.200 1156.030 2698.380 1157.210 ;
        RECT 2697.200 1154.430 2698.380 1155.610 ;
        RECT 2697.200 1152.830 2698.380 1154.010 ;
        RECT 2899.000 1165.630 2900.180 1166.810 ;
        RECT 2899.000 1164.030 2900.180 1165.210 ;
        RECT 2899.000 1162.430 2900.180 1163.610 ;
        RECT 2899.000 1160.830 2900.180 1162.010 ;
        RECT 2899.000 1159.230 2900.180 1160.410 ;
        RECT 2899.000 1157.630 2900.180 1158.810 ;
        RECT 2899.000 1156.030 2900.180 1157.210 ;
        RECT 2899.000 1154.430 2900.180 1155.610 ;
        RECT 2899.000 1152.830 2900.180 1154.010 ;
        RECT 2919.000 1165.630 2920.180 1166.810 ;
        RECT 2919.000 1164.030 2920.180 1165.210 ;
        RECT 2919.000 1162.430 2920.180 1163.610 ;
        RECT 2919.000 1160.830 2920.180 1162.010 ;
        RECT 2919.000 1159.230 2920.180 1160.410 ;
        RECT 2919.000 1157.630 2920.180 1158.810 ;
        RECT 2919.000 1156.030 2920.180 1157.210 ;
        RECT 2919.000 1154.430 2920.180 1155.610 ;
        RECT 2919.000 1152.830 2920.180 1154.010 ;
        RECT 2923.050 1048.975 2935.430 1061.355 ;
        RECT 2967.320 1048.975 2979.700 1061.355 ;
        RECT 3136.515 1048.790 3139.295 1061.170 ;
        RECT 3213.315 1048.790 3216.095 1061.170 ;
        RECT 3290.115 1048.790 3292.895 1061.170 ;
        RECT 256.155 1045.600 257.335 1046.780 ;
        RECT 256.155 1044.000 257.335 1045.180 ;
        RECT 256.155 995.600 257.335 996.780 ;
        RECT 256.155 994.000 257.335 995.180 ;
        RECT 2923.915 995.485 2934.695 998.265 ;
        RECT 2960.190 995.895 2961.370 997.075 ;
        RECT 2961.790 995.895 2962.970 997.075 ;
        RECT 2963.390 995.895 2964.570 997.075 ;
        RECT 256.155 945.600 257.335 946.780 ;
        RECT 256.155 944.000 257.335 945.180 ;
        RECT 2923.915 917.285 2934.695 920.065 ;
        RECT 2960.190 917.695 2961.370 918.875 ;
        RECT 2961.790 917.695 2962.970 918.875 ;
        RECT 2963.390 917.695 2964.570 918.875 ;
        RECT 256.155 895.600 257.335 896.780 ;
        RECT 256.155 894.000 257.335 895.180 ;
        RECT 210.435 868.545 227.615 882.525 ;
        RECT 212.465 844.850 213.645 846.030 ;
        RECT 214.065 844.850 215.245 846.030 ;
        RECT 215.665 844.850 216.845 846.030 ;
        RECT 217.265 844.850 218.445 846.030 ;
        RECT 218.865 844.850 220.045 846.030 ;
        RECT 220.465 844.850 221.645 846.030 ;
        RECT 222.065 844.850 223.245 846.030 ;
        RECT 223.665 844.850 224.845 846.030 ;
        RECT 225.265 844.850 226.445 846.030 ;
        RECT 256.155 845.600 257.335 846.780 ;
        RECT 256.155 844.000 257.335 845.180 ;
        RECT 2923.915 839.085 2934.695 841.865 ;
        RECT 2960.190 839.495 2961.370 840.675 ;
        RECT 2961.790 839.495 2962.970 840.675 ;
        RECT 2963.390 839.495 2964.570 840.675 ;
        RECT 212.465 794.850 213.645 796.030 ;
        RECT 214.065 794.850 215.245 796.030 ;
        RECT 215.665 794.850 216.845 796.030 ;
        RECT 217.265 794.850 218.445 796.030 ;
        RECT 218.865 794.850 220.045 796.030 ;
        RECT 220.465 794.850 221.645 796.030 ;
        RECT 222.065 794.850 223.245 796.030 ;
        RECT 223.665 794.850 224.845 796.030 ;
        RECT 225.265 794.850 226.445 796.030 ;
        RECT 256.155 795.600 257.335 796.780 ;
        RECT 256.155 794.000 257.335 795.180 ;
        RECT 2923.915 760.885 2934.695 763.665 ;
        RECT 2960.190 761.295 2961.370 762.475 ;
        RECT 2961.790 761.295 2962.970 762.475 ;
        RECT 2963.390 761.295 2964.570 762.475 ;
        RECT 212.465 744.850 213.645 746.030 ;
        RECT 214.065 744.850 215.245 746.030 ;
        RECT 215.665 744.850 216.845 746.030 ;
        RECT 217.265 744.850 218.445 746.030 ;
        RECT 218.865 744.850 220.045 746.030 ;
        RECT 220.465 744.850 221.645 746.030 ;
        RECT 222.065 744.850 223.245 746.030 ;
        RECT 223.665 744.850 224.845 746.030 ;
        RECT 225.265 744.850 226.445 746.030 ;
        RECT 256.155 745.600 257.335 746.780 ;
        RECT 256.155 744.000 257.335 745.180 ;
        RECT 212.465 694.850 213.645 696.030 ;
        RECT 214.065 694.850 215.245 696.030 ;
        RECT 215.665 694.850 216.845 696.030 ;
        RECT 217.265 694.850 218.445 696.030 ;
        RECT 218.865 694.850 220.045 696.030 ;
        RECT 220.465 694.850 221.645 696.030 ;
        RECT 222.065 694.850 223.245 696.030 ;
        RECT 223.665 694.850 224.845 696.030 ;
        RECT 225.265 694.850 226.445 696.030 ;
        RECT 256.155 695.600 257.335 696.780 ;
        RECT 256.155 694.000 257.335 695.180 ;
        RECT 2923.915 682.685 2934.695 685.465 ;
        RECT 2960.190 683.095 2961.370 684.275 ;
        RECT 2961.790 683.095 2962.970 684.275 ;
        RECT 2963.390 683.095 2964.570 684.275 ;
        RECT 212.465 644.850 213.645 646.030 ;
        RECT 214.065 644.850 215.245 646.030 ;
        RECT 215.665 644.850 216.845 646.030 ;
        RECT 217.265 644.850 218.445 646.030 ;
        RECT 218.865 644.850 220.045 646.030 ;
        RECT 220.465 644.850 221.645 646.030 ;
        RECT 222.065 644.850 223.245 646.030 ;
        RECT 223.665 644.850 224.845 646.030 ;
        RECT 225.265 644.850 226.445 646.030 ;
        RECT 256.155 645.600 257.335 646.780 ;
        RECT 256.155 644.000 257.335 645.180 ;
        RECT 2960.190 604.895 2961.370 606.075 ;
        RECT 2961.790 604.895 2962.970 606.075 ;
        RECT 2963.390 604.895 2964.570 606.075 ;
        RECT 2923.915 598.485 2934.695 601.265 ;
        RECT 212.465 594.850 213.645 596.030 ;
        RECT 214.065 594.850 215.245 596.030 ;
        RECT 215.665 594.850 216.845 596.030 ;
        RECT 217.265 594.850 218.445 596.030 ;
        RECT 218.865 594.850 220.045 596.030 ;
        RECT 220.465 594.850 221.645 596.030 ;
        RECT 222.065 594.850 223.245 596.030 ;
        RECT 223.665 594.850 224.845 596.030 ;
        RECT 225.265 594.850 226.445 596.030 ;
        RECT 256.155 595.600 257.335 596.780 ;
        RECT 256.155 594.000 257.335 595.180 ;
        RECT 212.465 544.850 213.645 546.030 ;
        RECT 214.065 544.850 215.245 546.030 ;
        RECT 215.665 544.850 216.845 546.030 ;
        RECT 217.265 544.850 218.445 546.030 ;
        RECT 218.865 544.850 220.045 546.030 ;
        RECT 220.465 544.850 221.645 546.030 ;
        RECT 222.065 544.850 223.245 546.030 ;
        RECT 223.665 544.850 224.845 546.030 ;
        RECT 225.265 544.850 226.445 546.030 ;
        RECT 256.155 545.600 257.335 546.780 ;
        RECT 256.155 544.000 257.335 545.180 ;
        RECT 2923.915 526.285 2934.695 529.065 ;
        RECT 2960.190 526.695 2961.370 527.875 ;
        RECT 2961.790 526.695 2962.970 527.875 ;
        RECT 2963.390 526.695 2964.570 527.875 ;
        RECT 212.465 494.850 213.645 496.030 ;
        RECT 214.065 494.850 215.245 496.030 ;
        RECT 215.665 494.850 216.845 496.030 ;
        RECT 217.265 494.850 218.445 496.030 ;
        RECT 218.865 494.850 220.045 496.030 ;
        RECT 220.465 494.850 221.645 496.030 ;
        RECT 222.065 494.850 223.245 496.030 ;
        RECT 223.665 494.850 224.845 496.030 ;
        RECT 225.265 494.850 226.445 496.030 ;
        RECT 256.155 495.600 257.335 496.780 ;
        RECT 256.155 494.000 257.335 495.180 ;
        RECT 212.465 444.850 213.645 446.030 ;
        RECT 214.065 444.850 215.245 446.030 ;
        RECT 215.665 444.850 216.845 446.030 ;
        RECT 217.265 444.850 218.445 446.030 ;
        RECT 218.865 444.850 220.045 446.030 ;
        RECT 220.465 444.850 221.645 446.030 ;
        RECT 222.065 444.850 223.245 446.030 ;
        RECT 223.665 444.850 224.845 446.030 ;
        RECT 225.265 444.850 226.445 446.030 ;
        RECT 256.155 445.600 257.335 446.780 ;
        RECT 256.155 444.000 257.335 445.180 ;
        RECT 210.455 391.380 227.635 413.360 ;
        RECT 256.155 395.600 257.335 396.780 ;
        RECT 256.155 394.000 257.335 395.180 ;
        RECT 3161.270 392.365 3164.050 403.145 ;
        RECT 3201.160 391.700 3203.940 404.080 ;
        RECT 3149.495 384.785 3150.675 385.965 ;
        RECT 3149.495 383.185 3150.675 384.365 ;
        RECT 3149.495 381.585 3150.675 382.765 ;
        RECT 3165.055 384.855 3166.235 386.035 ;
        RECT 3165.055 383.255 3166.235 384.435 ;
        RECT 3165.055 381.655 3166.235 382.835 ;
        RECT 3180.505 384.835 3181.685 386.015 ;
        RECT 3180.505 383.235 3181.685 384.415 ;
        RECT 3180.505 381.635 3181.685 382.815 ;
        RECT 3195.975 384.835 3197.155 386.015 ;
        RECT 3195.975 383.235 3197.155 384.415 ;
        RECT 3195.975 381.635 3197.155 382.815 ;
        RECT 3211.515 384.895 3212.695 386.075 ;
        RECT 3211.515 383.295 3212.695 384.475 ;
        RECT 3211.515 381.695 3212.695 382.875 ;
        RECT 210.335 341.860 227.515 363.840 ;
        RECT 256.155 345.600 257.335 346.780 ;
        RECT 256.155 344.000 257.335 345.180 ;
        RECT 3149.495 316.815 3150.675 317.995 ;
        RECT 3149.495 315.215 3150.675 316.395 ;
        RECT 3149.495 313.615 3150.675 314.795 ;
        RECT 3165.055 316.885 3166.235 318.065 ;
        RECT 3165.055 315.285 3166.235 316.465 ;
        RECT 3165.055 313.685 3166.235 314.865 ;
        RECT 3180.505 316.865 3181.685 318.045 ;
        RECT 3180.505 315.265 3181.685 316.445 ;
        RECT 3180.505 313.665 3181.685 314.845 ;
        RECT 3195.975 316.865 3197.155 318.045 ;
        RECT 3195.975 315.265 3197.155 316.445 ;
        RECT 3195.975 313.665 3197.155 314.845 ;
        RECT 3211.515 316.925 3212.695 318.105 ;
        RECT 3211.515 315.325 3212.695 316.505 ;
        RECT 3211.515 313.725 3212.695 314.905 ;
        RECT 212.465 294.750 213.645 295.930 ;
        RECT 214.065 294.750 215.245 295.930 ;
        RECT 215.665 294.750 216.845 295.930 ;
        RECT 217.265 294.750 218.445 295.930 ;
        RECT 218.865 294.750 220.045 295.930 ;
        RECT 220.465 294.750 221.645 295.930 ;
        RECT 222.065 294.750 223.245 295.930 ;
        RECT 223.665 294.750 224.845 295.930 ;
        RECT 225.265 294.750 226.445 295.930 ;
        RECT 256.155 295.600 257.335 296.780 ;
        RECT 256.155 294.000 257.335 295.180 ;
        RECT 210.400 242.390 227.580 259.570 ;
        RECT 273.250 242.220 290.430 259.400 ;
        RECT 717.115 250.180 723.095 252.960 ;
        RECT 3332.610 235.190 3333.790 236.370 ;
        RECT 3334.210 235.190 3335.390 236.370 ;
        RECT 3335.810 235.190 3336.990 236.370 ;
        RECT 3337.410 235.190 3338.590 236.370 ;
        RECT 3339.010 235.190 3340.190 236.370 ;
        RECT 3340.610 235.190 3341.790 236.370 ;
        RECT 3342.210 235.190 3343.390 236.370 ;
        RECT 3343.810 235.190 3344.990 236.370 ;
        RECT 3345.410 235.190 3346.590 236.370 ;
      LAYER met5 ;
        RECT 281.480 1152.330 2936.870 1167.330 ;
        RECT 255.920 1043.790 266.080 1046.990 ;
        RECT 2873.230 1043.790 2901.550 1046.990 ;
        RECT 2898.350 1037.390 2901.550 1043.790 ;
        RECT 2921.870 1037.390 2936.870 1152.330 ;
        RECT 3243.040 1129.360 3256.790 1130.960 ;
        RECT 3251.120 1110.960 3256.790 1129.360 ;
        RECT 3243.200 1109.360 3256.790 1110.960 ;
        RECT 3251.120 1062.520 3256.790 1109.360 ;
        RECT 2966.260 1047.520 3347.130 1062.520 ;
        RECT 2898.350 1034.210 2936.870 1037.390 ;
        RECT 2901.550 1034.190 2936.870 1034.210 ;
        RECT 2921.870 996.990 2936.870 1034.190 ;
        RECT 3332.130 997.300 3347.130 1047.520 ;
        RECT 255.920 993.790 266.080 996.990 ;
        RECT 2873.230 993.790 2936.870 996.990 ;
        RECT 2959.880 995.700 2967.970 997.300 ;
        RECT 3325.880 995.700 3347.130 997.300 ;
        RECT 2921.870 946.990 2936.870 993.790 ;
        RECT 255.920 943.790 266.080 946.990 ;
        RECT 2873.230 943.790 2936.870 946.990 ;
        RECT 2921.870 896.990 2936.870 943.790 ;
        RECT 3332.130 919.100 3347.130 995.700 ;
        RECT 2959.880 917.500 2967.970 919.100 ;
        RECT 3325.880 917.500 3347.130 919.100 ;
        RECT 255.920 893.790 266.080 896.990 ;
        RECT 2873.230 893.790 2936.870 896.990 ;
        RECT 208.840 240.370 228.840 884.370 ;
        RECT 2921.870 846.990 2936.870 893.790 ;
        RECT 255.920 843.790 266.080 846.990 ;
        RECT 2873.230 843.790 2936.870 846.990 ;
        RECT 2921.870 796.990 2936.870 843.790 ;
        RECT 3332.130 840.900 3347.130 917.500 ;
        RECT 2959.880 839.300 2967.970 840.900 ;
        RECT 3325.880 839.300 3347.130 840.900 ;
        RECT 255.920 793.790 266.080 796.990 ;
        RECT 2873.230 793.790 2936.870 796.990 ;
        RECT 2921.870 746.990 2936.870 793.790 ;
        RECT 3332.130 762.700 3347.130 839.300 ;
        RECT 2959.880 761.100 2967.970 762.700 ;
        RECT 3325.880 761.100 3347.130 762.700 ;
        RECT 255.920 743.790 266.080 746.990 ;
        RECT 2873.230 743.790 2936.870 746.990 ;
        RECT 2921.870 696.990 2936.870 743.790 ;
        RECT 255.920 693.790 266.080 696.990 ;
        RECT 2873.230 693.790 2936.870 696.990 ;
        RECT 2921.870 646.990 2936.870 693.790 ;
        RECT 3332.130 684.500 3347.130 761.100 ;
        RECT 2959.880 682.900 2967.970 684.500 ;
        RECT 3325.880 682.900 3347.130 684.500 ;
        RECT 255.920 643.790 266.080 646.990 ;
        RECT 2873.230 643.790 2936.870 646.990 ;
        RECT 2921.870 596.990 2936.870 643.790 ;
        RECT 3332.130 606.300 3347.130 682.900 ;
        RECT 2959.880 604.700 2967.970 606.300 ;
        RECT 3325.880 604.700 3347.130 606.300 ;
        RECT 255.920 593.790 266.080 596.990 ;
        RECT 2873.230 593.790 2936.870 596.990 ;
        RECT 2921.870 546.990 2936.870 593.790 ;
        RECT 255.920 543.790 266.080 546.990 ;
        RECT 2873.230 543.790 2936.870 546.990 ;
        RECT 2921.870 496.990 2936.870 543.790 ;
        RECT 3332.130 528.100 3347.130 604.700 ;
        RECT 2959.880 526.500 2967.970 528.100 ;
        RECT 3325.880 526.500 3347.130 528.100 ;
        RECT 255.920 493.790 266.080 496.990 ;
        RECT 2873.230 493.790 2936.870 496.990 ;
        RECT 2921.870 446.990 2936.870 493.790 ;
        RECT 3217.720 467.370 3232.720 467.940 ;
        RECT 3209.530 465.770 3232.720 467.370 ;
        RECT 3332.130 467.030 3347.130 526.500 ;
        RECT 255.920 443.790 266.080 446.990 ;
        RECT 2873.230 443.790 2936.870 446.990 ;
        RECT 2921.870 396.990 2936.870 443.790 ;
        RECT 3217.720 427.370 3232.720 465.770 ;
        RECT 3312.610 465.430 3347.130 467.030 ;
        RECT 3332.130 458.870 3347.130 465.430 ;
        RECT 3312.420 457.270 3347.130 458.870 ;
        RECT 3332.130 450.710 3347.130 457.270 ;
        RECT 3312.520 449.110 3347.130 450.710 ;
        RECT 3209.840 425.770 3232.720 427.370 ;
        RECT 3217.720 405.410 3232.720 425.770 ;
        RECT 3332.130 405.410 3347.130 449.110 ;
        RECT 255.920 393.790 266.080 396.990 ;
        RECT 2873.230 393.790 2936.870 396.990 ;
        RECT 2921.870 346.990 2936.870 393.790 ;
        RECT 3160.010 390.410 3347.130 405.410 ;
        RECT 3226.280 386.340 3235.420 390.410 ;
        RECT 3148.930 381.340 3235.420 386.340 ;
        RECT 3231.420 367.430 3235.420 381.340 ;
        RECT 3227.680 365.830 3235.420 367.430 ;
        RECT 3231.420 350.530 3235.420 365.830 ;
        RECT 3227.510 348.930 3235.420 350.530 ;
        RECT 255.920 343.790 266.080 346.990 ;
        RECT 2873.230 343.790 2936.870 346.990 ;
        RECT 2921.870 296.990 2936.870 343.790 ;
        RECT 3231.420 333.630 3235.420 348.930 ;
        RECT 3228.120 332.030 3235.420 333.630 ;
        RECT 3231.420 318.370 3235.420 332.030 ;
        RECT 3148.930 313.370 3235.420 318.370 ;
        RECT 255.920 293.790 266.080 296.990 ;
        RECT 2873.230 293.790 2936.870 296.990 ;
        RECT 2921.870 261.110 2936.870 293.790 ;
        RECT 271.870 241.110 2936.870 261.110 ;
        RECT 3332.130 234.890 3347.130 390.410 ;
    END
  END vccd_core
  PIN vssd_core
    PORT
      LAYER met1 ;
        RECT 3240.520 233.690 3248.350 235.940 ;
        RECT 3240.520 232.990 3250.800 233.690 ;
        RECT 3240.520 232.950 3248.350 232.990 ;
      LAYER via ;
        RECT 3240.945 233.370 3247.925 235.550 ;
      LAYER met2 ;
        RECT 3240.520 233.690 3248.350 235.940 ;
        RECT 3240.520 232.990 3250.800 233.690 ;
        RECT 3240.520 232.950 3248.350 232.990 ;
      LAYER via2 ;
        RECT 3240.895 233.320 3247.975 235.600 ;
      LAYER met3 ;
        RECT 3240.520 234.220 3248.350 235.940 ;
        RECT 1208.450 197.130 1230.245 233.430 ;
        RECT 1256.500 197.130 1278.510 233.430 ;
        RECT 3240.520 232.990 3250.790 234.220 ;
        RECT 3240.520 232.950 3248.350 232.990 ;
      LAYER via3 ;
        RECT 1208.755 214.285 1229.875 233.005 ;
        RECT 1257.015 214.355 1278.135 233.075 ;
        RECT 3240.875 233.300 3247.995 235.620 ;
      LAYER met4 ;
        RECT 238.930 1172.330 316.250 1187.330 ;
        RECT 702.220 1172.240 704.620 1187.370 ;
        RECT 777.620 1172.240 780.020 1187.370 ;
        RECT 852.870 1172.240 855.270 1187.370 ;
        RECT 927.920 1172.240 930.320 1187.370 ;
        RECT 1078.620 1172.240 1081.020 1187.370 ;
        RECT 1153.870 1172.240 1156.270 1187.370 ;
        RECT 1229.120 1172.240 1231.520 1187.370 ;
        RECT 1304.370 1172.240 1306.770 1187.370 ;
        RECT 1379.620 1172.240 1382.020 1187.370 ;
        RECT 1454.870 1172.240 1457.270 1187.370 ;
        RECT 1529.920 1172.240 1532.320 1187.370 ;
        RECT 1605.870 1172.240 1608.270 1187.370 ;
        RECT 1680.620 1172.240 1683.020 1187.370 ;
        RECT 1755.570 1172.240 1757.970 1187.370 ;
        RECT 1831.120 1172.240 1833.520 1187.370 ;
        RECT 1905.770 1172.240 1908.170 1187.370 ;
        RECT 1981.220 1172.240 1983.620 1187.370 ;
        RECT 2056.870 1172.240 2059.270 1187.370 ;
        RECT 2132.120 1172.240 2134.520 1187.370 ;
        RECT 2207.370 1172.240 2209.770 1187.370 ;
        RECT 2282.620 1172.240 2285.020 1187.370 ;
        RECT 2357.870 1172.240 2360.270 1187.370 ;
        RECT 2433.120 1172.240 2435.520 1187.370 ;
        RECT 2508.370 1172.240 2510.770 1187.370 ;
        RECT 2583.620 1172.240 2586.020 1187.370 ;
        RECT 2658.870 1172.240 2661.270 1187.370 ;
        RECT 2733.870 1172.240 2736.270 1187.370 ;
        RECT 2911.310 1039.310 2956.940 1042.510 ;
        RECT 2910.360 1005.310 2956.940 1008.510 ;
        RECT 2910.360 955.310 2956.940 958.510 ;
        RECT 2910.360 905.310 2956.940 908.510 ;
        RECT 2910.360 855.310 2956.940 858.510 ;
        RECT 2910.360 805.310 2956.940 808.510 ;
        RECT 2910.360 755.310 2956.940 758.510 ;
        RECT 2910.360 705.310 2956.940 708.510 ;
        RECT 2910.360 655.310 2956.940 658.510 ;
        RECT 2910.360 605.310 2956.940 608.510 ;
        RECT 2910.360 555.310 2956.940 558.510 ;
        RECT 2910.360 505.310 2956.940 508.510 ;
        RECT 2986.510 493.800 2988.110 511.580 ;
        RECT 3063.310 494.020 3064.910 511.190 ;
        RECT 3140.110 494.020 3141.710 511.190 ;
        RECT 3216.910 494.020 3218.510 511.190 ;
        RECT 3293.710 494.020 3295.310 510.650 ;
        RECT 2983.710 479.780 2990.760 493.800 ;
        RECT 3061.120 480.250 3067.710 494.020 ;
        RECT 3137.920 480.250 3144.510 494.020 ;
        RECT 3180.400 482.170 3184.970 493.790 ;
        RECT 3181.770 472.240 3183.370 482.170 ;
        RECT 3214.720 480.250 3221.310 494.020 ;
        RECT 3291.520 480.250 3297.965 494.020 ;
        RECT 2910.360 455.310 2956.940 458.510 ;
        RECT 2910.360 405.310 2956.940 408.510 ;
        RECT 3157.090 370.520 3158.690 386.870 ;
        RECT 3172.590 370.520 3174.190 386.870 ;
        RECT 3188.090 370.520 3189.690 386.870 ;
        RECT 3203.590 370.520 3205.190 386.870 ;
        RECT 3219.090 370.520 3220.690 386.870 ;
        RECT 2910.360 355.310 2956.940 358.510 ;
        RECT 2910.360 305.310 2956.940 308.510 ;
        RECT 3157.090 302.550 3158.690 318.900 ;
        RECT 3172.590 302.550 3174.190 318.900 ;
        RECT 3188.090 302.550 3189.690 318.900 ;
        RECT 3203.590 302.550 3205.190 318.900 ;
        RECT 3219.090 302.550 3220.690 318.900 ;
        RECT 712.800 226.980 713.700 236.280 ;
        RECT 708.880 226.970 714.330 226.980 ;
        RECT 706.880 220.650 714.330 226.970 ;
        RECT 1208.400 213.920 1230.280 233.460 ;
        RECT 1256.510 213.940 1278.500 233.420 ;
        RECT 3240.520 232.950 3248.350 235.940 ;
      LAYER via4 ;
        RECT 240.455 1173.695 252.835 1186.075 ;
        RECT 282.275 1173.725 315.455 1186.105 ;
        RECT 702.600 1185.625 703.780 1186.805 ;
        RECT 702.600 1184.025 703.780 1185.205 ;
        RECT 702.600 1182.425 703.780 1183.605 ;
        RECT 702.600 1180.825 703.780 1182.005 ;
        RECT 702.600 1179.225 703.780 1180.405 ;
        RECT 702.600 1177.625 703.780 1178.805 ;
        RECT 702.600 1176.025 703.780 1177.205 ;
        RECT 702.600 1174.425 703.780 1175.605 ;
        RECT 702.600 1172.825 703.780 1174.005 ;
        RECT 778.000 1185.625 779.180 1186.805 ;
        RECT 778.000 1184.025 779.180 1185.205 ;
        RECT 778.000 1182.425 779.180 1183.605 ;
        RECT 778.000 1180.825 779.180 1182.005 ;
        RECT 778.000 1179.225 779.180 1180.405 ;
        RECT 778.000 1177.625 779.180 1178.805 ;
        RECT 778.000 1176.025 779.180 1177.205 ;
        RECT 778.000 1174.425 779.180 1175.605 ;
        RECT 778.000 1172.825 779.180 1174.005 ;
        RECT 853.250 1185.625 854.430 1186.805 ;
        RECT 853.250 1184.025 854.430 1185.205 ;
        RECT 853.250 1182.425 854.430 1183.605 ;
        RECT 853.250 1180.825 854.430 1182.005 ;
        RECT 853.250 1179.225 854.430 1180.405 ;
        RECT 853.250 1177.625 854.430 1178.805 ;
        RECT 853.250 1176.025 854.430 1177.205 ;
        RECT 853.250 1174.425 854.430 1175.605 ;
        RECT 853.250 1172.825 854.430 1174.005 ;
        RECT 928.300 1185.625 929.480 1186.805 ;
        RECT 928.300 1184.025 929.480 1185.205 ;
        RECT 928.300 1182.425 929.480 1183.605 ;
        RECT 928.300 1180.825 929.480 1182.005 ;
        RECT 928.300 1179.225 929.480 1180.405 ;
        RECT 928.300 1177.625 929.480 1178.805 ;
        RECT 928.300 1176.025 929.480 1177.205 ;
        RECT 928.300 1174.425 929.480 1175.605 ;
        RECT 928.300 1172.825 929.480 1174.005 ;
        RECT 1079.000 1185.625 1080.180 1186.805 ;
        RECT 1079.000 1184.025 1080.180 1185.205 ;
        RECT 1079.000 1182.425 1080.180 1183.605 ;
        RECT 1079.000 1180.825 1080.180 1182.005 ;
        RECT 1079.000 1179.225 1080.180 1180.405 ;
        RECT 1079.000 1177.625 1080.180 1178.805 ;
        RECT 1079.000 1176.025 1080.180 1177.205 ;
        RECT 1079.000 1174.425 1080.180 1175.605 ;
        RECT 1079.000 1172.825 1080.180 1174.005 ;
        RECT 1154.250 1185.625 1155.430 1186.805 ;
        RECT 1154.250 1184.025 1155.430 1185.205 ;
        RECT 1154.250 1182.425 1155.430 1183.605 ;
        RECT 1154.250 1180.825 1155.430 1182.005 ;
        RECT 1154.250 1179.225 1155.430 1180.405 ;
        RECT 1154.250 1177.625 1155.430 1178.805 ;
        RECT 1154.250 1176.025 1155.430 1177.205 ;
        RECT 1154.250 1174.425 1155.430 1175.605 ;
        RECT 1154.250 1172.825 1155.430 1174.005 ;
        RECT 1229.500 1185.625 1230.680 1186.805 ;
        RECT 1229.500 1184.025 1230.680 1185.205 ;
        RECT 1229.500 1182.425 1230.680 1183.605 ;
        RECT 1229.500 1180.825 1230.680 1182.005 ;
        RECT 1229.500 1179.225 1230.680 1180.405 ;
        RECT 1229.500 1177.625 1230.680 1178.805 ;
        RECT 1229.500 1176.025 1230.680 1177.205 ;
        RECT 1229.500 1174.425 1230.680 1175.605 ;
        RECT 1229.500 1172.825 1230.680 1174.005 ;
        RECT 1304.750 1185.625 1305.930 1186.805 ;
        RECT 1304.750 1184.025 1305.930 1185.205 ;
        RECT 1304.750 1182.425 1305.930 1183.605 ;
        RECT 1304.750 1180.825 1305.930 1182.005 ;
        RECT 1304.750 1179.225 1305.930 1180.405 ;
        RECT 1304.750 1177.625 1305.930 1178.805 ;
        RECT 1304.750 1176.025 1305.930 1177.205 ;
        RECT 1304.750 1174.425 1305.930 1175.605 ;
        RECT 1304.750 1172.825 1305.930 1174.005 ;
        RECT 1380.000 1185.625 1381.180 1186.805 ;
        RECT 1380.000 1184.025 1381.180 1185.205 ;
        RECT 1380.000 1182.425 1381.180 1183.605 ;
        RECT 1380.000 1180.825 1381.180 1182.005 ;
        RECT 1380.000 1179.225 1381.180 1180.405 ;
        RECT 1380.000 1177.625 1381.180 1178.805 ;
        RECT 1380.000 1176.025 1381.180 1177.205 ;
        RECT 1380.000 1174.425 1381.180 1175.605 ;
        RECT 1380.000 1172.825 1381.180 1174.005 ;
        RECT 1455.250 1185.625 1456.430 1186.805 ;
        RECT 1455.250 1184.025 1456.430 1185.205 ;
        RECT 1455.250 1182.425 1456.430 1183.605 ;
        RECT 1455.250 1180.825 1456.430 1182.005 ;
        RECT 1455.250 1179.225 1456.430 1180.405 ;
        RECT 1455.250 1177.625 1456.430 1178.805 ;
        RECT 1455.250 1176.025 1456.430 1177.205 ;
        RECT 1455.250 1174.425 1456.430 1175.605 ;
        RECT 1455.250 1172.825 1456.430 1174.005 ;
        RECT 1530.300 1185.625 1531.480 1186.805 ;
        RECT 1530.300 1184.025 1531.480 1185.205 ;
        RECT 1530.300 1182.425 1531.480 1183.605 ;
        RECT 1530.300 1180.825 1531.480 1182.005 ;
        RECT 1530.300 1179.225 1531.480 1180.405 ;
        RECT 1530.300 1177.625 1531.480 1178.805 ;
        RECT 1530.300 1176.025 1531.480 1177.205 ;
        RECT 1530.300 1174.425 1531.480 1175.605 ;
        RECT 1530.300 1172.825 1531.480 1174.005 ;
        RECT 1606.250 1185.625 1607.430 1186.805 ;
        RECT 1606.250 1184.025 1607.430 1185.205 ;
        RECT 1606.250 1182.425 1607.430 1183.605 ;
        RECT 1606.250 1180.825 1607.430 1182.005 ;
        RECT 1606.250 1179.225 1607.430 1180.405 ;
        RECT 1606.250 1177.625 1607.430 1178.805 ;
        RECT 1606.250 1176.025 1607.430 1177.205 ;
        RECT 1606.250 1174.425 1607.430 1175.605 ;
        RECT 1606.250 1172.825 1607.430 1174.005 ;
        RECT 1681.000 1185.625 1682.180 1186.805 ;
        RECT 1681.000 1184.025 1682.180 1185.205 ;
        RECT 1681.000 1182.425 1682.180 1183.605 ;
        RECT 1681.000 1180.825 1682.180 1182.005 ;
        RECT 1681.000 1179.225 1682.180 1180.405 ;
        RECT 1681.000 1177.625 1682.180 1178.805 ;
        RECT 1681.000 1176.025 1682.180 1177.205 ;
        RECT 1681.000 1174.425 1682.180 1175.605 ;
        RECT 1681.000 1172.825 1682.180 1174.005 ;
        RECT 1755.950 1185.625 1757.130 1186.805 ;
        RECT 1755.950 1184.025 1757.130 1185.205 ;
        RECT 1755.950 1182.425 1757.130 1183.605 ;
        RECT 1755.950 1180.825 1757.130 1182.005 ;
        RECT 1755.950 1179.225 1757.130 1180.405 ;
        RECT 1755.950 1177.625 1757.130 1178.805 ;
        RECT 1755.950 1176.025 1757.130 1177.205 ;
        RECT 1755.950 1174.425 1757.130 1175.605 ;
        RECT 1755.950 1172.825 1757.130 1174.005 ;
        RECT 1831.500 1185.625 1832.680 1186.805 ;
        RECT 1831.500 1184.025 1832.680 1185.205 ;
        RECT 1831.500 1182.425 1832.680 1183.605 ;
        RECT 1831.500 1180.825 1832.680 1182.005 ;
        RECT 1831.500 1179.225 1832.680 1180.405 ;
        RECT 1831.500 1177.625 1832.680 1178.805 ;
        RECT 1831.500 1176.025 1832.680 1177.205 ;
        RECT 1831.500 1174.425 1832.680 1175.605 ;
        RECT 1831.500 1172.825 1832.680 1174.005 ;
        RECT 1906.150 1185.625 1907.330 1186.805 ;
        RECT 1906.150 1184.025 1907.330 1185.205 ;
        RECT 1906.150 1182.425 1907.330 1183.605 ;
        RECT 1906.150 1180.825 1907.330 1182.005 ;
        RECT 1906.150 1179.225 1907.330 1180.405 ;
        RECT 1906.150 1177.625 1907.330 1178.805 ;
        RECT 1906.150 1176.025 1907.330 1177.205 ;
        RECT 1906.150 1174.425 1907.330 1175.605 ;
        RECT 1906.150 1172.825 1907.330 1174.005 ;
        RECT 1981.600 1185.625 1982.780 1186.805 ;
        RECT 1981.600 1184.025 1982.780 1185.205 ;
        RECT 1981.600 1182.425 1982.780 1183.605 ;
        RECT 1981.600 1180.825 1982.780 1182.005 ;
        RECT 1981.600 1179.225 1982.780 1180.405 ;
        RECT 1981.600 1177.625 1982.780 1178.805 ;
        RECT 1981.600 1176.025 1982.780 1177.205 ;
        RECT 1981.600 1174.425 1982.780 1175.605 ;
        RECT 1981.600 1172.825 1982.780 1174.005 ;
        RECT 2057.250 1185.625 2058.430 1186.805 ;
        RECT 2057.250 1184.025 2058.430 1185.205 ;
        RECT 2057.250 1182.425 2058.430 1183.605 ;
        RECT 2057.250 1180.825 2058.430 1182.005 ;
        RECT 2057.250 1179.225 2058.430 1180.405 ;
        RECT 2057.250 1177.625 2058.430 1178.805 ;
        RECT 2057.250 1176.025 2058.430 1177.205 ;
        RECT 2057.250 1174.425 2058.430 1175.605 ;
        RECT 2057.250 1172.825 2058.430 1174.005 ;
        RECT 2132.500 1185.625 2133.680 1186.805 ;
        RECT 2132.500 1184.025 2133.680 1185.205 ;
        RECT 2132.500 1182.425 2133.680 1183.605 ;
        RECT 2132.500 1180.825 2133.680 1182.005 ;
        RECT 2132.500 1179.225 2133.680 1180.405 ;
        RECT 2132.500 1177.625 2133.680 1178.805 ;
        RECT 2132.500 1176.025 2133.680 1177.205 ;
        RECT 2132.500 1174.425 2133.680 1175.605 ;
        RECT 2132.500 1172.825 2133.680 1174.005 ;
        RECT 2207.750 1185.625 2208.930 1186.805 ;
        RECT 2207.750 1184.025 2208.930 1185.205 ;
        RECT 2207.750 1182.425 2208.930 1183.605 ;
        RECT 2207.750 1180.825 2208.930 1182.005 ;
        RECT 2207.750 1179.225 2208.930 1180.405 ;
        RECT 2207.750 1177.625 2208.930 1178.805 ;
        RECT 2207.750 1176.025 2208.930 1177.205 ;
        RECT 2207.750 1174.425 2208.930 1175.605 ;
        RECT 2207.750 1172.825 2208.930 1174.005 ;
        RECT 2283.000 1185.625 2284.180 1186.805 ;
        RECT 2283.000 1184.025 2284.180 1185.205 ;
        RECT 2283.000 1182.425 2284.180 1183.605 ;
        RECT 2283.000 1180.825 2284.180 1182.005 ;
        RECT 2283.000 1179.225 2284.180 1180.405 ;
        RECT 2283.000 1177.625 2284.180 1178.805 ;
        RECT 2283.000 1176.025 2284.180 1177.205 ;
        RECT 2283.000 1174.425 2284.180 1175.605 ;
        RECT 2283.000 1172.825 2284.180 1174.005 ;
        RECT 2358.250 1185.625 2359.430 1186.805 ;
        RECT 2358.250 1184.025 2359.430 1185.205 ;
        RECT 2358.250 1182.425 2359.430 1183.605 ;
        RECT 2358.250 1180.825 2359.430 1182.005 ;
        RECT 2358.250 1179.225 2359.430 1180.405 ;
        RECT 2358.250 1177.625 2359.430 1178.805 ;
        RECT 2358.250 1176.025 2359.430 1177.205 ;
        RECT 2358.250 1174.425 2359.430 1175.605 ;
        RECT 2358.250 1172.825 2359.430 1174.005 ;
        RECT 2433.500 1185.625 2434.680 1186.805 ;
        RECT 2433.500 1184.025 2434.680 1185.205 ;
        RECT 2433.500 1182.425 2434.680 1183.605 ;
        RECT 2433.500 1180.825 2434.680 1182.005 ;
        RECT 2433.500 1179.225 2434.680 1180.405 ;
        RECT 2433.500 1177.625 2434.680 1178.805 ;
        RECT 2433.500 1176.025 2434.680 1177.205 ;
        RECT 2433.500 1174.425 2434.680 1175.605 ;
        RECT 2433.500 1172.825 2434.680 1174.005 ;
        RECT 2508.750 1185.625 2509.930 1186.805 ;
        RECT 2508.750 1184.025 2509.930 1185.205 ;
        RECT 2508.750 1182.425 2509.930 1183.605 ;
        RECT 2508.750 1180.825 2509.930 1182.005 ;
        RECT 2508.750 1179.225 2509.930 1180.405 ;
        RECT 2508.750 1177.625 2509.930 1178.805 ;
        RECT 2508.750 1176.025 2509.930 1177.205 ;
        RECT 2508.750 1174.425 2509.930 1175.605 ;
        RECT 2508.750 1172.825 2509.930 1174.005 ;
        RECT 2584.000 1185.625 2585.180 1186.805 ;
        RECT 2584.000 1184.025 2585.180 1185.205 ;
        RECT 2584.000 1182.425 2585.180 1183.605 ;
        RECT 2584.000 1180.825 2585.180 1182.005 ;
        RECT 2584.000 1179.225 2585.180 1180.405 ;
        RECT 2584.000 1177.625 2585.180 1178.805 ;
        RECT 2584.000 1176.025 2585.180 1177.205 ;
        RECT 2584.000 1174.425 2585.180 1175.605 ;
        RECT 2584.000 1172.825 2585.180 1174.005 ;
        RECT 2659.250 1185.625 2660.430 1186.805 ;
        RECT 2659.250 1184.025 2660.430 1185.205 ;
        RECT 2659.250 1182.425 2660.430 1183.605 ;
        RECT 2659.250 1180.825 2660.430 1182.005 ;
        RECT 2659.250 1179.225 2660.430 1180.405 ;
        RECT 2659.250 1177.625 2660.430 1178.805 ;
        RECT 2659.250 1176.025 2660.430 1177.205 ;
        RECT 2659.250 1174.425 2660.430 1175.605 ;
        RECT 2659.250 1172.825 2660.430 1174.005 ;
        RECT 2734.250 1185.625 2735.430 1186.805 ;
        RECT 2734.250 1184.025 2735.430 1185.205 ;
        RECT 2734.250 1182.425 2735.430 1183.605 ;
        RECT 2734.250 1180.825 2735.430 1182.005 ;
        RECT 2734.250 1179.225 2735.430 1180.405 ;
        RECT 2734.250 1177.625 2735.430 1178.805 ;
        RECT 2734.250 1176.025 2735.430 1177.205 ;
        RECT 2734.250 1174.425 2735.430 1175.605 ;
        RECT 2734.250 1172.825 2735.430 1174.005 ;
        RECT 2912.000 1040.330 2913.180 1041.510 ;
        RECT 2913.600 1040.330 2914.780 1041.510 ;
        RECT 2915.200 1040.330 2916.380 1041.510 ;
        RECT 2916.800 1040.330 2917.980 1041.510 ;
        RECT 2942.465 1040.330 2943.645 1041.510 ;
        RECT 2944.065 1040.330 2945.245 1041.510 ;
        RECT 2945.665 1040.330 2946.845 1041.510 ;
        RECT 2947.265 1040.330 2948.445 1041.510 ;
        RECT 2948.865 1040.330 2950.045 1041.510 ;
        RECT 2950.465 1040.330 2951.645 1041.510 ;
        RECT 2952.065 1040.330 2953.245 1041.510 ;
        RECT 2953.665 1040.330 2954.845 1041.510 ;
        RECT 2955.265 1040.330 2956.445 1041.510 ;
        RECT 2911.020 1006.270 2912.200 1007.450 ;
        RECT 2912.620 1006.270 2913.800 1007.450 ;
        RECT 2942.465 1006.250 2943.645 1007.430 ;
        RECT 2944.065 1006.250 2945.245 1007.430 ;
        RECT 2945.665 1006.250 2946.845 1007.430 ;
        RECT 2947.265 1006.250 2948.445 1007.430 ;
        RECT 2948.865 1006.250 2950.045 1007.430 ;
        RECT 2950.465 1006.250 2951.645 1007.430 ;
        RECT 2952.065 1006.250 2953.245 1007.430 ;
        RECT 2953.665 1006.250 2954.845 1007.430 ;
        RECT 2955.265 1006.250 2956.445 1007.430 ;
        RECT 2911.020 956.270 2912.200 957.450 ;
        RECT 2912.620 956.270 2913.800 957.450 ;
        RECT 2942.465 956.250 2943.645 957.430 ;
        RECT 2944.065 956.250 2945.245 957.430 ;
        RECT 2945.665 956.250 2946.845 957.430 ;
        RECT 2947.265 956.250 2948.445 957.430 ;
        RECT 2948.865 956.250 2950.045 957.430 ;
        RECT 2950.465 956.250 2951.645 957.430 ;
        RECT 2952.065 956.250 2953.245 957.430 ;
        RECT 2953.665 956.250 2954.845 957.430 ;
        RECT 2955.265 956.250 2956.445 957.430 ;
        RECT 2911.020 906.270 2912.200 907.450 ;
        RECT 2912.620 906.270 2913.800 907.450 ;
        RECT 2942.465 906.250 2943.645 907.430 ;
        RECT 2944.065 906.250 2945.245 907.430 ;
        RECT 2945.665 906.250 2946.845 907.430 ;
        RECT 2947.265 906.250 2948.445 907.430 ;
        RECT 2948.865 906.250 2950.045 907.430 ;
        RECT 2950.465 906.250 2951.645 907.430 ;
        RECT 2952.065 906.250 2953.245 907.430 ;
        RECT 2953.665 906.250 2954.845 907.430 ;
        RECT 2955.265 906.250 2956.445 907.430 ;
        RECT 2911.020 856.270 2912.200 857.450 ;
        RECT 2912.620 856.270 2913.800 857.450 ;
        RECT 2942.465 856.250 2943.645 857.430 ;
        RECT 2944.065 856.250 2945.245 857.430 ;
        RECT 2945.665 856.250 2946.845 857.430 ;
        RECT 2947.265 856.250 2948.445 857.430 ;
        RECT 2948.865 856.250 2950.045 857.430 ;
        RECT 2950.465 856.250 2951.645 857.430 ;
        RECT 2952.065 856.250 2953.245 857.430 ;
        RECT 2953.665 856.250 2954.845 857.430 ;
        RECT 2955.265 856.250 2956.445 857.430 ;
        RECT 2911.020 806.270 2912.200 807.450 ;
        RECT 2912.620 806.270 2913.800 807.450 ;
        RECT 2942.465 806.250 2943.645 807.430 ;
        RECT 2944.065 806.250 2945.245 807.430 ;
        RECT 2945.665 806.250 2946.845 807.430 ;
        RECT 2947.265 806.250 2948.445 807.430 ;
        RECT 2948.865 806.250 2950.045 807.430 ;
        RECT 2950.465 806.250 2951.645 807.430 ;
        RECT 2952.065 806.250 2953.245 807.430 ;
        RECT 2953.665 806.250 2954.845 807.430 ;
        RECT 2955.265 806.250 2956.445 807.430 ;
        RECT 2911.020 756.270 2912.200 757.450 ;
        RECT 2912.620 756.270 2913.800 757.450 ;
        RECT 2942.465 756.250 2943.645 757.430 ;
        RECT 2944.065 756.250 2945.245 757.430 ;
        RECT 2945.665 756.250 2946.845 757.430 ;
        RECT 2947.265 756.250 2948.445 757.430 ;
        RECT 2948.865 756.250 2950.045 757.430 ;
        RECT 2950.465 756.250 2951.645 757.430 ;
        RECT 2952.065 756.250 2953.245 757.430 ;
        RECT 2953.665 756.250 2954.845 757.430 ;
        RECT 2955.265 756.250 2956.445 757.430 ;
        RECT 2911.020 706.270 2912.200 707.450 ;
        RECT 2912.620 706.270 2913.800 707.450 ;
        RECT 2942.465 706.250 2943.645 707.430 ;
        RECT 2944.065 706.250 2945.245 707.430 ;
        RECT 2945.665 706.250 2946.845 707.430 ;
        RECT 2947.265 706.250 2948.445 707.430 ;
        RECT 2948.865 706.250 2950.045 707.430 ;
        RECT 2950.465 706.250 2951.645 707.430 ;
        RECT 2952.065 706.250 2953.245 707.430 ;
        RECT 2953.665 706.250 2954.845 707.430 ;
        RECT 2955.265 706.250 2956.445 707.430 ;
        RECT 2911.020 656.270 2912.200 657.450 ;
        RECT 2912.620 656.270 2913.800 657.450 ;
        RECT 2942.465 656.250 2943.645 657.430 ;
        RECT 2944.065 656.250 2945.245 657.430 ;
        RECT 2945.665 656.250 2946.845 657.430 ;
        RECT 2947.265 656.250 2948.445 657.430 ;
        RECT 2948.865 656.250 2950.045 657.430 ;
        RECT 2950.465 656.250 2951.645 657.430 ;
        RECT 2952.065 656.250 2953.245 657.430 ;
        RECT 2953.665 656.250 2954.845 657.430 ;
        RECT 2955.265 656.250 2956.445 657.430 ;
        RECT 2911.020 606.270 2912.200 607.450 ;
        RECT 2912.620 606.270 2913.800 607.450 ;
        RECT 2942.465 606.250 2943.645 607.430 ;
        RECT 2944.065 606.250 2945.245 607.430 ;
        RECT 2945.665 606.250 2946.845 607.430 ;
        RECT 2947.265 606.250 2948.445 607.430 ;
        RECT 2948.865 606.250 2950.045 607.430 ;
        RECT 2950.465 606.250 2951.645 607.430 ;
        RECT 2952.065 606.250 2953.245 607.430 ;
        RECT 2953.665 606.250 2954.845 607.430 ;
        RECT 2955.265 606.250 2956.445 607.430 ;
        RECT 2911.020 556.270 2912.200 557.450 ;
        RECT 2912.620 556.270 2913.800 557.450 ;
        RECT 2942.465 556.250 2943.645 557.430 ;
        RECT 2944.065 556.250 2945.245 557.430 ;
        RECT 2945.665 556.250 2946.845 557.430 ;
        RECT 2947.265 556.250 2948.445 557.430 ;
        RECT 2948.865 556.250 2950.045 557.430 ;
        RECT 2950.465 556.250 2951.645 557.430 ;
        RECT 2952.065 556.250 2953.245 557.430 ;
        RECT 2953.665 556.250 2954.845 557.430 ;
        RECT 2955.265 556.250 2956.445 557.430 ;
        RECT 2911.020 506.270 2912.200 507.450 ;
        RECT 2912.620 506.270 2913.800 507.450 ;
        RECT 2942.465 506.250 2943.645 507.430 ;
        RECT 2944.065 506.250 2945.245 507.430 ;
        RECT 2945.665 506.250 2946.845 507.430 ;
        RECT 2947.265 506.250 2948.445 507.430 ;
        RECT 2948.865 506.250 2950.045 507.430 ;
        RECT 2950.465 506.250 2951.645 507.430 ;
        RECT 2952.065 506.250 2953.245 507.430 ;
        RECT 2953.665 506.250 2954.845 507.430 ;
        RECT 2955.265 506.250 2956.445 507.430 ;
        RECT 2985.060 480.635 2989.440 493.015 ;
        RECT 3062.315 480.945 3066.695 493.325 ;
        RECT 3139.115 480.945 3143.495 493.325 ;
        RECT 3181.295 483.425 3184.075 492.605 ;
        RECT 3215.915 480.945 3220.295 493.325 ;
        RECT 3292.715 480.945 3297.095 493.325 ;
        RECT 2911.020 456.270 2912.200 457.450 ;
        RECT 2912.620 456.270 2913.800 457.450 ;
        RECT 2942.465 456.250 2943.645 457.430 ;
        RECT 2944.065 456.250 2945.245 457.430 ;
        RECT 2945.665 456.250 2946.845 457.430 ;
        RECT 2947.265 456.250 2948.445 457.430 ;
        RECT 2948.865 456.250 2950.045 457.430 ;
        RECT 2950.465 456.250 2951.645 457.430 ;
        RECT 2952.065 456.250 2953.245 457.430 ;
        RECT 2953.665 456.250 2954.845 457.430 ;
        RECT 2955.265 456.250 2956.445 457.430 ;
        RECT 2911.020 406.270 2912.200 407.450 ;
        RECT 2912.620 406.270 2913.800 407.450 ;
        RECT 2942.465 406.250 2943.645 407.430 ;
        RECT 2944.065 406.250 2945.245 407.430 ;
        RECT 2945.665 406.250 2946.845 407.430 ;
        RECT 2947.265 406.250 2948.445 407.430 ;
        RECT 2948.865 406.250 2950.045 407.430 ;
        RECT 2950.465 406.250 2951.645 407.430 ;
        RECT 2952.065 406.250 2953.245 407.430 ;
        RECT 2953.665 406.250 2954.845 407.430 ;
        RECT 2955.265 406.250 2956.445 407.430 ;
        RECT 3157.255 377.775 3158.435 378.955 ;
        RECT 3157.255 376.175 3158.435 377.355 ;
        RECT 3157.255 374.575 3158.435 375.755 ;
        RECT 3172.725 377.795 3173.905 378.975 ;
        RECT 3172.725 376.195 3173.905 377.375 ;
        RECT 3172.725 374.595 3173.905 375.775 ;
        RECT 3188.265 377.815 3189.445 378.995 ;
        RECT 3188.265 376.215 3189.445 377.395 ;
        RECT 3188.265 374.615 3189.445 375.795 ;
        RECT 3203.785 377.775 3204.965 378.955 ;
        RECT 3203.785 376.175 3204.965 377.355 ;
        RECT 3203.785 374.575 3204.965 375.755 ;
        RECT 3219.295 377.905 3220.475 379.085 ;
        RECT 3219.295 376.305 3220.475 377.485 ;
        RECT 3219.295 374.705 3220.475 375.885 ;
        RECT 2911.020 356.270 2912.200 357.450 ;
        RECT 2912.620 356.270 2913.800 357.450 ;
        RECT 2942.465 356.250 2943.645 357.430 ;
        RECT 2944.065 356.250 2945.245 357.430 ;
        RECT 2945.665 356.250 2946.845 357.430 ;
        RECT 2947.265 356.250 2948.445 357.430 ;
        RECT 2948.865 356.250 2950.045 357.430 ;
        RECT 2950.465 356.250 2951.645 357.430 ;
        RECT 2952.065 356.250 2953.245 357.430 ;
        RECT 2953.665 356.250 2954.845 357.430 ;
        RECT 2955.265 356.250 2956.445 357.430 ;
        RECT 3157.255 309.805 3158.435 310.985 ;
        RECT 2911.020 306.270 2912.200 307.450 ;
        RECT 2912.620 306.270 2913.800 307.450 ;
        RECT 2942.465 306.250 2943.645 307.430 ;
        RECT 2944.065 306.250 2945.245 307.430 ;
        RECT 2945.665 306.250 2946.845 307.430 ;
        RECT 2947.265 306.250 2948.445 307.430 ;
        RECT 2948.865 306.250 2950.045 307.430 ;
        RECT 2950.465 306.250 2951.645 307.430 ;
        RECT 2952.065 306.250 2953.245 307.430 ;
        RECT 2953.665 306.250 2954.845 307.430 ;
        RECT 2955.265 306.250 2956.445 307.430 ;
        RECT 3157.255 308.205 3158.435 309.385 ;
        RECT 3157.255 306.605 3158.435 307.785 ;
        RECT 3172.725 309.825 3173.905 311.005 ;
        RECT 3172.725 308.225 3173.905 309.405 ;
        RECT 3172.725 306.625 3173.905 307.805 ;
        RECT 3188.265 309.845 3189.445 311.025 ;
        RECT 3188.265 308.245 3189.445 309.425 ;
        RECT 3188.265 306.645 3189.445 307.825 ;
        RECT 3203.785 309.805 3204.965 310.985 ;
        RECT 3203.785 308.205 3204.965 309.385 ;
        RECT 3203.785 306.605 3204.965 307.785 ;
        RECT 3219.295 309.935 3220.475 311.115 ;
        RECT 3219.295 308.335 3220.475 309.515 ;
        RECT 3219.295 306.735 3220.475 307.915 ;
        RECT 3241.445 233.870 3242.625 235.050 ;
        RECT 3243.045 233.870 3244.225 235.050 ;
        RECT 3244.645 233.870 3245.825 235.050 ;
        RECT 3246.245 233.870 3247.425 235.050 ;
        RECT 707.640 221.590 713.620 225.970 ;
        RECT 1209.125 214.255 1229.505 233.035 ;
        RECT 1257.385 214.325 1277.765 233.105 ;
      LAYER met5 ;
        RECT 239.180 1058.490 254.180 1188.060 ;
        RECT 281.440 1172.330 2956.950 1187.330 ;
        RECT 2941.950 1130.420 2956.950 1172.330 ;
        RECT 2941.950 1120.960 3201.830 1130.420 ;
        RECT 2941.950 1120.410 3209.990 1120.960 ;
        RECT 239.180 1055.290 266.160 1058.490 ;
        RECT 2873.230 1055.290 2914.550 1058.490 ;
        RECT 239.180 1008.490 254.180 1055.290 ;
        RECT 2911.350 1042.510 2914.550 1055.290 ;
        RECT 2911.350 1039.310 2918.710 1042.510 ;
        RECT 2941.950 1036.400 2956.950 1120.410 ;
        RECT 3197.330 1119.360 3209.990 1120.410 ;
        RECT 2941.950 1034.800 2967.970 1036.400 ;
        RECT 239.180 1005.290 266.160 1008.490 ;
        RECT 2873.230 1005.290 2914.550 1008.490 ;
        RECT 239.180 958.490 254.180 1005.290 ;
        RECT 239.180 955.290 266.160 958.490 ;
        RECT 2873.230 955.290 2914.550 958.490 ;
        RECT 2941.950 958.200 2956.950 1034.800 ;
        RECT 2941.950 956.600 2967.970 958.200 ;
        RECT 239.180 908.490 254.180 955.290 ;
        RECT 239.180 905.290 266.160 908.490 ;
        RECT 2873.230 905.290 2914.550 908.490 ;
        RECT 239.180 858.490 254.180 905.290 ;
        RECT 2941.950 880.000 2956.950 956.600 ;
        RECT 2941.950 878.400 2967.970 880.000 ;
        RECT 239.180 855.290 266.160 858.490 ;
        RECT 2873.230 855.290 2914.550 858.490 ;
        RECT 239.180 833.940 254.180 855.290 ;
        RECT 234.180 808.490 254.180 833.940 ;
        RECT 234.180 805.290 266.160 808.490 ;
        RECT 2873.230 805.290 2914.550 808.490 ;
        RECT 234.180 758.490 254.180 805.290 ;
        RECT 2941.950 801.800 2956.950 878.400 ;
        RECT 2941.950 800.200 2967.970 801.800 ;
        RECT 234.180 755.290 266.160 758.490 ;
        RECT 2873.230 755.290 2914.550 758.490 ;
        RECT 234.180 708.490 254.180 755.290 ;
        RECT 2941.950 723.600 2956.950 800.200 ;
        RECT 2941.950 722.000 2967.970 723.600 ;
        RECT 234.180 705.290 266.160 708.490 ;
        RECT 2873.230 705.290 2914.550 708.490 ;
        RECT 234.180 658.490 254.180 705.290 ;
        RECT 234.180 655.290 266.160 658.490 ;
        RECT 2873.230 655.290 2914.550 658.490 ;
        RECT 234.180 608.490 254.180 655.290 ;
        RECT 2941.950 645.400 2956.950 722.000 ;
        RECT 2941.950 643.800 2967.970 645.400 ;
        RECT 234.180 605.290 266.160 608.490 ;
        RECT 2873.230 605.290 2914.550 608.490 ;
        RECT 234.180 558.490 254.180 605.290 ;
        RECT 2941.950 567.200 2956.950 643.800 ;
        RECT 2941.950 565.600 2968.050 567.200 ;
        RECT 234.180 555.290 266.160 558.490 ;
        RECT 2873.230 555.290 2914.550 558.490 ;
        RECT 234.180 508.490 254.180 555.290 ;
        RECT 234.180 505.290 266.160 508.490 ;
        RECT 2873.230 505.290 2914.550 508.490 ;
        RECT 234.180 458.490 254.180 505.290 ;
        RECT 2941.950 494.780 2956.950 565.600 ;
        RECT 2941.950 479.780 3297.965 494.780 ;
        RECT 234.180 455.290 266.160 458.490 ;
        RECT 2873.230 455.290 2914.550 458.490 ;
        RECT 234.180 408.490 254.180 455.290 ;
        RECT 234.180 405.290 266.160 408.490 ;
        RECT 2873.230 405.290 2914.550 408.490 ;
        RECT 234.180 358.490 254.180 405.290 ;
        RECT 234.180 355.290 266.160 358.490 ;
        RECT 2873.230 355.290 2914.550 358.490 ;
        RECT 234.180 308.490 254.180 355.290 ;
        RECT 234.180 305.290 266.160 308.490 ;
        RECT 2873.230 305.290 2914.550 308.490 ;
        RECT 234.180 233.940 254.180 305.290 ;
        RECT 2941.950 235.940 2956.950 479.780 ;
        RECT 3124.120 447.370 3139.120 479.780 ;
        RECT 3254.970 462.950 3269.970 479.780 ;
        RECT 3254.970 461.350 3288.770 462.950 ;
        RECT 3254.970 454.790 3269.970 461.350 ;
        RECT 3254.970 453.190 3288.920 454.790 ;
        RECT 3254.970 452.610 3269.970 453.190 ;
        RECT 3124.120 445.770 3146.810 447.370 ;
        RECT 3124.120 445.060 3139.120 445.770 ;
        RECT 3128.090 379.340 3135.170 445.060 ;
        RECT 3128.090 374.340 3220.940 379.340 ;
        RECT 3128.090 358.980 3132.090 374.340 ;
        RECT 3128.090 357.380 3134.840 358.980 ;
        RECT 3128.090 342.080 3132.090 357.380 ;
        RECT 3128.090 340.480 3134.840 342.080 ;
        RECT 3128.090 311.370 3132.090 340.480 ;
        RECT 3128.090 306.370 3220.940 311.370 ;
        RECT 2941.950 233.940 3248.340 235.940 ;
        RECT 234.180 232.940 3248.340 233.940 ;
        RECT 234.180 213.940 2956.980 232.940 ;
    END
  END vssd_core
  PIN vccd2_core
    PORT
      LAYER met4 ;
        RECT 306.910 1342.690 310.010 1379.380 ;
        RECT 306.910 1339.590 326.260 1342.690 ;
        RECT 323.160 1207.330 326.260 1339.590 ;
        RECT 220.980 1192.330 326.260 1207.330 ;
        RECT 974.410 1192.330 976.070 1207.320 ;
        RECT 1025.010 1192.330 1026.670 1207.320 ;
        RECT 220.980 1172.330 234.010 1192.330 ;
        RECT 323.160 1192.000 326.260 1192.330 ;
        RECT 3262.690 1191.330 3265.790 1379.380 ;
      LAYER via4 ;
        RECT 222.040 1173.135 232.820 1206.315 ;
        RECT 282.830 1193.695 316.010 1206.075 ;
        RECT 324.065 1205.650 325.245 1206.830 ;
        RECT 324.065 1204.050 325.245 1205.230 ;
        RECT 324.065 1202.450 325.245 1203.630 ;
        RECT 324.065 1200.850 325.245 1202.030 ;
        RECT 324.065 1199.250 325.245 1200.430 ;
        RECT 324.065 1197.650 325.245 1198.830 ;
        RECT 324.065 1196.050 325.245 1197.230 ;
        RECT 324.065 1194.450 325.245 1195.630 ;
        RECT 324.065 1192.850 325.245 1194.030 ;
        RECT 974.650 1205.685 975.830 1206.865 ;
        RECT 974.650 1204.085 975.830 1205.265 ;
        RECT 974.650 1202.485 975.830 1203.665 ;
        RECT 974.650 1200.885 975.830 1202.065 ;
        RECT 974.650 1199.285 975.830 1200.465 ;
        RECT 974.650 1197.685 975.830 1198.865 ;
        RECT 974.650 1196.085 975.830 1197.265 ;
        RECT 974.650 1194.485 975.830 1195.665 ;
        RECT 974.650 1192.885 975.830 1194.065 ;
        RECT 1025.250 1205.685 1026.430 1206.865 ;
        RECT 1025.250 1204.085 1026.430 1205.265 ;
        RECT 1025.250 1202.485 1026.430 1203.665 ;
        RECT 1025.250 1200.885 1026.430 1202.065 ;
        RECT 1025.250 1199.285 1026.430 1200.465 ;
        RECT 1025.250 1197.685 1026.430 1198.865 ;
        RECT 1025.250 1196.085 1026.430 1197.265 ;
        RECT 1025.250 1194.485 1026.430 1195.665 ;
        RECT 1025.250 1192.885 1026.430 1194.065 ;
        RECT 3263.605 1205.675 3264.785 1206.855 ;
        RECT 3263.605 1204.075 3264.785 1205.255 ;
        RECT 3263.605 1202.475 3264.785 1203.655 ;
        RECT 3263.605 1200.875 3264.785 1202.055 ;
        RECT 3263.605 1199.275 3264.785 1200.455 ;
        RECT 3263.605 1197.675 3264.785 1198.855 ;
        RECT 3263.605 1196.075 3264.785 1197.255 ;
        RECT 3263.605 1194.475 3264.785 1195.655 ;
        RECT 3263.605 1192.875 3264.785 1194.055 ;
      LAYER met5 ;
        RECT 221.270 1172.660 233.590 1206.790 ;
        RECT 281.390 1192.330 3266.530 1207.330 ;
    END
  END vccd2_core
  PIN vssd2_core
    PORT
      LAYER met4 ;
        RECT 302.110 1337.890 305.210 1374.610 ;
        RECT 302.110 1334.790 321.460 1337.890 ;
        RECT 318.360 1227.330 321.460 1334.790 ;
        RECT 204.920 1212.330 321.460 1227.330 ;
        RECT 995.310 1212.330 996.970 1227.320 ;
        RECT 1045.610 1212.340 1047.270 1227.330 ;
        RECT 204.920 1191.330 218.060 1212.330 ;
        RECT 318.360 1211.790 321.460 1212.330 ;
        RECT 3267.490 1211.810 3270.590 1374.580 ;
      LAYER via4 ;
        RECT 206.100 1191.985 216.880 1226.765 ;
        RECT 282.755 1213.525 315.935 1225.905 ;
        RECT 319.315 1225.670 320.495 1226.850 ;
        RECT 319.315 1224.070 320.495 1225.250 ;
        RECT 319.315 1222.470 320.495 1223.650 ;
        RECT 319.315 1220.870 320.495 1222.050 ;
        RECT 319.315 1219.270 320.495 1220.450 ;
        RECT 319.315 1217.670 320.495 1218.850 ;
        RECT 319.315 1216.070 320.495 1217.250 ;
        RECT 319.315 1214.470 320.495 1215.650 ;
        RECT 319.315 1212.870 320.495 1214.050 ;
        RECT 995.550 1225.685 996.730 1226.865 ;
        RECT 995.550 1224.085 996.730 1225.265 ;
        RECT 995.550 1222.485 996.730 1223.665 ;
        RECT 995.550 1220.885 996.730 1222.065 ;
        RECT 995.550 1219.285 996.730 1220.465 ;
        RECT 995.550 1217.685 996.730 1218.865 ;
        RECT 995.550 1216.085 996.730 1217.265 ;
        RECT 995.550 1214.485 996.730 1215.665 ;
        RECT 995.550 1212.885 996.730 1214.065 ;
        RECT 1045.850 1225.695 1047.030 1226.875 ;
        RECT 1045.850 1224.095 1047.030 1225.275 ;
        RECT 1045.850 1222.495 1047.030 1223.675 ;
        RECT 1045.850 1220.895 1047.030 1222.075 ;
        RECT 1045.850 1219.295 1047.030 1220.475 ;
        RECT 1045.850 1217.695 1047.030 1218.875 ;
        RECT 1045.850 1216.095 1047.030 1217.275 ;
        RECT 1045.850 1214.495 1047.030 1215.675 ;
        RECT 1045.850 1212.895 1047.030 1214.075 ;
        RECT 3268.395 1225.685 3269.575 1226.865 ;
        RECT 3268.395 1224.085 3269.575 1225.265 ;
        RECT 3268.395 1222.485 3269.575 1223.665 ;
        RECT 3268.395 1220.885 3269.575 1222.065 ;
        RECT 3268.395 1219.285 3269.575 1220.465 ;
        RECT 3268.395 1217.685 3269.575 1218.865 ;
        RECT 3268.395 1216.085 3269.575 1217.265 ;
        RECT 3268.395 1214.485 3269.575 1215.665 ;
        RECT 3268.395 1212.885 3269.575 1214.065 ;
      LAYER met5 ;
        RECT 205.330 1191.810 217.650 1226.940 ;
        RECT 281.390 1212.330 3271.110 1227.330 ;
    END
  END vssd2_core
  PIN vdda2_core
    PORT
      LAYER met3 ;
        RECT 199.620 2465.390 261.460 2489.290 ;
        RECT 199.620 2415.495 261.460 2439.395 ;
      LAYER via3 ;
        RECT 251.980 2466.295 260.300 2488.615 ;
        RECT 251.920 2416.345 260.240 2438.665 ;
      LAYER met4 ;
        RECT 250.970 4943.680 282.170 4946.740 ;
        RECT 250.860 2465.420 260.980 2489.370 ;
        RECT 250.990 2415.470 261.110 2439.420 ;
        RECT 250.930 1363.190 260.990 1367.190 ;
        RECT 250.930 1360.130 282.030 1363.190 ;
        RECT 287.710 1323.490 290.810 1360.210 ;
        RECT 287.710 1320.390 307.060 1323.490 ;
        RECT 303.960 1287.330 307.060 1320.390 ;
        RECT 250.850 1272.330 307.060 1287.330 ;
        RECT 303.960 1272.110 307.060 1272.330 ;
        RECT 1922.930 1272.260 1928.540 1287.350 ;
        RECT 1998.430 1272.260 2004.040 1287.350 ;
        RECT 3281.890 1271.930 3284.990 1360.180 ;
      LAYER via4 ;
        RECT 251.400 4944.625 252.580 4945.805 ;
        RECT 253.000 4944.625 254.180 4945.805 ;
        RECT 254.600 4944.625 255.780 4945.805 ;
        RECT 256.200 4944.625 257.380 4945.805 ;
        RECT 257.800 4944.625 258.980 4945.805 ;
        RECT 259.400 4944.625 260.580 4945.805 ;
        RECT 279.165 4944.650 280.345 4945.830 ;
        RECT 280.765 4944.650 281.945 4945.830 ;
        RECT 252.350 2466.465 259.930 2488.445 ;
        RECT 252.290 2416.515 259.870 2438.495 ;
        RECT 251.365 1360.680 260.545 1366.660 ;
        RECT 279.010 1360.285 281.790 1363.065 ;
        RECT 252.355 1273.845 259.935 1286.225 ;
        RECT 282.820 1273.540 301.600 1285.920 ;
        RECT 304.900 1285.630 306.080 1286.810 ;
        RECT 304.900 1284.030 306.080 1285.210 ;
        RECT 304.900 1282.430 306.080 1283.610 ;
        RECT 304.900 1280.830 306.080 1282.010 ;
        RECT 304.900 1279.230 306.080 1280.410 ;
        RECT 304.900 1277.630 306.080 1278.810 ;
        RECT 304.900 1276.030 306.080 1277.210 ;
        RECT 304.900 1274.430 306.080 1275.610 ;
        RECT 304.900 1272.830 306.080 1274.010 ;
        RECT 1923.575 1272.850 1927.955 1286.830 ;
        RECT 1999.075 1272.850 2003.455 1286.830 ;
        RECT 3282.805 1285.595 3283.985 1286.775 ;
        RECT 3282.805 1283.995 3283.985 1285.175 ;
        RECT 3282.805 1282.395 3283.985 1283.575 ;
        RECT 3282.805 1280.795 3283.985 1281.975 ;
        RECT 3282.805 1279.195 3283.985 1280.375 ;
        RECT 3282.805 1277.595 3283.985 1278.775 ;
        RECT 3282.805 1275.995 3283.985 1277.175 ;
        RECT 3282.805 1274.395 3283.985 1275.575 ;
        RECT 3282.805 1272.795 3283.985 1273.975 ;
      LAYER met5 ;
        RECT 250.990 1272.490 260.990 4952.330 ;
        RECT 278.880 4943.640 287.760 4946.740 ;
        RECT 278.770 1360.120 287.730 1363.220 ;
        RECT 281.850 1272.330 3285.380 1287.330 ;
    END
  END vdda2_core
  PIN vssa2_core
    PORT
      LAYER met3 ;
        RECT 199.260 4188.390 250.010 4212.290 ;
        RECT 199.260 4138.495 250.010 4162.395 ;
      LAYER via3 ;
        RECT 239.645 4189.150 248.365 4211.470 ;
        RECT 239.645 4139.490 248.365 4161.810 ;
      LAYER met4 ;
        RECT 238.980 4948.460 282.910 4951.550 ;
        RECT 238.960 4188.290 249.110 4212.310 ;
        RECT 238.960 4138.510 249.110 4162.530 ;
        RECT 238.960 1355.410 283.080 1358.440 ;
        RECT 238.960 1355.290 286.010 1355.410 ;
        RECT 238.960 1351.290 249.010 1355.290 ;
        RECT 282.860 1307.330 286.010 1355.290 ;
        RECT 238.850 1292.330 297.350 1307.330 ;
        RECT 1959.720 1292.340 1964.230 1307.250 ;
        RECT 2035.320 1292.340 2039.830 1307.250 ;
        RECT 3286.690 1291.950 3289.790 1355.410 ;
      LAYER via4 ;
        RECT 239.370 4949.445 240.550 4950.625 ;
        RECT 240.970 4949.445 242.150 4950.625 ;
        RECT 242.570 4949.445 243.750 4950.625 ;
        RECT 244.170 4949.445 245.350 4950.625 ;
        RECT 245.770 4949.445 246.950 4950.625 ;
        RECT 247.370 4949.445 248.550 4950.625 ;
        RECT 279.145 4949.450 280.325 4950.630 ;
        RECT 280.745 4949.450 281.925 4950.630 ;
        RECT 240.215 4189.320 247.795 4211.300 ;
        RECT 240.215 4139.660 247.795 4161.640 ;
        RECT 239.395 1351.915 248.575 1357.895 ;
        RECT 279.280 1355.470 282.060 1358.250 ;
        RECT 240.355 1293.845 247.935 1306.225 ;
        RECT 282.775 1293.540 296.755 1305.920 ;
        RECT 1960.585 1293.565 1963.365 1305.945 ;
        RECT 2036.185 1293.565 2038.965 1305.945 ;
        RECT 3287.615 1305.685 3288.795 1306.865 ;
        RECT 3287.615 1304.085 3288.795 1305.265 ;
        RECT 3287.615 1302.485 3288.795 1303.665 ;
        RECT 3287.615 1300.885 3288.795 1302.065 ;
        RECT 3287.615 1299.285 3288.795 1300.465 ;
        RECT 3287.615 1297.685 3288.795 1298.865 ;
        RECT 3287.615 1296.085 3288.795 1297.265 ;
        RECT 3287.615 1294.485 3288.795 1295.665 ;
        RECT 3287.615 1292.885 3288.795 1294.065 ;
      LAYER met5 ;
        RECT 238.990 1292.420 248.990 4952.330 ;
        RECT 278.880 4948.440 282.980 4951.540 ;
        RECT 278.770 1355.320 282.950 1358.420 ;
        RECT 281.850 1292.330 3290.450 1307.330 ;
    END
  END vssa2_core
  PIN vssd1_core
    PORT
      LAYER met3 ;
        RECT 565.910 4977.510 571.910 5152.410 ;
        RECT 822.910 4977.510 828.910 5152.410 ;
        RECT 1079.910 4977.510 1085.910 5152.410 ;
        RECT 1336.910 4977.510 1342.910 5152.410 ;
        RECT 1594.910 4977.510 1600.910 5152.410 ;
        RECT 1846.910 4977.510 1852.910 5152.410 ;
        RECT 2183.910 4977.510 2189.910 5152.410 ;
        RECT 2568.910 4977.510 2574.910 5152.410 ;
        RECT 2825.910 4977.510 2831.910 5152.410 ;
        RECT 36.180 4740.910 283.050 4741.910 ;
        RECT 36.180 4735.910 314.720 4740.910 ;
        RECT 277.160 4734.910 314.720 4735.910 ;
        RECT 36.180 4106.910 314.720 4112.910 ;
        RECT 36.180 3890.910 314.720 3896.910 ;
        RECT 36.180 3674.910 314.720 3680.910 ;
        RECT 36.180 3458.910 314.720 3464.910 ;
        RECT 36.180 3242.910 314.720 3248.910 ;
        RECT 36.180 3026.910 314.720 3032.910 ;
        RECT 36.180 2810.910 314.720 2816.910 ;
        RECT 36.180 2172.910 314.720 2178.910 ;
        RECT 36.180 1956.910 314.720 1962.910 ;
        RECT 36.180 1740.910 314.720 1746.910 ;
        RECT 36.180 1524.910 314.720 1530.910 ;
        RECT 36.180 1308.910 269.080 1314.910 ;
        RECT 36.180 1092.910 269.080 1098.910 ;
      LAYER via3 ;
        RECT 566.140 5148.340 571.710 5151.840 ;
        RECT 566.150 4977.920 571.640 4983.330 ;
        RECT 823.140 5148.340 828.710 5151.840 ;
        RECT 823.150 4977.920 828.640 4983.330 ;
        RECT 1080.140 5148.340 1085.710 5151.840 ;
        RECT 1080.150 4977.920 1085.640 4983.330 ;
        RECT 1337.140 5148.340 1342.710 5151.840 ;
        RECT 1337.150 4977.920 1342.640 4983.330 ;
        RECT 1595.140 5148.340 1600.710 5151.840 ;
        RECT 1595.150 4977.920 1600.640 4983.330 ;
        RECT 1847.140 5148.340 1852.710 5151.840 ;
        RECT 1847.150 4977.920 1852.640 4983.330 ;
        RECT 2184.140 5148.340 2189.710 5151.840 ;
        RECT 2184.150 4977.920 2189.640 4983.330 ;
        RECT 2569.140 5148.340 2574.710 5151.840 ;
        RECT 2569.150 4977.920 2574.640 4983.330 ;
        RECT 2826.140 5148.340 2831.710 5151.840 ;
        RECT 2826.150 4977.920 2831.640 4983.330 ;
        RECT 36.750 4736.140 40.250 4741.710 ;
        RECT 263.260 4736.150 268.670 4741.640 ;
        RECT 312.055 4735.085 314.375 4740.605 ;
        RECT 36.750 4107.140 40.250 4112.710 ;
        RECT 263.260 4107.150 268.670 4112.640 ;
        RECT 312.055 4107.085 314.375 4112.605 ;
        RECT 36.750 3891.140 40.250 3896.710 ;
        RECT 263.260 3891.150 268.670 3896.640 ;
        RECT 312.055 3891.085 314.375 3896.605 ;
        RECT 36.750 3675.140 40.250 3680.710 ;
        RECT 263.260 3675.150 268.670 3680.640 ;
        RECT 312.055 3675.085 314.375 3680.605 ;
        RECT 36.750 3459.140 40.250 3464.710 ;
        RECT 263.260 3459.150 268.670 3464.640 ;
        RECT 312.055 3459.085 314.375 3464.605 ;
        RECT 36.750 3243.140 40.250 3248.710 ;
        RECT 263.260 3243.150 268.670 3248.640 ;
        RECT 312.055 3243.085 314.375 3248.605 ;
        RECT 36.750 3027.140 40.250 3032.710 ;
        RECT 263.260 3027.150 268.670 3032.640 ;
        RECT 312.055 3027.085 314.375 3032.605 ;
        RECT 36.750 2811.140 40.250 2816.710 ;
        RECT 263.260 2811.150 268.670 2816.640 ;
        RECT 312.055 2811.085 314.375 2816.605 ;
        RECT 36.750 2173.140 40.250 2178.710 ;
        RECT 263.260 2173.150 268.670 2178.640 ;
        RECT 312.055 2173.085 314.375 2178.605 ;
        RECT 36.750 1957.140 40.250 1962.710 ;
        RECT 263.260 1957.150 268.670 1962.640 ;
        RECT 312.055 1957.085 314.375 1962.605 ;
        RECT 36.750 1741.140 40.250 1746.710 ;
        RECT 263.260 1741.150 268.670 1746.640 ;
        RECT 312.055 1741.085 314.375 1746.605 ;
        RECT 36.750 1525.140 40.250 1530.710 ;
        RECT 263.260 1525.150 268.670 1530.640 ;
        RECT 312.055 1525.085 314.375 1530.605 ;
        RECT 36.750 1309.140 40.250 1314.710 ;
        RECT 263.260 1309.150 268.670 1314.640 ;
        RECT 36.750 1093.140 40.250 1098.710 ;
        RECT 263.260 1093.150 268.670 1098.640 ;
      LAYER met4 ;
        RECT 505.380 5148.060 572.210 5152.060 ;
        RECT 762.380 5148.060 829.210 5152.060 ;
        RECT 1019.380 5148.060 1086.210 5152.060 ;
        RECT 1276.380 5148.060 1343.210 5152.060 ;
        RECT 1534.380 5148.060 1601.210 5152.060 ;
        RECT 1786.380 5148.060 1853.210 5152.060 ;
        RECT 2123.380 5148.060 2190.210 5152.060 ;
        RECT 2508.380 5148.060 2575.210 5152.060 ;
        RECT 2765.380 5148.060 2832.210 5152.060 ;
        RECT 565.870 4977.660 571.940 4983.690 ;
        RECT 822.870 4977.660 828.940 4983.690 ;
        RECT 1079.870 4977.660 1085.940 4983.690 ;
        RECT 1336.870 4977.660 1342.940 4983.690 ;
        RECT 1594.870 4977.660 1600.940 4983.690 ;
        RECT 1846.870 4977.660 1852.940 4983.690 ;
        RECT 2183.870 4977.660 2189.940 4983.690 ;
        RECT 2568.870 4977.660 2574.940 4983.690 ;
        RECT 2825.870 4977.660 2831.940 4983.690 ;
        RECT 3354.080 4983.460 3367.130 4983.480 ;
        RECT 3354.040 4977.460 3383.270 4983.460 ;
        RECT 3354.080 4951.000 3367.130 4977.460 ;
        RECT 262.980 4919.640 282.020 4922.740 ;
        RECT 36.530 4675.380 40.530 4742.210 ;
        RECT 262.900 4735.870 268.930 4741.940 ;
        RECT 311.910 4735.070 314.520 4740.620 ;
        RECT 36.530 4046.380 40.530 4113.210 ;
        RECT 262.900 4106.870 268.930 4112.940 ;
        RECT 311.910 4107.070 314.520 4112.620 ;
        RECT 36.530 3830.380 40.530 3897.210 ;
        RECT 262.900 3890.870 268.930 3896.940 ;
        RECT 311.910 3891.070 314.520 3896.620 ;
        RECT 36.530 3614.380 40.530 3681.210 ;
        RECT 262.900 3674.870 268.930 3680.940 ;
        RECT 311.910 3675.070 314.520 3680.620 ;
        RECT 36.530 3398.380 40.530 3465.210 ;
        RECT 262.900 3458.870 268.930 3464.940 ;
        RECT 311.910 3459.070 314.520 3464.620 ;
        RECT 36.530 3182.380 40.530 3249.210 ;
        RECT 262.900 3242.870 268.930 3248.940 ;
        RECT 311.910 3243.070 314.520 3248.620 ;
        RECT 36.530 2966.380 40.530 3033.210 ;
        RECT 262.900 3026.870 268.930 3032.940 ;
        RECT 311.910 3027.070 314.520 3032.620 ;
        RECT 36.530 2750.380 40.530 2817.210 ;
        RECT 262.900 2810.870 268.930 2816.940 ;
        RECT 311.910 2811.070 314.520 2816.620 ;
        RECT 36.530 2112.380 40.530 2179.210 ;
        RECT 262.900 2172.870 268.930 2178.940 ;
        RECT 311.910 2173.070 314.520 2178.620 ;
        RECT 36.530 1896.380 40.530 1963.210 ;
        RECT 262.900 1956.870 268.930 1962.940 ;
        RECT 311.910 1957.070 314.520 1962.620 ;
        RECT 36.530 1680.380 40.530 1747.210 ;
        RECT 262.900 1740.870 268.930 1746.940 ;
        RECT 311.910 1741.070 314.520 1746.620 ;
        RECT 36.530 1464.380 40.530 1531.210 ;
        RECT 262.900 1524.870 268.930 1530.940 ;
        RECT 311.910 1525.070 314.520 1530.620 ;
        RECT 262.910 1387.230 269.000 1390.230 ;
        RECT 262.910 1384.110 282.080 1387.230 ;
        RECT 311.710 1347.490 314.810 1384.170 ;
        RECT 311.710 1344.390 331.060 1347.490 ;
        RECT 36.530 1248.380 40.530 1315.210 ;
        RECT 262.900 1308.870 268.930 1314.940 ;
        RECT 262.890 1252.330 316.460 1267.330 ;
        RECT 327.960 1251.930 331.060 1344.390 ;
        RECT 1383.610 1252.350 1386.300 1267.360 ;
        RECT 1458.610 1252.350 1461.300 1267.360 ;
        RECT 1533.810 1252.350 1536.500 1267.360 ;
        RECT 1609.410 1252.350 1612.100 1267.360 ;
        RECT 3257.890 1251.960 3260.990 1384.220 ;
        RECT 36.530 1032.380 40.530 1099.210 ;
        RECT 262.900 1092.870 268.930 1098.940 ;
      LAYER via4 ;
        RECT 505.640 5148.140 507.130 5152.010 ;
        RECT 522.590 5148.160 524.010 5151.990 ;
        RECT 539.470 5148.150 540.890 5151.980 ;
        RECT 762.640 5148.140 764.130 5152.010 ;
        RECT 779.590 5148.160 781.010 5151.990 ;
        RECT 796.470 5148.150 797.890 5151.980 ;
        RECT 1019.640 5148.140 1021.130 5152.010 ;
        RECT 1036.590 5148.160 1038.010 5151.990 ;
        RECT 1053.470 5148.150 1054.890 5151.980 ;
        RECT 1276.640 5148.140 1278.130 5152.010 ;
        RECT 1293.590 5148.160 1295.010 5151.990 ;
        RECT 1310.470 5148.150 1311.890 5151.980 ;
        RECT 1534.640 5148.140 1536.130 5152.010 ;
        RECT 1551.590 5148.160 1553.010 5151.990 ;
        RECT 1568.470 5148.150 1569.890 5151.980 ;
        RECT 1786.640 5148.140 1788.130 5152.010 ;
        RECT 1803.590 5148.160 1805.010 5151.990 ;
        RECT 1820.470 5148.150 1821.890 5151.980 ;
        RECT 2123.640 5148.140 2125.130 5152.010 ;
        RECT 2140.590 5148.160 2142.010 5151.990 ;
        RECT 2157.470 5148.150 2158.890 5151.980 ;
        RECT 2508.640 5148.140 2510.130 5152.010 ;
        RECT 2525.590 5148.160 2527.010 5151.990 ;
        RECT 2542.470 5148.150 2543.890 5151.980 ;
        RECT 2765.640 5148.140 2767.130 5152.010 ;
        RECT 2782.590 5148.160 2784.010 5151.990 ;
        RECT 2799.470 5148.150 2800.890 5151.980 ;
        RECT 566.150 4977.920 571.640 4983.330 ;
        RECT 823.150 4977.920 828.640 4983.330 ;
        RECT 1080.150 4977.920 1085.640 4983.330 ;
        RECT 1337.150 4977.920 1342.640 4983.330 ;
        RECT 1595.150 4977.920 1600.640 4983.330 ;
        RECT 1847.150 4977.920 1852.640 4983.330 ;
        RECT 2184.150 4977.920 2189.640 4983.330 ;
        RECT 2569.150 4977.920 2574.640 4983.330 ;
        RECT 2826.150 4977.920 2831.640 4983.330 ;
        RECT 3355.180 4978.340 3381.960 4982.720 ;
        RECT 3355.210 4951.820 3365.990 4962.600 ;
        RECT 263.795 4920.605 264.975 4921.785 ;
        RECT 265.395 4920.605 266.575 4921.785 ;
        RECT 266.995 4920.605 268.175 4921.785 ;
        RECT 279.055 4919.805 281.835 4922.585 ;
        RECT 263.260 4736.150 268.670 4741.640 ;
        RECT 36.590 4709.440 40.460 4710.930 ;
        RECT 36.600 4692.590 40.460 4693.980 ;
        RECT 36.580 4675.640 40.450 4677.130 ;
        RECT 263.260 4107.150 268.670 4112.640 ;
        RECT 36.590 4080.440 40.460 4081.930 ;
        RECT 36.600 4063.590 40.460 4064.980 ;
        RECT 36.580 4046.640 40.450 4048.130 ;
        RECT 263.260 3891.150 268.670 3896.640 ;
        RECT 36.590 3864.440 40.460 3865.930 ;
        RECT 36.600 3847.590 40.460 3848.980 ;
        RECT 36.580 3830.640 40.450 3832.130 ;
        RECT 263.260 3675.150 268.670 3680.640 ;
        RECT 36.590 3648.440 40.460 3649.930 ;
        RECT 36.600 3631.590 40.460 3632.980 ;
        RECT 36.580 3614.640 40.450 3616.130 ;
        RECT 263.260 3459.150 268.670 3464.640 ;
        RECT 36.590 3432.440 40.460 3433.930 ;
        RECT 36.600 3415.590 40.460 3416.980 ;
        RECT 36.580 3398.640 40.450 3400.130 ;
        RECT 263.260 3243.150 268.670 3248.640 ;
        RECT 36.590 3216.440 40.460 3217.930 ;
        RECT 36.600 3199.590 40.460 3200.980 ;
        RECT 36.580 3182.640 40.450 3184.130 ;
        RECT 263.260 3027.150 268.670 3032.640 ;
        RECT 36.590 3000.440 40.460 3001.930 ;
        RECT 36.600 2983.590 40.460 2984.980 ;
        RECT 36.580 2966.640 40.450 2968.130 ;
        RECT 263.260 2811.150 268.670 2816.640 ;
        RECT 36.590 2784.440 40.460 2785.930 ;
        RECT 36.600 2767.590 40.460 2768.980 ;
        RECT 36.580 2750.640 40.450 2752.130 ;
        RECT 263.260 2173.150 268.670 2178.640 ;
        RECT 36.590 2146.440 40.460 2147.930 ;
        RECT 36.600 2129.590 40.460 2130.980 ;
        RECT 36.580 2112.640 40.450 2114.130 ;
        RECT 263.260 1957.150 268.670 1962.640 ;
        RECT 36.590 1930.440 40.460 1931.930 ;
        RECT 36.600 1913.590 40.460 1914.980 ;
        RECT 36.580 1896.640 40.450 1898.130 ;
        RECT 263.260 1741.150 268.670 1746.640 ;
        RECT 36.590 1714.440 40.460 1715.930 ;
        RECT 36.600 1697.590 40.460 1698.980 ;
        RECT 36.580 1680.640 40.450 1682.130 ;
        RECT 263.260 1525.150 268.670 1530.640 ;
        RECT 36.590 1498.440 40.460 1499.930 ;
        RECT 36.600 1481.590 40.460 1482.980 ;
        RECT 36.580 1464.640 40.450 1466.130 ;
        RECT 263.765 1385.050 268.145 1389.430 ;
        RECT 279.030 1384.295 281.810 1387.075 ;
        RECT 263.260 1309.150 268.670 1314.640 ;
        RECT 36.590 1282.440 40.460 1283.930 ;
        RECT 36.600 1265.590 40.460 1266.980 ;
        RECT 263.810 1252.860 268.190 1266.840 ;
        RECT 281.160 1252.870 315.940 1266.850 ;
        RECT 328.875 1265.610 330.055 1266.790 ;
        RECT 328.875 1264.010 330.055 1265.190 ;
        RECT 328.875 1262.410 330.055 1263.590 ;
        RECT 328.875 1260.810 330.055 1261.990 ;
        RECT 328.875 1259.210 330.055 1260.390 ;
        RECT 328.875 1257.610 330.055 1258.790 ;
        RECT 328.875 1256.010 330.055 1257.190 ;
        RECT 328.875 1254.410 330.055 1255.590 ;
        RECT 328.875 1252.810 330.055 1253.990 ;
        RECT 1384.135 1265.700 1385.315 1266.880 ;
        RECT 1384.135 1264.100 1385.315 1265.280 ;
        RECT 1384.135 1262.500 1385.315 1263.680 ;
        RECT 1384.135 1260.900 1385.315 1262.080 ;
        RECT 1384.135 1259.300 1385.315 1260.480 ;
        RECT 1384.135 1257.700 1385.315 1258.880 ;
        RECT 1384.135 1256.100 1385.315 1257.280 ;
        RECT 1384.135 1254.500 1385.315 1255.680 ;
        RECT 1384.135 1252.900 1385.315 1254.080 ;
        RECT 1459.135 1265.700 1460.315 1266.880 ;
        RECT 1459.135 1264.100 1460.315 1265.280 ;
        RECT 1459.135 1262.500 1460.315 1263.680 ;
        RECT 1459.135 1260.900 1460.315 1262.080 ;
        RECT 1459.135 1259.300 1460.315 1260.480 ;
        RECT 1459.135 1257.700 1460.315 1258.880 ;
        RECT 1459.135 1256.100 1460.315 1257.280 ;
        RECT 1459.135 1254.500 1460.315 1255.680 ;
        RECT 1459.135 1252.900 1460.315 1254.080 ;
        RECT 1534.335 1265.700 1535.515 1266.880 ;
        RECT 1534.335 1264.100 1535.515 1265.280 ;
        RECT 1534.335 1262.500 1535.515 1263.680 ;
        RECT 1534.335 1260.900 1535.515 1262.080 ;
        RECT 1534.335 1259.300 1535.515 1260.480 ;
        RECT 1534.335 1257.700 1535.515 1258.880 ;
        RECT 1534.335 1256.100 1535.515 1257.280 ;
        RECT 1534.335 1254.500 1535.515 1255.680 ;
        RECT 1534.335 1252.900 1535.515 1254.080 ;
        RECT 1609.935 1265.700 1611.115 1266.880 ;
        RECT 1609.935 1264.100 1611.115 1265.280 ;
        RECT 1609.935 1262.500 1611.115 1263.680 ;
        RECT 1609.935 1260.900 1611.115 1262.080 ;
        RECT 1609.935 1259.300 1611.115 1260.480 ;
        RECT 1609.935 1257.700 1611.115 1258.880 ;
        RECT 1609.935 1256.100 1611.115 1257.280 ;
        RECT 1609.935 1254.500 1611.115 1255.680 ;
        RECT 1609.935 1252.900 1611.115 1254.080 ;
        RECT 3258.070 1252.805 3260.850 1266.785 ;
        RECT 36.580 1248.640 40.450 1250.130 ;
        RECT 263.260 1093.150 268.670 1098.640 ;
        RECT 36.590 1066.440 40.460 1067.930 ;
        RECT 36.600 1049.590 40.460 1050.980 ;
        RECT 36.580 1032.640 40.450 1034.130 ;
      LAYER met5 ;
        RECT 505.510 5147.980 507.260 5152.140 ;
        RECT 505.590 5145.520 507.190 5147.980 ;
        RECT 522.400 5147.940 524.130 5152.320 ;
        RECT 539.340 5147.970 541.070 5152.350 ;
        RECT 762.510 5147.980 764.260 5152.140 ;
        RECT 522.490 5145.680 524.090 5147.940 ;
        RECT 539.390 5145.680 540.990 5147.970 ;
        RECT 762.590 5145.520 764.190 5147.980 ;
        RECT 779.400 5147.940 781.130 5152.320 ;
        RECT 796.340 5147.970 798.070 5152.350 ;
        RECT 1019.510 5147.980 1021.260 5152.140 ;
        RECT 779.490 5145.680 781.090 5147.940 ;
        RECT 796.390 5145.680 797.990 5147.970 ;
        RECT 1019.590 5145.520 1021.190 5147.980 ;
        RECT 1036.400 5147.940 1038.130 5152.320 ;
        RECT 1053.340 5147.970 1055.070 5152.350 ;
        RECT 1276.510 5147.980 1278.260 5152.140 ;
        RECT 1036.490 5145.680 1038.090 5147.940 ;
        RECT 1053.390 5145.680 1054.990 5147.970 ;
        RECT 1276.590 5145.520 1278.190 5147.980 ;
        RECT 1293.400 5147.940 1295.130 5152.320 ;
        RECT 1310.340 5147.970 1312.070 5152.350 ;
        RECT 1534.510 5147.980 1536.260 5152.140 ;
        RECT 1293.490 5145.680 1295.090 5147.940 ;
        RECT 1310.390 5145.680 1311.990 5147.970 ;
        RECT 1534.590 5145.520 1536.190 5147.980 ;
        RECT 1551.400 5147.940 1553.130 5152.320 ;
        RECT 1568.340 5147.970 1570.070 5152.350 ;
        RECT 1786.510 5147.980 1788.260 5152.140 ;
        RECT 1551.490 5145.680 1553.090 5147.940 ;
        RECT 1568.390 5145.680 1569.990 5147.970 ;
        RECT 1786.590 5145.520 1788.190 5147.980 ;
        RECT 1803.400 5147.940 1805.130 5152.320 ;
        RECT 1820.340 5147.970 1822.070 5152.350 ;
        RECT 2123.510 5147.980 2125.260 5152.140 ;
        RECT 1803.490 5145.680 1805.090 5147.940 ;
        RECT 1820.390 5145.680 1821.990 5147.970 ;
        RECT 2123.590 5145.520 2125.190 5147.980 ;
        RECT 2140.400 5147.940 2142.130 5152.320 ;
        RECT 2157.340 5147.970 2159.070 5152.350 ;
        RECT 2508.510 5147.980 2510.260 5152.140 ;
        RECT 2140.490 5145.680 2142.090 5147.940 ;
        RECT 2157.390 5145.680 2158.990 5147.970 ;
        RECT 2508.590 5145.520 2510.190 5147.980 ;
        RECT 2525.400 5147.940 2527.130 5152.320 ;
        RECT 2542.340 5147.970 2544.070 5152.350 ;
        RECT 2765.510 5147.980 2767.260 5152.140 ;
        RECT 2525.490 5145.680 2527.090 5147.940 ;
        RECT 2542.390 5145.680 2543.990 5147.970 ;
        RECT 2765.590 5145.520 2767.190 5147.980 ;
        RECT 2782.400 5147.940 2784.130 5152.320 ;
        RECT 2799.340 5147.970 2801.070 5152.350 ;
        RECT 2782.490 5145.680 2784.090 5147.940 ;
        RECT 2799.390 5145.680 2800.990 5147.970 ;
        RECT 262.990 4977.510 3383.300 4983.510 ;
        RECT 36.395 4710.990 40.590 4711.095 ;
        RECT 36.300 4709.390 42.910 4710.990 ;
        RECT 36.395 4709.290 40.590 4709.390 ;
        RECT 36.485 4694.090 40.680 4694.205 ;
        RECT 36.330 4692.490 42.910 4694.090 ;
        RECT 36.485 4692.400 40.680 4692.490 ;
        RECT 36.385 4677.190 40.860 4677.265 ;
        RECT 36.385 4675.590 43.070 4677.190 ;
        RECT 36.385 4675.510 40.860 4675.590 ;
        RECT 36.395 4081.990 40.590 4082.095 ;
        RECT 36.300 4080.390 42.910 4081.990 ;
        RECT 36.395 4080.290 40.590 4080.390 ;
        RECT 36.485 4065.090 40.680 4065.205 ;
        RECT 36.330 4063.490 42.910 4065.090 ;
        RECT 36.485 4063.400 40.680 4063.490 ;
        RECT 36.385 4048.190 40.860 4048.265 ;
        RECT 36.385 4046.590 43.070 4048.190 ;
        RECT 36.385 4046.510 40.860 4046.590 ;
        RECT 36.395 3865.990 40.590 3866.095 ;
        RECT 36.300 3864.390 42.910 3865.990 ;
        RECT 36.395 3864.290 40.590 3864.390 ;
        RECT 36.485 3849.090 40.680 3849.205 ;
        RECT 36.330 3847.490 42.910 3849.090 ;
        RECT 36.485 3847.400 40.680 3847.490 ;
        RECT 36.385 3832.190 40.860 3832.265 ;
        RECT 36.385 3830.590 43.070 3832.190 ;
        RECT 36.385 3830.510 40.860 3830.590 ;
        RECT 36.395 3649.990 40.590 3650.095 ;
        RECT 36.300 3648.390 42.910 3649.990 ;
        RECT 36.395 3648.290 40.590 3648.390 ;
        RECT 36.485 3633.090 40.680 3633.205 ;
        RECT 36.330 3631.490 42.910 3633.090 ;
        RECT 36.485 3631.400 40.680 3631.490 ;
        RECT 36.385 3616.190 40.860 3616.265 ;
        RECT 36.385 3614.590 43.070 3616.190 ;
        RECT 36.385 3614.510 40.860 3614.590 ;
        RECT 36.395 3433.990 40.590 3434.095 ;
        RECT 36.300 3432.390 42.910 3433.990 ;
        RECT 36.395 3432.290 40.590 3432.390 ;
        RECT 36.485 3417.090 40.680 3417.205 ;
        RECT 36.330 3415.490 42.910 3417.090 ;
        RECT 36.485 3415.400 40.680 3415.490 ;
        RECT 36.385 3400.190 40.860 3400.265 ;
        RECT 36.385 3398.590 43.070 3400.190 ;
        RECT 36.385 3398.510 40.860 3398.590 ;
        RECT 36.395 3217.990 40.590 3218.095 ;
        RECT 36.300 3216.390 42.910 3217.990 ;
        RECT 36.395 3216.290 40.590 3216.390 ;
        RECT 36.485 3201.090 40.680 3201.205 ;
        RECT 36.330 3199.490 42.910 3201.090 ;
        RECT 36.485 3199.400 40.680 3199.490 ;
        RECT 36.385 3184.190 40.860 3184.265 ;
        RECT 36.385 3182.590 43.070 3184.190 ;
        RECT 36.385 3182.510 40.860 3182.590 ;
        RECT 36.395 3001.990 40.590 3002.095 ;
        RECT 36.300 3000.390 42.910 3001.990 ;
        RECT 36.395 3000.290 40.590 3000.390 ;
        RECT 36.485 2985.090 40.680 2985.205 ;
        RECT 36.330 2983.490 42.910 2985.090 ;
        RECT 36.485 2983.400 40.680 2983.490 ;
        RECT 36.385 2968.190 40.860 2968.265 ;
        RECT 36.385 2966.590 43.070 2968.190 ;
        RECT 36.385 2966.510 40.860 2966.590 ;
        RECT 36.395 2785.990 40.590 2786.095 ;
        RECT 36.300 2784.390 42.910 2785.990 ;
        RECT 36.395 2784.290 40.590 2784.390 ;
        RECT 36.485 2769.090 40.680 2769.205 ;
        RECT 36.330 2767.490 42.910 2769.090 ;
        RECT 36.485 2767.400 40.680 2767.490 ;
        RECT 36.385 2752.190 40.860 2752.265 ;
        RECT 36.385 2750.590 43.070 2752.190 ;
        RECT 36.385 2750.510 40.860 2750.590 ;
        RECT 36.395 2147.990 40.590 2148.095 ;
        RECT 36.300 2146.390 42.910 2147.990 ;
        RECT 36.395 2146.290 40.590 2146.390 ;
        RECT 36.485 2131.090 40.680 2131.205 ;
        RECT 36.330 2129.490 42.910 2131.090 ;
        RECT 36.485 2129.400 40.680 2129.490 ;
        RECT 36.385 2114.190 40.860 2114.265 ;
        RECT 36.385 2112.590 43.070 2114.190 ;
        RECT 36.385 2112.510 40.860 2112.590 ;
        RECT 36.395 1931.990 40.590 1932.095 ;
        RECT 36.300 1930.390 42.910 1931.990 ;
        RECT 36.395 1930.290 40.590 1930.390 ;
        RECT 36.485 1915.090 40.680 1915.205 ;
        RECT 36.330 1913.490 42.910 1915.090 ;
        RECT 36.485 1913.400 40.680 1913.490 ;
        RECT 36.385 1898.190 40.860 1898.265 ;
        RECT 36.385 1896.590 43.070 1898.190 ;
        RECT 36.385 1896.510 40.860 1896.590 ;
        RECT 36.395 1715.990 40.590 1716.095 ;
        RECT 36.300 1714.390 42.910 1715.990 ;
        RECT 36.395 1714.290 40.590 1714.390 ;
        RECT 36.485 1699.090 40.680 1699.205 ;
        RECT 36.330 1697.490 42.910 1699.090 ;
        RECT 36.485 1697.400 40.680 1697.490 ;
        RECT 36.385 1682.190 40.860 1682.265 ;
        RECT 36.385 1680.590 43.070 1682.190 ;
        RECT 36.385 1680.510 40.860 1680.590 ;
        RECT 36.395 1499.990 40.590 1500.095 ;
        RECT 36.300 1498.390 42.910 1499.990 ;
        RECT 36.395 1498.290 40.590 1498.390 ;
        RECT 36.485 1483.090 40.680 1483.205 ;
        RECT 36.330 1481.490 42.910 1483.090 ;
        RECT 36.485 1481.400 40.680 1481.490 ;
        RECT 36.385 1466.190 40.860 1466.265 ;
        RECT 36.385 1464.590 43.070 1466.190 ;
        RECT 36.385 1464.510 40.860 1464.590 ;
        RECT 36.395 1283.990 40.590 1284.095 ;
        RECT 36.300 1282.390 42.910 1283.990 ;
        RECT 36.395 1282.290 40.590 1282.390 ;
        RECT 36.485 1267.090 40.680 1267.205 ;
        RECT 36.330 1265.490 42.910 1267.090 ;
        RECT 36.485 1265.400 40.680 1265.490 ;
        RECT 36.385 1250.190 40.860 1250.265 ;
        RECT 36.385 1248.590 43.070 1250.190 ;
        RECT 36.385 1248.510 40.860 1248.590 ;
        RECT 262.990 1088.710 268.990 4977.510 ;
        RECT 3354.880 4951.770 3366.320 4962.650 ;
        RECT 278.880 4919.640 311.790 4922.740 ;
        RECT 278.770 1384.120 311.760 1387.220 ;
        RECT 280.630 1252.330 3354.930 1267.330 ;
        RECT 36.395 1067.990 40.590 1068.095 ;
        RECT 36.300 1066.390 42.910 1067.990 ;
        RECT 36.395 1066.290 40.590 1066.390 ;
        RECT 36.485 1051.090 40.680 1051.205 ;
        RECT 36.330 1049.490 42.910 1051.090 ;
        RECT 36.485 1049.400 40.680 1049.490 ;
        RECT 36.385 1034.190 40.860 1034.265 ;
        RECT 36.385 1032.590 43.070 1034.190 ;
        RECT 36.385 1032.510 40.860 1032.590 ;
    END
  END vssd1_core
  PIN vccd1_core
    PORT
      LAYER met3 ;
        RECT 573.910 4969.290 579.910 5158.480 ;
        RECT 830.910 4969.290 836.910 5158.480 ;
        RECT 1087.910 4969.290 1093.910 5158.480 ;
        RECT 1344.910 4969.290 1350.910 5158.480 ;
        RECT 1602.910 4969.290 1608.910 5158.480 ;
        RECT 1854.910 4969.290 1860.910 5158.480 ;
        RECT 2191.910 4969.290 2197.910 5158.480 ;
        RECT 2576.910 4969.290 2582.910 5158.480 ;
        RECT 2833.910 4969.290 2839.910 5158.480 ;
        RECT 30.110 4748.410 291.090 4749.910 ;
        RECT 30.110 4743.910 319.610 4748.410 ;
        RECT 285.190 4742.410 319.610 4743.910 ;
        RECT 30.110 4114.910 319.610 4120.910 ;
        RECT 280.390 3904.910 319.610 3910.910 ;
        RECT 30.110 3898.910 286.850 3904.910 ;
        RECT 30.110 3682.910 319.610 3688.910 ;
        RECT 30.110 3466.910 319.610 3472.910 ;
        RECT 30.110 3250.910 319.610 3256.910 ;
        RECT 30.110 3034.910 319.610 3040.910 ;
        RECT 30.110 2818.910 319.610 2824.910 ;
        RECT 30.110 2180.910 319.610 2186.910 ;
        RECT 30.110 1964.910 319.610 1970.910 ;
        RECT 279.840 1754.910 319.610 1758.910 ;
        RECT 30.110 1752.910 319.610 1754.910 ;
        RECT 30.110 1748.910 286.320 1752.910 ;
        RECT 30.110 1532.910 319.610 1538.910 ;
        RECT 30.110 1316.910 277.300 1322.910 ;
        RECT 30.110 1100.910 277.300 1106.910 ;
      LAYER via3 ;
        RECT 574.120 5154.330 579.690 5157.830 ;
        RECT 574.240 4969.950 579.730 4975.360 ;
        RECT 831.120 5154.330 836.690 5157.830 ;
        RECT 831.240 4969.950 836.730 4975.360 ;
        RECT 1088.120 5154.330 1093.690 5157.830 ;
        RECT 1088.240 4969.950 1093.730 4975.360 ;
        RECT 1345.120 5154.330 1350.690 5157.830 ;
        RECT 1345.240 4969.950 1350.730 4975.360 ;
        RECT 1603.120 5154.330 1608.690 5157.830 ;
        RECT 1603.240 4969.950 1608.730 4975.360 ;
        RECT 1855.120 5154.330 1860.690 5157.830 ;
        RECT 1855.240 4969.950 1860.730 4975.360 ;
        RECT 2192.120 5154.330 2197.690 5157.830 ;
        RECT 2192.240 4969.950 2197.730 4975.360 ;
        RECT 2577.120 5154.330 2582.690 5157.830 ;
        RECT 2577.240 4969.950 2582.730 4975.360 ;
        RECT 2834.120 5154.330 2839.690 5157.830 ;
        RECT 2834.240 4969.950 2839.730 4975.360 ;
        RECT 30.760 4744.120 34.260 4749.690 ;
        RECT 271.230 4744.240 276.640 4749.730 ;
        RECT 316.895 4742.625 319.215 4748.145 ;
        RECT 30.760 4115.120 34.260 4120.690 ;
        RECT 271.230 4115.240 276.640 4120.730 ;
        RECT 316.895 4115.125 319.215 4120.645 ;
        RECT 316.895 3905.125 319.215 3910.645 ;
        RECT 30.760 3899.120 34.260 3904.690 ;
        RECT 271.230 3899.240 276.640 3904.730 ;
        RECT 30.760 3683.120 34.260 3688.690 ;
        RECT 271.230 3683.240 276.640 3688.730 ;
        RECT 316.895 3683.125 319.215 3688.645 ;
        RECT 30.760 3467.120 34.260 3472.690 ;
        RECT 271.230 3467.240 276.640 3472.730 ;
        RECT 316.895 3467.125 319.215 3472.645 ;
        RECT 30.760 3251.120 34.260 3256.690 ;
        RECT 271.230 3251.240 276.640 3256.730 ;
        RECT 316.895 3251.125 319.215 3256.645 ;
        RECT 30.760 3035.120 34.260 3040.690 ;
        RECT 271.230 3035.240 276.640 3040.730 ;
        RECT 316.895 3035.125 319.215 3040.645 ;
        RECT 30.760 2819.120 34.260 2824.690 ;
        RECT 271.230 2819.240 276.640 2824.730 ;
        RECT 316.895 2819.125 319.215 2824.645 ;
        RECT 30.760 2181.120 34.260 2186.690 ;
        RECT 271.230 2181.240 276.640 2186.730 ;
        RECT 316.895 2181.125 319.215 2186.645 ;
        RECT 30.760 1965.120 34.260 1970.690 ;
        RECT 271.230 1965.240 276.640 1970.730 ;
        RECT 316.895 1965.125 319.215 1970.645 ;
        RECT 30.760 1749.120 34.260 1754.690 ;
        RECT 271.230 1749.240 276.640 1754.730 ;
        RECT 316.895 1753.125 319.215 1758.645 ;
        RECT 30.760 1533.120 34.260 1538.690 ;
        RECT 271.230 1533.240 276.640 1538.730 ;
        RECT 316.895 1533.125 319.215 1538.645 ;
        RECT 30.760 1317.120 34.260 1322.690 ;
        RECT 271.230 1317.240 276.640 1322.730 ;
        RECT 30.760 1101.120 34.260 1106.690 ;
        RECT 271.230 1101.240 276.640 1106.730 ;
      LAYER met4 ;
        RECT 496.730 5154.060 580.350 5158.060 ;
        RECT 753.730 5154.060 837.350 5158.060 ;
        RECT 1010.730 5154.060 1094.350 5158.060 ;
        RECT 1267.730 5154.060 1351.350 5158.060 ;
        RECT 1525.730 5154.060 1609.350 5158.060 ;
        RECT 1777.730 5154.060 1861.350 5158.060 ;
        RECT 2114.730 5154.060 2198.350 5158.060 ;
        RECT 2499.730 5154.060 2583.350 5158.060 ;
        RECT 2756.730 5154.060 2840.350 5158.060 ;
        RECT 573.870 4969.640 579.940 4975.670 ;
        RECT 830.870 4969.640 836.940 4975.670 ;
        RECT 1087.870 4969.640 1093.940 4975.670 ;
        RECT 1344.870 4969.640 1350.940 4975.670 ;
        RECT 1602.870 4969.640 1608.940 4975.670 ;
        RECT 1854.870 4969.640 1860.940 4975.670 ;
        RECT 2191.870 4969.640 2197.940 4975.670 ;
        RECT 2576.870 4969.640 2582.940 4975.670 ;
        RECT 2833.870 4969.640 2839.940 4975.670 ;
        RECT 30.530 4666.730 34.530 4750.350 ;
        RECT 270.920 4743.870 276.950 4749.940 ;
        RECT 316.750 4742.610 319.360 4748.160 ;
        RECT 30.530 4037.730 34.530 4121.350 ;
        RECT 270.920 4114.870 276.950 4120.940 ;
        RECT 316.750 4115.110 319.360 4120.660 ;
        RECT 30.530 3821.730 34.530 3905.350 ;
        RECT 316.750 3905.110 319.360 3910.660 ;
        RECT 270.920 3898.870 276.950 3904.940 ;
        RECT 30.530 3605.730 34.530 3689.350 ;
        RECT 270.920 3682.870 276.950 3688.940 ;
        RECT 316.750 3683.110 319.360 3688.660 ;
        RECT 30.530 3389.730 34.530 3473.350 ;
        RECT 270.920 3466.870 276.950 3472.940 ;
        RECT 316.750 3467.110 319.360 3472.660 ;
        RECT 30.530 3173.730 34.530 3257.350 ;
        RECT 270.920 3250.870 276.950 3256.940 ;
        RECT 316.750 3251.110 319.360 3256.660 ;
        RECT 30.530 2957.730 34.530 3041.350 ;
        RECT 270.920 3034.870 276.950 3040.940 ;
        RECT 316.750 3035.110 319.360 3040.660 ;
        RECT 30.530 2741.730 34.530 2825.350 ;
        RECT 270.920 2818.870 276.950 2824.940 ;
        RECT 316.750 2819.110 319.360 2824.660 ;
        RECT 30.530 2103.730 34.530 2187.350 ;
        RECT 270.920 2180.870 276.950 2186.940 ;
        RECT 316.750 2181.110 319.360 2186.660 ;
        RECT 30.530 1887.730 34.530 1971.350 ;
        RECT 270.920 1964.870 276.950 1970.940 ;
        RECT 316.750 1965.110 319.360 1970.660 ;
        RECT 30.530 1671.730 34.530 1755.350 ;
        RECT 270.920 1748.870 276.950 1754.940 ;
        RECT 316.750 1753.110 319.360 1758.660 ;
        RECT 30.530 1455.730 34.530 1539.350 ;
        RECT 270.920 1532.870 276.950 1538.940 ;
        RECT 316.750 1533.110 319.360 1538.660 ;
        RECT 316.510 1352.290 319.610 1388.960 ;
        RECT 316.510 1349.190 335.860 1352.290 ;
        RECT 30.530 1239.730 34.530 1323.350 ;
        RECT 270.920 1316.870 276.950 1322.940 ;
        RECT 332.760 1231.740 335.860 1349.190 ;
        RECT 1346.820 1232.340 1349.060 1246.620 ;
        RECT 1421.770 1232.340 1424.010 1246.620 ;
        RECT 1496.770 1232.340 1499.010 1246.620 ;
        RECT 1573.070 1232.340 1575.310 1246.620 ;
        RECT 3253.090 1231.480 3256.190 1388.990 ;
        RECT 3334.450 1232.330 3383.350 1247.380 ;
        RECT 30.530 1023.730 34.530 1107.350 ;
        RECT 270.920 1100.870 276.950 1106.940 ;
      LAYER via4 ;
        RECT 497.200 5154.110 498.690 5157.980 ;
        RECT 514.180 5154.130 515.580 5158.000 ;
        RECT 531.020 5154.140 532.440 5157.970 ;
        RECT 754.200 5154.110 755.690 5157.980 ;
        RECT 771.180 5154.130 772.580 5158.000 ;
        RECT 788.020 5154.140 789.440 5157.970 ;
        RECT 1011.200 5154.110 1012.690 5157.980 ;
        RECT 1028.180 5154.130 1029.580 5158.000 ;
        RECT 1045.020 5154.140 1046.440 5157.970 ;
        RECT 1268.200 5154.110 1269.690 5157.980 ;
        RECT 1285.180 5154.130 1286.580 5158.000 ;
        RECT 1302.020 5154.140 1303.440 5157.970 ;
        RECT 1526.200 5154.110 1527.690 5157.980 ;
        RECT 1543.180 5154.130 1544.580 5158.000 ;
        RECT 1560.020 5154.140 1561.440 5157.970 ;
        RECT 1778.200 5154.110 1779.690 5157.980 ;
        RECT 1795.180 5154.130 1796.580 5158.000 ;
        RECT 1812.020 5154.140 1813.440 5157.970 ;
        RECT 2115.200 5154.110 2116.690 5157.980 ;
        RECT 2132.180 5154.130 2133.580 5158.000 ;
        RECT 2149.020 5154.140 2150.440 5157.970 ;
        RECT 2500.200 5154.110 2501.690 5157.980 ;
        RECT 2517.180 5154.130 2518.580 5158.000 ;
        RECT 2534.020 5154.140 2535.440 5157.970 ;
        RECT 2757.200 5154.110 2758.690 5157.980 ;
        RECT 2774.180 5154.130 2775.580 5158.000 ;
        RECT 2791.020 5154.140 2792.440 5157.970 ;
        RECT 574.240 4969.950 579.730 4975.360 ;
        RECT 831.240 4969.950 836.730 4975.360 ;
        RECT 1088.240 4969.950 1093.730 4975.360 ;
        RECT 1345.240 4969.950 1350.730 4975.360 ;
        RECT 1603.240 4969.950 1608.730 4975.360 ;
        RECT 1855.240 4969.950 1860.730 4975.360 ;
        RECT 2192.240 4969.950 2197.730 4975.360 ;
        RECT 2577.240 4969.950 2582.730 4975.360 ;
        RECT 2834.240 4969.950 2839.730 4975.360 ;
        RECT 271.230 4744.240 276.640 4749.730 ;
        RECT 30.580 4701.030 34.440 4702.420 ;
        RECT 30.600 4684.200 34.480 4685.590 ;
        RECT 30.610 4667.200 34.480 4668.690 ;
        RECT 271.230 4115.240 276.640 4120.730 ;
        RECT 30.580 4072.030 34.440 4073.420 ;
        RECT 30.600 4055.200 34.480 4056.590 ;
        RECT 30.610 4038.200 34.480 4039.690 ;
        RECT 271.230 3899.240 276.640 3904.730 ;
        RECT 30.580 3856.030 34.440 3857.420 ;
        RECT 30.600 3839.200 34.480 3840.590 ;
        RECT 30.610 3822.200 34.480 3823.690 ;
        RECT 271.230 3683.240 276.640 3688.730 ;
        RECT 30.580 3640.030 34.440 3641.420 ;
        RECT 30.600 3623.200 34.480 3624.590 ;
        RECT 30.610 3606.200 34.480 3607.690 ;
        RECT 271.230 3467.240 276.640 3472.730 ;
        RECT 30.580 3424.030 34.440 3425.420 ;
        RECT 30.600 3407.200 34.480 3408.590 ;
        RECT 30.610 3390.200 34.480 3391.690 ;
        RECT 271.230 3251.240 276.640 3256.730 ;
        RECT 30.580 3208.030 34.440 3209.420 ;
        RECT 30.600 3191.200 34.480 3192.590 ;
        RECT 30.610 3174.200 34.480 3175.690 ;
        RECT 271.230 3035.240 276.640 3040.730 ;
        RECT 30.580 2992.030 34.440 2993.420 ;
        RECT 30.600 2975.200 34.480 2976.590 ;
        RECT 30.610 2958.200 34.480 2959.690 ;
        RECT 271.230 2819.240 276.640 2824.730 ;
        RECT 30.580 2776.030 34.440 2777.420 ;
        RECT 30.600 2759.200 34.480 2760.590 ;
        RECT 30.610 2742.200 34.480 2743.690 ;
        RECT 271.230 2181.240 276.640 2186.730 ;
        RECT 30.580 2138.030 34.440 2139.420 ;
        RECT 30.600 2121.200 34.480 2122.590 ;
        RECT 30.610 2104.200 34.480 2105.690 ;
        RECT 271.230 1965.240 276.640 1970.730 ;
        RECT 30.580 1922.030 34.440 1923.420 ;
        RECT 30.600 1905.200 34.480 1906.590 ;
        RECT 30.610 1888.200 34.480 1889.690 ;
        RECT 271.230 1749.240 276.640 1754.730 ;
        RECT 30.580 1706.030 34.440 1707.420 ;
        RECT 30.600 1689.200 34.480 1690.590 ;
        RECT 30.610 1672.200 34.480 1673.690 ;
        RECT 271.230 1533.240 276.640 1538.730 ;
        RECT 30.580 1490.030 34.440 1491.420 ;
        RECT 30.600 1473.200 34.480 1474.590 ;
        RECT 30.610 1456.200 34.480 1457.690 ;
        RECT 271.230 1317.240 276.640 1322.730 ;
        RECT 30.580 1274.030 34.440 1275.420 ;
        RECT 30.600 1257.200 34.480 1258.590 ;
        RECT 30.610 1240.200 34.480 1241.690 ;
        RECT 333.695 1245.670 334.875 1246.850 ;
        RECT 333.695 1244.070 334.875 1245.250 ;
        RECT 333.695 1242.470 334.875 1243.650 ;
        RECT 333.695 1240.870 334.875 1242.050 ;
        RECT 333.695 1239.270 334.875 1240.450 ;
        RECT 333.695 1237.670 334.875 1238.850 ;
        RECT 333.695 1236.070 334.875 1237.250 ;
        RECT 333.695 1234.470 334.875 1235.650 ;
        RECT 333.695 1232.870 334.875 1234.050 ;
        RECT 1347.350 1244.705 1348.530 1245.885 ;
        RECT 1347.350 1243.105 1348.530 1244.285 ;
        RECT 1347.350 1241.505 1348.530 1242.685 ;
        RECT 1347.350 1239.905 1348.530 1241.085 ;
        RECT 1347.350 1238.305 1348.530 1239.485 ;
        RECT 1347.350 1236.705 1348.530 1237.885 ;
        RECT 1347.350 1235.105 1348.530 1236.285 ;
        RECT 1347.350 1233.505 1348.530 1234.685 ;
        RECT 1422.300 1244.705 1423.480 1245.885 ;
        RECT 1422.300 1243.105 1423.480 1244.285 ;
        RECT 1422.300 1241.505 1423.480 1242.685 ;
        RECT 1422.300 1239.905 1423.480 1241.085 ;
        RECT 1422.300 1238.305 1423.480 1239.485 ;
        RECT 1422.300 1236.705 1423.480 1237.885 ;
        RECT 1422.300 1235.105 1423.480 1236.285 ;
        RECT 1422.300 1233.505 1423.480 1234.685 ;
        RECT 1497.300 1244.705 1498.480 1245.885 ;
        RECT 1497.300 1243.105 1498.480 1244.285 ;
        RECT 1497.300 1241.505 1498.480 1242.685 ;
        RECT 1497.300 1239.905 1498.480 1241.085 ;
        RECT 1497.300 1238.305 1498.480 1239.485 ;
        RECT 1497.300 1236.705 1498.480 1237.885 ;
        RECT 1497.300 1235.105 1498.480 1236.285 ;
        RECT 1497.300 1233.505 1498.480 1234.685 ;
        RECT 1573.600 1244.705 1574.780 1245.885 ;
        RECT 1573.600 1243.105 1574.780 1244.285 ;
        RECT 1573.600 1241.505 1574.780 1242.685 ;
        RECT 1573.600 1239.905 1574.780 1241.085 ;
        RECT 1573.600 1238.305 1574.780 1239.485 ;
        RECT 1573.600 1236.705 1574.780 1237.885 ;
        RECT 1573.600 1235.105 1574.780 1236.285 ;
        RECT 1573.600 1233.505 1574.780 1234.685 ;
        RECT 3253.240 1232.895 3256.020 1246.875 ;
        RECT 3335.560 1233.685 3347.940 1246.065 ;
        RECT 3371.130 1233.590 3381.910 1245.970 ;
        RECT 271.230 1101.240 276.640 1106.730 ;
        RECT 30.580 1058.030 34.440 1059.420 ;
        RECT 30.600 1041.200 34.480 1042.590 ;
        RECT 30.610 1024.200 34.480 1025.690 ;
      LAYER met5 ;
        RECT 497.060 5153.970 498.810 5158.130 ;
        RECT 514.010 5154.010 515.740 5158.390 ;
        RECT 497.140 5145.520 498.740 5153.970 ;
        RECT 514.040 5145.680 515.640 5154.010 ;
        RECT 530.830 5153.990 532.560 5158.370 ;
        RECT 530.940 5145.680 532.540 5153.990 ;
        RECT 754.060 5153.970 755.810 5158.130 ;
        RECT 771.010 5154.010 772.740 5158.390 ;
        RECT 754.140 5145.520 755.740 5153.970 ;
        RECT 771.040 5145.680 772.640 5154.010 ;
        RECT 787.830 5153.990 789.560 5158.370 ;
        RECT 787.940 5145.680 789.540 5153.990 ;
        RECT 1011.060 5153.970 1012.810 5158.130 ;
        RECT 1028.010 5154.010 1029.740 5158.390 ;
        RECT 1011.140 5145.520 1012.740 5153.970 ;
        RECT 1028.040 5145.680 1029.640 5154.010 ;
        RECT 1044.830 5153.990 1046.560 5158.370 ;
        RECT 1044.940 5145.680 1046.540 5153.990 ;
        RECT 1268.060 5153.970 1269.810 5158.130 ;
        RECT 1285.010 5154.010 1286.740 5158.390 ;
        RECT 1268.140 5145.520 1269.740 5153.970 ;
        RECT 1285.040 5145.680 1286.640 5154.010 ;
        RECT 1301.830 5153.990 1303.560 5158.370 ;
        RECT 1301.940 5145.680 1303.540 5153.990 ;
        RECT 1526.060 5153.970 1527.810 5158.130 ;
        RECT 1543.010 5154.010 1544.740 5158.390 ;
        RECT 1526.140 5145.520 1527.740 5153.970 ;
        RECT 1543.040 5145.680 1544.640 5154.010 ;
        RECT 1559.830 5153.990 1561.560 5158.370 ;
        RECT 1559.940 5145.680 1561.540 5153.990 ;
        RECT 1778.060 5153.970 1779.810 5158.130 ;
        RECT 1795.010 5154.010 1796.740 5158.390 ;
        RECT 1778.140 5145.520 1779.740 5153.970 ;
        RECT 1795.040 5145.680 1796.640 5154.010 ;
        RECT 1811.830 5153.990 1813.560 5158.370 ;
        RECT 1811.940 5145.680 1813.540 5153.990 ;
        RECT 2115.060 5153.970 2116.810 5158.130 ;
        RECT 2132.010 5154.010 2133.740 5158.390 ;
        RECT 2115.140 5145.520 2116.740 5153.970 ;
        RECT 2132.040 5145.680 2133.640 5154.010 ;
        RECT 2148.830 5153.990 2150.560 5158.370 ;
        RECT 2148.940 5145.680 2150.540 5153.990 ;
        RECT 2500.060 5153.970 2501.810 5158.130 ;
        RECT 2517.010 5154.010 2518.740 5158.390 ;
        RECT 2500.140 5145.520 2501.740 5153.970 ;
        RECT 2517.040 5145.680 2518.640 5154.010 ;
        RECT 2533.830 5153.990 2535.560 5158.370 ;
        RECT 2533.940 5145.680 2535.540 5153.990 ;
        RECT 2757.060 5153.970 2758.810 5158.130 ;
        RECT 2774.010 5154.010 2775.740 5158.390 ;
        RECT 2757.140 5145.520 2758.740 5153.970 ;
        RECT 2774.040 5145.680 2775.640 5154.010 ;
        RECT 2790.830 5153.990 2792.560 5158.370 ;
        RECT 2790.940 5145.680 2792.540 5153.990 ;
        RECT 270.990 4969.510 3383.100 4975.510 ;
        RECT 270.990 4917.940 276.990 4969.510 ;
        RECT 3370.100 4963.480 3383.100 4969.510 ;
        RECT 270.990 4914.840 316.580 4917.940 ;
        RECT 30.440 4702.540 34.635 4702.700 ;
        RECT 30.240 4700.940 42.910 4702.540 ;
        RECT 30.440 4700.895 34.635 4700.940 ;
        RECT 30.170 4685.640 34.645 4685.770 ;
        RECT 30.170 4684.040 42.910 4685.640 ;
        RECT 30.170 4684.030 34.645 4684.040 ;
        RECT 30.425 4668.740 34.900 4668.850 ;
        RECT 30.425 4667.140 43.070 4668.740 ;
        RECT 30.425 4667.040 34.900 4667.140 ;
        RECT 30.440 4073.540 34.635 4073.700 ;
        RECT 30.240 4071.940 42.910 4073.540 ;
        RECT 30.440 4071.895 34.635 4071.940 ;
        RECT 30.170 4056.640 34.645 4056.770 ;
        RECT 30.170 4055.040 42.910 4056.640 ;
        RECT 30.170 4055.030 34.645 4055.040 ;
        RECT 30.425 4039.740 34.900 4039.850 ;
        RECT 30.425 4038.140 43.070 4039.740 ;
        RECT 30.425 4038.040 34.900 4038.140 ;
        RECT 30.440 3857.540 34.635 3857.700 ;
        RECT 30.240 3855.940 42.910 3857.540 ;
        RECT 30.440 3855.895 34.635 3855.940 ;
        RECT 30.170 3840.640 34.645 3840.770 ;
        RECT 30.170 3839.040 42.910 3840.640 ;
        RECT 30.170 3839.030 34.645 3839.040 ;
        RECT 30.425 3823.740 34.900 3823.850 ;
        RECT 30.425 3822.140 43.070 3823.740 ;
        RECT 30.425 3822.040 34.900 3822.140 ;
        RECT 30.440 3641.540 34.635 3641.700 ;
        RECT 30.240 3639.940 42.910 3641.540 ;
        RECT 30.440 3639.895 34.635 3639.940 ;
        RECT 30.170 3624.640 34.645 3624.770 ;
        RECT 30.170 3623.040 42.910 3624.640 ;
        RECT 30.170 3623.030 34.645 3623.040 ;
        RECT 30.425 3607.740 34.900 3607.850 ;
        RECT 30.425 3606.140 43.070 3607.740 ;
        RECT 30.425 3606.040 34.900 3606.140 ;
        RECT 30.440 3425.540 34.635 3425.700 ;
        RECT 30.240 3423.940 42.910 3425.540 ;
        RECT 30.440 3423.895 34.635 3423.940 ;
        RECT 30.170 3408.640 34.645 3408.770 ;
        RECT 30.170 3407.040 42.910 3408.640 ;
        RECT 30.170 3407.030 34.645 3407.040 ;
        RECT 30.425 3391.740 34.900 3391.850 ;
        RECT 30.425 3390.140 43.070 3391.740 ;
        RECT 30.425 3390.040 34.900 3390.140 ;
        RECT 30.440 3209.540 34.635 3209.700 ;
        RECT 30.240 3207.940 42.910 3209.540 ;
        RECT 30.440 3207.895 34.635 3207.940 ;
        RECT 30.170 3192.640 34.645 3192.770 ;
        RECT 30.170 3191.040 42.910 3192.640 ;
        RECT 30.170 3191.030 34.645 3191.040 ;
        RECT 30.425 3175.740 34.900 3175.850 ;
        RECT 30.425 3174.140 43.070 3175.740 ;
        RECT 30.425 3174.040 34.900 3174.140 ;
        RECT 30.440 2993.540 34.635 2993.700 ;
        RECT 30.240 2991.940 42.910 2993.540 ;
        RECT 30.440 2991.895 34.635 2991.940 ;
        RECT 30.170 2976.640 34.645 2976.770 ;
        RECT 30.170 2975.040 42.910 2976.640 ;
        RECT 30.170 2975.030 34.645 2975.040 ;
        RECT 30.425 2959.740 34.900 2959.850 ;
        RECT 30.425 2958.140 43.070 2959.740 ;
        RECT 30.425 2958.040 34.900 2958.140 ;
        RECT 30.440 2777.540 34.635 2777.700 ;
        RECT 30.240 2775.940 42.910 2777.540 ;
        RECT 30.440 2775.895 34.635 2775.940 ;
        RECT 30.170 2760.640 34.645 2760.770 ;
        RECT 30.170 2759.040 42.910 2760.640 ;
        RECT 30.170 2759.030 34.645 2759.040 ;
        RECT 30.425 2743.740 34.900 2743.850 ;
        RECT 30.425 2742.140 43.070 2743.740 ;
        RECT 30.425 2742.040 34.900 2742.140 ;
        RECT 30.440 2139.540 34.635 2139.700 ;
        RECT 30.240 2137.940 42.910 2139.540 ;
        RECT 30.440 2137.895 34.635 2137.940 ;
        RECT 30.170 2122.640 34.645 2122.770 ;
        RECT 30.170 2121.040 42.910 2122.640 ;
        RECT 30.170 2121.030 34.645 2121.040 ;
        RECT 30.425 2105.740 34.900 2105.850 ;
        RECT 30.425 2104.140 43.070 2105.740 ;
        RECT 30.425 2104.040 34.900 2104.140 ;
        RECT 30.440 1923.540 34.635 1923.700 ;
        RECT 30.240 1921.940 42.910 1923.540 ;
        RECT 30.440 1921.895 34.635 1921.940 ;
        RECT 30.170 1906.640 34.645 1906.770 ;
        RECT 30.170 1905.040 42.910 1906.640 ;
        RECT 30.170 1905.030 34.645 1905.040 ;
        RECT 30.425 1889.740 34.900 1889.850 ;
        RECT 30.425 1888.140 43.070 1889.740 ;
        RECT 30.425 1888.040 34.900 1888.140 ;
        RECT 30.440 1707.540 34.635 1707.700 ;
        RECT 30.240 1705.940 42.910 1707.540 ;
        RECT 30.440 1705.895 34.635 1705.940 ;
        RECT 30.170 1690.640 34.645 1690.770 ;
        RECT 30.170 1689.040 42.910 1690.640 ;
        RECT 30.170 1689.030 34.645 1689.040 ;
        RECT 30.425 1673.740 34.900 1673.850 ;
        RECT 30.425 1672.140 43.070 1673.740 ;
        RECT 30.425 1672.040 34.900 1672.140 ;
        RECT 30.440 1491.540 34.635 1491.700 ;
        RECT 30.240 1489.940 42.910 1491.540 ;
        RECT 30.440 1489.895 34.635 1489.940 ;
        RECT 30.170 1474.640 34.645 1474.770 ;
        RECT 30.170 1473.040 42.910 1474.640 ;
        RECT 30.170 1473.030 34.645 1473.040 ;
        RECT 30.425 1457.740 34.900 1457.850 ;
        RECT 30.425 1456.140 43.070 1457.740 ;
        RECT 30.425 1456.040 34.900 1456.140 ;
        RECT 270.990 1392.020 276.990 4914.840 ;
        RECT 270.990 1388.920 316.560 1392.020 ;
        RECT 30.440 1275.540 34.635 1275.700 ;
        RECT 30.240 1273.940 42.910 1275.540 ;
        RECT 30.440 1273.895 34.635 1273.940 ;
        RECT 30.170 1258.640 34.645 1258.770 ;
        RECT 30.170 1257.040 42.910 1258.640 ;
        RECT 30.170 1257.030 34.645 1257.040 ;
        RECT 270.990 1247.330 276.990 1388.920 ;
        RECT 30.425 1241.740 34.900 1241.850 ;
        RECT 30.425 1240.140 43.070 1241.740 ;
        RECT 30.425 1240.040 34.900 1240.140 ;
        RECT 270.990 1232.330 3349.450 1247.330 ;
        RECT 3370.780 1233.080 3382.260 1246.480 ;
        RECT 270.990 1096.710 276.990 1232.330 ;
        RECT 30.440 1059.540 34.635 1059.700 ;
        RECT 30.240 1057.940 42.910 1059.540 ;
        RECT 30.440 1057.895 34.635 1057.940 ;
        RECT 30.170 1042.640 34.645 1042.770 ;
        RECT 30.170 1041.040 42.910 1042.640 ;
        RECT 30.170 1041.030 34.645 1041.040 ;
        RECT 30.425 1025.740 34.900 1025.850 ;
        RECT 30.425 1024.140 43.070 1025.740 ;
        RECT 30.425 1024.040 34.900 1024.140 ;
    END
  END vccd1_core
  PIN vssa1_core
    PORT
      LAYER met3 ;
        RECT 2878.500 4975.160 2902.395 4988.390 ;
        RECT 2928.390 4975.160 2952.290 4988.390 ;
        RECT 3319.570 2128.740 3388.560 2152.505 ;
        RECT 3319.570 2127.810 3335.550 2128.740 ;
        RECT 3319.570 2078.710 3388.560 2102.610 ;
      LAYER via3 ;
        RECT 2879.070 4975.715 2901.790 4985.235 ;
        RECT 2928.920 4975.745 2951.640 4985.265 ;
        RECT 3320.725 2128.425 3332.645 2151.945 ;
        RECT 3320.640 2079.435 3332.560 2102.155 ;
      LAYER met4 ;
        RECT 2878.400 4953.940 2902.390 4985.650 ;
        RECT 2928.350 4954.010 2952.340 4985.720 ;
        RECT 3320.040 2127.860 3333.060 2152.450 ;
        RECT 3320.090 2078.800 3333.170 2102.620 ;
        RECT 292.510 1332.040 295.610 1364.960 ;
        RECT 1953.860 1332.370 1957.790 1347.350 ;
        RECT 2029.110 1332.370 2033.040 1347.350 ;
        RECT 1956.870 1311.040 1957.770 1332.370 ;
        RECT 2032.120 1311.040 2033.020 1332.370 ;
        RECT 3277.090 1331.930 3280.190 1365.020 ;
      LAYER via4 ;
        RECT 2879.375 4955.105 2901.355 4965.885 ;
        RECT 2929.355 4955.175 2951.335 4965.955 ;
        RECT 3321.295 2129.195 3332.075 2151.175 ;
        RECT 3321.210 2079.805 3331.990 2101.785 ;
        RECT 293.445 1345.640 294.625 1346.820 ;
        RECT 293.445 1344.040 294.625 1345.220 ;
        RECT 293.445 1342.440 294.625 1343.620 ;
        RECT 293.445 1340.840 294.625 1342.020 ;
        RECT 293.445 1339.240 294.625 1340.420 ;
        RECT 293.445 1337.640 294.625 1338.820 ;
        RECT 293.445 1336.040 294.625 1337.220 ;
        RECT 293.445 1334.440 294.625 1335.620 ;
        RECT 293.445 1332.840 294.625 1334.020 ;
        RECT 1954.455 1332.825 1957.235 1346.805 ;
        RECT 2029.705 1332.825 2032.485 1346.805 ;
        RECT 3278.035 1345.625 3279.215 1346.805 ;
        RECT 3278.035 1344.025 3279.215 1345.205 ;
        RECT 3278.035 1342.425 3279.215 1343.605 ;
        RECT 3278.035 1340.825 3279.215 1342.005 ;
        RECT 3278.035 1339.225 3279.215 1340.405 ;
        RECT 3278.035 1337.625 3279.215 1338.805 ;
        RECT 3278.035 1336.025 3279.215 1337.205 ;
        RECT 3278.035 1334.425 3279.215 1335.605 ;
        RECT 3278.035 1332.825 3279.215 1334.005 ;
      LAYER met5 ;
        RECT 2878.200 4953.980 3333.100 4966.980 ;
        RECT 3320.100 4941.940 3333.100 4953.980 ;
        RECT 3280.190 4938.840 3333.100 4941.940 ;
        RECT 3320.100 1368.020 3333.100 4938.840 ;
        RECT 3280.130 1364.920 3333.100 1368.020 ;
        RECT 3320.100 1347.330 3333.100 1364.920 ;
        RECT 291.940 1332.330 3333.100 1347.330 ;
    END
  END vssa1_core
  PIN vdda1_core
    PORT
      LAYER met3 ;
        RECT 3335.860 4142.605 3389.090 4166.505 ;
        RECT 3335.860 4092.710 3389.090 4116.610 ;
        RECT 3335.310 2569.605 3388.500 2593.505 ;
        RECT 3335.310 2519.710 3388.500 2543.610 ;
      LAYER via3 ;
        RECT 3336.580 4143.230 3348.500 4165.950 ;
        RECT 3336.510 4093.260 3348.430 4115.980 ;
        RECT 3336.845 2570.435 3348.365 2592.755 ;
        RECT 3336.915 2520.485 3348.435 2542.805 ;
      LAYER met4 ;
        RECT 3291.900 4934.060 3349.130 4937.180 ;
        RECT 3336.010 4142.600 3349.010 4166.550 ;
        RECT 3336.070 4092.730 3349.070 4116.680 ;
        RECT 3336.030 2569.600 3349.070 2593.480 ;
        RECT 3336.090 2519.750 3349.130 2543.630 ;
        RECT 297.310 1333.090 300.410 1369.760 ;
        RECT 297.310 1329.990 316.660 1333.090 ;
        RECT 313.560 1312.010 316.660 1329.990 ;
        RECT 1919.970 1327.310 1920.870 1327.380 ;
        RECT 1995.220 1327.310 1996.120 1327.380 ;
        RECT 1916.830 1314.270 1920.870 1327.310 ;
        RECT 1992.080 1314.270 1996.120 1327.310 ;
        RECT 1919.970 1311.220 1920.870 1314.270 ;
        RECT 1995.220 1311.220 1996.120 1314.270 ;
        RECT 3272.290 1311.810 3275.390 1369.780 ;
        RECT 3294.750 1369.690 3349.060 1372.870 ;
        RECT 3336.080 1365.690 3349.060 1369.690 ;
      LAYER via4 ;
        RECT 3292.885 4935.030 3294.065 4936.210 ;
        RECT 3294.485 4935.030 3295.665 4936.210 ;
        RECT 3296.085 4935.030 3297.265 4936.210 ;
        RECT 3297.685 4935.030 3298.865 4936.210 ;
        RECT 3299.285 4935.030 3300.465 4936.210 ;
        RECT 3300.885 4935.030 3302.065 4936.210 ;
        RECT 3302.485 4935.030 3303.665 4936.210 ;
        RECT 3304.085 4935.030 3305.265 4936.210 ;
        RECT 3305.685 4935.030 3306.865 4936.210 ;
        RECT 3307.285 4935.030 3308.465 4936.210 ;
        RECT 3308.885 4935.030 3310.065 4936.210 ;
        RECT 3310.485 4935.030 3311.665 4936.210 ;
        RECT 3312.085 4935.030 3313.265 4936.210 ;
        RECT 3313.685 4935.030 3314.865 4936.210 ;
        RECT 3336.405 4935.055 3337.585 4936.235 ;
        RECT 3338.005 4935.055 3339.185 4936.235 ;
        RECT 3339.605 4935.055 3340.785 4936.235 ;
        RECT 3341.205 4935.055 3342.385 4936.235 ;
        RECT 3342.805 4935.055 3343.985 4936.235 ;
        RECT 3344.405 4935.055 3345.585 4936.235 ;
        RECT 3346.005 4935.055 3347.185 4936.235 ;
        RECT 3347.605 4935.055 3348.785 4936.235 ;
        RECT 3337.150 4143.600 3347.930 4165.580 ;
        RECT 3337.080 4093.630 3347.860 4115.610 ;
        RECT 3337.215 2570.605 3347.995 2592.585 ;
        RECT 3337.285 2520.655 3348.065 2542.635 ;
        RECT 3295.925 1370.645 3297.105 1371.825 ;
        RECT 3297.525 1370.645 3298.705 1371.825 ;
        RECT 3299.125 1370.645 3300.305 1371.825 ;
        RECT 3300.725 1370.645 3301.905 1371.825 ;
        RECT 3302.325 1370.645 3303.505 1371.825 ;
        RECT 3303.925 1370.645 3305.105 1371.825 ;
        RECT 3305.525 1370.645 3306.705 1371.825 ;
        RECT 3307.125 1370.645 3308.305 1371.825 ;
        RECT 3308.725 1370.645 3309.905 1371.825 ;
        RECT 3310.325 1370.645 3311.505 1371.825 ;
        RECT 3311.925 1370.645 3313.105 1371.825 ;
        RECT 3313.525 1370.645 3314.705 1371.825 ;
        RECT 314.485 1325.620 315.665 1326.800 ;
        RECT 314.485 1324.020 315.665 1325.200 ;
        RECT 314.485 1322.420 315.665 1323.600 ;
        RECT 314.485 1320.820 315.665 1322.000 ;
        RECT 314.485 1319.220 315.665 1320.400 ;
        RECT 314.485 1317.620 315.665 1318.800 ;
        RECT 314.485 1316.020 315.665 1317.200 ;
        RECT 314.485 1314.420 315.665 1315.600 ;
        RECT 1917.435 1315.260 1920.215 1326.040 ;
        RECT 1992.685 1315.260 1995.465 1326.040 ;
        RECT 314.485 1312.820 315.665 1314.000 ;
        RECT 3337.240 1366.280 3348.020 1372.260 ;
        RECT 3273.245 1325.615 3274.425 1326.795 ;
        RECT 3273.245 1324.015 3274.425 1325.195 ;
        RECT 3273.245 1322.415 3274.425 1323.595 ;
        RECT 3273.245 1320.815 3274.425 1321.995 ;
        RECT 3273.245 1319.215 3274.425 1320.395 ;
        RECT 3273.245 1317.615 3274.425 1318.795 ;
        RECT 3273.245 1316.015 3274.425 1317.195 ;
        RECT 3273.245 1314.415 3274.425 1315.595 ;
        RECT 3273.245 1312.815 3274.425 1313.995 ;
      LAYER met5 ;
        RECT 3275.390 4934.040 3315.890 4937.140 ;
        RECT 3275.300 1369.720 3315.790 1372.820 ;
        RECT 3336.100 1327.330 3349.100 4937.830 ;
        RECT 312.670 1312.330 3349.100 1327.330 ;
    END
  END vdda1_core
  OBS
      LAYER met2 ;
        RECT 2208.095 203.885 2209.960 211.885 ;
        RECT 2208.015 202.820 2210.045 203.885 ;
      LAYER via2 ;
        RECT 2208.095 202.910 2209.960 203.810 ;
      LAYER met3 ;
        RECT 549.500 4996.630 555.500 5093.480 ;
        RECT 557.500 5029.580 563.500 5099.450 ;
        RECT 806.500 4996.630 812.500 5093.480 ;
        RECT 814.500 5029.580 820.500 5099.450 ;
        RECT 842.905 4986.595 844.770 5034.235 ;
        RECT 848.895 4985.700 850.745 5001.540 ;
        RECT 1063.500 4996.630 1069.500 5093.480 ;
        RECT 1071.500 5029.580 1077.500 5099.450 ;
        RECT 1320.500 4996.630 1326.500 5093.480 ;
        RECT 1328.500 5029.580 1334.500 5099.450 ;
        RECT 1578.500 4996.630 1584.500 5093.480 ;
        RECT 1586.500 5029.580 1592.500 5099.450 ;
        RECT 1830.500 4996.630 1836.500 5093.480 ;
        RECT 1838.500 5029.580 1844.500 5099.450 ;
        RECT 2085.090 4986.595 2086.955 5034.235 ;
        RECT 2091.080 4985.695 2092.930 5001.535 ;
        RECT 2167.500 4996.630 2173.500 5093.480 ;
        RECT 2175.500 5029.580 2181.500 5099.450 ;
        RECT 2552.500 4996.630 2558.500 5093.480 ;
        RECT 2560.500 5029.580 2566.500 5099.450 ;
        RECT 2809.500 4996.630 2815.500 5093.480 ;
        RECT 2817.500 5029.580 2823.500 5099.450 ;
        RECT 3318.140 4986.595 3320.005 5034.235 ;
        RECT 3324.130 4985.695 3325.980 5001.535 ;
        RECT 220.990 4759.620 309.980 4765.620 ;
        RECT 204.920 4751.620 305.160 4757.620 ;
        RECT 89.140 4727.500 158.310 4733.500 ;
        RECT 3253.080 4725.910 3559.020 4731.910 ;
        RECT 95.110 4719.500 191.260 4725.500 ;
        RECT 3257.900 4717.910 3552.950 4723.910 ;
        RECT 3429.570 4709.500 3499.990 4715.500 ;
        RECT 3396.620 4701.500 3494.020 4707.500 ;
        RECT 3253.080 4499.910 3379.150 4505.910 ;
        RECT 3257.900 4491.910 3363.380 4497.910 ;
        RECT 153.765 4446.875 202.365 4448.740 ;
        RECT 186.465 4440.905 202.345 4442.755 ;
        RECT 3253.080 4274.910 3376.320 4280.910 ;
        RECT 3257.900 4266.910 3363.540 4272.910 ;
        RECT 220.990 4130.620 309.980 4136.620 ;
        RECT 204.920 4122.620 305.160 4128.620 ;
        RECT 89.140 4098.500 158.310 4104.500 ;
        RECT 95.110 4090.500 191.260 4096.500 ;
        RECT 220.990 3922.620 309.980 3928.620 ;
        RECT 204.920 3914.620 305.160 3920.620 ;
        RECT 89.140 3882.500 158.310 3888.500 ;
        RECT 95.110 3874.500 191.260 3880.500 ;
        RECT 3253.080 3833.910 3559.070 3839.910 ;
        RECT 3257.900 3825.910 3553.000 3831.910 ;
        RECT 3429.620 3817.500 3500.040 3823.500 ;
        RECT 3396.670 3809.500 3494.070 3815.500 ;
        RECT 220.990 3698.620 309.980 3704.620 ;
        RECT 204.920 3690.620 305.160 3696.620 ;
        RECT 89.140 3666.500 158.310 3672.500 ;
        RECT 95.110 3658.500 191.260 3664.500 ;
        RECT 3386.595 3622.445 3434.235 3624.310 ;
        RECT 3385.695 3616.470 3401.535 3618.320 ;
        RECT 3253.080 3608.910 3559.070 3614.910 ;
        RECT 3257.900 3600.910 3553.000 3606.910 ;
        RECT 3429.620 3592.500 3500.040 3598.500 ;
        RECT 3396.670 3584.500 3494.070 3590.500 ;
        RECT 220.990 3482.620 309.980 3488.620 ;
        RECT 204.920 3474.620 305.160 3480.620 ;
        RECT 89.140 3450.500 158.310 3456.500 ;
        RECT 95.110 3442.500 191.260 3448.500 ;
        RECT 3253.080 3382.910 3559.070 3388.910 ;
        RECT 3257.900 3374.910 3553.000 3380.910 ;
        RECT 3429.620 3366.500 3500.040 3372.500 ;
        RECT 3396.670 3358.500 3494.070 3364.500 ;
        RECT 220.990 3266.620 309.980 3272.620 ;
        RECT 204.920 3258.620 305.160 3264.620 ;
        RECT 89.140 3234.500 158.310 3240.500 ;
        RECT 95.110 3226.500 191.260 3232.500 ;
        RECT 3253.080 3157.910 3559.070 3163.910 ;
        RECT 3296.550 3149.910 3553.000 3155.910 ;
        RECT 3257.900 3143.910 3303.000 3149.910 ;
        RECT 3429.620 3141.500 3500.040 3147.500 ;
        RECT 3396.670 3133.500 3494.070 3139.500 ;
        RECT 220.990 3055.920 309.980 3061.920 ;
        RECT 204.920 3047.920 305.160 3053.920 ;
        RECT 153.865 3024.500 202.150 3024.870 ;
        RECT 89.140 3023.005 202.150 3024.500 ;
        RECT 89.140 3018.500 158.310 3023.005 ;
        RECT 188.000 3017.035 201.990 3018.885 ;
        RECT 188.000 3016.500 191.260 3017.035 ;
        RECT 95.110 3010.500 191.260 3016.500 ;
        RECT 3253.080 2931.910 3559.070 2937.910 ;
        RECT 3257.900 2923.910 3553.000 2929.910 ;
        RECT 3429.620 2915.500 3500.040 2921.500 ;
        RECT 3396.670 2907.500 3494.070 2913.500 ;
        RECT 220.990 2834.620 309.980 2840.620 ;
        RECT 204.920 2826.620 305.160 2832.620 ;
        RECT 89.140 2802.500 158.310 2808.500 ;
        RECT 95.110 2794.500 191.260 2800.500 ;
        RECT 3253.080 2706.910 3559.070 2712.910 ;
        RECT 3257.900 2698.910 3553.000 2704.910 ;
        RECT 3429.620 2690.500 3500.040 2696.500 ;
        RECT 3396.670 2682.500 3494.070 2688.500 ;
        RECT 3253.080 2492.910 3298.790 2495.910 ;
        RECT 3253.080 2489.910 3559.070 2492.910 ;
        RECT 3292.840 2486.910 3559.070 2489.910 ;
        RECT 3257.900 2478.910 3553.000 2484.910 ;
        RECT 3429.620 2470.500 3500.040 2476.500 ;
        RECT 3396.670 2462.500 3494.070 2468.500 ;
        RECT 3386.595 2240.440 3434.235 2242.305 ;
        RECT 3385.695 2234.465 3401.535 2236.315 ;
        RECT 220.990 2196.620 309.980 2202.620 ;
        RECT 204.920 2188.620 305.160 2194.620 ;
        RECT 89.140 2164.500 158.310 2170.500 ;
        RECT 95.110 2156.500 191.260 2162.500 ;
        RECT 3253.080 2045.910 3559.070 2051.910 ;
        RECT 3257.900 2037.910 3553.000 2043.910 ;
        RECT 3429.620 2029.500 3500.040 2035.500 ;
        RECT 3396.670 2021.500 3494.070 2027.500 ;
        RECT 220.990 1980.620 309.980 1986.620 ;
        RECT 204.920 1972.620 305.160 1978.620 ;
        RECT 89.140 1948.500 158.310 1954.500 ;
        RECT 95.110 1940.500 191.260 1946.500 ;
        RECT 3253.080 1826.910 3328.320 1832.910 ;
        RECT 3322.320 1825.910 3328.320 1826.910 ;
        RECT 3322.320 1819.910 3559.070 1825.910 ;
        RECT 3257.900 1811.910 3553.000 1817.910 ;
        RECT 3429.620 1803.500 3500.040 1809.500 ;
        RECT 3396.670 1795.500 3494.070 1801.500 ;
        RECT 220.990 1769.620 309.980 1775.620 ;
        RECT 204.920 1761.620 305.160 1767.620 ;
        RECT 89.140 1736.615 158.310 1738.500 ;
        RECT 89.140 1734.750 202.545 1736.615 ;
        RECT 89.140 1732.500 158.310 1734.750 ;
        RECT 186.465 1730.500 203.595 1730.630 ;
        RECT 95.110 1728.780 203.595 1730.500 ;
        RECT 95.110 1724.500 191.260 1728.780 ;
        RECT 3253.080 1594.910 3559.070 1600.910 ;
        RECT 3257.900 1586.910 3553.000 1592.910 ;
        RECT 3429.620 1578.500 3500.040 1584.500 ;
        RECT 3396.670 1570.500 3494.070 1576.500 ;
        RECT 220.990 1548.620 309.980 1554.620 ;
        RECT 204.920 1540.620 305.160 1546.620 ;
        RECT 89.140 1516.500 158.310 1522.500 ;
        RECT 95.110 1508.500 191.260 1514.500 ;
        RECT 3376.380 1369.910 3559.070 1375.910 ;
        RECT 3358.100 1361.910 3553.000 1367.910 ;
        RECT 3429.620 1353.500 3500.040 1359.500 ;
        RECT 3396.670 1345.500 3494.070 1351.500 ;
        RECT 89.140 1300.500 158.310 1306.500 ;
        RECT 95.110 1292.500 191.260 1298.500 ;
        RECT 3376.380 1143.910 3559.070 1149.910 ;
        RECT 3358.100 1135.910 3553.000 1141.910 ;
        RECT 3429.620 1127.500 3500.040 1133.500 ;
        RECT 3396.670 1119.500 3494.070 1125.500 ;
        RECT 89.140 1084.500 158.310 1090.500 ;
        RECT 95.110 1076.500 191.260 1082.500 ;
        RECT 3376.380 918.910 3559.070 924.910 ;
        RECT 3358.100 910.910 3553.000 916.910 ;
        RECT 3429.620 902.500 3500.040 908.500 ;
        RECT 3396.670 894.500 3494.070 900.500 ;
        RECT 3376.380 692.910 3559.070 698.910 ;
        RECT 3358.100 684.910 3553.000 690.910 ;
        RECT 3429.620 676.500 3500.040 682.500 ;
        RECT 3396.670 668.500 3494.070 674.500 ;
        RECT 730.965 209.380 732.815 211.400 ;
        RECT 736.940 209.835 746.570 210.455 ;
        RECT 2202.265 209.980 2202.585 210.300 ;
        RECT 2202.665 209.980 2202.985 210.300 ;
        RECT 2203.065 209.980 2203.385 210.300 ;
        RECT 2203.465 209.980 2203.785 210.300 ;
        RECT 643.050 169.500 647.340 208.000 ;
        RECT 730.965 207.390 740.895 209.380 ;
        RECT 650.710 175.570 655.000 204.610 ;
        RECT 738.975 186.505 740.900 203.515 ;
        RECT 2130.090 154.030 2131.995 203.810 ;
        RECT 2135.095 186.700 2137.000 205.790 ;
        RECT 2208.015 202.820 2210.045 203.885 ;
        RECT 2281.685 186.700 2283.590 203.810 ;
        RECT 2286.695 154.030 2288.600 203.810 ;
        RECT 3209.770 169.600 3218.470 220.130 ;
        RECT 3267.310 179.040 3284.550 225.780 ;
      LAYER via3 ;
        RECT 557.680 5095.410 563.340 5099.160 ;
        RECT 549.690 5089.390 555.350 5093.140 ;
        RECT 814.680 5095.410 820.340 5099.160 ;
        RECT 557.770 5030.020 563.160 5033.790 ;
        RECT 806.690 5089.390 812.350 5093.140 ;
        RECT 549.900 4997.290 555.320 5001.100 ;
        RECT 1071.680 5095.410 1077.340 5099.160 ;
        RECT 1063.690 5089.390 1069.350 5093.140 ;
        RECT 814.770 5030.020 820.160 5033.790 ;
        RECT 843.255 5029.885 844.375 5033.405 ;
        RECT 806.900 4997.290 812.320 5001.100 ;
        RECT 849.235 4997.440 850.355 5000.960 ;
        RECT 1328.680 5095.410 1334.340 5099.160 ;
        RECT 1071.770 5030.020 1077.160 5033.790 ;
        RECT 1320.690 5089.390 1326.350 5093.140 ;
        RECT 1063.900 4997.290 1069.320 5001.100 ;
        RECT 1586.680 5095.410 1592.340 5099.160 ;
        RECT 1328.770 5030.020 1334.160 5033.790 ;
        RECT 1578.690 5089.390 1584.350 5093.140 ;
        RECT 1320.900 4997.290 1326.320 5001.100 ;
        RECT 1838.680 5095.410 1844.340 5099.160 ;
        RECT 1586.770 5030.020 1592.160 5033.790 ;
        RECT 1830.690 5089.390 1836.350 5093.140 ;
        RECT 1578.900 4997.290 1584.320 5001.100 ;
        RECT 2175.680 5095.410 2181.340 5099.160 ;
        RECT 2167.690 5089.390 2173.350 5093.140 ;
        RECT 1838.770 5030.020 1844.160 5033.790 ;
        RECT 2085.440 5029.885 2086.560 5033.405 ;
        RECT 1830.900 4997.290 1836.320 5001.100 ;
        RECT 2091.420 4997.435 2092.540 5000.955 ;
        RECT 2560.680 5095.410 2566.340 5099.160 ;
        RECT 2175.770 5030.020 2181.160 5033.790 ;
        RECT 2552.690 5089.390 2558.350 5093.140 ;
        RECT 2167.900 4997.290 2173.320 5001.100 ;
        RECT 2817.680 5095.410 2823.340 5099.160 ;
        RECT 2560.770 5030.020 2566.160 5033.790 ;
        RECT 2809.690 5089.390 2815.350 5093.140 ;
        RECT 2552.900 4997.290 2558.320 5001.100 ;
        RECT 2817.770 5030.020 2823.160 5033.790 ;
        RECT 3318.490 5029.885 3319.610 5033.405 ;
        RECT 2809.900 4997.290 2815.320 5001.100 ;
        RECT 3324.470 4997.435 3325.590 5000.955 ;
        RECT 221.570 4759.955 233.490 4765.075 ;
        RECT 307.305 4759.840 309.625 4765.360 ;
        RECT 205.520 4752.045 217.440 4757.165 ;
        RECT 302.485 4751.880 304.805 4757.400 ;
        RECT 89.430 4727.680 93.180 4733.340 ;
        RECT 154.100 4727.770 157.870 4733.160 ;
        RECT 3253.280 4726.165 3256.000 4731.685 ;
        RECT 3376.990 4726.240 3382.400 4731.730 ;
        RECT 3554.870 4726.120 3558.370 4731.690 ;
        RECT 95.450 4719.690 99.200 4725.350 ;
        RECT 186.790 4719.900 190.600 4725.320 ;
        RECT 3258.070 4718.145 3260.790 4723.665 ;
        RECT 3358.460 4718.150 3363.870 4723.640 ;
        RECT 3548.880 4718.140 3552.380 4723.710 ;
        RECT 3430.010 4709.770 3433.780 4715.160 ;
        RECT 3495.950 4709.680 3499.700 4715.340 ;
        RECT 3397.280 4701.900 3401.090 4707.320 ;
        RECT 3489.930 4701.690 3493.680 4707.350 ;
        RECT 3253.280 4500.165 3256.000 4505.685 ;
        RECT 3373.825 4500.405 3378.545 4505.525 ;
        RECT 3258.070 4492.145 3260.790 4497.665 ;
        RECT 3357.845 4492.365 3362.965 4497.485 ;
        RECT 154.235 4447.440 157.755 4448.560 ;
        RECT 186.935 4441.455 190.455 4442.575 ;
        RECT 3253.280 4275.165 3256.000 4280.685 ;
        RECT 3370.680 4275.360 3375.800 4280.480 ;
        RECT 3258.070 4267.145 3260.790 4272.665 ;
        RECT 3357.960 4267.350 3363.080 4272.470 ;
        RECT 221.570 4130.955 233.490 4136.075 ;
        RECT 307.305 4130.840 309.625 4136.360 ;
        RECT 205.520 4123.045 217.440 4128.165 ;
        RECT 302.485 4122.880 304.805 4128.400 ;
        RECT 89.430 4098.680 93.180 4104.340 ;
        RECT 154.100 4098.770 157.870 4104.160 ;
        RECT 95.450 4090.690 99.200 4096.350 ;
        RECT 186.790 4090.900 190.600 4096.320 ;
        RECT 221.570 3922.955 233.490 3928.075 ;
        RECT 307.305 3922.840 309.625 3928.360 ;
        RECT 205.520 3915.045 217.440 3920.165 ;
        RECT 302.485 3914.880 304.805 3920.400 ;
        RECT 89.430 3882.680 93.180 3888.340 ;
        RECT 154.100 3882.770 157.870 3888.160 ;
        RECT 95.450 3874.690 99.200 3880.350 ;
        RECT 186.790 3874.900 190.600 3880.320 ;
        RECT 3253.280 3834.165 3256.000 3839.685 ;
        RECT 3377.040 3834.240 3382.450 3839.730 ;
        RECT 3554.920 3834.120 3558.420 3839.690 ;
        RECT 3258.070 3826.145 3260.790 3831.665 ;
        RECT 3358.510 3826.150 3363.920 3831.640 ;
        RECT 3548.930 3826.140 3552.430 3831.710 ;
        RECT 3430.060 3817.770 3433.830 3823.160 ;
        RECT 3496.000 3817.680 3499.750 3823.340 ;
        RECT 3397.330 3809.900 3401.140 3815.320 ;
        RECT 3489.980 3809.690 3493.730 3815.350 ;
        RECT 221.570 3698.955 233.490 3704.075 ;
        RECT 307.305 3698.840 309.625 3704.360 ;
        RECT 205.520 3691.045 217.440 3696.165 ;
        RECT 302.485 3690.880 304.805 3696.400 ;
        RECT 89.430 3666.680 93.180 3672.340 ;
        RECT 154.100 3666.770 157.870 3672.160 ;
        RECT 95.450 3658.690 99.200 3664.350 ;
        RECT 186.790 3658.900 190.600 3664.320 ;
        RECT 3429.885 3622.840 3433.405 3623.960 ;
        RECT 3397.435 3616.860 3400.955 3617.980 ;
        RECT 3253.280 3609.165 3256.000 3614.685 ;
        RECT 3377.040 3609.240 3382.450 3614.730 ;
        RECT 3554.920 3609.120 3558.420 3614.690 ;
        RECT 3258.070 3601.145 3260.790 3606.665 ;
        RECT 3358.510 3601.150 3363.920 3606.640 ;
        RECT 3548.930 3601.140 3552.430 3606.710 ;
        RECT 3430.060 3592.770 3433.830 3598.160 ;
        RECT 3496.000 3592.680 3499.750 3598.340 ;
        RECT 3397.330 3584.900 3401.140 3590.320 ;
        RECT 3489.980 3584.690 3493.730 3590.350 ;
        RECT 221.570 3482.955 233.490 3488.075 ;
        RECT 307.305 3482.840 309.625 3488.360 ;
        RECT 205.520 3475.045 217.440 3480.165 ;
        RECT 302.485 3474.880 304.805 3480.400 ;
        RECT 89.430 3450.680 93.180 3456.340 ;
        RECT 154.100 3450.770 157.870 3456.160 ;
        RECT 95.450 3442.690 99.200 3448.350 ;
        RECT 186.790 3442.900 190.600 3448.320 ;
        RECT 3253.280 3383.165 3256.000 3388.685 ;
        RECT 3377.040 3383.240 3382.450 3388.730 ;
        RECT 3554.920 3383.120 3558.420 3388.690 ;
        RECT 3258.070 3375.145 3260.790 3380.665 ;
        RECT 3358.510 3375.150 3363.920 3380.640 ;
        RECT 3548.930 3375.140 3552.430 3380.710 ;
        RECT 3430.060 3366.770 3433.830 3372.160 ;
        RECT 3496.000 3366.680 3499.750 3372.340 ;
        RECT 3397.330 3358.900 3401.140 3364.320 ;
        RECT 3489.980 3358.690 3493.730 3364.350 ;
        RECT 221.570 3266.955 233.490 3272.075 ;
        RECT 307.305 3266.840 309.625 3272.360 ;
        RECT 205.520 3259.045 217.440 3264.165 ;
        RECT 302.485 3258.880 304.805 3264.400 ;
        RECT 89.430 3234.680 93.180 3240.340 ;
        RECT 154.100 3234.770 157.870 3240.160 ;
        RECT 95.450 3226.690 99.200 3232.350 ;
        RECT 186.790 3226.900 190.600 3232.320 ;
        RECT 3253.280 3158.165 3256.000 3163.685 ;
        RECT 3377.040 3158.240 3382.450 3163.730 ;
        RECT 3554.920 3158.120 3558.420 3163.690 ;
        RECT 3358.510 3150.150 3363.920 3155.640 ;
        RECT 3548.930 3150.140 3552.430 3155.710 ;
        RECT 3258.070 3144.145 3260.790 3149.665 ;
        RECT 3430.060 3141.770 3433.830 3147.160 ;
        RECT 3496.000 3141.680 3499.750 3147.340 ;
        RECT 3397.330 3133.900 3401.140 3139.320 ;
        RECT 3489.980 3133.690 3493.730 3139.350 ;
        RECT 221.570 3056.255 233.490 3061.375 ;
        RECT 307.305 3056.140 309.625 3061.660 ;
        RECT 205.520 3048.345 217.440 3053.465 ;
        RECT 302.485 3048.180 304.805 3053.700 ;
        RECT 89.430 3018.680 93.180 3024.340 ;
        RECT 154.100 3018.770 157.870 3024.160 ;
        RECT 95.450 3010.690 99.200 3016.350 ;
        RECT 186.790 3010.900 190.600 3016.320 ;
        RECT 3253.280 2932.165 3256.000 2937.685 ;
        RECT 3377.040 2932.240 3382.450 2937.730 ;
        RECT 3554.920 2932.120 3558.420 2937.690 ;
        RECT 3258.070 2924.145 3260.790 2929.665 ;
        RECT 3358.510 2924.150 3363.920 2929.640 ;
        RECT 3548.930 2924.140 3552.430 2929.710 ;
        RECT 3430.060 2915.770 3433.830 2921.160 ;
        RECT 3496.000 2915.680 3499.750 2921.340 ;
        RECT 3397.330 2907.900 3401.140 2913.320 ;
        RECT 3489.980 2907.690 3493.730 2913.350 ;
        RECT 221.570 2834.955 233.490 2840.075 ;
        RECT 307.305 2834.840 309.625 2840.360 ;
        RECT 205.520 2827.045 217.440 2832.165 ;
        RECT 302.485 2826.880 304.805 2832.400 ;
        RECT 89.430 2802.680 93.180 2808.340 ;
        RECT 154.100 2802.770 157.870 2808.160 ;
        RECT 95.450 2794.690 99.200 2800.350 ;
        RECT 186.790 2794.900 190.600 2800.320 ;
        RECT 3253.280 2707.165 3256.000 2712.685 ;
        RECT 3377.040 2707.240 3382.450 2712.730 ;
        RECT 3554.920 2707.120 3558.420 2712.690 ;
        RECT 3258.070 2699.145 3260.790 2704.665 ;
        RECT 3358.510 2699.150 3363.920 2704.640 ;
        RECT 3548.930 2699.140 3552.430 2704.710 ;
        RECT 3430.060 2690.770 3433.830 2696.160 ;
        RECT 3496.000 2690.680 3499.750 2696.340 ;
        RECT 3397.330 2682.900 3401.140 2688.320 ;
        RECT 3489.980 2682.690 3493.730 2688.350 ;
        RECT 3253.280 2490.165 3256.000 2495.685 ;
        RECT 3377.040 2487.240 3382.450 2492.730 ;
        RECT 3554.920 2487.120 3558.420 2492.690 ;
        RECT 3258.070 2479.145 3260.790 2484.665 ;
        RECT 3358.510 2479.150 3363.920 2484.640 ;
        RECT 3548.930 2479.140 3552.430 2484.710 ;
        RECT 3430.060 2470.770 3433.830 2476.160 ;
        RECT 3496.000 2470.680 3499.750 2476.340 ;
        RECT 3397.330 2462.900 3401.140 2468.320 ;
        RECT 3489.980 2462.690 3493.730 2468.350 ;
        RECT 3429.885 2240.835 3433.405 2241.955 ;
        RECT 3397.435 2234.855 3400.955 2235.975 ;
        RECT 221.570 2196.955 233.490 2202.075 ;
        RECT 307.305 2196.840 309.625 2202.360 ;
        RECT 205.520 2189.045 217.440 2194.165 ;
        RECT 302.485 2188.880 304.805 2194.400 ;
        RECT 89.430 2164.680 93.180 2170.340 ;
        RECT 154.100 2164.770 157.870 2170.160 ;
        RECT 95.450 2156.690 99.200 2162.350 ;
        RECT 186.790 2156.900 190.600 2162.320 ;
        RECT 3253.280 2046.165 3256.000 2051.685 ;
        RECT 3377.040 2046.240 3382.450 2051.730 ;
        RECT 3554.920 2046.120 3558.420 2051.690 ;
        RECT 3258.070 2038.145 3260.790 2043.665 ;
        RECT 3358.510 2038.150 3363.920 2043.640 ;
        RECT 3548.930 2038.140 3552.430 2043.710 ;
        RECT 3430.060 2029.770 3433.830 2035.160 ;
        RECT 3496.000 2029.680 3499.750 2035.340 ;
        RECT 3397.330 2021.900 3401.140 2027.320 ;
        RECT 3489.980 2021.690 3493.730 2027.350 ;
        RECT 221.570 1980.955 233.490 1986.075 ;
        RECT 307.305 1980.840 309.625 1986.360 ;
        RECT 205.520 1973.045 217.440 1978.165 ;
        RECT 302.485 1972.880 304.805 1978.400 ;
        RECT 89.430 1948.680 93.180 1954.340 ;
        RECT 154.100 1948.770 157.870 1954.160 ;
        RECT 95.450 1940.690 99.200 1946.350 ;
        RECT 186.790 1940.900 190.600 1946.320 ;
        RECT 3253.280 1827.165 3256.000 1832.685 ;
        RECT 3377.040 1820.240 3382.450 1825.730 ;
        RECT 3554.920 1820.120 3558.420 1825.690 ;
        RECT 3258.070 1812.145 3260.790 1817.665 ;
        RECT 3358.510 1812.150 3363.920 1817.640 ;
        RECT 3548.930 1812.140 3552.430 1817.710 ;
        RECT 3430.060 1803.770 3433.830 1809.160 ;
        RECT 3496.000 1803.680 3499.750 1809.340 ;
        RECT 3397.330 1795.900 3401.140 1801.320 ;
        RECT 3489.980 1795.690 3493.730 1801.350 ;
        RECT 221.570 1769.955 233.490 1775.075 ;
        RECT 307.305 1769.840 309.625 1775.360 ;
        RECT 205.520 1762.045 217.440 1767.165 ;
        RECT 302.485 1761.880 304.805 1767.400 ;
        RECT 89.430 1732.680 93.180 1738.340 ;
        RECT 154.100 1732.770 157.870 1738.160 ;
        RECT 95.450 1724.690 99.200 1730.350 ;
        RECT 186.790 1724.900 190.600 1730.320 ;
        RECT 3253.280 1595.165 3256.000 1600.685 ;
        RECT 3377.040 1595.240 3382.450 1600.730 ;
        RECT 3554.920 1595.120 3558.420 1600.690 ;
        RECT 3258.070 1587.145 3260.790 1592.665 ;
        RECT 3358.510 1587.150 3363.920 1592.640 ;
        RECT 3548.930 1587.140 3552.430 1592.710 ;
        RECT 3430.060 1578.770 3433.830 1584.160 ;
        RECT 3496.000 1578.680 3499.750 1584.340 ;
        RECT 3397.330 1570.900 3401.140 1576.320 ;
        RECT 3489.980 1570.690 3493.730 1576.350 ;
        RECT 221.570 1548.955 233.490 1554.075 ;
        RECT 307.305 1548.840 309.625 1554.360 ;
        RECT 205.520 1541.045 217.440 1546.165 ;
        RECT 302.485 1540.880 304.805 1546.400 ;
        RECT 89.430 1516.680 93.180 1522.340 ;
        RECT 154.100 1516.770 157.870 1522.160 ;
        RECT 95.450 1508.690 99.200 1514.350 ;
        RECT 186.790 1508.900 190.600 1514.320 ;
        RECT 3377.040 1370.240 3382.450 1375.730 ;
        RECT 3554.920 1370.120 3558.420 1375.690 ;
        RECT 3358.510 1362.150 3363.920 1367.640 ;
        RECT 3548.930 1362.140 3552.430 1367.710 ;
        RECT 3430.060 1353.770 3433.830 1359.160 ;
        RECT 3496.000 1353.680 3499.750 1359.340 ;
        RECT 3397.330 1345.900 3401.140 1351.320 ;
        RECT 3489.980 1345.690 3493.730 1351.350 ;
        RECT 89.430 1300.680 93.180 1306.340 ;
        RECT 154.100 1300.770 157.870 1306.160 ;
        RECT 95.450 1292.690 99.200 1298.350 ;
        RECT 186.790 1292.900 190.600 1298.320 ;
        RECT 3377.040 1144.240 3382.450 1149.730 ;
        RECT 3554.920 1144.120 3558.420 1149.690 ;
        RECT 3358.510 1136.150 3363.920 1141.640 ;
        RECT 3548.930 1136.140 3552.430 1141.710 ;
        RECT 3430.060 1127.770 3433.830 1133.160 ;
        RECT 3496.000 1127.680 3499.750 1133.340 ;
        RECT 3397.330 1119.900 3401.140 1125.320 ;
        RECT 3489.980 1119.690 3493.730 1125.350 ;
        RECT 89.430 1084.680 93.180 1090.340 ;
        RECT 154.100 1084.770 157.870 1090.160 ;
        RECT 95.450 1076.690 99.200 1082.350 ;
        RECT 186.790 1076.900 190.600 1082.320 ;
        RECT 3377.040 919.240 3382.450 924.730 ;
        RECT 3554.920 919.120 3558.420 924.690 ;
        RECT 3358.510 911.150 3363.920 916.640 ;
        RECT 3548.930 911.140 3552.430 916.710 ;
        RECT 3430.060 902.770 3433.830 908.160 ;
        RECT 3496.000 902.680 3499.750 908.340 ;
        RECT 3397.330 894.900 3401.140 900.320 ;
        RECT 3489.980 894.690 3493.730 900.350 ;
        RECT 3377.040 693.240 3382.450 698.730 ;
        RECT 3554.920 693.120 3558.420 698.690 ;
        RECT 3358.510 685.150 3363.920 690.640 ;
        RECT 3548.930 685.140 3552.430 690.710 ;
        RECT 3430.060 676.770 3433.830 682.160 ;
        RECT 3496.000 676.680 3499.750 682.340 ;
        RECT 3397.330 668.900 3401.140 674.320 ;
        RECT 3489.980 668.690 3493.730 674.350 ;
        RECT 3209.975 211.105 3218.295 219.825 ;
        RECT 745.760 210.055 746.080 210.375 ;
        RECT 746.160 210.055 746.480 210.375 ;
        RECT 643.235 206.790 647.155 207.910 ;
        RECT 739.075 207.520 740.805 209.280 ;
        RECT 2135.295 204.980 2136.815 205.700 ;
        RECT 650.895 203.000 654.815 204.120 ;
        RECT 739.060 200.390 740.800 203.425 ;
        RECT 739.085 186.710 740.800 190.915 ;
        RECT 2130.290 203.000 2131.810 203.720 ;
        RECT 650.910 175.945 654.830 179.865 ;
        RECT 643.260 169.905 647.180 173.825 ;
        RECT 2208.095 202.910 2209.960 203.810 ;
        RECT 2135.285 187.050 2136.805 190.570 ;
        RECT 2281.885 200.080 2283.405 203.600 ;
        RECT 2281.885 187.050 2283.405 190.570 ;
        RECT 2286.890 200.080 2288.410 203.600 ;
        RECT 2130.280 154.380 2131.800 157.900 ;
        RECT 3267.915 213.190 3283.835 225.110 ;
        RECT 3210.190 170.110 3218.110 173.630 ;
        RECT 2286.890 154.380 2288.410 157.900 ;
      LAYER met4 ;
        RECT 500.110 5095.240 563.550 5099.240 ;
        RECT 757.110 5095.240 820.550 5099.240 ;
        RECT 1014.110 5095.240 1077.550 5099.240 ;
        RECT 1271.110 5095.240 1334.550 5099.240 ;
        RECT 1529.110 5095.240 1592.550 5099.240 ;
        RECT 1781.110 5095.240 1844.550 5099.240 ;
        RECT 2118.110 5095.240 2181.550 5099.240 ;
        RECT 2503.110 5095.240 2566.550 5099.240 ;
        RECT 2760.110 5095.240 2823.550 5099.240 ;
        RECT 491.740 5089.240 556.660 5093.240 ;
        RECT 748.740 5089.240 813.660 5093.240 ;
        RECT 1005.740 5089.240 1070.660 5093.240 ;
        RECT 1262.740 5089.240 1327.660 5093.240 ;
        RECT 1520.740 5089.240 1585.660 5093.240 ;
        RECT 1772.740 5089.240 1837.660 5093.240 ;
        RECT 2109.740 5089.240 2174.660 5093.240 ;
        RECT 2494.740 5089.240 2559.660 5093.240 ;
        RECT 2751.740 5089.240 2816.660 5093.240 ;
        RECT 557.770 5030.020 563.160 5033.790 ;
        RECT 814.770 5030.020 820.160 5033.790 ;
        RECT 843.255 5029.885 844.375 5033.405 ;
        RECT 1071.770 5030.020 1077.160 5033.790 ;
        RECT 1328.770 5030.020 1334.160 5033.790 ;
        RECT 1586.770 5030.020 1592.160 5033.790 ;
        RECT 1838.770 5030.020 1844.160 5033.790 ;
        RECT 2085.440 5029.885 2086.560 5033.405 ;
        RECT 2175.770 5030.020 2181.160 5033.790 ;
        RECT 2560.770 5030.020 2566.160 5033.790 ;
        RECT 2817.770 5030.020 2823.160 5033.790 ;
        RECT 3318.490 5029.885 3319.610 5033.405 ;
        RECT 549.900 4997.290 555.320 5001.100 ;
        RECT 806.900 4997.290 812.320 5001.100 ;
        RECT 849.235 4997.440 850.355 5000.960 ;
        RECT 1063.900 4997.290 1069.320 5001.100 ;
        RECT 1320.900 4997.290 1326.320 5001.100 ;
        RECT 1578.900 4997.290 1584.320 5001.100 ;
        RECT 1830.900 4997.290 1836.320 5001.100 ;
        RECT 2091.420 4997.435 2092.540 5000.955 ;
        RECT 2167.900 4997.290 2173.320 5001.100 ;
        RECT 2552.900 4997.290 2558.320 5001.100 ;
        RECT 2809.900 4997.290 2815.320 5001.100 ;
        RECT 3324.470 4997.435 3325.590 5000.955 ;
        RECT 204.965 4929.270 282.070 4932.340 ;
        RECT 221.000 4924.370 282.200 4927.630 ;
        RECT 3291.580 4919.640 3367.150 4922.850 ;
        RECT 3291.440 4914.800 3383.120 4918.010 ;
        RECT 221.000 4759.610 233.960 4765.630 ;
        RECT 307.120 4759.800 309.810 4765.400 ;
        RECT 204.970 4751.630 217.940 4757.610 ;
        RECT 302.300 4751.840 304.990 4757.440 ;
        RECT 89.350 4670.110 93.350 4733.550 ;
        RECT 154.100 4727.770 157.870 4733.160 ;
        RECT 95.350 4661.740 99.350 4726.660 ;
        RECT 3253.270 4726.120 3256.010 4731.730 ;
        RECT 3376.680 4725.870 3382.710 4731.940 ;
        RECT 186.790 4719.900 190.600 4725.320 ;
        RECT 3258.010 4718.060 3260.850 4723.750 ;
        RECT 3358.200 4717.870 3364.230 4723.940 ;
        RECT 3430.010 4709.770 3433.780 4715.160 ;
        RECT 3397.280 4701.900 3401.090 4707.320 ;
        RECT 3489.780 4643.740 3493.780 4708.660 ;
        RECT 3495.780 4652.110 3499.780 4715.550 ;
        RECT 3548.600 4657.380 3552.600 4724.210 ;
        RECT 3554.600 4648.730 3558.600 4732.350 ;
        RECT 3253.270 4500.120 3256.010 4505.730 ;
        RECT 3373.150 4499.910 3379.150 4505.910 ;
        RECT 3258.010 4492.060 3260.850 4497.750 ;
        RECT 3357.380 4491.910 3363.380 4497.910 ;
        RECT 154.235 4447.440 157.755 4448.560 ;
        RECT 186.935 4441.455 190.455 4442.575 ;
        RECT 3253.270 4275.120 3256.010 4280.730 ;
        RECT 3370.270 4274.910 3376.270 4280.910 ;
        RECT 3258.010 4267.060 3260.850 4272.750 ;
        RECT 3357.540 4266.910 3363.540 4272.910 ;
        RECT 221.000 4130.610 233.960 4136.630 ;
        RECT 307.120 4130.800 309.810 4136.400 ;
        RECT 204.970 4122.630 217.940 4128.610 ;
        RECT 302.300 4122.840 304.990 4128.440 ;
        RECT 89.350 4041.110 93.350 4104.550 ;
        RECT 154.100 4098.770 157.870 4104.160 ;
        RECT 95.350 4032.740 99.350 4097.660 ;
        RECT 186.790 4090.900 190.600 4096.320 ;
        RECT 221.000 3922.610 233.960 3928.630 ;
        RECT 307.120 3922.800 309.810 3928.400 ;
        RECT 204.970 3914.630 217.940 3920.610 ;
        RECT 302.300 3914.840 304.990 3920.440 ;
        RECT 89.350 3825.110 93.350 3888.550 ;
        RECT 154.100 3882.770 157.870 3888.160 ;
        RECT 95.350 3816.740 99.350 3881.660 ;
        RECT 186.790 3874.900 190.600 3880.320 ;
        RECT 3253.270 3834.120 3256.010 3839.730 ;
        RECT 3376.730 3833.870 3382.760 3839.940 ;
        RECT 3258.010 3826.060 3260.850 3831.750 ;
        RECT 3358.250 3825.870 3364.280 3831.940 ;
        RECT 3430.060 3817.770 3433.830 3823.160 ;
        RECT 3397.330 3809.900 3401.140 3815.320 ;
        RECT 3489.830 3751.740 3493.830 3816.660 ;
        RECT 3495.830 3760.110 3499.830 3823.550 ;
        RECT 3548.650 3765.380 3552.650 3832.210 ;
        RECT 3554.650 3756.730 3558.650 3840.350 ;
        RECT 221.000 3698.610 233.960 3704.630 ;
        RECT 307.120 3698.800 309.810 3704.400 ;
        RECT 204.970 3690.630 217.940 3696.610 ;
        RECT 302.300 3690.840 304.990 3696.440 ;
        RECT 89.350 3609.110 93.350 3672.550 ;
        RECT 154.100 3666.770 157.870 3672.160 ;
        RECT 95.350 3600.740 99.350 3665.660 ;
        RECT 186.790 3658.900 190.600 3664.320 ;
        RECT 3429.885 3622.840 3433.405 3623.960 ;
        RECT 3397.435 3616.860 3400.955 3617.980 ;
        RECT 3253.270 3609.120 3256.010 3614.730 ;
        RECT 3376.730 3608.870 3382.760 3614.940 ;
        RECT 3258.010 3601.060 3260.850 3606.750 ;
        RECT 3358.250 3600.870 3364.280 3606.940 ;
        RECT 3430.060 3592.770 3433.830 3598.160 ;
        RECT 3397.330 3584.900 3401.140 3590.320 ;
        RECT 3489.830 3526.740 3493.830 3591.660 ;
        RECT 3495.830 3535.110 3499.830 3598.550 ;
        RECT 3548.650 3540.380 3552.650 3607.210 ;
        RECT 3554.650 3531.730 3558.650 3615.350 ;
        RECT 221.000 3482.610 233.960 3488.630 ;
        RECT 307.120 3482.800 309.810 3488.400 ;
        RECT 204.970 3474.630 217.940 3480.610 ;
        RECT 302.300 3474.840 304.990 3480.440 ;
        RECT 89.350 3393.110 93.350 3456.550 ;
        RECT 154.100 3450.770 157.870 3456.160 ;
        RECT 95.350 3384.740 99.350 3449.660 ;
        RECT 186.790 3442.900 190.600 3448.320 ;
        RECT 3253.270 3383.120 3256.010 3388.730 ;
        RECT 3376.730 3382.870 3382.760 3388.940 ;
        RECT 3258.010 3375.060 3260.850 3380.750 ;
        RECT 3358.250 3374.870 3364.280 3380.940 ;
        RECT 3430.060 3366.770 3433.830 3372.160 ;
        RECT 3397.330 3358.900 3401.140 3364.320 ;
        RECT 3489.830 3300.740 3493.830 3365.660 ;
        RECT 3495.830 3309.110 3499.830 3372.550 ;
        RECT 3548.650 3314.380 3552.650 3381.210 ;
        RECT 3554.650 3305.730 3558.650 3389.350 ;
        RECT 221.000 3266.610 233.960 3272.630 ;
        RECT 307.120 3266.800 309.810 3272.400 ;
        RECT 204.970 3258.630 217.940 3264.610 ;
        RECT 302.300 3258.840 304.990 3264.440 ;
        RECT 89.350 3177.110 93.350 3240.550 ;
        RECT 154.100 3234.770 157.870 3240.160 ;
        RECT 95.350 3168.740 99.350 3233.660 ;
        RECT 186.790 3226.900 190.600 3232.320 ;
        RECT 3253.270 3158.120 3256.010 3163.730 ;
        RECT 3376.730 3157.870 3382.760 3163.940 ;
        RECT 3358.250 3149.870 3364.280 3155.940 ;
        RECT 3258.010 3144.060 3260.850 3149.750 ;
        RECT 3430.060 3141.770 3433.830 3147.160 ;
        RECT 3397.330 3133.900 3401.140 3139.320 ;
        RECT 3489.830 3075.740 3493.830 3140.660 ;
        RECT 3495.830 3084.110 3499.830 3147.550 ;
        RECT 3548.650 3089.380 3552.650 3156.210 ;
        RECT 3554.650 3080.730 3558.650 3164.350 ;
        RECT 221.000 3055.910 233.960 3061.930 ;
        RECT 307.120 3056.100 309.810 3061.700 ;
        RECT 204.970 3047.930 217.940 3053.910 ;
        RECT 302.300 3048.140 304.990 3053.740 ;
        RECT 89.350 2961.110 93.350 3024.550 ;
        RECT 154.100 3018.770 157.870 3024.160 ;
        RECT 95.350 2952.740 99.350 3017.660 ;
        RECT 186.790 3010.900 190.600 3016.320 ;
        RECT 3253.270 2932.120 3256.010 2937.730 ;
        RECT 3376.730 2931.870 3382.760 2937.940 ;
        RECT 3258.010 2924.060 3260.850 2929.750 ;
        RECT 3358.250 2923.870 3364.280 2929.940 ;
        RECT 3430.060 2915.770 3433.830 2921.160 ;
        RECT 3397.330 2907.900 3401.140 2913.320 ;
        RECT 3489.830 2849.740 3493.830 2914.660 ;
        RECT 3495.830 2858.110 3499.830 2921.550 ;
        RECT 3548.650 2863.380 3552.650 2930.210 ;
        RECT 3554.650 2854.730 3558.650 2938.350 ;
        RECT 221.000 2834.610 233.960 2840.630 ;
        RECT 307.120 2834.800 309.810 2840.400 ;
        RECT 204.970 2826.630 217.940 2832.610 ;
        RECT 302.300 2826.840 304.990 2832.440 ;
        RECT 89.350 2745.110 93.350 2808.550 ;
        RECT 154.100 2802.770 157.870 2808.160 ;
        RECT 95.350 2736.740 99.350 2801.660 ;
        RECT 186.790 2794.900 190.600 2800.320 ;
        RECT 3253.270 2707.120 3256.010 2712.730 ;
        RECT 3376.730 2706.870 3382.760 2712.940 ;
        RECT 3258.010 2699.060 3260.850 2704.750 ;
        RECT 3358.250 2698.870 3364.280 2704.940 ;
        RECT 3430.060 2690.770 3433.830 2696.160 ;
        RECT 3397.330 2682.900 3401.140 2688.320 ;
        RECT 3489.830 2624.740 3493.830 2689.660 ;
        RECT 3495.830 2633.110 3499.830 2696.550 ;
        RECT 3548.650 2638.380 3552.650 2705.210 ;
        RECT 3554.650 2629.730 3558.650 2713.350 ;
        RECT 3253.270 2490.120 3256.010 2495.730 ;
        RECT 3376.730 2486.870 3382.760 2492.940 ;
        RECT 3258.010 2479.060 3260.850 2484.750 ;
        RECT 3358.250 2478.870 3364.280 2484.940 ;
        RECT 3430.060 2470.770 3433.830 2476.160 ;
        RECT 3397.330 2462.900 3401.140 2468.320 ;
        RECT 3489.830 2404.740 3493.830 2469.660 ;
        RECT 3495.830 2413.110 3499.830 2476.550 ;
        RECT 3548.650 2418.380 3552.650 2485.210 ;
        RECT 3554.650 2409.730 3558.650 2493.350 ;
        RECT 3429.885 2240.835 3433.405 2241.955 ;
        RECT 3397.435 2234.855 3400.955 2235.975 ;
        RECT 221.000 2196.610 233.960 2202.630 ;
        RECT 307.120 2196.800 309.810 2202.400 ;
        RECT 204.970 2188.630 217.940 2194.610 ;
        RECT 302.300 2188.840 304.990 2194.440 ;
        RECT 89.350 2107.110 93.350 2170.550 ;
        RECT 154.100 2164.770 157.870 2170.160 ;
        RECT 95.350 2098.740 99.350 2163.660 ;
        RECT 186.790 2156.900 190.600 2162.320 ;
        RECT 3253.270 2046.120 3256.010 2051.730 ;
        RECT 3376.730 2045.870 3382.760 2051.940 ;
        RECT 3258.010 2038.060 3260.850 2043.750 ;
        RECT 3358.250 2037.870 3364.280 2043.940 ;
        RECT 3430.060 2029.770 3433.830 2035.160 ;
        RECT 3397.330 2021.900 3401.140 2027.320 ;
        RECT 221.000 1980.610 233.960 1986.630 ;
        RECT 307.120 1980.800 309.810 1986.400 ;
        RECT 204.970 1972.630 217.940 1978.610 ;
        RECT 302.300 1972.840 304.990 1978.440 ;
        RECT 3489.830 1963.740 3493.830 2028.660 ;
        RECT 3495.830 1972.110 3499.830 2035.550 ;
        RECT 3548.650 1977.380 3552.650 2044.210 ;
        RECT 3554.650 1968.730 3558.650 2052.350 ;
        RECT 89.350 1891.110 93.350 1954.550 ;
        RECT 154.100 1948.770 157.870 1954.160 ;
        RECT 95.350 1882.740 99.350 1947.660 ;
        RECT 186.790 1940.900 190.600 1946.320 ;
        RECT 3253.270 1827.120 3256.010 1832.730 ;
        RECT 3376.730 1819.870 3382.760 1825.940 ;
        RECT 3258.010 1812.060 3260.850 1817.750 ;
        RECT 3358.250 1811.870 3364.280 1817.940 ;
        RECT 3430.060 1803.770 3433.830 1809.160 ;
        RECT 3397.330 1795.900 3401.140 1801.320 ;
        RECT 221.000 1769.610 233.960 1775.630 ;
        RECT 307.120 1769.800 309.810 1775.400 ;
        RECT 204.970 1761.630 217.940 1767.610 ;
        RECT 302.300 1761.840 304.990 1767.440 ;
        RECT 89.350 1675.110 93.350 1738.550 ;
        RECT 154.100 1732.770 157.870 1738.160 ;
        RECT 3489.830 1737.740 3493.830 1802.660 ;
        RECT 3495.830 1746.110 3499.830 1809.550 ;
        RECT 3548.650 1751.380 3552.650 1818.210 ;
        RECT 3554.650 1742.730 3558.650 1826.350 ;
        RECT 95.350 1666.740 99.350 1731.660 ;
        RECT 186.790 1724.900 190.600 1730.320 ;
        RECT 3253.270 1595.120 3256.010 1600.730 ;
        RECT 3376.730 1594.870 3382.760 1600.940 ;
        RECT 3258.010 1587.060 3260.850 1592.750 ;
        RECT 3358.250 1586.870 3364.280 1592.940 ;
        RECT 3430.060 1578.770 3433.830 1584.160 ;
        RECT 3397.330 1570.900 3401.140 1576.320 ;
        RECT 221.000 1548.610 233.960 1554.630 ;
        RECT 307.120 1548.800 309.810 1554.400 ;
        RECT 204.970 1540.630 217.940 1546.610 ;
        RECT 302.300 1540.840 304.990 1546.440 ;
        RECT 89.350 1459.110 93.350 1522.550 ;
        RECT 154.100 1516.770 157.870 1522.160 ;
        RECT 95.350 1450.740 99.350 1515.660 ;
        RECT 186.790 1508.900 190.600 1514.320 ;
        RECT 3489.830 1512.740 3493.830 1577.660 ;
        RECT 3495.830 1521.110 3499.830 1584.550 ;
        RECT 3548.650 1526.380 3552.650 1593.210 ;
        RECT 3554.650 1517.730 3558.650 1601.350 ;
        RECT 3294.410 1388.870 3383.140 1392.030 ;
        RECT 220.975 1382.420 234.010 1386.420 ;
        RECT 3294.280 1384.080 3367.250 1387.280 ;
        RECT 220.975 1379.290 282.160 1382.420 ;
        RECT 3354.090 1380.080 3367.250 1384.080 ;
        RECT 3370.080 1383.870 3383.140 1388.870 ;
        RECT 213.730 1374.530 282.240 1377.660 ;
        RECT 213.730 1346.390 218.050 1374.530 ;
        RECT 3376.730 1369.870 3382.760 1375.940 ;
        RECT 3358.250 1361.870 3364.280 1367.940 ;
        RECT 3430.060 1353.770 3433.830 1359.160 ;
        RECT 3397.330 1345.900 3401.140 1351.320 ;
        RECT 89.350 1243.110 93.350 1306.550 ;
        RECT 154.100 1300.770 157.870 1306.160 ;
        RECT 95.350 1234.740 99.350 1299.660 ;
        RECT 186.790 1292.900 190.600 1298.320 ;
        RECT 3489.830 1287.740 3493.830 1352.660 ;
        RECT 3495.830 1296.110 3499.830 1359.550 ;
        RECT 3548.650 1301.380 3552.650 1368.210 ;
        RECT 3554.650 1292.730 3558.650 1376.350 ;
        RECT 3376.730 1143.870 3382.760 1149.940 ;
        RECT 3358.250 1135.870 3364.280 1141.940 ;
        RECT 3430.060 1127.770 3433.830 1133.160 ;
        RECT 3397.330 1119.900 3401.140 1125.320 ;
        RECT 89.350 1027.110 93.350 1090.550 ;
        RECT 154.100 1084.770 157.870 1090.160 ;
        RECT 95.350 1018.740 99.350 1083.660 ;
        RECT 186.790 1076.900 190.600 1082.320 ;
        RECT 3489.830 1061.740 3493.830 1126.660 ;
        RECT 3495.830 1070.110 3499.830 1133.550 ;
        RECT 3548.650 1075.380 3552.650 1142.210 ;
        RECT 3554.650 1066.730 3558.650 1150.350 ;
        RECT 3376.730 918.870 3382.760 924.940 ;
        RECT 3358.250 910.870 3364.280 916.940 ;
        RECT 3430.060 902.770 3433.830 908.160 ;
        RECT 3397.330 894.900 3401.140 900.320 ;
        RECT 3489.830 836.740 3493.830 901.660 ;
        RECT 3495.830 845.110 3499.830 908.550 ;
        RECT 3548.650 850.380 3552.650 917.210 ;
        RECT 3554.650 841.730 3558.650 925.350 ;
        RECT 3376.730 692.870 3382.760 698.940 ;
        RECT 3358.250 684.870 3364.280 690.940 ;
        RECT 3430.060 676.770 3433.830 682.160 ;
        RECT 3397.330 668.900 3401.140 674.320 ;
        RECT 3489.830 610.740 3493.830 675.660 ;
        RECT 3495.830 619.110 3499.830 682.550 ;
        RECT 3548.650 624.380 3552.650 691.210 ;
        RECT 3554.650 615.730 3558.650 699.350 ;
        RECT 2281.685 243.200 2299.120 245.200 ;
        RECT 717.200 208.000 718.100 236.480 ;
        RECT 643.050 206.310 647.340 208.000 ;
        RECT 716.450 206.310 718.230 208.000 ;
        RECT 723.700 204.610 724.600 236.700 ;
        RECT 745.670 209.380 746.570 210.455 ;
        RECT 650.710 202.910 655.000 204.610 ;
        RECT 722.950 202.910 724.725 204.610 ;
        RECT 738.970 200.290 740.895 209.380 ;
        RECT 2202.120 205.790 2203.970 210.390 ;
        RECT 2135.095 204.890 2203.970 205.790 ;
        RECT 2208.015 203.810 2210.045 203.885 ;
        RECT 2130.090 202.910 2210.045 203.810 ;
        RECT 2208.015 202.820 2210.045 202.910 ;
        RECT 2281.685 199.890 2283.590 243.200 ;
        RECT 2302.000 241.200 2303.600 245.200 ;
        RECT 2286.695 239.200 2303.600 241.200 ;
        RECT 2286.695 199.890 2288.600 239.200 ;
        RECT 3209.680 238.135 3251.010 240.135 ;
        RECT 3209.680 210.820 3218.590 238.135 ;
        RECT 3267.160 212.440 3284.560 235.270 ;
        RECT 739.085 186.710 740.800 190.915 ;
        RECT 2135.225 186.860 2136.865 190.765 ;
        RECT 2281.825 186.860 2283.465 190.765 ;
        RECT 650.860 175.830 654.880 179.980 ;
        RECT 643.210 169.790 647.230 173.940 ;
        RECT 3210.130 169.940 3218.170 173.800 ;
        RECT 2130.220 154.190 2131.860 158.095 ;
        RECT 2286.830 154.190 2288.470 158.095 ;
      LAYER via4 ;
        RECT 500.410 5095.320 501.850 5099.180 ;
        RECT 517.320 5095.330 518.760 5099.190 ;
        RECT 534.230 5095.300 535.670 5099.160 ;
        RECT 558.280 5095.360 559.690 5099.140 ;
        RECT 757.410 5095.320 758.850 5099.180 ;
        RECT 774.320 5095.330 775.760 5099.190 ;
        RECT 791.230 5095.300 792.670 5099.160 ;
        RECT 815.280 5095.360 816.690 5099.140 ;
        RECT 1014.410 5095.320 1015.850 5099.180 ;
        RECT 1031.320 5095.330 1032.760 5099.190 ;
        RECT 1048.230 5095.300 1049.670 5099.160 ;
        RECT 1072.280 5095.360 1073.690 5099.140 ;
        RECT 1271.410 5095.320 1272.850 5099.180 ;
        RECT 1288.320 5095.330 1289.760 5099.190 ;
        RECT 1305.230 5095.300 1306.670 5099.160 ;
        RECT 1329.280 5095.360 1330.690 5099.140 ;
        RECT 1529.410 5095.320 1530.850 5099.180 ;
        RECT 1546.320 5095.330 1547.760 5099.190 ;
        RECT 1563.230 5095.300 1564.670 5099.160 ;
        RECT 1587.280 5095.360 1588.690 5099.140 ;
        RECT 1781.410 5095.320 1782.850 5099.180 ;
        RECT 1798.320 5095.330 1799.760 5099.190 ;
        RECT 1815.230 5095.300 1816.670 5099.160 ;
        RECT 1839.280 5095.360 1840.690 5099.140 ;
        RECT 2118.410 5095.320 2119.850 5099.180 ;
        RECT 2135.320 5095.330 2136.760 5099.190 ;
        RECT 2152.230 5095.300 2153.670 5099.160 ;
        RECT 2176.280 5095.360 2177.690 5099.140 ;
        RECT 2503.410 5095.320 2504.850 5099.180 ;
        RECT 2520.320 5095.330 2521.760 5099.190 ;
        RECT 2537.230 5095.300 2538.670 5099.160 ;
        RECT 2561.280 5095.360 2562.690 5099.140 ;
        RECT 2760.410 5095.320 2761.850 5099.180 ;
        RECT 2777.320 5095.330 2778.760 5099.190 ;
        RECT 2794.230 5095.300 2795.670 5099.160 ;
        RECT 2818.280 5095.360 2819.690 5099.140 ;
        RECT 491.980 5089.300 493.420 5093.160 ;
        RECT 508.880 5089.300 510.320 5093.160 ;
        RECT 525.780 5089.320 527.220 5093.180 ;
        RECT 554.760 5089.360 556.170 5093.140 ;
        RECT 748.980 5089.300 750.420 5093.160 ;
        RECT 765.880 5089.300 767.320 5093.160 ;
        RECT 782.780 5089.320 784.220 5093.180 ;
        RECT 811.760 5089.360 813.170 5093.140 ;
        RECT 1005.980 5089.300 1007.420 5093.160 ;
        RECT 1022.880 5089.300 1024.320 5093.160 ;
        RECT 1039.780 5089.320 1041.220 5093.180 ;
        RECT 1068.760 5089.360 1070.170 5093.140 ;
        RECT 1262.980 5089.300 1264.420 5093.160 ;
        RECT 1279.880 5089.300 1281.320 5093.160 ;
        RECT 1296.780 5089.320 1298.220 5093.180 ;
        RECT 1325.760 5089.360 1327.170 5093.140 ;
        RECT 1520.980 5089.300 1522.420 5093.160 ;
        RECT 1537.880 5089.300 1539.320 5093.160 ;
        RECT 1554.780 5089.320 1556.220 5093.180 ;
        RECT 1583.760 5089.360 1585.170 5093.140 ;
        RECT 1772.980 5089.300 1774.420 5093.160 ;
        RECT 1789.880 5089.300 1791.320 5093.160 ;
        RECT 1806.780 5089.320 1808.220 5093.180 ;
        RECT 1835.760 5089.360 1837.170 5093.140 ;
        RECT 2109.980 5089.300 2111.420 5093.160 ;
        RECT 2126.880 5089.300 2128.320 5093.160 ;
        RECT 2143.780 5089.320 2145.220 5093.180 ;
        RECT 2172.760 5089.360 2174.170 5093.140 ;
        RECT 2494.980 5089.300 2496.420 5093.160 ;
        RECT 2511.880 5089.300 2513.320 5093.160 ;
        RECT 2528.780 5089.320 2530.220 5093.180 ;
        RECT 2557.760 5089.360 2559.170 5093.140 ;
        RECT 2751.980 5089.300 2753.420 5093.160 ;
        RECT 2768.880 5089.300 2770.320 5093.160 ;
        RECT 2785.780 5089.320 2787.220 5093.180 ;
        RECT 2814.760 5089.360 2816.170 5093.140 ;
        RECT 205.330 4929.425 217.710 4932.205 ;
        RECT 279.065 4930.215 280.245 4931.395 ;
        RECT 280.665 4930.215 281.845 4931.395 ;
        RECT 221.345 4924.650 233.725 4927.430 ;
        RECT 279.140 4924.595 281.920 4927.375 ;
        RECT 3291.955 4920.600 3293.135 4921.780 ;
        RECT 3293.555 4920.600 3294.735 4921.780 ;
        RECT 3295.155 4920.600 3296.335 4921.780 ;
        RECT 3296.755 4920.600 3297.935 4921.780 ;
        RECT 3298.355 4920.600 3299.535 4921.780 ;
        RECT 3299.955 4920.600 3301.135 4921.780 ;
        RECT 3301.555 4920.600 3302.735 4921.780 ;
        RECT 3303.155 4920.600 3304.335 4921.780 ;
        RECT 3304.755 4920.600 3305.935 4921.780 ;
        RECT 3306.355 4920.600 3307.535 4921.780 ;
        RECT 3307.955 4920.600 3309.135 4921.780 ;
        RECT 3309.555 4920.600 3310.735 4921.780 ;
        RECT 3311.155 4920.600 3312.335 4921.780 ;
        RECT 3312.755 4920.600 3313.935 4921.780 ;
        RECT 3314.355 4920.600 3315.535 4921.780 ;
        RECT 3354.415 4919.825 3366.795 4922.605 ;
        RECT 3291.865 4915.820 3293.045 4917.000 ;
        RECT 3293.465 4915.820 3294.645 4917.000 ;
        RECT 3295.065 4915.820 3296.245 4917.000 ;
        RECT 3296.665 4915.820 3297.845 4917.000 ;
        RECT 3298.265 4915.820 3299.445 4917.000 ;
        RECT 3299.865 4915.820 3301.045 4917.000 ;
        RECT 3301.465 4915.820 3302.645 4917.000 ;
        RECT 3303.065 4915.820 3304.245 4917.000 ;
        RECT 3304.665 4915.820 3305.845 4917.000 ;
        RECT 3306.265 4915.820 3307.445 4917.000 ;
        RECT 3307.865 4915.820 3309.045 4917.000 ;
        RECT 3309.465 4915.820 3310.645 4917.000 ;
        RECT 3311.065 4915.820 3312.245 4917.000 ;
        RECT 3312.665 4915.820 3313.845 4917.000 ;
        RECT 3314.265 4915.820 3315.445 4917.000 ;
        RECT 3370.405 4915.015 3382.785 4917.795 ;
        RECT 222.140 4760.325 232.920 4764.705 ;
        RECT 206.090 4752.415 216.870 4756.795 ;
        RECT 89.450 4728.280 93.230 4729.690 ;
        RECT 89.430 4704.230 93.290 4705.670 ;
        RECT 89.400 4687.320 93.260 4688.760 ;
        RECT 89.410 4670.410 93.270 4671.850 ;
        RECT 95.450 4724.760 99.230 4726.170 ;
        RECT 3376.990 4726.240 3382.400 4731.730 ;
        RECT 3358.460 4718.150 3363.870 4723.640 ;
        RECT 3495.900 4710.280 3499.680 4711.690 ;
        RECT 3489.900 4706.760 3493.680 4708.170 ;
        RECT 95.410 4695.780 99.270 4697.220 ;
        RECT 95.430 4678.880 99.290 4680.320 ;
        RECT 95.430 4661.980 99.290 4663.420 ;
        RECT 3489.860 4677.780 3493.720 4679.220 ;
        RECT 3489.840 4660.880 3493.700 4662.320 ;
        RECT 3495.840 4686.230 3499.700 4687.670 ;
        RECT 3495.870 4669.320 3499.730 4670.760 ;
        RECT 3548.680 4691.500 3552.510 4692.850 ;
        RECT 3548.690 4674.580 3552.520 4675.930 ;
        RECT 3548.680 4657.640 3552.550 4659.130 ;
        RECT 3554.690 4683.020 3558.520 4684.370 ;
        RECT 3554.660 4666.220 3558.490 4667.570 ;
        RECT 3495.860 4652.410 3499.720 4653.850 ;
        RECT 3554.650 4649.200 3558.520 4650.690 ;
        RECT 3489.840 4643.980 3493.700 4645.420 ;
        RECT 3373.995 4500.775 3378.375 4505.155 ;
        RECT 3358.215 4492.735 3362.595 4497.115 ;
        RECT 3371.050 4275.730 3375.430 4280.110 ;
        RECT 3358.330 4267.720 3362.710 4272.100 ;
        RECT 222.140 4131.325 232.920 4135.705 ;
        RECT 206.090 4123.415 216.870 4127.795 ;
        RECT 89.450 4099.280 93.230 4100.690 ;
        RECT 89.430 4075.230 93.290 4076.670 ;
        RECT 89.400 4058.320 93.260 4059.760 ;
        RECT 89.410 4041.410 93.270 4042.850 ;
        RECT 95.450 4095.760 99.230 4097.170 ;
        RECT 95.410 4066.780 99.270 4068.220 ;
        RECT 95.430 4049.880 99.290 4051.320 ;
        RECT 95.430 4032.980 99.290 4034.420 ;
        RECT 222.140 3923.325 232.920 3927.705 ;
        RECT 206.090 3915.415 216.870 3919.795 ;
        RECT 89.450 3883.280 93.230 3884.690 ;
        RECT 89.430 3859.230 93.290 3860.670 ;
        RECT 89.400 3842.320 93.260 3843.760 ;
        RECT 89.410 3825.410 93.270 3826.850 ;
        RECT 95.450 3879.760 99.230 3881.170 ;
        RECT 95.410 3850.780 99.270 3852.220 ;
        RECT 95.430 3833.880 99.290 3835.320 ;
        RECT 3377.040 3834.240 3382.450 3839.730 ;
        RECT 3358.510 3826.150 3363.920 3831.640 ;
        RECT 95.430 3816.980 99.290 3818.420 ;
        RECT 3495.950 3818.280 3499.730 3819.690 ;
        RECT 3489.950 3814.760 3493.730 3816.170 ;
        RECT 3489.910 3785.780 3493.770 3787.220 ;
        RECT 3489.890 3768.880 3493.750 3770.320 ;
        RECT 3495.890 3794.230 3499.750 3795.670 ;
        RECT 3495.920 3777.320 3499.780 3778.760 ;
        RECT 3548.730 3799.500 3552.560 3800.850 ;
        RECT 3548.740 3782.580 3552.570 3783.930 ;
        RECT 3548.730 3765.640 3552.600 3767.130 ;
        RECT 3554.740 3791.020 3558.570 3792.370 ;
        RECT 3554.710 3774.220 3558.540 3775.570 ;
        RECT 3495.910 3760.410 3499.770 3761.850 ;
        RECT 3554.700 3757.200 3558.570 3758.690 ;
        RECT 3489.890 3751.980 3493.750 3753.420 ;
        RECT 222.140 3699.325 232.920 3703.705 ;
        RECT 206.090 3691.415 216.870 3695.795 ;
        RECT 89.450 3667.280 93.230 3668.690 ;
        RECT 89.430 3643.230 93.290 3644.670 ;
        RECT 89.400 3626.320 93.260 3627.760 ;
        RECT 89.410 3609.410 93.270 3610.850 ;
        RECT 95.450 3663.760 99.230 3665.170 ;
        RECT 95.410 3634.780 99.270 3636.220 ;
        RECT 95.430 3617.880 99.290 3619.320 ;
        RECT 3377.040 3609.240 3382.450 3614.730 ;
        RECT 95.430 3600.980 99.290 3602.420 ;
        RECT 3358.510 3601.150 3363.920 3606.640 ;
        RECT 3495.950 3593.280 3499.730 3594.690 ;
        RECT 3489.950 3589.760 3493.730 3591.170 ;
        RECT 3489.910 3560.780 3493.770 3562.220 ;
        RECT 3489.890 3543.880 3493.750 3545.320 ;
        RECT 3495.890 3569.230 3499.750 3570.670 ;
        RECT 3495.920 3552.320 3499.780 3553.760 ;
        RECT 3548.730 3574.500 3552.560 3575.850 ;
        RECT 3548.740 3557.580 3552.570 3558.930 ;
        RECT 3548.730 3540.640 3552.600 3542.130 ;
        RECT 3554.740 3566.020 3558.570 3567.370 ;
        RECT 3554.710 3549.220 3558.540 3550.570 ;
        RECT 3495.910 3535.410 3499.770 3536.850 ;
        RECT 3554.700 3532.200 3558.570 3533.690 ;
        RECT 3489.890 3526.980 3493.750 3528.420 ;
        RECT 222.140 3483.325 232.920 3487.705 ;
        RECT 206.090 3475.415 216.870 3479.795 ;
        RECT 89.450 3451.280 93.230 3452.690 ;
        RECT 89.430 3427.230 93.290 3428.670 ;
        RECT 89.400 3410.320 93.260 3411.760 ;
        RECT 89.410 3393.410 93.270 3394.850 ;
        RECT 95.450 3447.760 99.230 3449.170 ;
        RECT 95.410 3418.780 99.270 3420.220 ;
        RECT 95.430 3401.880 99.290 3403.320 ;
        RECT 95.430 3384.980 99.290 3386.420 ;
        RECT 3377.040 3383.240 3382.450 3388.730 ;
        RECT 3358.510 3375.150 3363.920 3380.640 ;
        RECT 3495.950 3367.280 3499.730 3368.690 ;
        RECT 3489.950 3363.760 3493.730 3365.170 ;
        RECT 3489.910 3334.780 3493.770 3336.220 ;
        RECT 3489.890 3317.880 3493.750 3319.320 ;
        RECT 3495.890 3343.230 3499.750 3344.670 ;
        RECT 3495.920 3326.320 3499.780 3327.760 ;
        RECT 3548.730 3348.500 3552.560 3349.850 ;
        RECT 3548.740 3331.580 3552.570 3332.930 ;
        RECT 3548.730 3314.640 3552.600 3316.130 ;
        RECT 3554.740 3340.020 3558.570 3341.370 ;
        RECT 3554.710 3323.220 3558.540 3324.570 ;
        RECT 3495.910 3309.410 3499.770 3310.850 ;
        RECT 3554.700 3306.200 3558.570 3307.690 ;
        RECT 3489.890 3300.980 3493.750 3302.420 ;
        RECT 222.140 3267.325 232.920 3271.705 ;
        RECT 206.090 3259.415 216.870 3263.795 ;
        RECT 89.450 3235.280 93.230 3236.690 ;
        RECT 89.430 3211.230 93.290 3212.670 ;
        RECT 89.400 3194.320 93.260 3195.760 ;
        RECT 89.410 3177.410 93.270 3178.850 ;
        RECT 95.450 3231.760 99.230 3233.170 ;
        RECT 95.410 3202.780 99.270 3204.220 ;
        RECT 95.430 3185.880 99.290 3187.320 ;
        RECT 95.430 3168.980 99.290 3170.420 ;
        RECT 3377.040 3158.240 3382.450 3163.730 ;
        RECT 3358.510 3150.150 3363.920 3155.640 ;
        RECT 3495.950 3142.280 3499.730 3143.690 ;
        RECT 3489.950 3138.760 3493.730 3140.170 ;
        RECT 3489.910 3109.780 3493.770 3111.220 ;
        RECT 3489.890 3092.880 3493.750 3094.320 ;
        RECT 3495.890 3118.230 3499.750 3119.670 ;
        RECT 3495.920 3101.320 3499.780 3102.760 ;
        RECT 3548.730 3123.500 3552.560 3124.850 ;
        RECT 3548.740 3106.580 3552.570 3107.930 ;
        RECT 3548.730 3089.640 3552.600 3091.130 ;
        RECT 3554.740 3115.020 3558.570 3116.370 ;
        RECT 3554.710 3098.220 3558.540 3099.570 ;
        RECT 3495.910 3084.410 3499.770 3085.850 ;
        RECT 3554.700 3081.200 3558.570 3082.690 ;
        RECT 3489.890 3075.980 3493.750 3077.420 ;
        RECT 222.140 3056.625 232.920 3061.005 ;
        RECT 206.090 3048.715 216.870 3053.095 ;
        RECT 89.450 3019.280 93.230 3020.690 ;
        RECT 89.430 2995.230 93.290 2996.670 ;
        RECT 89.400 2978.320 93.260 2979.760 ;
        RECT 89.410 2961.410 93.270 2962.850 ;
        RECT 95.450 3015.760 99.230 3017.170 ;
        RECT 95.410 2986.780 99.270 2988.220 ;
        RECT 95.430 2969.880 99.290 2971.320 ;
        RECT 95.430 2952.980 99.290 2954.420 ;
        RECT 3377.040 2932.240 3382.450 2937.730 ;
        RECT 3358.510 2924.150 3363.920 2929.640 ;
        RECT 3495.950 2916.280 3499.730 2917.690 ;
        RECT 3489.950 2912.760 3493.730 2914.170 ;
        RECT 3489.910 2883.780 3493.770 2885.220 ;
        RECT 3489.890 2866.880 3493.750 2868.320 ;
        RECT 3495.890 2892.230 3499.750 2893.670 ;
        RECT 3495.920 2875.320 3499.780 2876.760 ;
        RECT 3548.730 2897.500 3552.560 2898.850 ;
        RECT 3548.740 2880.580 3552.570 2881.930 ;
        RECT 3548.730 2863.640 3552.600 2865.130 ;
        RECT 3554.740 2889.020 3558.570 2890.370 ;
        RECT 3554.710 2872.220 3558.540 2873.570 ;
        RECT 3495.910 2858.410 3499.770 2859.850 ;
        RECT 3554.700 2855.200 3558.570 2856.690 ;
        RECT 3489.890 2849.980 3493.750 2851.420 ;
        RECT 222.140 2835.325 232.920 2839.705 ;
        RECT 206.090 2827.415 216.870 2831.795 ;
        RECT 89.450 2803.280 93.230 2804.690 ;
        RECT 89.430 2779.230 93.290 2780.670 ;
        RECT 89.400 2762.320 93.260 2763.760 ;
        RECT 89.410 2745.410 93.270 2746.850 ;
        RECT 95.450 2799.760 99.230 2801.170 ;
        RECT 95.410 2770.780 99.270 2772.220 ;
        RECT 95.430 2753.880 99.290 2755.320 ;
        RECT 95.430 2736.980 99.290 2738.420 ;
        RECT 3377.040 2707.240 3382.450 2712.730 ;
        RECT 3358.510 2699.150 3363.920 2704.640 ;
        RECT 3495.950 2691.280 3499.730 2692.690 ;
        RECT 3489.950 2687.760 3493.730 2689.170 ;
        RECT 3489.910 2658.780 3493.770 2660.220 ;
        RECT 3489.890 2641.880 3493.750 2643.320 ;
        RECT 3495.890 2667.230 3499.750 2668.670 ;
        RECT 3495.920 2650.320 3499.780 2651.760 ;
        RECT 3548.730 2672.500 3552.560 2673.850 ;
        RECT 3548.740 2655.580 3552.570 2656.930 ;
        RECT 3548.730 2638.640 3552.600 2640.130 ;
        RECT 3554.740 2664.020 3558.570 2665.370 ;
        RECT 3554.710 2647.220 3558.540 2648.570 ;
        RECT 3495.910 2633.410 3499.770 2634.850 ;
        RECT 3554.700 2630.200 3558.570 2631.690 ;
        RECT 3489.890 2624.980 3493.750 2626.420 ;
        RECT 3377.040 2487.240 3382.450 2492.730 ;
        RECT 3358.510 2479.150 3363.920 2484.640 ;
        RECT 3495.950 2471.280 3499.730 2472.690 ;
        RECT 3489.950 2467.760 3493.730 2469.170 ;
        RECT 3489.910 2438.780 3493.770 2440.220 ;
        RECT 3489.890 2421.880 3493.750 2423.320 ;
        RECT 3495.890 2447.230 3499.750 2448.670 ;
        RECT 3495.920 2430.320 3499.780 2431.760 ;
        RECT 3548.730 2452.500 3552.560 2453.850 ;
        RECT 3548.740 2435.580 3552.570 2436.930 ;
        RECT 3548.730 2418.640 3552.600 2420.130 ;
        RECT 3554.740 2444.020 3558.570 2445.370 ;
        RECT 3554.710 2427.220 3558.540 2428.570 ;
        RECT 3495.910 2413.410 3499.770 2414.850 ;
        RECT 3554.700 2410.200 3558.570 2411.690 ;
        RECT 3489.890 2404.980 3493.750 2406.420 ;
        RECT 222.140 2197.325 232.920 2201.705 ;
        RECT 206.090 2189.415 216.870 2193.795 ;
        RECT 89.450 2165.280 93.230 2166.690 ;
        RECT 89.430 2141.230 93.290 2142.670 ;
        RECT 89.400 2124.320 93.260 2125.760 ;
        RECT 89.410 2107.410 93.270 2108.850 ;
        RECT 95.450 2161.760 99.230 2163.170 ;
        RECT 95.410 2132.780 99.270 2134.220 ;
        RECT 95.430 2115.880 99.290 2117.320 ;
        RECT 95.430 2098.980 99.290 2100.420 ;
        RECT 3377.040 2046.240 3382.450 2051.730 ;
        RECT 3358.510 2038.150 3363.920 2043.640 ;
        RECT 3495.950 2030.280 3499.730 2031.690 ;
        RECT 3489.950 2026.760 3493.730 2028.170 ;
        RECT 3489.910 1997.780 3493.770 1999.220 ;
        RECT 222.140 1981.325 232.920 1985.705 ;
        RECT 3489.890 1980.880 3493.750 1982.320 ;
        RECT 206.090 1973.415 216.870 1977.795 ;
        RECT 3495.890 2006.230 3499.750 2007.670 ;
        RECT 3495.920 1989.320 3499.780 1990.760 ;
        RECT 3548.730 2011.500 3552.560 2012.850 ;
        RECT 3548.740 1994.580 3552.570 1995.930 ;
        RECT 3548.730 1977.640 3552.600 1979.130 ;
        RECT 3554.740 2003.020 3558.570 2004.370 ;
        RECT 3554.710 1986.220 3558.540 1987.570 ;
        RECT 3495.910 1972.410 3499.770 1973.850 ;
        RECT 3554.700 1969.200 3558.570 1970.690 ;
        RECT 3489.890 1963.980 3493.750 1965.420 ;
        RECT 89.450 1949.280 93.230 1950.690 ;
        RECT 89.430 1925.230 93.290 1926.670 ;
        RECT 89.400 1908.320 93.260 1909.760 ;
        RECT 89.410 1891.410 93.270 1892.850 ;
        RECT 95.450 1945.760 99.230 1947.170 ;
        RECT 95.410 1916.780 99.270 1918.220 ;
        RECT 95.430 1899.880 99.290 1901.320 ;
        RECT 95.430 1882.980 99.290 1884.420 ;
        RECT 3377.040 1820.240 3382.450 1825.730 ;
        RECT 3358.510 1812.150 3363.920 1817.640 ;
        RECT 3495.950 1804.280 3499.730 1805.690 ;
        RECT 3489.950 1800.760 3493.730 1802.170 ;
        RECT 222.140 1770.325 232.920 1774.705 ;
        RECT 3489.910 1771.780 3493.770 1773.220 ;
        RECT 206.090 1762.415 216.870 1766.795 ;
        RECT 3489.890 1754.880 3493.750 1756.320 ;
        RECT 3495.890 1780.230 3499.750 1781.670 ;
        RECT 3495.920 1763.320 3499.780 1764.760 ;
        RECT 3548.730 1785.500 3552.560 1786.850 ;
        RECT 3548.740 1768.580 3552.570 1769.930 ;
        RECT 3548.730 1751.640 3552.600 1753.130 ;
        RECT 3554.740 1777.020 3558.570 1778.370 ;
        RECT 3554.710 1760.220 3558.540 1761.570 ;
        RECT 3495.910 1746.410 3499.770 1747.850 ;
        RECT 3554.700 1743.200 3558.570 1744.690 ;
        RECT 89.450 1733.280 93.230 1734.690 ;
        RECT 3489.890 1737.980 3493.750 1739.420 ;
        RECT 89.430 1709.230 93.290 1710.670 ;
        RECT 89.400 1692.320 93.260 1693.760 ;
        RECT 89.410 1675.410 93.270 1676.850 ;
        RECT 95.450 1729.760 99.230 1731.170 ;
        RECT 95.410 1700.780 99.270 1702.220 ;
        RECT 95.430 1683.880 99.290 1685.320 ;
        RECT 95.430 1666.980 99.290 1668.420 ;
        RECT 3377.040 1595.240 3382.450 1600.730 ;
        RECT 3358.510 1587.150 3363.920 1592.640 ;
        RECT 3495.950 1579.280 3499.730 1580.690 ;
        RECT 3489.950 1575.760 3493.730 1577.170 ;
        RECT 222.140 1549.325 232.920 1553.705 ;
        RECT 3489.910 1546.780 3493.770 1548.220 ;
        RECT 206.090 1541.415 216.870 1545.795 ;
        RECT 3489.890 1529.880 3493.750 1531.320 ;
        RECT 89.450 1517.280 93.230 1518.690 ;
        RECT 89.430 1493.230 93.290 1494.670 ;
        RECT 89.400 1476.320 93.260 1477.760 ;
        RECT 89.410 1459.410 93.270 1460.850 ;
        RECT 95.450 1513.760 99.230 1515.170 ;
        RECT 3495.890 1555.230 3499.750 1556.670 ;
        RECT 3495.920 1538.320 3499.780 1539.760 ;
        RECT 3548.730 1560.500 3552.560 1561.850 ;
        RECT 3548.740 1543.580 3552.570 1544.930 ;
        RECT 3548.730 1526.640 3552.600 1528.130 ;
        RECT 3554.740 1552.020 3558.570 1553.370 ;
        RECT 3554.710 1535.220 3558.540 1536.570 ;
        RECT 3495.910 1521.410 3499.770 1522.850 ;
        RECT 3554.700 1518.200 3558.570 1519.690 ;
        RECT 3489.890 1512.980 3493.750 1514.420 ;
        RECT 95.410 1484.780 99.270 1486.220 ;
        RECT 95.430 1467.880 99.290 1469.320 ;
        RECT 95.430 1450.980 99.290 1452.420 ;
        RECT 3294.920 1389.875 3296.100 1391.055 ;
        RECT 3296.520 1389.875 3297.700 1391.055 ;
        RECT 3298.120 1389.875 3299.300 1391.055 ;
        RECT 3299.720 1389.875 3300.900 1391.055 ;
        RECT 3301.320 1389.875 3302.500 1391.055 ;
        RECT 3302.920 1389.875 3304.100 1391.055 ;
        RECT 3304.520 1389.875 3305.700 1391.055 ;
        RECT 3306.120 1389.875 3307.300 1391.055 ;
        RECT 3307.720 1389.875 3308.900 1391.055 ;
        RECT 3309.320 1389.875 3310.500 1391.055 ;
        RECT 3310.920 1389.875 3312.100 1391.055 ;
        RECT 3312.520 1389.875 3313.700 1391.055 ;
        RECT 3314.120 1389.875 3315.300 1391.055 ;
        RECT 221.285 1379.885 233.665 1385.865 ;
        RECT 3294.825 1385.150 3296.005 1386.330 ;
        RECT 3296.425 1385.150 3297.605 1386.330 ;
        RECT 3298.025 1385.150 3299.205 1386.330 ;
        RECT 3299.625 1385.150 3300.805 1386.330 ;
        RECT 3301.225 1385.150 3302.405 1386.330 ;
        RECT 3302.825 1385.150 3304.005 1386.330 ;
        RECT 3304.425 1385.150 3305.605 1386.330 ;
        RECT 3306.025 1385.150 3307.205 1386.330 ;
        RECT 3307.625 1385.150 3308.805 1386.330 ;
        RECT 3309.225 1385.150 3310.405 1386.330 ;
        RECT 3310.825 1385.150 3312.005 1386.330 ;
        RECT 3312.425 1385.150 3313.605 1386.330 ;
        RECT 3314.025 1385.150 3315.205 1386.330 ;
        RECT 279.080 1380.260 280.260 1381.440 ;
        RECT 280.680 1380.260 281.860 1381.440 ;
        RECT 3354.430 1380.720 3366.810 1386.700 ;
        RECT 3370.430 1384.150 3382.810 1391.730 ;
        RECT 214.505 1347.100 217.285 1377.080 ;
        RECT 279.120 1375.490 280.300 1376.670 ;
        RECT 280.720 1375.490 281.900 1376.670 ;
        RECT 3377.040 1370.240 3382.450 1375.730 ;
        RECT 3358.510 1362.150 3363.920 1367.640 ;
        RECT 3495.950 1354.280 3499.730 1355.690 ;
        RECT 3489.950 1350.760 3493.730 1352.170 ;
        RECT 3489.910 1321.780 3493.770 1323.220 ;
        RECT 89.450 1301.280 93.230 1302.690 ;
        RECT 3489.890 1304.880 3493.750 1306.320 ;
        RECT 89.430 1277.230 93.290 1278.670 ;
        RECT 89.400 1260.320 93.260 1261.760 ;
        RECT 89.410 1243.410 93.270 1244.850 ;
        RECT 95.450 1297.760 99.230 1299.170 ;
        RECT 3495.890 1330.230 3499.750 1331.670 ;
        RECT 3495.920 1313.320 3499.780 1314.760 ;
        RECT 3548.730 1335.500 3552.560 1336.850 ;
        RECT 3548.740 1318.580 3552.570 1319.930 ;
        RECT 3548.730 1301.640 3552.600 1303.130 ;
        RECT 3554.740 1327.020 3558.570 1328.370 ;
        RECT 3554.710 1310.220 3558.540 1311.570 ;
        RECT 3495.910 1296.410 3499.770 1297.850 ;
        RECT 3554.700 1293.200 3558.570 1294.690 ;
        RECT 3489.890 1287.980 3493.750 1289.420 ;
        RECT 95.410 1268.780 99.270 1270.220 ;
        RECT 95.430 1251.880 99.290 1253.320 ;
        RECT 95.430 1234.980 99.290 1236.420 ;
        RECT 3377.040 1144.240 3382.450 1149.730 ;
        RECT 3358.510 1136.150 3363.920 1141.640 ;
        RECT 3495.950 1128.280 3499.730 1129.690 ;
        RECT 3489.950 1124.760 3493.730 1126.170 ;
        RECT 3489.910 1095.780 3493.770 1097.220 ;
        RECT 89.450 1085.280 93.230 1086.690 ;
        RECT 89.430 1061.230 93.290 1062.670 ;
        RECT 89.400 1044.320 93.260 1045.760 ;
        RECT 89.410 1027.410 93.270 1028.850 ;
        RECT 95.450 1081.760 99.230 1083.170 ;
        RECT 3489.890 1078.880 3493.750 1080.320 ;
        RECT 3495.890 1104.230 3499.750 1105.670 ;
        RECT 3495.920 1087.320 3499.780 1088.760 ;
        RECT 3548.730 1109.500 3552.560 1110.850 ;
        RECT 3548.740 1092.580 3552.570 1093.930 ;
        RECT 3548.730 1075.640 3552.600 1077.130 ;
        RECT 3554.740 1101.020 3558.570 1102.370 ;
        RECT 3554.710 1084.220 3558.540 1085.570 ;
        RECT 3495.910 1070.410 3499.770 1071.850 ;
        RECT 3554.700 1067.200 3558.570 1068.690 ;
        RECT 3489.890 1061.980 3493.750 1063.420 ;
        RECT 95.410 1052.780 99.270 1054.220 ;
        RECT 95.430 1035.880 99.290 1037.320 ;
        RECT 95.430 1018.980 99.290 1020.420 ;
        RECT 3377.040 919.240 3382.450 924.730 ;
        RECT 3358.510 911.150 3363.920 916.640 ;
        RECT 3495.950 903.280 3499.730 904.690 ;
        RECT 3489.950 899.760 3493.730 901.170 ;
        RECT 3489.910 870.780 3493.770 872.220 ;
        RECT 3489.890 853.880 3493.750 855.320 ;
        RECT 3495.890 879.230 3499.750 880.670 ;
        RECT 3495.920 862.320 3499.780 863.760 ;
        RECT 3548.730 884.500 3552.560 885.850 ;
        RECT 3548.740 867.580 3552.570 868.930 ;
        RECT 3548.730 850.640 3552.600 852.130 ;
        RECT 3554.740 876.020 3558.570 877.370 ;
        RECT 3554.710 859.220 3558.540 860.570 ;
        RECT 3495.910 845.410 3499.770 846.850 ;
        RECT 3554.700 842.200 3558.570 843.690 ;
        RECT 3489.890 836.980 3493.750 838.420 ;
        RECT 3377.040 693.240 3382.450 698.730 ;
        RECT 3358.510 685.150 3363.920 690.640 ;
        RECT 3495.950 677.280 3499.730 678.690 ;
        RECT 3489.950 673.760 3493.730 675.170 ;
        RECT 3489.910 644.780 3493.770 646.220 ;
        RECT 3489.890 627.880 3493.750 629.320 ;
        RECT 3495.890 653.230 3499.750 654.670 ;
        RECT 3495.920 636.320 3499.780 637.760 ;
        RECT 3548.730 658.500 3552.560 659.850 ;
        RECT 3548.740 641.580 3552.570 642.930 ;
        RECT 3548.730 624.640 3552.600 626.130 ;
        RECT 3554.740 650.020 3558.570 651.370 ;
        RECT 3554.710 633.220 3558.540 634.570 ;
        RECT 3495.910 619.410 3499.770 620.850 ;
        RECT 3554.700 616.200 3558.570 617.690 ;
        RECT 3489.890 610.980 3493.750 612.420 ;
        RECT 643.800 206.700 644.980 207.880 ;
        RECT 645.405 206.700 646.585 207.880 ;
        RECT 716.920 206.700 718.100 207.880 ;
        RECT 651.460 203.310 652.640 204.490 ;
        RECT 653.065 203.310 654.245 204.490 ;
        RECT 723.420 203.310 724.600 204.490 ;
      LAYER met5 ;
        RECT 491.900 5093.460 493.500 5101.470 ;
        RECT 500.350 5099.450 501.950 5101.470 ;
        RECT 500.280 5095.070 502.010 5099.450 ;
        RECT 508.800 5093.470 510.400 5101.470 ;
        RECT 517.250 5099.530 518.850 5101.470 ;
        RECT 517.140 5095.150 518.900 5099.530 ;
        RECT 525.700 5093.480 527.300 5101.470 ;
        RECT 534.150 5099.390 535.750 5101.470 ;
        RECT 534.110 5095.010 535.840 5099.390 ;
        RECT 491.840 5089.080 493.570 5093.460 ;
        RECT 508.740 5089.090 510.470 5093.470 ;
        RECT 525.620 5089.100 527.350 5093.480 ;
        RECT 554.650 5093.350 556.250 5117.040 ;
        RECT 558.150 5099.610 559.750 5117.040 ;
        RECT 558.130 5095.230 559.860 5099.610 ;
        RECT 748.900 5093.460 750.500 5101.470 ;
        RECT 757.350 5099.450 758.950 5101.470 ;
        RECT 757.280 5095.070 759.010 5099.450 ;
        RECT 765.800 5093.470 767.400 5101.470 ;
        RECT 774.250 5099.530 775.850 5101.470 ;
        RECT 774.140 5095.150 775.900 5099.530 ;
        RECT 782.700 5093.480 784.300 5101.470 ;
        RECT 791.150 5099.390 792.750 5101.470 ;
        RECT 791.110 5095.010 792.840 5099.390 ;
        RECT 525.700 5089.090 527.300 5089.100 ;
        RECT 554.620 5088.970 556.350 5093.350 ;
        RECT 748.840 5089.080 750.570 5093.460 ;
        RECT 765.740 5089.090 767.470 5093.470 ;
        RECT 782.620 5089.100 784.350 5093.480 ;
        RECT 811.650 5093.350 813.250 5117.040 ;
        RECT 815.150 5099.610 816.750 5117.040 ;
        RECT 815.130 5095.230 816.860 5099.610 ;
        RECT 1005.900 5093.460 1007.500 5101.470 ;
        RECT 1014.350 5099.450 1015.950 5101.470 ;
        RECT 1014.280 5095.070 1016.010 5099.450 ;
        RECT 1022.800 5093.470 1024.400 5101.470 ;
        RECT 1031.250 5099.530 1032.850 5101.470 ;
        RECT 1031.140 5095.150 1032.900 5099.530 ;
        RECT 1039.700 5093.480 1041.300 5101.470 ;
        RECT 1048.150 5099.390 1049.750 5101.470 ;
        RECT 1048.110 5095.010 1049.840 5099.390 ;
        RECT 782.700 5089.090 784.300 5089.100 ;
        RECT 811.620 5088.970 813.350 5093.350 ;
        RECT 1005.840 5089.080 1007.570 5093.460 ;
        RECT 1022.740 5089.090 1024.470 5093.470 ;
        RECT 1039.620 5089.100 1041.350 5093.480 ;
        RECT 1068.650 5093.350 1070.250 5117.040 ;
        RECT 1072.150 5099.610 1073.750 5117.040 ;
        RECT 1072.130 5095.230 1073.860 5099.610 ;
        RECT 1262.900 5093.460 1264.500 5101.470 ;
        RECT 1271.350 5099.450 1272.950 5101.470 ;
        RECT 1271.280 5095.070 1273.010 5099.450 ;
        RECT 1279.800 5093.470 1281.400 5101.470 ;
        RECT 1288.250 5099.530 1289.850 5101.470 ;
        RECT 1288.140 5095.150 1289.900 5099.530 ;
        RECT 1296.700 5093.480 1298.300 5101.470 ;
        RECT 1305.150 5099.390 1306.750 5101.470 ;
        RECT 1305.110 5095.010 1306.840 5099.390 ;
        RECT 1039.700 5089.090 1041.300 5089.100 ;
        RECT 1068.620 5088.970 1070.350 5093.350 ;
        RECT 1262.840 5089.080 1264.570 5093.460 ;
        RECT 1279.740 5089.090 1281.470 5093.470 ;
        RECT 1296.620 5089.100 1298.350 5093.480 ;
        RECT 1325.650 5093.350 1327.250 5117.040 ;
        RECT 1329.150 5099.610 1330.750 5117.040 ;
        RECT 1329.130 5095.230 1330.860 5099.610 ;
        RECT 1520.900 5093.460 1522.500 5101.470 ;
        RECT 1529.350 5099.450 1530.950 5101.470 ;
        RECT 1529.280 5095.070 1531.010 5099.450 ;
        RECT 1537.800 5093.470 1539.400 5101.470 ;
        RECT 1546.250 5099.530 1547.850 5101.470 ;
        RECT 1546.140 5095.150 1547.900 5099.530 ;
        RECT 1554.700 5093.480 1556.300 5101.470 ;
        RECT 1563.150 5099.390 1564.750 5101.470 ;
        RECT 1563.110 5095.010 1564.840 5099.390 ;
        RECT 1296.700 5089.090 1298.300 5089.100 ;
        RECT 1325.620 5088.970 1327.350 5093.350 ;
        RECT 1520.840 5089.080 1522.570 5093.460 ;
        RECT 1537.740 5089.090 1539.470 5093.470 ;
        RECT 1554.620 5089.100 1556.350 5093.480 ;
        RECT 1583.650 5093.350 1585.250 5117.040 ;
        RECT 1587.150 5099.610 1588.750 5117.040 ;
        RECT 1587.130 5095.230 1588.860 5099.610 ;
        RECT 1772.900 5093.460 1774.500 5101.470 ;
        RECT 1781.350 5099.450 1782.950 5101.470 ;
        RECT 1781.280 5095.070 1783.010 5099.450 ;
        RECT 1789.800 5093.470 1791.400 5101.470 ;
        RECT 1798.250 5099.530 1799.850 5101.470 ;
        RECT 1798.140 5095.150 1799.900 5099.530 ;
        RECT 1806.700 5093.480 1808.300 5101.470 ;
        RECT 1815.150 5099.390 1816.750 5101.470 ;
        RECT 1815.110 5095.010 1816.840 5099.390 ;
        RECT 1554.700 5089.090 1556.300 5089.100 ;
        RECT 1583.620 5088.970 1585.350 5093.350 ;
        RECT 1772.840 5089.080 1774.570 5093.460 ;
        RECT 1789.740 5089.090 1791.470 5093.470 ;
        RECT 1806.620 5089.100 1808.350 5093.480 ;
        RECT 1835.650 5093.350 1837.250 5117.040 ;
        RECT 1839.150 5099.610 1840.750 5117.040 ;
        RECT 1839.130 5095.230 1840.860 5099.610 ;
        RECT 2109.900 5093.460 2111.500 5101.470 ;
        RECT 2118.350 5099.450 2119.950 5101.470 ;
        RECT 2118.280 5095.070 2120.010 5099.450 ;
        RECT 2126.800 5093.470 2128.400 5101.470 ;
        RECT 2135.250 5099.530 2136.850 5101.470 ;
        RECT 2135.140 5095.150 2136.900 5099.530 ;
        RECT 2143.700 5093.480 2145.300 5101.470 ;
        RECT 2152.150 5099.390 2153.750 5101.470 ;
        RECT 2152.110 5095.010 2153.840 5099.390 ;
        RECT 1806.700 5089.090 1808.300 5089.100 ;
        RECT 1835.620 5088.970 1837.350 5093.350 ;
        RECT 2109.840 5089.080 2111.570 5093.460 ;
        RECT 2126.740 5089.090 2128.470 5093.470 ;
        RECT 2143.620 5089.100 2145.350 5093.480 ;
        RECT 2172.650 5093.350 2174.250 5117.040 ;
        RECT 2176.150 5099.610 2177.750 5117.040 ;
        RECT 2176.130 5095.230 2177.860 5099.610 ;
        RECT 2494.900 5093.460 2496.500 5101.470 ;
        RECT 2503.350 5099.450 2504.950 5101.470 ;
        RECT 2503.280 5095.070 2505.010 5099.450 ;
        RECT 2511.800 5093.470 2513.400 5101.470 ;
        RECT 2520.250 5099.530 2521.850 5101.470 ;
        RECT 2520.140 5095.150 2521.900 5099.530 ;
        RECT 2528.700 5093.480 2530.300 5101.470 ;
        RECT 2537.150 5099.390 2538.750 5101.470 ;
        RECT 2537.110 5095.010 2538.840 5099.390 ;
        RECT 2143.700 5089.090 2145.300 5089.100 ;
        RECT 2172.620 5088.970 2174.350 5093.350 ;
        RECT 2494.840 5089.080 2496.570 5093.460 ;
        RECT 2511.740 5089.090 2513.470 5093.470 ;
        RECT 2528.620 5089.100 2530.350 5093.480 ;
        RECT 2557.650 5093.350 2559.250 5117.040 ;
        RECT 2561.150 5099.610 2562.750 5117.040 ;
        RECT 2561.130 5095.230 2562.860 5099.610 ;
        RECT 2751.900 5093.460 2753.500 5101.470 ;
        RECT 2760.350 5099.450 2761.950 5101.470 ;
        RECT 2760.280 5095.070 2762.010 5099.450 ;
        RECT 2768.800 5093.470 2770.400 5101.470 ;
        RECT 2777.250 5099.530 2778.850 5101.470 ;
        RECT 2777.140 5095.150 2778.900 5099.530 ;
        RECT 2785.700 5093.480 2787.300 5101.470 ;
        RECT 2794.150 5099.390 2795.750 5101.470 ;
        RECT 2794.110 5095.010 2795.840 5099.390 ;
        RECT 2528.700 5089.090 2530.300 5089.100 ;
        RECT 2557.620 5088.970 2559.350 5093.350 ;
        RECT 2751.840 5089.080 2753.570 5093.460 ;
        RECT 2768.740 5089.090 2770.470 5093.470 ;
        RECT 2785.620 5089.100 2787.350 5093.480 ;
        RECT 2814.650 5093.350 2816.250 5117.040 ;
        RECT 2818.150 5099.610 2819.750 5117.040 ;
        RECT 2818.130 5095.230 2819.860 5099.610 ;
        RECT 2785.700 5089.090 2787.300 5089.100 ;
        RECT 2814.620 5088.970 2816.350 5093.350 ;
        RECT 205.170 4929.390 217.870 4932.240 ;
        RECT 278.880 4929.240 302.180 4932.340 ;
        RECT 221.210 4924.590 233.860 4927.490 ;
        RECT 278.880 4924.440 306.990 4927.540 ;
        RECT 3260.900 4919.640 3315.890 4922.740 ;
        RECT 3354.290 4919.750 3366.920 4922.680 ;
        RECT 3256.140 4914.840 3315.890 4917.940 ;
        RECT 3370.280 4914.940 3382.910 4917.870 ;
        RECT 221.390 4759.880 233.670 4765.150 ;
        RECT 205.340 4751.970 217.620 4757.240 ;
        RECT 89.230 4729.780 93.425 4729.895 ;
        RECT 71.550 4728.180 93.425 4729.780 ;
        RECT 89.230 4728.090 93.425 4728.180 ;
        RECT 95.260 4726.280 99.455 4726.350 ;
        RECT 71.550 4724.680 99.610 4726.280 ;
        RECT 3376.990 4726.240 3382.400 4731.730 ;
        RECT 95.260 4724.545 99.455 4724.680 ;
        RECT 3358.460 4718.150 3363.870 4723.640 ;
        RECT 3495.740 4711.780 3499.870 4711.840 ;
        RECT 3495.740 4710.180 3517.580 4711.780 ;
        RECT 3495.740 4710.125 3499.870 4710.180 ;
        RECT 3489.685 4708.280 3493.815 4708.355 ;
        RECT 3489.520 4706.680 3517.580 4708.280 ;
        RECT 3489.685 4706.640 3493.815 4706.680 ;
        RECT 89.245 4705.750 93.455 4705.840 ;
        RECT 87.120 4704.150 93.540 4705.750 ;
        RECT 89.245 4704.040 93.455 4704.150 ;
        RECT 95.280 4697.300 99.490 4697.365 ;
        RECT 87.120 4695.700 99.500 4697.300 ;
        RECT 95.280 4695.620 99.490 4695.700 ;
        RECT 3548.530 4692.990 3552.715 4693.075 ;
        RECT 3546.220 4691.390 3552.830 4692.990 ;
        RECT 3548.530 4691.300 3552.715 4691.390 ;
        RECT 89.285 4688.850 93.495 4688.890 ;
        RECT 87.120 4687.250 93.495 4688.850 ;
        RECT 89.285 4687.145 93.495 4687.250 ;
        RECT 3495.580 4687.750 3499.905 4687.850 ;
        RECT 3495.580 4686.150 3502.010 4687.750 ;
        RECT 3495.580 4686.080 3499.905 4686.150 ;
        RECT 3554.535 4684.540 3558.720 4684.620 ;
        RECT 3546.220 4682.940 3558.890 4684.540 ;
        RECT 3554.535 4682.845 3558.720 4682.940 ;
        RECT 95.265 4680.400 99.475 4680.475 ;
        RECT 87.120 4678.800 99.500 4680.400 ;
        RECT 3489.595 4679.300 3493.920 4679.360 ;
        RECT 95.265 4678.730 99.475 4678.800 ;
        RECT 3489.595 4677.700 3502.010 4679.300 ;
        RECT 3489.595 4677.590 3493.920 4677.700 ;
        RECT 3548.505 4676.090 3552.690 4676.205 ;
        RECT 3546.220 4674.490 3552.800 4676.090 ;
        RECT 3548.505 4674.430 3552.690 4674.490 ;
        RECT 89.265 4671.950 93.475 4672.025 ;
        RECT 87.120 4670.350 93.510 4671.950 ;
        RECT 3495.695 4670.850 3500.020 4670.935 ;
        RECT 89.265 4670.280 93.475 4670.350 ;
        RECT 3495.695 4669.250 3502.010 4670.850 ;
        RECT 3495.695 4669.165 3500.020 4669.250 ;
        RECT 3554.480 4667.640 3558.890 4667.750 ;
        RECT 3546.220 4666.140 3558.890 4667.640 ;
        RECT 3546.220 4666.060 3558.885 4666.140 ;
        RECT 3546.220 4666.040 3558.880 4666.060 ;
        RECT 95.310 4663.500 99.520 4663.575 ;
        RECT 87.120 4661.900 99.520 4663.500 ;
        RECT 95.310 4661.830 99.520 4661.900 ;
        RECT 3489.600 4662.400 3493.925 4662.460 ;
        RECT 3489.600 4660.800 3502.010 4662.400 ;
        RECT 3489.600 4660.690 3493.925 4660.800 ;
        RECT 3548.510 4659.190 3552.690 4659.280 ;
        RECT 3546.060 4657.590 3552.690 4659.190 ;
        RECT 3548.510 4657.480 3552.690 4657.590 ;
        RECT 3495.600 4653.950 3499.925 4654.055 ;
        RECT 3495.600 4652.350 3502.010 4653.950 ;
        RECT 3495.600 4652.285 3499.925 4652.350 ;
        RECT 3554.475 4650.740 3558.660 4650.820 ;
        RECT 3546.060 4649.140 3558.660 4650.740 ;
        RECT 3554.475 4649.045 3558.660 4649.140 ;
        RECT 3489.630 4645.500 3493.955 4645.600 ;
        RECT 3489.630 4643.900 3502.010 4645.500 ;
        RECT 3489.630 4643.830 3493.955 4643.900 ;
        RECT 3373.670 4500.370 3378.700 4505.560 ;
        RECT 3357.830 4492.330 3362.980 4497.520 ;
        RECT 3370.580 4275.260 3375.900 4280.580 ;
        RECT 3357.850 4267.210 3363.190 4272.610 ;
        RECT 221.390 4130.880 233.670 4136.150 ;
        RECT 205.340 4122.970 217.620 4128.240 ;
        RECT 89.230 4100.780 93.425 4100.895 ;
        RECT 71.550 4099.180 93.425 4100.780 ;
        RECT 89.230 4099.090 93.425 4099.180 ;
        RECT 95.260 4097.280 99.455 4097.350 ;
        RECT 71.550 4095.680 99.610 4097.280 ;
        RECT 95.260 4095.545 99.455 4095.680 ;
        RECT 89.245 4076.750 93.455 4076.840 ;
        RECT 87.120 4075.150 93.540 4076.750 ;
        RECT 89.245 4075.040 93.455 4075.150 ;
        RECT 95.280 4068.300 99.490 4068.365 ;
        RECT 87.120 4066.700 99.500 4068.300 ;
        RECT 95.280 4066.620 99.490 4066.700 ;
        RECT 89.285 4059.850 93.495 4059.890 ;
        RECT 87.120 4058.250 93.495 4059.850 ;
        RECT 89.285 4058.145 93.495 4058.250 ;
        RECT 95.265 4051.400 99.475 4051.475 ;
        RECT 87.120 4049.800 99.500 4051.400 ;
        RECT 95.265 4049.730 99.475 4049.800 ;
        RECT 89.265 4042.950 93.475 4043.025 ;
        RECT 87.120 4041.350 93.510 4042.950 ;
        RECT 89.265 4041.280 93.475 4041.350 ;
        RECT 95.310 4034.500 99.520 4034.575 ;
        RECT 87.120 4032.900 99.520 4034.500 ;
        RECT 95.310 4032.830 99.520 4032.900 ;
        RECT 221.390 3922.880 233.670 3928.150 ;
        RECT 205.340 3914.970 217.620 3920.240 ;
        RECT 89.230 3884.780 93.425 3884.895 ;
        RECT 71.550 3883.180 93.425 3884.780 ;
        RECT 89.230 3883.090 93.425 3883.180 ;
        RECT 95.260 3881.280 99.455 3881.350 ;
        RECT 71.550 3879.680 99.610 3881.280 ;
        RECT 95.260 3879.545 99.455 3879.680 ;
        RECT 89.245 3860.750 93.455 3860.840 ;
        RECT 87.120 3859.150 93.540 3860.750 ;
        RECT 89.245 3859.040 93.455 3859.150 ;
        RECT 95.280 3852.300 99.490 3852.365 ;
        RECT 87.120 3850.700 99.500 3852.300 ;
        RECT 95.280 3850.620 99.490 3850.700 ;
        RECT 89.285 3843.850 93.495 3843.890 ;
        RECT 87.120 3842.250 93.495 3843.850 ;
        RECT 89.285 3842.145 93.495 3842.250 ;
        RECT 95.265 3835.400 99.475 3835.475 ;
        RECT 87.120 3833.800 99.500 3835.400 ;
        RECT 3377.040 3834.240 3382.450 3839.730 ;
        RECT 95.265 3833.730 99.475 3833.800 ;
        RECT 89.265 3826.950 93.475 3827.025 ;
        RECT 87.120 3825.350 93.510 3826.950 ;
        RECT 3358.510 3826.150 3363.920 3831.640 ;
        RECT 89.265 3825.280 93.475 3825.350 ;
        RECT 3495.790 3819.780 3499.920 3819.840 ;
        RECT 95.310 3818.500 99.520 3818.575 ;
        RECT 87.120 3816.900 99.520 3818.500 ;
        RECT 3495.790 3818.180 3517.630 3819.780 ;
        RECT 3495.790 3818.125 3499.920 3818.180 ;
        RECT 95.310 3816.830 99.520 3816.900 ;
        RECT 3489.735 3816.280 3493.865 3816.355 ;
        RECT 3489.570 3814.680 3517.630 3816.280 ;
        RECT 3489.735 3814.640 3493.865 3814.680 ;
        RECT 3548.580 3800.990 3552.765 3801.075 ;
        RECT 3546.270 3799.390 3552.880 3800.990 ;
        RECT 3548.580 3799.300 3552.765 3799.390 ;
        RECT 3495.630 3795.750 3499.955 3795.850 ;
        RECT 3495.630 3794.150 3502.060 3795.750 ;
        RECT 3495.630 3794.080 3499.955 3794.150 ;
        RECT 3554.585 3792.540 3558.770 3792.620 ;
        RECT 3546.270 3790.940 3558.940 3792.540 ;
        RECT 3554.585 3790.845 3558.770 3790.940 ;
        RECT 3489.645 3787.300 3493.970 3787.360 ;
        RECT 3489.645 3785.700 3502.060 3787.300 ;
        RECT 3489.645 3785.590 3493.970 3785.700 ;
        RECT 3548.555 3784.090 3552.740 3784.205 ;
        RECT 3546.270 3782.490 3552.850 3784.090 ;
        RECT 3548.555 3782.430 3552.740 3782.490 ;
        RECT 3495.745 3778.850 3500.070 3778.935 ;
        RECT 3495.745 3777.250 3502.060 3778.850 ;
        RECT 3495.745 3777.165 3500.070 3777.250 ;
        RECT 3554.530 3775.640 3558.940 3775.750 ;
        RECT 3546.270 3774.140 3558.940 3775.640 ;
        RECT 3546.270 3774.060 3558.935 3774.140 ;
        RECT 3546.270 3774.040 3558.930 3774.060 ;
        RECT 3489.650 3770.400 3493.975 3770.460 ;
        RECT 3489.650 3768.800 3502.060 3770.400 ;
        RECT 3489.650 3768.690 3493.975 3768.800 ;
        RECT 3548.560 3767.190 3552.740 3767.280 ;
        RECT 3546.110 3765.590 3552.740 3767.190 ;
        RECT 3548.560 3765.480 3552.740 3765.590 ;
        RECT 3495.650 3761.950 3499.975 3762.055 ;
        RECT 3495.650 3760.350 3502.060 3761.950 ;
        RECT 3495.650 3760.285 3499.975 3760.350 ;
        RECT 3554.525 3758.740 3558.710 3758.820 ;
        RECT 3546.110 3757.140 3558.710 3758.740 ;
        RECT 3554.525 3757.045 3558.710 3757.140 ;
        RECT 3489.680 3753.500 3494.005 3753.600 ;
        RECT 3489.680 3751.900 3502.060 3753.500 ;
        RECT 3489.680 3751.830 3494.005 3751.900 ;
        RECT 221.390 3698.880 233.670 3704.150 ;
        RECT 205.340 3690.970 217.620 3696.240 ;
        RECT 89.230 3668.780 93.425 3668.895 ;
        RECT 71.550 3667.180 93.425 3668.780 ;
        RECT 89.230 3667.090 93.425 3667.180 ;
        RECT 95.260 3665.280 99.455 3665.350 ;
        RECT 71.550 3663.680 99.610 3665.280 ;
        RECT 95.260 3663.545 99.455 3663.680 ;
        RECT 89.245 3644.750 93.455 3644.840 ;
        RECT 87.120 3643.150 93.540 3644.750 ;
        RECT 89.245 3643.040 93.455 3643.150 ;
        RECT 95.280 3636.300 99.490 3636.365 ;
        RECT 87.120 3634.700 99.500 3636.300 ;
        RECT 95.280 3634.620 99.490 3634.700 ;
        RECT 89.285 3627.850 93.495 3627.890 ;
        RECT 87.120 3626.250 93.495 3627.850 ;
        RECT 89.285 3626.145 93.495 3626.250 ;
        RECT 95.265 3619.400 99.475 3619.475 ;
        RECT 87.120 3617.800 99.500 3619.400 ;
        RECT 95.265 3617.730 99.475 3617.800 ;
        RECT 89.265 3610.950 93.475 3611.025 ;
        RECT 87.120 3609.350 93.510 3610.950 ;
        RECT 89.265 3609.280 93.475 3609.350 ;
        RECT 3377.040 3609.240 3382.450 3614.730 ;
        RECT 95.310 3602.500 99.520 3602.575 ;
        RECT 87.120 3600.900 99.520 3602.500 ;
        RECT 3358.510 3601.150 3363.920 3606.640 ;
        RECT 95.310 3600.830 99.520 3600.900 ;
        RECT 3495.790 3594.780 3499.920 3594.840 ;
        RECT 3495.790 3593.180 3517.630 3594.780 ;
        RECT 3495.790 3593.125 3499.920 3593.180 ;
        RECT 3489.735 3591.280 3493.865 3591.355 ;
        RECT 3489.570 3589.680 3517.630 3591.280 ;
        RECT 3489.735 3589.640 3493.865 3589.680 ;
        RECT 3548.580 3575.990 3552.765 3576.075 ;
        RECT 3546.270 3574.390 3552.880 3575.990 ;
        RECT 3548.580 3574.300 3552.765 3574.390 ;
        RECT 3495.630 3570.750 3499.955 3570.850 ;
        RECT 3495.630 3569.150 3502.060 3570.750 ;
        RECT 3495.630 3569.080 3499.955 3569.150 ;
        RECT 3554.585 3567.540 3558.770 3567.620 ;
        RECT 3546.270 3565.940 3558.940 3567.540 ;
        RECT 3554.585 3565.845 3558.770 3565.940 ;
        RECT 3489.645 3562.300 3493.970 3562.360 ;
        RECT 3489.645 3560.700 3502.060 3562.300 ;
        RECT 3489.645 3560.590 3493.970 3560.700 ;
        RECT 3548.555 3559.090 3552.740 3559.205 ;
        RECT 3546.270 3557.490 3552.850 3559.090 ;
        RECT 3548.555 3557.430 3552.740 3557.490 ;
        RECT 3495.745 3553.850 3500.070 3553.935 ;
        RECT 3495.745 3552.250 3502.060 3553.850 ;
        RECT 3495.745 3552.165 3500.070 3552.250 ;
        RECT 3554.530 3550.640 3558.940 3550.750 ;
        RECT 3546.270 3549.140 3558.940 3550.640 ;
        RECT 3546.270 3549.060 3558.935 3549.140 ;
        RECT 3546.270 3549.040 3558.930 3549.060 ;
        RECT 3489.650 3545.400 3493.975 3545.460 ;
        RECT 3489.650 3543.800 3502.060 3545.400 ;
        RECT 3489.650 3543.690 3493.975 3543.800 ;
        RECT 3548.560 3542.190 3552.740 3542.280 ;
        RECT 3546.110 3540.590 3552.740 3542.190 ;
        RECT 3548.560 3540.480 3552.740 3540.590 ;
        RECT 3495.650 3536.950 3499.975 3537.055 ;
        RECT 3495.650 3535.350 3502.060 3536.950 ;
        RECT 3495.650 3535.285 3499.975 3535.350 ;
        RECT 3554.525 3533.740 3558.710 3533.820 ;
        RECT 3546.110 3532.140 3558.710 3533.740 ;
        RECT 3554.525 3532.045 3558.710 3532.140 ;
        RECT 3489.680 3528.500 3494.005 3528.600 ;
        RECT 3489.680 3526.900 3502.060 3528.500 ;
        RECT 3489.680 3526.830 3494.005 3526.900 ;
        RECT 221.390 3482.880 233.670 3488.150 ;
        RECT 205.340 3474.970 217.620 3480.240 ;
        RECT 89.230 3452.780 93.425 3452.895 ;
        RECT 71.550 3451.180 93.425 3452.780 ;
        RECT 89.230 3451.090 93.425 3451.180 ;
        RECT 95.260 3449.280 99.455 3449.350 ;
        RECT 71.550 3447.680 99.610 3449.280 ;
        RECT 95.260 3447.545 99.455 3447.680 ;
        RECT 89.245 3428.750 93.455 3428.840 ;
        RECT 87.120 3427.150 93.540 3428.750 ;
        RECT 89.245 3427.040 93.455 3427.150 ;
        RECT 95.280 3420.300 99.490 3420.365 ;
        RECT 87.120 3418.700 99.500 3420.300 ;
        RECT 95.280 3418.620 99.490 3418.700 ;
        RECT 89.285 3411.850 93.495 3411.890 ;
        RECT 87.120 3410.250 93.495 3411.850 ;
        RECT 89.285 3410.145 93.495 3410.250 ;
        RECT 95.265 3403.400 99.475 3403.475 ;
        RECT 87.120 3401.800 99.500 3403.400 ;
        RECT 95.265 3401.730 99.475 3401.800 ;
        RECT 89.265 3394.950 93.475 3395.025 ;
        RECT 87.120 3393.350 93.510 3394.950 ;
        RECT 89.265 3393.280 93.475 3393.350 ;
        RECT 95.310 3386.500 99.520 3386.575 ;
        RECT 87.120 3384.900 99.520 3386.500 ;
        RECT 95.310 3384.830 99.520 3384.900 ;
        RECT 3377.040 3383.240 3382.450 3388.730 ;
        RECT 3358.510 3375.150 3363.920 3380.640 ;
        RECT 3495.790 3368.780 3499.920 3368.840 ;
        RECT 3495.790 3367.180 3517.630 3368.780 ;
        RECT 3495.790 3367.125 3499.920 3367.180 ;
        RECT 3489.735 3365.280 3493.865 3365.355 ;
        RECT 3489.570 3363.680 3517.630 3365.280 ;
        RECT 3489.735 3363.640 3493.865 3363.680 ;
        RECT 3548.580 3349.990 3552.765 3350.075 ;
        RECT 3546.270 3348.390 3552.880 3349.990 ;
        RECT 3548.580 3348.300 3552.765 3348.390 ;
        RECT 3495.630 3344.750 3499.955 3344.850 ;
        RECT 3495.630 3343.150 3502.060 3344.750 ;
        RECT 3495.630 3343.080 3499.955 3343.150 ;
        RECT 3554.585 3341.540 3558.770 3341.620 ;
        RECT 3546.270 3339.940 3558.940 3341.540 ;
        RECT 3554.585 3339.845 3558.770 3339.940 ;
        RECT 3489.645 3336.300 3493.970 3336.360 ;
        RECT 3489.645 3334.700 3502.060 3336.300 ;
        RECT 3489.645 3334.590 3493.970 3334.700 ;
        RECT 3548.555 3333.090 3552.740 3333.205 ;
        RECT 3546.270 3331.490 3552.850 3333.090 ;
        RECT 3548.555 3331.430 3552.740 3331.490 ;
        RECT 3495.745 3327.850 3500.070 3327.935 ;
        RECT 3495.745 3326.250 3502.060 3327.850 ;
        RECT 3495.745 3326.165 3500.070 3326.250 ;
        RECT 3554.530 3324.640 3558.940 3324.750 ;
        RECT 3546.270 3323.140 3558.940 3324.640 ;
        RECT 3546.270 3323.060 3558.935 3323.140 ;
        RECT 3546.270 3323.040 3558.930 3323.060 ;
        RECT 3489.650 3319.400 3493.975 3319.460 ;
        RECT 3489.650 3317.800 3502.060 3319.400 ;
        RECT 3489.650 3317.690 3493.975 3317.800 ;
        RECT 3548.560 3316.190 3552.740 3316.280 ;
        RECT 3546.110 3314.590 3552.740 3316.190 ;
        RECT 3548.560 3314.480 3552.740 3314.590 ;
        RECT 3495.650 3310.950 3499.975 3311.055 ;
        RECT 3495.650 3309.350 3502.060 3310.950 ;
        RECT 3495.650 3309.285 3499.975 3309.350 ;
        RECT 3554.525 3307.740 3558.710 3307.820 ;
        RECT 3546.110 3306.140 3558.710 3307.740 ;
        RECT 3554.525 3306.045 3558.710 3306.140 ;
        RECT 3489.680 3302.500 3494.005 3302.600 ;
        RECT 3489.680 3300.900 3502.060 3302.500 ;
        RECT 3489.680 3300.830 3494.005 3300.900 ;
        RECT 221.390 3266.880 233.670 3272.150 ;
        RECT 205.340 3258.970 217.620 3264.240 ;
        RECT 89.230 3236.780 93.425 3236.895 ;
        RECT 71.550 3235.180 93.425 3236.780 ;
        RECT 89.230 3235.090 93.425 3235.180 ;
        RECT 95.260 3233.280 99.455 3233.350 ;
        RECT 71.550 3231.680 99.610 3233.280 ;
        RECT 95.260 3231.545 99.455 3231.680 ;
        RECT 89.245 3212.750 93.455 3212.840 ;
        RECT 87.120 3211.150 93.540 3212.750 ;
        RECT 89.245 3211.040 93.455 3211.150 ;
        RECT 95.280 3204.300 99.490 3204.365 ;
        RECT 87.120 3202.700 99.500 3204.300 ;
        RECT 95.280 3202.620 99.490 3202.700 ;
        RECT 89.285 3195.850 93.495 3195.890 ;
        RECT 87.120 3194.250 93.495 3195.850 ;
        RECT 89.285 3194.145 93.495 3194.250 ;
        RECT 95.265 3187.400 99.475 3187.475 ;
        RECT 87.120 3185.800 99.500 3187.400 ;
        RECT 95.265 3185.730 99.475 3185.800 ;
        RECT 89.265 3178.950 93.475 3179.025 ;
        RECT 87.120 3177.350 93.510 3178.950 ;
        RECT 89.265 3177.280 93.475 3177.350 ;
        RECT 95.310 3170.500 99.520 3170.575 ;
        RECT 87.120 3168.900 99.520 3170.500 ;
        RECT 95.310 3168.830 99.520 3168.900 ;
        RECT 3377.040 3158.240 3382.450 3163.730 ;
        RECT 3358.510 3150.150 3363.920 3155.640 ;
        RECT 3495.790 3143.780 3499.920 3143.840 ;
        RECT 3495.790 3142.180 3517.630 3143.780 ;
        RECT 3495.790 3142.125 3499.920 3142.180 ;
        RECT 3489.735 3140.280 3493.865 3140.355 ;
        RECT 3489.570 3138.680 3517.630 3140.280 ;
        RECT 3489.735 3138.640 3493.865 3138.680 ;
        RECT 3548.580 3124.990 3552.765 3125.075 ;
        RECT 3546.270 3123.390 3552.880 3124.990 ;
        RECT 3548.580 3123.300 3552.765 3123.390 ;
        RECT 3495.630 3119.750 3499.955 3119.850 ;
        RECT 3495.630 3118.150 3502.060 3119.750 ;
        RECT 3495.630 3118.080 3499.955 3118.150 ;
        RECT 3554.585 3116.540 3558.770 3116.620 ;
        RECT 3546.270 3114.940 3558.940 3116.540 ;
        RECT 3554.585 3114.845 3558.770 3114.940 ;
        RECT 3489.645 3111.300 3493.970 3111.360 ;
        RECT 3489.645 3109.700 3502.060 3111.300 ;
        RECT 3489.645 3109.590 3493.970 3109.700 ;
        RECT 3548.555 3108.090 3552.740 3108.205 ;
        RECT 3546.270 3106.490 3552.850 3108.090 ;
        RECT 3548.555 3106.430 3552.740 3106.490 ;
        RECT 3495.745 3102.850 3500.070 3102.935 ;
        RECT 3495.745 3101.250 3502.060 3102.850 ;
        RECT 3495.745 3101.165 3500.070 3101.250 ;
        RECT 3554.530 3099.640 3558.940 3099.750 ;
        RECT 3546.270 3098.140 3558.940 3099.640 ;
        RECT 3546.270 3098.060 3558.935 3098.140 ;
        RECT 3546.270 3098.040 3558.930 3098.060 ;
        RECT 3489.650 3094.400 3493.975 3094.460 ;
        RECT 3489.650 3092.800 3502.060 3094.400 ;
        RECT 3489.650 3092.690 3493.975 3092.800 ;
        RECT 3548.560 3091.190 3552.740 3091.280 ;
        RECT 3546.110 3089.590 3552.740 3091.190 ;
        RECT 3548.560 3089.480 3552.740 3089.590 ;
        RECT 3495.650 3085.950 3499.975 3086.055 ;
        RECT 3495.650 3084.350 3502.060 3085.950 ;
        RECT 3495.650 3084.285 3499.975 3084.350 ;
        RECT 3554.525 3082.740 3558.710 3082.820 ;
        RECT 3546.110 3081.140 3558.710 3082.740 ;
        RECT 3554.525 3081.045 3558.710 3081.140 ;
        RECT 3489.680 3077.500 3494.005 3077.600 ;
        RECT 3489.680 3075.900 3502.060 3077.500 ;
        RECT 3489.680 3075.830 3494.005 3075.900 ;
        RECT 221.390 3056.180 233.670 3061.450 ;
        RECT 205.340 3048.270 217.620 3053.540 ;
        RECT 89.230 3020.780 93.425 3020.895 ;
        RECT 71.550 3019.180 93.425 3020.780 ;
        RECT 89.230 3019.090 93.425 3019.180 ;
        RECT 95.260 3017.280 99.455 3017.350 ;
        RECT 71.550 3015.680 99.610 3017.280 ;
        RECT 95.260 3015.545 99.455 3015.680 ;
        RECT 89.245 2996.750 93.455 2996.840 ;
        RECT 87.120 2995.150 93.540 2996.750 ;
        RECT 89.245 2995.040 93.455 2995.150 ;
        RECT 95.280 2988.300 99.490 2988.365 ;
        RECT 87.120 2986.700 99.500 2988.300 ;
        RECT 95.280 2986.620 99.490 2986.700 ;
        RECT 89.285 2979.850 93.495 2979.890 ;
        RECT 87.120 2978.250 93.495 2979.850 ;
        RECT 89.285 2978.145 93.495 2978.250 ;
        RECT 95.265 2971.400 99.475 2971.475 ;
        RECT 87.120 2969.800 99.500 2971.400 ;
        RECT 95.265 2969.730 99.475 2969.800 ;
        RECT 89.265 2962.950 93.475 2963.025 ;
        RECT 87.120 2961.350 93.510 2962.950 ;
        RECT 89.265 2961.280 93.475 2961.350 ;
        RECT 95.310 2954.500 99.520 2954.575 ;
        RECT 87.120 2952.900 99.520 2954.500 ;
        RECT 95.310 2952.830 99.520 2952.900 ;
        RECT 3377.040 2932.240 3382.450 2937.730 ;
        RECT 3358.510 2924.150 3363.920 2929.640 ;
        RECT 3495.790 2917.780 3499.920 2917.840 ;
        RECT 3495.790 2916.180 3517.630 2917.780 ;
        RECT 3495.790 2916.125 3499.920 2916.180 ;
        RECT 3489.735 2914.280 3493.865 2914.355 ;
        RECT 3489.570 2912.680 3517.630 2914.280 ;
        RECT 3489.735 2912.640 3493.865 2912.680 ;
        RECT 3548.580 2898.990 3552.765 2899.075 ;
        RECT 3546.270 2897.390 3552.880 2898.990 ;
        RECT 3548.580 2897.300 3552.765 2897.390 ;
        RECT 3495.630 2893.750 3499.955 2893.850 ;
        RECT 3495.630 2892.150 3502.060 2893.750 ;
        RECT 3495.630 2892.080 3499.955 2892.150 ;
        RECT 3554.585 2890.540 3558.770 2890.620 ;
        RECT 3546.270 2888.940 3558.940 2890.540 ;
        RECT 3554.585 2888.845 3558.770 2888.940 ;
        RECT 3489.645 2885.300 3493.970 2885.360 ;
        RECT 3489.645 2883.700 3502.060 2885.300 ;
        RECT 3489.645 2883.590 3493.970 2883.700 ;
        RECT 3548.555 2882.090 3552.740 2882.205 ;
        RECT 3546.270 2880.490 3552.850 2882.090 ;
        RECT 3548.555 2880.430 3552.740 2880.490 ;
        RECT 3495.745 2876.850 3500.070 2876.935 ;
        RECT 3495.745 2875.250 3502.060 2876.850 ;
        RECT 3495.745 2875.165 3500.070 2875.250 ;
        RECT 3554.530 2873.640 3558.940 2873.750 ;
        RECT 3546.270 2872.140 3558.940 2873.640 ;
        RECT 3546.270 2872.060 3558.935 2872.140 ;
        RECT 3546.270 2872.040 3558.930 2872.060 ;
        RECT 3489.650 2868.400 3493.975 2868.460 ;
        RECT 3489.650 2866.800 3502.060 2868.400 ;
        RECT 3489.650 2866.690 3493.975 2866.800 ;
        RECT 3548.560 2865.190 3552.740 2865.280 ;
        RECT 3546.110 2863.590 3552.740 2865.190 ;
        RECT 3548.560 2863.480 3552.740 2863.590 ;
        RECT 3495.650 2859.950 3499.975 2860.055 ;
        RECT 3495.650 2858.350 3502.060 2859.950 ;
        RECT 3495.650 2858.285 3499.975 2858.350 ;
        RECT 3554.525 2856.740 3558.710 2856.820 ;
        RECT 3546.110 2855.140 3558.710 2856.740 ;
        RECT 3554.525 2855.045 3558.710 2855.140 ;
        RECT 3489.680 2851.500 3494.005 2851.600 ;
        RECT 3489.680 2849.900 3502.060 2851.500 ;
        RECT 3489.680 2849.830 3494.005 2849.900 ;
        RECT 221.390 2834.880 233.670 2840.150 ;
        RECT 205.340 2826.970 217.620 2832.240 ;
        RECT 89.230 2804.780 93.425 2804.895 ;
        RECT 71.550 2803.180 93.425 2804.780 ;
        RECT 89.230 2803.090 93.425 2803.180 ;
        RECT 95.260 2801.280 99.455 2801.350 ;
        RECT 71.550 2799.680 99.610 2801.280 ;
        RECT 95.260 2799.545 99.455 2799.680 ;
        RECT 89.245 2780.750 93.455 2780.840 ;
        RECT 87.120 2779.150 93.540 2780.750 ;
        RECT 89.245 2779.040 93.455 2779.150 ;
        RECT 95.280 2772.300 99.490 2772.365 ;
        RECT 87.120 2770.700 99.500 2772.300 ;
        RECT 95.280 2770.620 99.490 2770.700 ;
        RECT 89.285 2763.850 93.495 2763.890 ;
        RECT 87.120 2762.250 93.495 2763.850 ;
        RECT 89.285 2762.145 93.495 2762.250 ;
        RECT 95.265 2755.400 99.475 2755.475 ;
        RECT 87.120 2753.800 99.500 2755.400 ;
        RECT 95.265 2753.730 99.475 2753.800 ;
        RECT 89.265 2746.950 93.475 2747.025 ;
        RECT 87.120 2745.350 93.510 2746.950 ;
        RECT 89.265 2745.280 93.475 2745.350 ;
        RECT 95.310 2738.500 99.520 2738.575 ;
        RECT 87.120 2736.900 99.520 2738.500 ;
        RECT 95.310 2736.830 99.520 2736.900 ;
        RECT 3377.040 2707.240 3382.450 2712.730 ;
        RECT 3358.510 2699.150 3363.920 2704.640 ;
        RECT 3495.790 2692.780 3499.920 2692.840 ;
        RECT 3495.790 2691.180 3517.630 2692.780 ;
        RECT 3495.790 2691.125 3499.920 2691.180 ;
        RECT 3489.735 2689.280 3493.865 2689.355 ;
        RECT 3489.570 2687.680 3517.630 2689.280 ;
        RECT 3489.735 2687.640 3493.865 2687.680 ;
        RECT 3548.580 2673.990 3552.765 2674.075 ;
        RECT 3546.270 2672.390 3552.880 2673.990 ;
        RECT 3548.580 2672.300 3552.765 2672.390 ;
        RECT 3495.630 2668.750 3499.955 2668.850 ;
        RECT 3495.630 2667.150 3502.060 2668.750 ;
        RECT 3495.630 2667.080 3499.955 2667.150 ;
        RECT 3554.585 2665.540 3558.770 2665.620 ;
        RECT 3546.270 2663.940 3558.940 2665.540 ;
        RECT 3554.585 2663.845 3558.770 2663.940 ;
        RECT 3489.645 2660.300 3493.970 2660.360 ;
        RECT 3489.645 2658.700 3502.060 2660.300 ;
        RECT 3489.645 2658.590 3493.970 2658.700 ;
        RECT 3548.555 2657.090 3552.740 2657.205 ;
        RECT 3546.270 2655.490 3552.850 2657.090 ;
        RECT 3548.555 2655.430 3552.740 2655.490 ;
        RECT 3495.745 2651.850 3500.070 2651.935 ;
        RECT 3495.745 2650.250 3502.060 2651.850 ;
        RECT 3495.745 2650.165 3500.070 2650.250 ;
        RECT 3554.530 2648.640 3558.940 2648.750 ;
        RECT 3546.270 2647.140 3558.940 2648.640 ;
        RECT 3546.270 2647.060 3558.935 2647.140 ;
        RECT 3546.270 2647.040 3558.930 2647.060 ;
        RECT 3489.650 2643.400 3493.975 2643.460 ;
        RECT 3489.650 2641.800 3502.060 2643.400 ;
        RECT 3489.650 2641.690 3493.975 2641.800 ;
        RECT 3548.560 2640.190 3552.740 2640.280 ;
        RECT 3546.110 2638.590 3552.740 2640.190 ;
        RECT 3548.560 2638.480 3552.740 2638.590 ;
        RECT 3495.650 2634.950 3499.975 2635.055 ;
        RECT 3495.650 2633.350 3502.060 2634.950 ;
        RECT 3495.650 2633.285 3499.975 2633.350 ;
        RECT 3554.525 2631.740 3558.710 2631.820 ;
        RECT 3546.110 2630.140 3558.710 2631.740 ;
        RECT 3554.525 2630.045 3558.710 2630.140 ;
        RECT 3489.680 2626.500 3494.005 2626.600 ;
        RECT 3489.680 2624.900 3502.060 2626.500 ;
        RECT 3489.680 2624.830 3494.005 2624.900 ;
        RECT 3377.040 2487.240 3382.450 2492.730 ;
        RECT 3358.510 2479.150 3363.920 2484.640 ;
        RECT 3495.790 2472.780 3499.920 2472.840 ;
        RECT 3495.790 2471.180 3517.630 2472.780 ;
        RECT 3495.790 2471.125 3499.920 2471.180 ;
        RECT 3489.735 2469.280 3493.865 2469.355 ;
        RECT 3489.570 2467.680 3517.630 2469.280 ;
        RECT 3489.735 2467.640 3493.865 2467.680 ;
        RECT 3548.580 2453.990 3552.765 2454.075 ;
        RECT 3546.270 2452.390 3552.880 2453.990 ;
        RECT 3548.580 2452.300 3552.765 2452.390 ;
        RECT 3495.630 2448.750 3499.955 2448.850 ;
        RECT 3495.630 2447.150 3502.060 2448.750 ;
        RECT 3495.630 2447.080 3499.955 2447.150 ;
        RECT 3554.585 2445.540 3558.770 2445.620 ;
        RECT 3546.270 2443.940 3558.940 2445.540 ;
        RECT 3554.585 2443.845 3558.770 2443.940 ;
        RECT 3489.645 2440.300 3493.970 2440.360 ;
        RECT 3489.645 2438.700 3502.060 2440.300 ;
        RECT 3489.645 2438.590 3493.970 2438.700 ;
        RECT 3548.555 2437.090 3552.740 2437.205 ;
        RECT 3546.270 2435.490 3552.850 2437.090 ;
        RECT 3548.555 2435.430 3552.740 2435.490 ;
        RECT 3495.745 2431.850 3500.070 2431.935 ;
        RECT 3495.745 2430.250 3502.060 2431.850 ;
        RECT 3495.745 2430.165 3500.070 2430.250 ;
        RECT 3554.530 2428.640 3558.940 2428.750 ;
        RECT 3546.270 2427.140 3558.940 2428.640 ;
        RECT 3546.270 2427.060 3558.935 2427.140 ;
        RECT 3546.270 2427.040 3558.930 2427.060 ;
        RECT 3489.650 2423.400 3493.975 2423.460 ;
        RECT 3489.650 2421.800 3502.060 2423.400 ;
        RECT 3489.650 2421.690 3493.975 2421.800 ;
        RECT 3548.560 2420.190 3552.740 2420.280 ;
        RECT 3546.110 2418.590 3552.740 2420.190 ;
        RECT 3548.560 2418.480 3552.740 2418.590 ;
        RECT 3495.650 2414.950 3499.975 2415.055 ;
        RECT 3495.650 2413.350 3502.060 2414.950 ;
        RECT 3495.650 2413.285 3499.975 2413.350 ;
        RECT 3554.525 2411.740 3558.710 2411.820 ;
        RECT 3546.110 2410.140 3558.710 2411.740 ;
        RECT 3554.525 2410.045 3558.710 2410.140 ;
        RECT 3489.680 2406.500 3494.005 2406.600 ;
        RECT 3489.680 2404.900 3502.060 2406.500 ;
        RECT 3489.680 2404.830 3494.005 2404.900 ;
        RECT 221.390 2196.880 233.670 2202.150 ;
        RECT 205.340 2188.970 217.620 2194.240 ;
        RECT 89.230 2166.780 93.425 2166.895 ;
        RECT 71.550 2165.180 93.425 2166.780 ;
        RECT 89.230 2165.090 93.425 2165.180 ;
        RECT 95.260 2163.280 99.455 2163.350 ;
        RECT 71.550 2161.680 99.610 2163.280 ;
        RECT 95.260 2161.545 99.455 2161.680 ;
        RECT 89.245 2142.750 93.455 2142.840 ;
        RECT 87.120 2141.150 93.540 2142.750 ;
        RECT 89.245 2141.040 93.455 2141.150 ;
        RECT 95.280 2134.300 99.490 2134.365 ;
        RECT 87.120 2132.700 99.500 2134.300 ;
        RECT 95.280 2132.620 99.490 2132.700 ;
        RECT 89.285 2125.850 93.495 2125.890 ;
        RECT 87.120 2124.250 93.495 2125.850 ;
        RECT 89.285 2124.145 93.495 2124.250 ;
        RECT 95.265 2117.400 99.475 2117.475 ;
        RECT 87.120 2115.800 99.500 2117.400 ;
        RECT 95.265 2115.730 99.475 2115.800 ;
        RECT 89.265 2108.950 93.475 2109.025 ;
        RECT 87.120 2107.350 93.510 2108.950 ;
        RECT 89.265 2107.280 93.475 2107.350 ;
        RECT 95.310 2100.500 99.520 2100.575 ;
        RECT 87.120 2098.900 99.520 2100.500 ;
        RECT 95.310 2098.830 99.520 2098.900 ;
        RECT 3377.040 2046.240 3382.450 2051.730 ;
        RECT 3358.510 2038.150 3363.920 2043.640 ;
        RECT 3495.790 2031.780 3499.920 2031.840 ;
        RECT 3495.790 2030.180 3517.630 2031.780 ;
        RECT 3495.790 2030.125 3499.920 2030.180 ;
        RECT 3489.735 2028.280 3493.865 2028.355 ;
        RECT 3489.570 2026.680 3517.630 2028.280 ;
        RECT 3489.735 2026.640 3493.865 2026.680 ;
        RECT 3548.580 2012.990 3552.765 2013.075 ;
        RECT 3546.270 2011.390 3552.880 2012.990 ;
        RECT 3548.580 2011.300 3552.765 2011.390 ;
        RECT 3495.630 2007.750 3499.955 2007.850 ;
        RECT 3495.630 2006.150 3502.060 2007.750 ;
        RECT 3495.630 2006.080 3499.955 2006.150 ;
        RECT 3554.585 2004.540 3558.770 2004.620 ;
        RECT 3546.270 2002.940 3558.940 2004.540 ;
        RECT 3554.585 2002.845 3558.770 2002.940 ;
        RECT 3489.645 1999.300 3493.970 1999.360 ;
        RECT 3489.645 1997.700 3502.060 1999.300 ;
        RECT 3489.645 1997.590 3493.970 1997.700 ;
        RECT 3548.555 1996.090 3552.740 1996.205 ;
        RECT 3546.270 1994.490 3552.850 1996.090 ;
        RECT 3548.555 1994.430 3552.740 1994.490 ;
        RECT 3495.745 1990.850 3500.070 1990.935 ;
        RECT 3495.745 1989.250 3502.060 1990.850 ;
        RECT 3495.745 1989.165 3500.070 1989.250 ;
        RECT 3554.530 1987.640 3558.940 1987.750 ;
        RECT 221.390 1980.880 233.670 1986.150 ;
        RECT 3546.270 1986.140 3558.940 1987.640 ;
        RECT 3546.270 1986.060 3558.935 1986.140 ;
        RECT 3546.270 1986.040 3558.930 1986.060 ;
        RECT 3489.650 1982.400 3493.975 1982.460 ;
        RECT 3489.650 1980.800 3502.060 1982.400 ;
        RECT 3489.650 1980.690 3493.975 1980.800 ;
        RECT 3548.560 1979.190 3552.740 1979.280 ;
        RECT 205.340 1972.970 217.620 1978.240 ;
        RECT 3546.110 1977.590 3552.740 1979.190 ;
        RECT 3548.560 1977.480 3552.740 1977.590 ;
        RECT 3495.650 1973.950 3499.975 1974.055 ;
        RECT 3495.650 1972.350 3502.060 1973.950 ;
        RECT 3495.650 1972.285 3499.975 1972.350 ;
        RECT 3554.525 1970.740 3558.710 1970.820 ;
        RECT 3546.110 1969.140 3558.710 1970.740 ;
        RECT 3554.525 1969.045 3558.710 1969.140 ;
        RECT 3489.680 1965.500 3494.005 1965.600 ;
        RECT 3489.680 1963.900 3502.060 1965.500 ;
        RECT 3489.680 1963.830 3494.005 1963.900 ;
        RECT 89.230 1950.780 93.425 1950.895 ;
        RECT 71.550 1949.180 93.425 1950.780 ;
        RECT 89.230 1949.090 93.425 1949.180 ;
        RECT 95.260 1947.280 99.455 1947.350 ;
        RECT 71.550 1945.680 99.610 1947.280 ;
        RECT 95.260 1945.545 99.455 1945.680 ;
        RECT 89.245 1926.750 93.455 1926.840 ;
        RECT 87.120 1925.150 93.540 1926.750 ;
        RECT 89.245 1925.040 93.455 1925.150 ;
        RECT 95.280 1918.300 99.490 1918.365 ;
        RECT 87.120 1916.700 99.500 1918.300 ;
        RECT 95.280 1916.620 99.490 1916.700 ;
        RECT 89.285 1909.850 93.495 1909.890 ;
        RECT 87.120 1908.250 93.495 1909.850 ;
        RECT 89.285 1908.145 93.495 1908.250 ;
        RECT 95.265 1901.400 99.475 1901.475 ;
        RECT 87.120 1899.800 99.500 1901.400 ;
        RECT 95.265 1899.730 99.475 1899.800 ;
        RECT 89.265 1892.950 93.475 1893.025 ;
        RECT 87.120 1891.350 93.510 1892.950 ;
        RECT 89.265 1891.280 93.475 1891.350 ;
        RECT 95.310 1884.500 99.520 1884.575 ;
        RECT 87.120 1882.900 99.520 1884.500 ;
        RECT 95.310 1882.830 99.520 1882.900 ;
        RECT 3377.040 1820.240 3382.450 1825.730 ;
        RECT 3358.510 1812.150 3363.920 1817.640 ;
        RECT 3495.790 1805.780 3499.920 1805.840 ;
        RECT 3495.790 1804.180 3517.630 1805.780 ;
        RECT 3495.790 1804.125 3499.920 1804.180 ;
        RECT 3489.735 1802.280 3493.865 1802.355 ;
        RECT 3489.570 1800.680 3517.630 1802.280 ;
        RECT 3489.735 1800.640 3493.865 1800.680 ;
        RECT 3548.580 1786.990 3552.765 1787.075 ;
        RECT 3546.270 1785.390 3552.880 1786.990 ;
        RECT 3548.580 1785.300 3552.765 1785.390 ;
        RECT 3495.630 1781.750 3499.955 1781.850 ;
        RECT 3495.630 1780.150 3502.060 1781.750 ;
        RECT 3495.630 1780.080 3499.955 1780.150 ;
        RECT 3554.585 1778.540 3558.770 1778.620 ;
        RECT 3546.270 1776.940 3558.940 1778.540 ;
        RECT 3554.585 1776.845 3558.770 1776.940 ;
        RECT 221.390 1769.880 233.670 1775.150 ;
        RECT 3489.645 1773.300 3493.970 1773.360 ;
        RECT 3489.645 1771.700 3502.060 1773.300 ;
        RECT 3489.645 1771.590 3493.970 1771.700 ;
        RECT 3548.555 1770.090 3552.740 1770.205 ;
        RECT 3546.270 1768.490 3552.850 1770.090 ;
        RECT 3548.555 1768.430 3552.740 1768.490 ;
        RECT 205.340 1761.970 217.620 1767.240 ;
        RECT 3495.745 1764.850 3500.070 1764.935 ;
        RECT 3495.745 1763.250 3502.060 1764.850 ;
        RECT 3495.745 1763.165 3500.070 1763.250 ;
        RECT 3554.530 1761.640 3558.940 1761.750 ;
        RECT 3546.270 1760.140 3558.940 1761.640 ;
        RECT 3546.270 1760.060 3558.935 1760.140 ;
        RECT 3546.270 1760.040 3558.930 1760.060 ;
        RECT 3489.650 1756.400 3493.975 1756.460 ;
        RECT 3489.650 1754.800 3502.060 1756.400 ;
        RECT 3489.650 1754.690 3493.975 1754.800 ;
        RECT 3548.560 1753.190 3552.740 1753.280 ;
        RECT 3546.110 1751.590 3552.740 1753.190 ;
        RECT 3548.560 1751.480 3552.740 1751.590 ;
        RECT 3495.650 1747.950 3499.975 1748.055 ;
        RECT 3495.650 1746.350 3502.060 1747.950 ;
        RECT 3495.650 1746.285 3499.975 1746.350 ;
        RECT 3554.525 1744.740 3558.710 1744.820 ;
        RECT 3546.110 1743.140 3558.710 1744.740 ;
        RECT 3554.525 1743.045 3558.710 1743.140 ;
        RECT 3489.680 1739.500 3494.005 1739.600 ;
        RECT 3489.680 1737.900 3502.060 1739.500 ;
        RECT 3489.680 1737.830 3494.005 1737.900 ;
        RECT 89.230 1734.780 93.425 1734.895 ;
        RECT 71.550 1733.180 93.425 1734.780 ;
        RECT 89.230 1733.090 93.425 1733.180 ;
        RECT 95.260 1731.280 99.455 1731.350 ;
        RECT 71.550 1729.680 99.610 1731.280 ;
        RECT 95.260 1729.545 99.455 1729.680 ;
        RECT 89.245 1710.750 93.455 1710.840 ;
        RECT 87.120 1709.150 93.540 1710.750 ;
        RECT 89.245 1709.040 93.455 1709.150 ;
        RECT 95.280 1702.300 99.490 1702.365 ;
        RECT 87.120 1700.700 99.500 1702.300 ;
        RECT 95.280 1700.620 99.490 1700.700 ;
        RECT 89.285 1693.850 93.495 1693.890 ;
        RECT 87.120 1692.250 93.495 1693.850 ;
        RECT 89.285 1692.145 93.495 1692.250 ;
        RECT 95.265 1685.400 99.475 1685.475 ;
        RECT 87.120 1683.800 99.500 1685.400 ;
        RECT 95.265 1683.730 99.475 1683.800 ;
        RECT 89.265 1676.950 93.475 1677.025 ;
        RECT 87.120 1675.350 93.510 1676.950 ;
        RECT 89.265 1675.280 93.475 1675.350 ;
        RECT 95.310 1668.500 99.520 1668.575 ;
        RECT 87.120 1666.900 99.520 1668.500 ;
        RECT 95.310 1666.830 99.520 1666.900 ;
        RECT 3377.040 1595.240 3382.450 1600.730 ;
        RECT 3358.510 1587.150 3363.920 1592.640 ;
        RECT 3495.790 1580.780 3499.920 1580.840 ;
        RECT 3495.790 1579.180 3517.630 1580.780 ;
        RECT 3495.790 1579.125 3499.920 1579.180 ;
        RECT 3489.735 1577.280 3493.865 1577.355 ;
        RECT 3489.570 1575.680 3517.630 1577.280 ;
        RECT 3489.735 1575.640 3493.865 1575.680 ;
        RECT 3548.580 1561.990 3552.765 1562.075 ;
        RECT 3546.270 1560.390 3552.880 1561.990 ;
        RECT 3548.580 1560.300 3552.765 1560.390 ;
        RECT 3495.630 1556.750 3499.955 1556.850 ;
        RECT 3495.630 1555.150 3502.060 1556.750 ;
        RECT 3495.630 1555.080 3499.955 1555.150 ;
        RECT 221.390 1548.880 233.670 1554.150 ;
        RECT 3554.585 1553.540 3558.770 1553.620 ;
        RECT 3546.270 1551.940 3558.940 1553.540 ;
        RECT 3554.585 1551.845 3558.770 1551.940 ;
        RECT 3489.645 1548.300 3493.970 1548.360 ;
        RECT 3489.645 1546.700 3502.060 1548.300 ;
        RECT 3489.645 1546.590 3493.970 1546.700 ;
        RECT 205.340 1540.970 217.620 1546.240 ;
        RECT 3548.555 1545.090 3552.740 1545.205 ;
        RECT 3546.270 1543.490 3552.850 1545.090 ;
        RECT 3548.555 1543.430 3552.740 1543.490 ;
        RECT 3495.745 1539.850 3500.070 1539.935 ;
        RECT 3495.745 1538.250 3502.060 1539.850 ;
        RECT 3495.745 1538.165 3500.070 1538.250 ;
        RECT 3554.530 1536.640 3558.940 1536.750 ;
        RECT 3546.270 1535.140 3558.940 1536.640 ;
        RECT 3546.270 1535.060 3558.935 1535.140 ;
        RECT 3546.270 1535.040 3558.930 1535.060 ;
        RECT 3489.650 1531.400 3493.975 1531.460 ;
        RECT 3489.650 1529.800 3502.060 1531.400 ;
        RECT 3489.650 1529.690 3493.975 1529.800 ;
        RECT 3548.560 1528.190 3552.740 1528.280 ;
        RECT 3546.110 1526.590 3552.740 1528.190 ;
        RECT 3548.560 1526.480 3552.740 1526.590 ;
        RECT 3495.650 1522.950 3499.975 1523.055 ;
        RECT 3495.650 1521.350 3502.060 1522.950 ;
        RECT 3495.650 1521.285 3499.975 1521.350 ;
        RECT 3554.525 1519.740 3558.710 1519.820 ;
        RECT 89.230 1518.780 93.425 1518.895 ;
        RECT 71.550 1517.180 93.425 1518.780 ;
        RECT 3546.110 1518.140 3558.710 1519.740 ;
        RECT 3554.525 1518.045 3558.710 1518.140 ;
        RECT 89.230 1517.090 93.425 1517.180 ;
        RECT 95.260 1515.280 99.455 1515.350 ;
        RECT 71.550 1513.680 99.610 1515.280 ;
        RECT 3489.680 1514.500 3494.005 1514.600 ;
        RECT 95.260 1513.545 99.455 1513.680 ;
        RECT 3489.680 1512.900 3502.060 1514.500 ;
        RECT 3489.680 1512.830 3494.005 1512.900 ;
        RECT 89.245 1494.750 93.455 1494.840 ;
        RECT 87.120 1493.150 93.540 1494.750 ;
        RECT 89.245 1493.040 93.455 1493.150 ;
        RECT 95.280 1486.300 99.490 1486.365 ;
        RECT 87.120 1484.700 99.500 1486.300 ;
        RECT 95.280 1484.620 99.490 1484.700 ;
        RECT 89.285 1477.850 93.495 1477.890 ;
        RECT 87.120 1476.250 93.495 1477.850 ;
        RECT 89.285 1476.145 93.495 1476.250 ;
        RECT 95.265 1469.400 99.475 1469.475 ;
        RECT 87.120 1467.800 99.500 1469.400 ;
        RECT 95.265 1467.730 99.475 1467.800 ;
        RECT 89.265 1460.950 93.475 1461.025 ;
        RECT 87.120 1459.350 93.510 1460.950 ;
        RECT 89.265 1459.280 93.475 1459.350 ;
        RECT 95.310 1452.500 99.520 1452.575 ;
        RECT 87.120 1450.900 99.520 1452.500 ;
        RECT 95.310 1450.830 99.520 1450.900 ;
        RECT 3256.130 1388.920 3315.790 1392.020 ;
        RECT 221.140 1379.440 233.810 1386.310 ;
        RECT 3260.940 1384.120 3315.790 1387.220 ;
        RECT 278.770 1379.320 306.940 1382.420 ;
        RECT 3354.420 1380.370 3366.820 1387.050 ;
        RECT 3370.420 1384.100 3382.820 1391.780 ;
        RECT 214.150 1346.890 217.640 1377.290 ;
        RECT 278.770 1374.520 302.140 1377.620 ;
        RECT 3377.040 1370.240 3382.450 1375.730 ;
        RECT 3358.510 1362.150 3363.920 1367.640 ;
        RECT 3495.790 1355.780 3499.920 1355.840 ;
        RECT 3495.790 1354.180 3517.630 1355.780 ;
        RECT 3495.790 1354.125 3499.920 1354.180 ;
        RECT 3489.735 1352.280 3493.865 1352.355 ;
        RECT 3489.570 1350.680 3517.630 1352.280 ;
        RECT 3489.735 1350.640 3493.865 1350.680 ;
        RECT 3548.580 1336.990 3552.765 1337.075 ;
        RECT 3546.270 1335.390 3552.880 1336.990 ;
        RECT 3548.580 1335.300 3552.765 1335.390 ;
        RECT 3495.630 1331.750 3499.955 1331.850 ;
        RECT 3495.630 1330.150 3502.060 1331.750 ;
        RECT 3495.630 1330.080 3499.955 1330.150 ;
        RECT 3554.585 1328.540 3558.770 1328.620 ;
        RECT 3546.270 1326.940 3558.940 1328.540 ;
        RECT 3554.585 1326.845 3558.770 1326.940 ;
        RECT 3489.645 1323.300 3493.970 1323.360 ;
        RECT 3489.645 1321.700 3502.060 1323.300 ;
        RECT 3489.645 1321.590 3493.970 1321.700 ;
        RECT 3548.555 1320.090 3552.740 1320.205 ;
        RECT 3546.270 1318.490 3552.850 1320.090 ;
        RECT 3548.555 1318.430 3552.740 1318.490 ;
        RECT 3495.745 1314.850 3500.070 1314.935 ;
        RECT 3495.745 1313.250 3502.060 1314.850 ;
        RECT 3495.745 1313.165 3500.070 1313.250 ;
        RECT 3554.530 1311.640 3558.940 1311.750 ;
        RECT 3546.270 1310.140 3558.940 1311.640 ;
        RECT 3546.270 1310.060 3558.935 1310.140 ;
        RECT 3546.270 1310.040 3558.930 1310.060 ;
        RECT 3489.650 1306.400 3493.975 1306.460 ;
        RECT 3489.650 1304.800 3502.060 1306.400 ;
        RECT 3489.650 1304.690 3493.975 1304.800 ;
        RECT 3548.560 1303.190 3552.740 1303.280 ;
        RECT 89.230 1302.780 93.425 1302.895 ;
        RECT 71.550 1301.180 93.425 1302.780 ;
        RECT 3546.110 1301.590 3552.740 1303.190 ;
        RECT 3548.560 1301.480 3552.740 1301.590 ;
        RECT 89.230 1301.090 93.425 1301.180 ;
        RECT 95.260 1299.280 99.455 1299.350 ;
        RECT 71.550 1297.680 99.610 1299.280 ;
        RECT 3495.650 1297.950 3499.975 1298.055 ;
        RECT 95.260 1297.545 99.455 1297.680 ;
        RECT 3495.650 1296.350 3502.060 1297.950 ;
        RECT 3495.650 1296.285 3499.975 1296.350 ;
        RECT 3554.525 1294.740 3558.710 1294.820 ;
        RECT 3546.110 1293.140 3558.710 1294.740 ;
        RECT 3554.525 1293.045 3558.710 1293.140 ;
        RECT 3489.680 1289.500 3494.005 1289.600 ;
        RECT 3489.680 1287.900 3502.060 1289.500 ;
        RECT 3489.680 1287.830 3494.005 1287.900 ;
        RECT 89.245 1278.750 93.455 1278.840 ;
        RECT 87.120 1277.150 93.540 1278.750 ;
        RECT 89.245 1277.040 93.455 1277.150 ;
        RECT 95.280 1270.300 99.490 1270.365 ;
        RECT 87.120 1268.700 99.500 1270.300 ;
        RECT 95.280 1268.620 99.490 1268.700 ;
        RECT 89.285 1261.850 93.495 1261.890 ;
        RECT 87.120 1260.250 93.495 1261.850 ;
        RECT 89.285 1260.145 93.495 1260.250 ;
        RECT 95.265 1253.400 99.475 1253.475 ;
        RECT 87.120 1251.800 99.500 1253.400 ;
        RECT 95.265 1251.730 99.475 1251.800 ;
        RECT 89.265 1244.950 93.475 1245.025 ;
        RECT 87.120 1243.350 93.510 1244.950 ;
        RECT 89.265 1243.280 93.475 1243.350 ;
        RECT 95.310 1236.500 99.520 1236.575 ;
        RECT 87.120 1234.900 99.520 1236.500 ;
        RECT 95.310 1234.830 99.520 1234.900 ;
        RECT 3377.040 1144.240 3382.450 1149.730 ;
        RECT 3358.510 1136.150 3363.920 1141.640 ;
        RECT 3495.790 1129.780 3499.920 1129.840 ;
        RECT 3495.790 1128.180 3517.630 1129.780 ;
        RECT 3495.790 1128.125 3499.920 1128.180 ;
        RECT 3489.735 1126.280 3493.865 1126.355 ;
        RECT 3489.570 1124.680 3517.630 1126.280 ;
        RECT 3489.735 1124.640 3493.865 1124.680 ;
        RECT 3548.580 1110.990 3552.765 1111.075 ;
        RECT 3546.270 1109.390 3552.880 1110.990 ;
        RECT 3548.580 1109.300 3552.765 1109.390 ;
        RECT 3495.630 1105.750 3499.955 1105.850 ;
        RECT 3495.630 1104.150 3502.060 1105.750 ;
        RECT 3495.630 1104.080 3499.955 1104.150 ;
        RECT 3554.585 1102.540 3558.770 1102.620 ;
        RECT 3546.270 1100.940 3558.940 1102.540 ;
        RECT 3554.585 1100.845 3558.770 1100.940 ;
        RECT 3489.645 1097.300 3493.970 1097.360 ;
        RECT 3489.645 1095.700 3502.060 1097.300 ;
        RECT 3489.645 1095.590 3493.970 1095.700 ;
        RECT 3548.555 1094.090 3552.740 1094.205 ;
        RECT 3546.270 1092.490 3552.850 1094.090 ;
        RECT 3548.555 1092.430 3552.740 1092.490 ;
        RECT 3495.745 1088.850 3500.070 1088.935 ;
        RECT 3495.745 1087.250 3502.060 1088.850 ;
        RECT 3495.745 1087.165 3500.070 1087.250 ;
        RECT 89.230 1086.780 93.425 1086.895 ;
        RECT 71.550 1085.180 93.425 1086.780 ;
        RECT 3554.530 1085.640 3558.940 1085.750 ;
        RECT 89.230 1085.090 93.425 1085.180 ;
        RECT 3546.270 1084.140 3558.940 1085.640 ;
        RECT 3546.270 1084.060 3558.935 1084.140 ;
        RECT 3546.270 1084.040 3558.930 1084.060 ;
        RECT 95.260 1083.280 99.455 1083.350 ;
        RECT 71.550 1081.680 99.610 1083.280 ;
        RECT 95.260 1081.545 99.455 1081.680 ;
        RECT 3489.650 1080.400 3493.975 1080.460 ;
        RECT 3489.650 1078.800 3502.060 1080.400 ;
        RECT 3489.650 1078.690 3493.975 1078.800 ;
        RECT 3548.560 1077.190 3552.740 1077.280 ;
        RECT 3546.110 1075.590 3552.740 1077.190 ;
        RECT 3548.560 1075.480 3552.740 1075.590 ;
        RECT 3495.650 1071.950 3499.975 1072.055 ;
        RECT 3495.650 1070.350 3502.060 1071.950 ;
        RECT 3495.650 1070.285 3499.975 1070.350 ;
        RECT 3554.525 1068.740 3558.710 1068.820 ;
        RECT 3546.110 1067.140 3558.710 1068.740 ;
        RECT 3554.525 1067.045 3558.710 1067.140 ;
        RECT 3489.680 1063.500 3494.005 1063.600 ;
        RECT 89.245 1062.750 93.455 1062.840 ;
        RECT 87.120 1061.150 93.540 1062.750 ;
        RECT 3489.680 1061.900 3502.060 1063.500 ;
        RECT 3489.680 1061.830 3494.005 1061.900 ;
        RECT 89.245 1061.040 93.455 1061.150 ;
        RECT 95.280 1054.300 99.490 1054.365 ;
        RECT 87.120 1052.700 99.500 1054.300 ;
        RECT 95.280 1052.620 99.490 1052.700 ;
        RECT 89.285 1045.850 93.495 1045.890 ;
        RECT 87.120 1044.250 93.495 1045.850 ;
        RECT 89.285 1044.145 93.495 1044.250 ;
        RECT 95.265 1037.400 99.475 1037.475 ;
        RECT 87.120 1035.800 99.500 1037.400 ;
        RECT 95.265 1035.730 99.475 1035.800 ;
        RECT 89.265 1028.950 93.475 1029.025 ;
        RECT 87.120 1027.350 93.510 1028.950 ;
        RECT 89.265 1027.280 93.475 1027.350 ;
        RECT 95.310 1020.500 99.520 1020.575 ;
        RECT 87.120 1018.900 99.520 1020.500 ;
        RECT 95.310 1018.830 99.520 1018.900 ;
        RECT 3377.040 919.240 3382.450 924.730 ;
        RECT 3358.510 911.150 3363.920 916.640 ;
        RECT 3495.790 904.780 3499.920 904.840 ;
        RECT 3495.790 903.180 3517.630 904.780 ;
        RECT 3495.790 903.125 3499.920 903.180 ;
        RECT 3489.735 901.280 3493.865 901.355 ;
        RECT 3489.570 899.680 3517.630 901.280 ;
        RECT 3489.735 899.640 3493.865 899.680 ;
        RECT 3548.580 885.990 3552.765 886.075 ;
        RECT 3546.270 884.390 3552.880 885.990 ;
        RECT 3548.580 884.300 3552.765 884.390 ;
        RECT 3495.630 880.750 3499.955 880.850 ;
        RECT 3495.630 879.150 3502.060 880.750 ;
        RECT 3495.630 879.080 3499.955 879.150 ;
        RECT 3554.585 877.540 3558.770 877.620 ;
        RECT 3546.270 875.940 3558.940 877.540 ;
        RECT 3554.585 875.845 3558.770 875.940 ;
        RECT 3489.645 872.300 3493.970 872.360 ;
        RECT 3489.645 870.700 3502.060 872.300 ;
        RECT 3489.645 870.590 3493.970 870.700 ;
        RECT 3548.555 869.090 3552.740 869.205 ;
        RECT 3546.270 867.490 3552.850 869.090 ;
        RECT 3548.555 867.430 3552.740 867.490 ;
        RECT 3495.745 863.850 3500.070 863.935 ;
        RECT 3495.745 862.250 3502.060 863.850 ;
        RECT 3495.745 862.165 3500.070 862.250 ;
        RECT 3554.530 860.640 3558.940 860.750 ;
        RECT 3546.270 859.140 3558.940 860.640 ;
        RECT 3546.270 859.060 3558.935 859.140 ;
        RECT 3546.270 859.040 3558.930 859.060 ;
        RECT 3489.650 855.400 3493.975 855.460 ;
        RECT 3489.650 853.800 3502.060 855.400 ;
        RECT 3489.650 853.690 3493.975 853.800 ;
        RECT 3548.560 852.190 3552.740 852.280 ;
        RECT 3546.110 850.590 3552.740 852.190 ;
        RECT 3548.560 850.480 3552.740 850.590 ;
        RECT 3495.650 846.950 3499.975 847.055 ;
        RECT 3495.650 845.350 3502.060 846.950 ;
        RECT 3495.650 845.285 3499.975 845.350 ;
        RECT 3554.525 843.740 3558.710 843.820 ;
        RECT 3546.110 842.140 3558.710 843.740 ;
        RECT 3554.525 842.045 3558.710 842.140 ;
        RECT 3489.680 838.500 3494.005 838.600 ;
        RECT 3489.680 836.900 3502.060 838.500 ;
        RECT 3489.680 836.830 3494.005 836.900 ;
        RECT 3377.040 693.240 3382.450 698.730 ;
        RECT 3358.510 685.150 3363.920 690.640 ;
        RECT 3495.790 678.780 3499.920 678.840 ;
        RECT 3495.790 677.180 3517.630 678.780 ;
        RECT 3495.790 677.125 3499.920 677.180 ;
        RECT 3489.735 675.280 3493.865 675.355 ;
        RECT 3489.570 673.680 3517.630 675.280 ;
        RECT 3489.735 673.640 3493.865 673.680 ;
        RECT 3548.580 659.990 3552.765 660.075 ;
        RECT 3546.270 658.390 3552.880 659.990 ;
        RECT 3548.580 658.300 3552.765 658.390 ;
        RECT 3495.630 654.750 3499.955 654.850 ;
        RECT 3495.630 653.150 3502.060 654.750 ;
        RECT 3495.630 653.080 3499.955 653.150 ;
        RECT 3554.585 651.540 3558.770 651.620 ;
        RECT 3546.270 649.940 3558.940 651.540 ;
        RECT 3554.585 649.845 3558.770 649.940 ;
        RECT 3489.645 646.300 3493.970 646.360 ;
        RECT 3489.645 644.700 3502.060 646.300 ;
        RECT 3489.645 644.590 3493.970 644.700 ;
        RECT 3548.555 643.090 3552.740 643.205 ;
        RECT 3546.270 641.490 3552.850 643.090 ;
        RECT 3548.555 641.430 3552.740 641.490 ;
        RECT 3495.745 637.850 3500.070 637.935 ;
        RECT 3495.745 636.250 3502.060 637.850 ;
        RECT 3495.745 636.165 3500.070 636.250 ;
        RECT 3554.530 634.640 3558.940 634.750 ;
        RECT 3546.270 633.140 3558.940 634.640 ;
        RECT 3546.270 633.060 3558.935 633.140 ;
        RECT 3546.270 633.040 3558.930 633.060 ;
        RECT 3489.650 629.400 3493.975 629.460 ;
        RECT 3489.650 627.800 3502.060 629.400 ;
        RECT 3489.650 627.690 3493.975 627.800 ;
        RECT 3548.560 626.190 3552.740 626.280 ;
        RECT 3546.110 624.590 3552.740 626.190 ;
        RECT 3548.560 624.480 3552.740 624.590 ;
        RECT 3495.650 620.950 3499.975 621.055 ;
        RECT 3495.650 619.350 3502.060 620.950 ;
        RECT 3495.650 619.285 3499.975 619.350 ;
        RECT 3554.525 617.740 3558.710 617.820 ;
        RECT 3546.110 616.140 3558.710 617.740 ;
        RECT 3554.525 616.045 3558.710 616.140 ;
        RECT 3489.680 612.500 3494.005 612.600 ;
        RECT 3489.680 610.900 3502.060 612.500 ;
        RECT 3489.680 610.830 3494.005 610.900 ;
        RECT 643.050 206.310 718.230 208.000 ;
        RECT 650.710 202.910 724.725 204.610 ;
  END
END caravel_power_routing
END LIBRARY

